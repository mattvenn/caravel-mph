VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2183.690 89.660 2184.010 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2183.690 89.520 2899.310 89.660 ;
        RECT 2183.690 89.460 2184.010 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2183.720 89.460 2183.980 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2183.710 601.955 2183.990 602.325 ;
        RECT 2183.780 89.750 2183.920 601.955 ;
        RECT 2183.720 89.430 2183.980 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2183.710 602.000 2183.990 602.280 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2166.000 604.800 2170.000 605.400 ;
        RECT 2169.670 602.290 2169.970 604.800 ;
        RECT 2183.685 602.290 2184.015 602.305 ;
        RECT 2169.670 601.990 2184.015 602.290 ;
        RECT 2183.685 601.975 2184.015 601.990 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2191.050 2429.200 2191.370 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 2191.050 2429.060 2901.150 2429.200 ;
        RECT 2191.050 2429.000 2191.370 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 2180.470 710.500 2180.790 710.560 ;
        RECT 2191.050 710.500 2191.370 710.560 ;
        RECT 2180.470 710.360 2191.370 710.500 ;
        RECT 2180.470 710.300 2180.790 710.360 ;
        RECT 2191.050 710.300 2191.370 710.360 ;
      LAYER via ;
        RECT 2191.080 2429.000 2191.340 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 2180.500 710.300 2180.760 710.560 ;
        RECT 2191.080 710.300 2191.340 710.560 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 2191.080 2428.970 2191.340 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 2191.140 710.590 2191.280 2428.970 ;
        RECT 2180.500 710.445 2180.760 710.590 ;
        RECT 2180.490 710.075 2180.770 710.445 ;
        RECT 2191.080 710.270 2191.340 710.590 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 2180.490 710.120 2180.770 710.400 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2180.465 710.410 2180.795 710.425 ;
        RECT 2169.670 710.120 2180.795 710.410 ;
        RECT 2166.000 710.110 2180.795 710.120 ;
        RECT 2166.000 709.520 2170.000 710.110 ;
        RECT 2180.465 710.095 2180.795 710.110 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2570.090 2663.800 2570.410 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 2570.090 2663.660 2901.150 2663.800 ;
        RECT 2570.090 2663.600 2570.410 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 2185.070 724.440 2185.390 724.500 ;
        RECT 2570.090 724.440 2570.410 724.500 ;
        RECT 2185.070 724.300 2570.410 724.440 ;
        RECT 2185.070 724.240 2185.390 724.300 ;
        RECT 2570.090 724.240 2570.410 724.300 ;
      LAYER via ;
        RECT 2570.120 2663.600 2570.380 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 2185.100 724.240 2185.360 724.500 ;
        RECT 2570.120 724.240 2570.380 724.500 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 2570.120 2663.570 2570.380 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 2570.180 724.530 2570.320 2663.570 ;
        RECT 2185.100 724.210 2185.360 724.530 ;
        RECT 2570.120 724.210 2570.380 724.530 ;
        RECT 2185.160 722.685 2185.300 724.210 ;
        RECT 2185.090 722.315 2185.370 722.685 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
        RECT 2185.090 722.360 2185.370 722.640 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2185.065 722.650 2185.395 722.665 ;
        RECT 2169.670 722.350 2185.395 722.650 ;
        RECT 2169.670 721.000 2169.970 722.350 ;
        RECT 2185.065 722.335 2185.395 722.350 ;
        RECT 2166.000 720.400 2170.000 721.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2211.290 2898.400 2211.610 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2211.290 2898.260 2901.150 2898.400 ;
        RECT 2211.290 2898.200 2211.610 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2186.910 730.900 2187.230 730.960 ;
        RECT 2211.290 730.900 2211.610 730.960 ;
        RECT 2186.910 730.760 2211.610 730.900 ;
        RECT 2186.910 730.700 2187.230 730.760 ;
        RECT 2211.290 730.700 2211.610 730.760 ;
      LAYER via ;
        RECT 2211.320 2898.200 2211.580 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2186.940 730.700 2187.200 730.960 ;
        RECT 2211.320 730.700 2211.580 730.960 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2211.320 2898.170 2211.580 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2186.930 731.155 2187.210 731.525 ;
        RECT 2187.000 730.990 2187.140 731.155 ;
        RECT 2211.380 730.990 2211.520 2898.170 ;
        RECT 2186.940 730.670 2187.200 730.990 ;
        RECT 2211.320 730.670 2211.580 730.990 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 2186.930 731.200 2187.210 731.480 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2186.905 731.490 2187.235 731.505 ;
        RECT 2169.670 731.200 2187.235 731.490 ;
        RECT 2166.000 731.190 2187.235 731.200 ;
        RECT 2166.000 730.600 2170.000 731.190 ;
        RECT 2186.905 731.175 2187.235 731.190 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2225.090 3133.000 2225.410 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2225.090 3132.860 2901.150 3133.000 ;
        RECT 2225.090 3132.800 2225.410 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 2180.470 745.180 2180.790 745.240 ;
        RECT 2225.090 745.180 2225.410 745.240 ;
        RECT 2180.470 745.040 2225.410 745.180 ;
        RECT 2180.470 744.980 2180.790 745.040 ;
        RECT 2225.090 744.980 2225.410 745.040 ;
      LAYER via ;
        RECT 2225.120 3132.800 2225.380 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 2180.500 744.980 2180.760 745.240 ;
        RECT 2225.120 744.980 2225.380 745.240 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2225.120 3132.770 2225.380 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 2225.180 745.270 2225.320 3132.770 ;
        RECT 2180.500 744.950 2180.760 745.270 ;
        RECT 2225.120 744.950 2225.380 745.270 ;
        RECT 2180.560 743.765 2180.700 744.950 ;
        RECT 2180.490 743.395 2180.770 743.765 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 2180.490 743.440 2180.770 743.720 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2180.465 743.730 2180.795 743.745 ;
        RECT 2169.670 743.430 2180.795 743.730 ;
        RECT 2169.670 742.080 2169.970 743.430 ;
        RECT 2180.465 743.415 2180.795 743.430 ;
        RECT 2166.000 741.480 2170.000 742.080 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2231.990 3367.600 2232.310 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2231.990 3367.460 2901.150 3367.600 ;
        RECT 2231.990 3367.400 2232.310 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 2186.910 751.980 2187.230 752.040 ;
        RECT 2231.990 751.980 2232.310 752.040 ;
        RECT 2186.910 751.840 2232.310 751.980 ;
        RECT 2186.910 751.780 2187.230 751.840 ;
        RECT 2231.990 751.780 2232.310 751.840 ;
      LAYER via ;
        RECT 2232.020 3367.400 2232.280 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 2186.940 751.780 2187.200 752.040 ;
        RECT 2232.020 751.780 2232.280 752.040 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2232.020 3367.370 2232.280 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 2232.080 752.070 2232.220 3367.370 ;
        RECT 2186.940 751.750 2187.200 752.070 ;
        RECT 2232.020 751.750 2232.280 752.070 ;
        RECT 2187.000 751.245 2187.140 751.750 ;
        RECT 2186.930 750.875 2187.210 751.245 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 2186.930 750.920 2187.210 751.200 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2166.000 751.680 2170.000 752.280 ;
        RECT 2169.670 751.210 2169.970 751.680 ;
        RECT 2186.905 751.210 2187.235 751.225 ;
        RECT 2169.670 750.910 2187.235 751.210 ;
        RECT 2186.905 750.895 2187.235 750.910 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2238.890 3501.560 2239.210 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 2238.890 3501.420 2798.570 3501.560 ;
        RECT 2238.890 3501.360 2239.210 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
        RECT 2186.910 765.920 2187.230 765.980 ;
        RECT 2238.890 765.920 2239.210 765.980 ;
        RECT 2186.910 765.780 2239.210 765.920 ;
        RECT 2186.910 765.720 2187.230 765.780 ;
        RECT 2238.890 765.720 2239.210 765.780 ;
      LAYER via ;
        RECT 2238.920 3501.360 2239.180 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
        RECT 2186.940 765.720 2187.200 765.980 ;
        RECT 2238.920 765.720 2239.180 765.980 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 2238.920 3501.330 2239.180 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 2238.980 766.010 2239.120 3501.330 ;
        RECT 2186.940 765.690 2187.200 766.010 ;
        RECT 2238.920 765.690 2239.180 766.010 ;
        RECT 2187.000 764.165 2187.140 765.690 ;
        RECT 2186.930 763.795 2187.210 764.165 ;
      LAYER via2 ;
        RECT 2186.930 763.840 2187.210 764.120 ;
      LAYER met3 ;
        RECT 2186.905 764.130 2187.235 764.145 ;
        RECT 2169.670 763.830 2187.235 764.130 ;
        RECT 2169.670 763.160 2169.970 763.830 ;
        RECT 2186.905 763.815 2187.235 763.830 ;
        RECT 2166.000 762.560 2170.000 763.160 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2190.590 3502.240 2190.910 3502.300 ;
        RECT 2473.950 3502.240 2474.270 3502.300 ;
        RECT 2190.590 3502.100 2474.270 3502.240 ;
        RECT 2190.590 3502.040 2190.910 3502.100 ;
        RECT 2473.950 3502.040 2474.270 3502.100 ;
        RECT 2180.470 776.120 2180.790 776.180 ;
        RECT 2190.590 776.120 2190.910 776.180 ;
        RECT 2180.470 775.980 2190.910 776.120 ;
        RECT 2180.470 775.920 2180.790 775.980 ;
        RECT 2190.590 775.920 2190.910 775.980 ;
      LAYER via ;
        RECT 2190.620 3502.040 2190.880 3502.300 ;
        RECT 2473.980 3502.040 2474.240 3502.300 ;
        RECT 2180.500 775.920 2180.760 776.180 ;
        RECT 2190.620 775.920 2190.880 776.180 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3502.330 2474.180 3517.600 ;
        RECT 2190.620 3502.010 2190.880 3502.330 ;
        RECT 2473.980 3502.010 2474.240 3502.330 ;
        RECT 2190.680 776.210 2190.820 3502.010 ;
        RECT 2180.500 775.890 2180.760 776.210 ;
        RECT 2190.620 775.890 2190.880 776.210 ;
        RECT 2180.560 775.725 2180.700 775.890 ;
        RECT 2180.490 775.355 2180.770 775.725 ;
      LAYER via2 ;
        RECT 2180.490 775.400 2180.770 775.680 ;
      LAYER met3 ;
        RECT 2180.465 775.690 2180.795 775.705 ;
        RECT 2169.670 775.390 2180.795 775.690 ;
        RECT 2169.670 773.360 2169.970 775.390 ;
        RECT 2180.465 775.375 2180.795 775.390 ;
        RECT 2166.000 772.760 2170.000 773.360 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2149.190 3498.500 2149.510 3498.560 ;
        RECT 2169.430 3498.500 2169.750 3498.560 ;
        RECT 2149.190 3498.360 2169.750 3498.500 ;
        RECT 2149.190 3498.300 2149.510 3498.360 ;
        RECT 2169.430 3498.300 2169.750 3498.360 ;
      LAYER via ;
        RECT 2149.220 3498.300 2149.480 3498.560 ;
        RECT 2169.460 3498.300 2169.720 3498.560 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3498.590 2149.420 3517.600 ;
        RECT 2149.220 3498.270 2149.480 3498.590 ;
        RECT 2169.460 3498.270 2169.720 3498.590 ;
        RECT 2169.520 786.605 2169.660 3498.270 ;
        RECT 2169.450 786.235 2169.730 786.605 ;
      LAYER via2 ;
        RECT 2169.450 786.280 2169.730 786.560 ;
      LAYER met3 ;
        RECT 2169.425 786.570 2169.755 786.585 ;
        RECT 2169.425 786.255 2169.970 786.570 ;
        RECT 2169.670 784.240 2169.970 786.255 ;
        RECT 2166.000 783.640 2170.000 784.240 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3503.600 1825.210 3503.660 ;
        RECT 2169.890 3503.600 2170.210 3503.660 ;
        RECT 1824.890 3503.460 2170.210 3503.600 ;
        RECT 1824.890 3503.400 1825.210 3503.460 ;
        RECT 2169.890 3503.400 2170.210 3503.460 ;
      LAYER via ;
        RECT 1824.920 3503.400 1825.180 3503.660 ;
        RECT 2169.920 3503.400 2170.180 3503.660 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3503.690 1825.120 3517.600 ;
        RECT 1824.920 3503.370 1825.180 3503.690 ;
        RECT 2169.920 3503.370 2170.180 3503.690 ;
        RECT 2169.980 796.805 2170.120 3503.370 ;
        RECT 2169.910 796.435 2170.190 796.805 ;
      LAYER via2 ;
        RECT 2169.910 796.480 2170.190 796.760 ;
      LAYER met3 ;
        RECT 2169.885 796.770 2170.215 796.785 ;
        RECT 2169.670 796.455 2170.215 796.770 ;
        RECT 2169.670 794.440 2169.970 796.455 ;
        RECT 2166.000 793.840 2170.000 794.440 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3504.620 1500.910 3504.680 ;
        RECT 2170.350 3504.620 2170.670 3504.680 ;
        RECT 1500.590 3504.480 2170.670 3504.620 ;
        RECT 1500.590 3504.420 1500.910 3504.480 ;
        RECT 2170.350 3504.420 2170.670 3504.480 ;
      LAYER via ;
        RECT 1500.620 3504.420 1500.880 3504.680 ;
        RECT 2170.380 3504.420 2170.640 3504.680 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3504.710 1500.820 3517.600 ;
        RECT 1500.620 3504.390 1500.880 3504.710 ;
        RECT 2170.380 3504.390 2170.640 3504.710 ;
        RECT 2170.440 806.325 2170.580 3504.390 ;
        RECT 2170.370 805.955 2170.650 806.325 ;
      LAYER via2 ;
        RECT 2170.370 806.000 2170.650 806.280 ;
      LAYER met3 ;
        RECT 2170.345 806.290 2170.675 806.305 ;
        RECT 2169.670 805.990 2170.675 806.290 ;
        RECT 2169.670 805.320 2169.970 805.990 ;
        RECT 2170.345 805.975 2170.675 805.990 ;
        RECT 2166.000 804.720 2170.000 805.320 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2184.150 324.260 2184.470 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2184.150 324.120 2899.310 324.260 ;
        RECT 2184.150 324.060 2184.470 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2184.180 324.060 2184.440 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2184.170 614.195 2184.450 614.565 ;
        RECT 2184.240 324.350 2184.380 614.195 ;
        RECT 2184.180 324.030 2184.440 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2184.170 614.240 2184.450 614.520 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2166.000 615.000 2170.000 615.600 ;
        RECT 2169.670 614.530 2169.970 615.000 ;
        RECT 2184.145 614.530 2184.475 614.545 ;
        RECT 2169.670 614.230 2184.475 614.530 ;
        RECT 2184.145 614.215 2184.475 614.230 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3503.940 1176.150 3504.000 ;
        RECT 2170.810 3503.940 2171.130 3504.000 ;
        RECT 1175.830 3503.800 2171.130 3503.940 ;
        RECT 1175.830 3503.740 1176.150 3503.800 ;
        RECT 2170.810 3503.740 2171.130 3503.800 ;
      LAYER via ;
        RECT 1175.860 3503.740 1176.120 3504.000 ;
        RECT 2170.840 3503.740 2171.100 3504.000 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3504.030 1176.060 3517.600 ;
        RECT 1175.860 3503.710 1176.120 3504.030 ;
        RECT 2170.840 3503.710 2171.100 3504.030 ;
        RECT 2170.900 817.885 2171.040 3503.710 ;
        RECT 2170.830 817.515 2171.110 817.885 ;
      LAYER via2 ;
        RECT 2170.830 817.560 2171.110 817.840 ;
      LAYER met3 ;
        RECT 2170.805 817.850 2171.135 817.865 ;
        RECT 2169.670 817.550 2171.135 817.850 ;
        RECT 2169.670 815.520 2169.970 817.550 ;
        RECT 2170.805 817.535 2171.135 817.550 ;
        RECT 2166.000 814.920 2170.000 815.520 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3503.260 851.850 3503.320 ;
        RECT 2171.730 3503.260 2172.050 3503.320 ;
        RECT 851.530 3503.120 2172.050 3503.260 ;
        RECT 851.530 3503.060 851.850 3503.120 ;
        RECT 2171.730 3503.060 2172.050 3503.120 ;
      LAYER via ;
        RECT 851.560 3503.060 851.820 3503.320 ;
        RECT 2171.760 3503.060 2172.020 3503.320 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3503.350 851.760 3517.600 ;
        RECT 851.560 3503.030 851.820 3503.350 ;
        RECT 2171.760 3503.030 2172.020 3503.350 ;
        RECT 2171.820 828.085 2171.960 3503.030 ;
        RECT 2171.750 827.715 2172.030 828.085 ;
      LAYER via2 ;
        RECT 2171.750 827.760 2172.030 828.040 ;
      LAYER met3 ;
        RECT 2171.725 828.050 2172.055 828.065 ;
        RECT 2169.670 827.750 2172.055 828.050 ;
        RECT 2169.670 825.720 2169.970 827.750 ;
        RECT 2171.725 827.735 2172.055 827.750 ;
        RECT 2166.000 825.120 2170.000 825.720 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3502.240 527.550 3502.300 ;
        RECT 2172.190 3502.240 2172.510 3502.300 ;
        RECT 527.230 3502.100 2172.510 3502.240 ;
        RECT 527.230 3502.040 527.550 3502.100 ;
        RECT 2172.190 3502.040 2172.510 3502.100 ;
      LAYER via ;
        RECT 527.260 3502.040 527.520 3502.300 ;
        RECT 2172.220 3502.040 2172.480 3502.300 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3502.330 527.460 3517.600 ;
        RECT 527.260 3502.010 527.520 3502.330 ;
        RECT 2172.220 3502.010 2172.480 3502.330 ;
        RECT 2172.280 838.965 2172.420 3502.010 ;
        RECT 2172.210 838.595 2172.490 838.965 ;
      LAYER via2 ;
        RECT 2172.210 838.640 2172.490 838.920 ;
      LAYER met3 ;
        RECT 2172.185 838.930 2172.515 838.945 ;
        RECT 2169.670 838.630 2172.515 838.930 ;
        RECT 2169.670 836.600 2169.970 838.630 ;
        RECT 2172.185 838.615 2172.515 838.630 ;
        RECT 2166.000 836.000 2170.000 836.600 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.560 202.790 3501.620 ;
        RECT 2171.270 3501.560 2171.590 3501.620 ;
        RECT 202.470 3501.420 2171.590 3501.560 ;
        RECT 202.470 3501.360 202.790 3501.420 ;
        RECT 2171.270 3501.360 2171.590 3501.420 ;
      LAYER via ;
        RECT 202.500 3501.360 202.760 3501.620 ;
        RECT 2171.300 3501.360 2171.560 3501.620 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.650 202.700 3517.600 ;
        RECT 202.500 3501.330 202.760 3501.650 ;
        RECT 2171.300 3501.330 2171.560 3501.650 ;
        RECT 2171.360 848.485 2171.500 3501.330 ;
        RECT 2171.290 848.115 2171.570 848.485 ;
      LAYER via2 ;
        RECT 2171.290 848.160 2171.570 848.440 ;
      LAYER met3 ;
        RECT 2171.265 848.450 2171.595 848.465 ;
        RECT 2169.670 848.150 2171.595 848.450 ;
        RECT 2169.670 846.800 2169.970 848.150 ;
        RECT 2171.265 848.135 2171.595 848.150 ;
        RECT 2166.000 846.200 2170.000 846.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 2173.570 3408.740 2173.890 3408.800 ;
        RECT 17.550 3408.600 2173.890 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 2173.570 3408.540 2173.890 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 2173.600 3408.540 2173.860 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 2173.600 3408.510 2173.860 3408.830 ;
        RECT 2173.660 860.045 2173.800 3408.510 ;
        RECT 2173.590 859.675 2173.870 860.045 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
        RECT 2173.590 859.720 2173.870 860.000 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
        RECT 2173.565 860.010 2173.895 860.025 ;
        RECT 2169.670 859.710 2173.895 860.010 ;
        RECT 2169.670 857.680 2169.970 859.710 ;
        RECT 2173.565 859.695 2173.895 859.710 ;
        RECT 2166.000 857.080 2170.000 857.680 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3119.060 17.410 3119.120 ;
        RECT 2174.030 3119.060 2174.350 3119.120 ;
        RECT 17.090 3118.920 2174.350 3119.060 ;
        RECT 17.090 3118.860 17.410 3118.920 ;
        RECT 2174.030 3118.860 2174.350 3118.920 ;
      LAYER via ;
        RECT 17.120 3118.860 17.380 3119.120 ;
        RECT 2174.060 3118.860 2174.320 3119.120 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.150 17.320 3124.075 ;
        RECT 17.120 3118.830 17.380 3119.150 ;
        RECT 2174.060 3118.830 2174.320 3119.150 ;
        RECT 2174.120 869.565 2174.260 3118.830 ;
        RECT 2174.050 869.195 2174.330 869.565 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
        RECT 2174.050 869.240 2174.330 869.520 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
        RECT 2174.025 869.530 2174.355 869.545 ;
        RECT 2169.670 869.230 2174.355 869.530 ;
        RECT 2169.670 867.880 2169.970 869.230 ;
        RECT 2174.025 869.215 2174.355 869.230 ;
        RECT 2166.000 867.280 2170.000 867.880 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1004.940 17.410 1005.000 ;
        RECT 2181.850 1004.940 2182.170 1005.000 ;
        RECT 17.090 1004.800 2182.170 1004.940 ;
        RECT 17.090 1004.740 17.410 1004.800 ;
        RECT 2181.850 1004.740 2182.170 1004.800 ;
      LAYER via ;
        RECT 17.120 1004.740 17.380 1005.000 ;
        RECT 2181.880 1004.740 2182.140 1005.000 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 1005.030 17.320 2836.435 ;
        RECT 17.120 1004.710 17.380 1005.030 ;
        RECT 2181.880 1004.710 2182.140 1005.030 ;
        RECT 2181.940 881.125 2182.080 1004.710 ;
        RECT 2181.870 880.755 2182.150 881.125 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
        RECT 2181.870 880.800 2182.150 881.080 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
        RECT 2181.845 881.090 2182.175 881.105 ;
        RECT 2169.670 880.790 2182.175 881.090 ;
        RECT 2169.670 878.760 2169.970 880.790 ;
        RECT 2181.845 880.775 2182.175 880.790 ;
        RECT 2166.000 878.160 2170.000 878.760 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 1005.280 18.330 1005.340 ;
        RECT 2182.310 1005.280 2182.630 1005.340 ;
        RECT 18.010 1005.140 2182.630 1005.280 ;
        RECT 18.010 1005.080 18.330 1005.140 ;
        RECT 2182.310 1005.080 2182.630 1005.140 ;
      LAYER via ;
        RECT 18.040 1005.080 18.300 1005.340 ;
        RECT 2182.340 1005.080 2182.600 1005.340 ;
      LAYER met2 ;
        RECT 18.030 2549.475 18.310 2549.845 ;
        RECT 18.100 1005.370 18.240 2549.475 ;
        RECT 18.040 1005.050 18.300 1005.370 ;
        RECT 2182.340 1005.050 2182.600 1005.370 ;
        RECT 2182.400 889.965 2182.540 1005.050 ;
        RECT 2182.330 889.595 2182.610 889.965 ;
      LAYER via2 ;
        RECT 18.030 2549.520 18.310 2549.800 ;
        RECT 2182.330 889.640 2182.610 889.920 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 18.005 2549.810 18.335 2549.825 ;
        RECT -4.800 2549.510 18.335 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 18.005 2549.495 18.335 2549.510 ;
        RECT 2182.305 889.930 2182.635 889.945 ;
        RECT 2169.670 889.630 2182.635 889.930 ;
        RECT 2169.670 888.960 2169.970 889.630 ;
        RECT 2182.305 889.615 2182.635 889.630 ;
        RECT 2166.000 888.360 2170.000 888.960 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 2256.820 15.570 2256.880 ;
        RECT 1336.370 2256.820 1336.690 2256.880 ;
        RECT 15.250 2256.680 1336.690 2256.820 ;
        RECT 15.250 2256.620 15.570 2256.680 ;
        RECT 1336.370 2256.620 1336.690 2256.680 ;
        RECT 1336.370 1928.380 1336.690 1928.440 ;
        RECT 2180.470 1928.380 2180.790 1928.440 ;
        RECT 1336.370 1928.240 2180.790 1928.380 ;
        RECT 1336.370 1928.180 1336.690 1928.240 ;
        RECT 2180.470 1928.180 2180.790 1928.240 ;
      LAYER via ;
        RECT 15.280 2256.620 15.540 2256.880 ;
        RECT 1336.400 2256.620 1336.660 2256.880 ;
        RECT 1336.400 1928.180 1336.660 1928.440 ;
        RECT 2180.500 1928.180 2180.760 1928.440 ;
      LAYER met2 ;
        RECT 15.270 2261.835 15.550 2262.205 ;
        RECT 15.340 2256.910 15.480 2261.835 ;
        RECT 15.280 2256.590 15.540 2256.910 ;
        RECT 1336.400 2256.590 1336.660 2256.910 ;
        RECT 1336.460 1928.470 1336.600 2256.590 ;
        RECT 1336.400 1928.150 1336.660 1928.470 ;
        RECT 2180.500 1928.150 2180.760 1928.470 ;
        RECT 2180.560 901.525 2180.700 1928.150 ;
        RECT 2180.490 901.155 2180.770 901.525 ;
      LAYER via2 ;
        RECT 15.270 2261.880 15.550 2262.160 ;
        RECT 2180.490 901.200 2180.770 901.480 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 15.245 2262.170 15.575 2262.185 ;
        RECT -4.800 2261.870 15.575 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 15.245 2261.855 15.575 2261.870 ;
        RECT 2180.465 901.490 2180.795 901.505 ;
        RECT 2169.670 901.190 2180.795 901.490 ;
        RECT 2169.670 899.840 2169.970 901.190 ;
        RECT 2180.465 901.175 2180.795 901.190 ;
        RECT 2166.000 899.240 2170.000 899.840 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 1005.620 19.710 1005.680 ;
        RECT 2182.770 1005.620 2183.090 1005.680 ;
        RECT 19.390 1005.480 2183.090 1005.620 ;
        RECT 19.390 1005.420 19.710 1005.480 ;
        RECT 2182.770 1005.420 2183.090 1005.480 ;
      LAYER via ;
        RECT 19.420 1005.420 19.680 1005.680 ;
        RECT 2182.800 1005.420 2183.060 1005.680 ;
      LAYER met2 ;
        RECT 19.410 1974.875 19.690 1975.245 ;
        RECT 19.480 1005.710 19.620 1974.875 ;
        RECT 19.420 1005.390 19.680 1005.710 ;
        RECT 2182.800 1005.390 2183.060 1005.710 ;
        RECT 2182.860 910.365 2183.000 1005.390 ;
        RECT 2182.790 909.995 2183.070 910.365 ;
      LAYER via2 ;
        RECT 19.410 1974.920 19.690 1975.200 ;
        RECT 2182.790 910.040 2183.070 910.320 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 19.385 1975.210 19.715 1975.225 ;
        RECT -4.800 1974.910 19.715 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 19.385 1974.895 19.715 1974.910 ;
        RECT 2182.765 910.330 2183.095 910.345 ;
        RECT 2169.670 910.040 2183.095 910.330 ;
        RECT 2166.000 910.030 2183.095 910.040 ;
        RECT 2166.000 909.440 2170.000 910.030 ;
        RECT 2182.765 910.015 2183.095 910.030 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2184.610 558.860 2184.930 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2184.610 558.720 2899.310 558.860 ;
        RECT 2184.610 558.660 2184.930 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2184.640 558.660 2184.900 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2184.630 622.355 2184.910 622.725 ;
        RECT 2184.700 558.950 2184.840 622.355 ;
        RECT 2184.640 558.630 2184.900 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2184.630 622.400 2184.910 622.680 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2166.000 625.200 2170.000 625.800 ;
        RECT 2169.670 622.690 2169.970 625.200 ;
        RECT 2184.605 622.690 2184.935 622.705 ;
        RECT 2169.670 622.390 2184.935 622.690 ;
        RECT 2184.605 622.375 2184.935 622.390 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 14.790 1683.920 15.110 1683.980 ;
        RECT 2174.490 1683.920 2174.810 1683.980 ;
        RECT 14.790 1683.780 2174.810 1683.920 ;
        RECT 14.790 1683.720 15.110 1683.780 ;
        RECT 2174.490 1683.720 2174.810 1683.780 ;
      LAYER via ;
        RECT 14.820 1683.720 15.080 1683.980 ;
        RECT 2174.520 1683.720 2174.780 1683.980 ;
      LAYER met2 ;
        RECT 14.810 1687.235 15.090 1687.605 ;
        RECT 14.880 1684.010 15.020 1687.235 ;
        RECT 14.820 1683.690 15.080 1684.010 ;
        RECT 2174.520 1683.690 2174.780 1684.010 ;
        RECT 2174.580 923.285 2174.720 1683.690 ;
        RECT 2174.510 922.915 2174.790 923.285 ;
      LAYER via2 ;
        RECT 14.810 1687.280 15.090 1687.560 ;
        RECT 2174.510 922.960 2174.790 923.240 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 14.785 1687.570 15.115 1687.585 ;
        RECT -4.800 1687.270 15.115 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 14.785 1687.255 15.115 1687.270 ;
        RECT 2174.485 923.250 2174.815 923.265 ;
        RECT 2169.670 922.950 2174.815 923.250 ;
        RECT 2169.670 920.920 2169.970 922.950 ;
        RECT 2174.485 922.935 2174.815 922.950 ;
        RECT 2166.000 920.320 2170.000 920.920 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 1470.060 16.950 1470.120 ;
        RECT 2172.650 1470.060 2172.970 1470.120 ;
        RECT 16.630 1469.920 2172.970 1470.060 ;
        RECT 16.630 1469.860 16.950 1469.920 ;
        RECT 2172.650 1469.860 2172.970 1469.920 ;
      LAYER via ;
        RECT 16.660 1469.860 16.920 1470.120 ;
        RECT 2172.680 1469.860 2172.940 1470.120 ;
      LAYER met2 ;
        RECT 16.650 1471.675 16.930 1472.045 ;
        RECT 16.720 1470.150 16.860 1471.675 ;
        RECT 16.660 1469.830 16.920 1470.150 ;
        RECT 2172.680 1469.830 2172.940 1470.150 ;
        RECT 2172.740 931.445 2172.880 1469.830 ;
        RECT 2172.670 931.075 2172.950 931.445 ;
      LAYER via2 ;
        RECT 16.650 1471.720 16.930 1472.000 ;
        RECT 2172.670 931.120 2172.950 931.400 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 16.625 1472.010 16.955 1472.025 ;
        RECT -4.800 1471.710 16.955 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 16.625 1471.695 16.955 1471.710 ;
        RECT 2172.645 931.410 2172.975 931.425 ;
        RECT 2169.670 931.120 2172.975 931.410 ;
        RECT 2166.000 931.110 2172.975 931.120 ;
        RECT 2166.000 930.520 2170.000 931.110 ;
        RECT 2172.645 931.095 2172.975 931.110 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 1256.200 16.950 1256.260 ;
        RECT 2175.410 1256.200 2175.730 1256.260 ;
        RECT 16.630 1256.060 2175.730 1256.200 ;
        RECT 16.630 1256.000 16.950 1256.060 ;
        RECT 2175.410 1256.000 2175.730 1256.060 ;
      LAYER via ;
        RECT 16.660 1256.000 16.920 1256.260 ;
        RECT 2175.440 1256.000 2175.700 1256.260 ;
      LAYER met2 ;
        RECT 16.650 1256.115 16.930 1256.485 ;
        RECT 16.660 1255.970 16.920 1256.115 ;
        RECT 2175.440 1255.970 2175.700 1256.290 ;
        RECT 2175.500 944.365 2175.640 1255.970 ;
        RECT 2175.430 943.995 2175.710 944.365 ;
      LAYER via2 ;
        RECT 16.650 1256.160 16.930 1256.440 ;
        RECT 2175.430 944.040 2175.710 944.320 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 16.625 1256.450 16.955 1256.465 ;
        RECT -4.800 1256.150 16.955 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 16.625 1256.135 16.955 1256.150 ;
        RECT 2175.405 944.330 2175.735 944.345 ;
        RECT 2169.670 944.030 2175.735 944.330 ;
        RECT 2169.670 942.000 2169.970 944.030 ;
        RECT 2175.405 944.015 2175.735 944.030 ;
        RECT 2166.000 941.400 2170.000 942.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 14.790 1035.200 15.110 1035.260 ;
        RECT 2175.870 1035.200 2176.190 1035.260 ;
        RECT 14.790 1035.060 2176.190 1035.200 ;
        RECT 14.790 1035.000 15.110 1035.060 ;
        RECT 2175.870 1035.000 2176.190 1035.060 ;
      LAYER via ;
        RECT 14.820 1035.000 15.080 1035.260 ;
        RECT 2175.900 1035.000 2176.160 1035.260 ;
      LAYER met2 ;
        RECT 14.810 1040.555 15.090 1040.925 ;
        RECT 14.880 1035.290 15.020 1040.555 ;
        RECT 14.820 1034.970 15.080 1035.290 ;
        RECT 2175.900 1034.970 2176.160 1035.290 ;
        RECT 2175.960 951.165 2176.100 1034.970 ;
        RECT 2175.890 950.795 2176.170 951.165 ;
      LAYER via2 ;
        RECT 14.810 1040.600 15.090 1040.880 ;
        RECT 2175.890 950.840 2176.170 951.120 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 14.785 1040.890 15.115 1040.905 ;
        RECT -4.800 1040.590 15.115 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 14.785 1040.575 15.115 1040.590 ;
        RECT 2166.000 951.600 2170.000 952.200 ;
        RECT 2169.670 951.130 2169.970 951.600 ;
        RECT 2175.865 951.130 2176.195 951.145 ;
        RECT 2169.670 950.830 2176.195 951.130 ;
        RECT 2175.865 950.815 2176.195 950.830 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 1000.860 16.490 1000.920 ;
        RECT 2183.230 1000.860 2183.550 1000.920 ;
        RECT 16.170 1000.720 2183.550 1000.860 ;
        RECT 16.170 1000.660 16.490 1000.720 ;
        RECT 2183.230 1000.660 2183.550 1000.720 ;
      LAYER via ;
        RECT 16.200 1000.660 16.460 1000.920 ;
        RECT 2183.260 1000.660 2183.520 1000.920 ;
      LAYER met2 ;
        RECT 16.200 1000.630 16.460 1000.950 ;
        RECT 2183.260 1000.630 2183.520 1000.950 ;
        RECT 16.260 825.365 16.400 1000.630 ;
        RECT 2183.320 965.445 2183.460 1000.630 ;
        RECT 2183.250 965.075 2183.530 965.445 ;
        RECT 16.190 824.995 16.470 825.365 ;
      LAYER via2 ;
        RECT 2183.250 965.120 2183.530 965.400 ;
        RECT 16.190 825.040 16.470 825.320 ;
      LAYER met3 ;
        RECT 2183.225 965.410 2183.555 965.425 ;
        RECT 2169.670 965.110 2183.555 965.410 ;
        RECT 2169.670 963.080 2169.970 965.110 ;
        RECT 2183.225 965.095 2183.555 965.110 ;
        RECT 2166.000 962.480 2170.000 963.080 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 16.165 825.330 16.495 825.345 ;
        RECT -4.800 825.030 16.495 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 16.165 825.015 16.495 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 603.060 16.950 603.120 ;
        RECT 2181.390 603.060 2181.710 603.120 ;
        RECT 16.630 602.920 2181.710 603.060 ;
        RECT 16.630 602.860 16.950 602.920 ;
        RECT 2181.390 602.860 2181.710 602.920 ;
      LAYER via ;
        RECT 16.660 602.860 16.920 603.120 ;
        RECT 2181.420 602.860 2181.680 603.120 ;
      LAYER met2 ;
        RECT 2181.410 969.835 2181.690 970.205 ;
        RECT 16.650 610.115 16.930 610.485 ;
        RECT 16.720 603.150 16.860 610.115 ;
        RECT 2181.480 603.150 2181.620 969.835 ;
        RECT 16.660 602.830 16.920 603.150 ;
        RECT 2181.420 602.830 2181.680 603.150 ;
      LAYER via2 ;
        RECT 2181.410 969.880 2181.690 970.160 ;
        RECT 16.650 610.160 16.930 610.440 ;
      LAYER met3 ;
        RECT 2166.000 972.680 2170.000 973.280 ;
        RECT 2169.670 970.170 2169.970 972.680 ;
        RECT 2181.385 970.170 2181.715 970.185 ;
        RECT 2169.670 969.870 2181.715 970.170 ;
        RECT 2181.385 969.855 2181.715 969.870 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 16.625 610.450 16.955 610.465 ;
        RECT -4.800 610.150 16.955 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 16.625 610.135 16.955 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 675.440 400.280 705.020 400.420 ;
        RECT 16.170 400.080 16.490 400.140 ;
        RECT 675.440 400.080 675.580 400.280 ;
        RECT 16.170 399.940 675.580 400.080 ;
        RECT 704.880 400.080 705.020 400.280 ;
        RECT 2037.500 400.280 2076.280 400.420 ;
        RECT 2037.500 400.080 2037.640 400.280 ;
        RECT 704.880 399.940 1068.880 400.080 ;
        RECT 16.170 399.880 16.490 399.940 ;
        RECT 1068.740 399.740 1068.880 399.940 ;
        RECT 1084.840 399.940 2037.640 400.080 ;
        RECT 2076.140 400.080 2076.280 400.280 ;
        RECT 2174.950 400.080 2175.270 400.140 ;
        RECT 2076.140 399.940 2175.270 400.080 ;
        RECT 1084.840 399.740 1084.980 399.940 ;
        RECT 2174.950 399.880 2175.270 399.940 ;
        RECT 1068.740 399.600 1084.980 399.740 ;
      LAYER via ;
        RECT 16.200 399.880 16.460 400.140 ;
        RECT 2174.980 399.880 2175.240 400.140 ;
      LAYER met2 ;
        RECT 2174.970 980.715 2175.250 981.085 ;
        RECT 2175.040 400.170 2175.180 980.715 ;
        RECT 16.200 399.850 16.460 400.170 ;
        RECT 2174.980 399.850 2175.240 400.170 ;
        RECT 16.260 394.925 16.400 399.850 ;
        RECT 16.190 394.555 16.470 394.925 ;
      LAYER via2 ;
        RECT 2174.970 980.760 2175.250 981.040 ;
        RECT 16.190 394.600 16.470 394.880 ;
      LAYER met3 ;
        RECT 2166.000 983.560 2170.000 984.160 ;
        RECT 2169.670 981.050 2169.970 983.560 ;
        RECT 2174.945 981.050 2175.275 981.065 ;
        RECT 2169.670 980.750 2175.275 981.050 ;
        RECT 2174.945 980.735 2175.275 980.750 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 16.165 394.890 16.495 394.905 ;
        RECT -4.800 394.590 16.495 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 16.165 394.575 16.495 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 2180.930 179.420 2181.250 179.480 ;
        RECT 17.090 179.280 2181.250 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 2180.930 179.220 2181.250 179.280 ;
      LAYER via ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 2180.960 179.220 2181.220 179.480 ;
      LAYER met2 ;
        RECT 2180.950 994.315 2181.230 994.685 ;
        RECT 2181.020 179.510 2181.160 994.315 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 2180.960 179.190 2181.220 179.510 ;
      LAYER via2 ;
        RECT 2180.950 994.360 2181.230 994.640 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 2180.925 994.650 2181.255 994.665 ;
        RECT 2169.670 994.360 2181.255 994.650 ;
        RECT 2166.000 994.350 2181.255 994.360 ;
        RECT 2166.000 993.760 2170.000 994.350 ;
        RECT 2180.925 994.335 2181.255 994.350 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2184.150 787.000 2184.470 787.060 ;
        RECT 2900.830 787.000 2901.150 787.060 ;
        RECT 2184.150 786.860 2901.150 787.000 ;
        RECT 2184.150 786.800 2184.470 786.860 ;
        RECT 2900.830 786.800 2901.150 786.860 ;
      LAYER via ;
        RECT 2184.180 786.800 2184.440 787.060 ;
        RECT 2900.860 786.800 2901.120 787.060 ;
      LAYER met2 ;
        RECT 2900.850 791.675 2901.130 792.045 ;
        RECT 2900.920 787.090 2901.060 791.675 ;
        RECT 2184.180 786.770 2184.440 787.090 ;
        RECT 2900.860 786.770 2901.120 787.090 ;
        RECT 2184.240 639.045 2184.380 786.770 ;
        RECT 2184.170 638.675 2184.450 639.045 ;
      LAYER via2 ;
        RECT 2900.850 791.720 2901.130 792.000 ;
        RECT 2184.170 638.720 2184.450 639.000 ;
      LAYER met3 ;
        RECT 2900.825 792.010 2901.155 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2900.825 791.710 2924.800 792.010 ;
        RECT 2900.825 791.695 2901.155 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2184.145 639.010 2184.475 639.025 ;
        RECT 2169.670 638.710 2184.475 639.010 ;
        RECT 2169.670 636.680 2169.970 638.710 ;
        RECT 2184.145 638.695 2184.475 638.710 ;
        RECT 2166.000 636.080 2170.000 636.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 648.620 2187.230 648.680 ;
        RECT 2904.050 648.620 2904.370 648.680 ;
        RECT 2186.910 648.480 2904.370 648.620 ;
        RECT 2186.910 648.420 2187.230 648.480 ;
        RECT 2904.050 648.420 2904.370 648.480 ;
      LAYER via ;
        RECT 2186.940 648.420 2187.200 648.680 ;
        RECT 2904.080 648.420 2904.340 648.680 ;
      LAYER met2 ;
        RECT 2904.070 1026.275 2904.350 1026.645 ;
        RECT 2904.140 648.710 2904.280 1026.275 ;
        RECT 2186.940 648.390 2187.200 648.710 ;
        RECT 2904.080 648.390 2904.340 648.710 ;
        RECT 2187.000 647.885 2187.140 648.390 ;
        RECT 2186.930 647.515 2187.210 647.885 ;
      LAYER via2 ;
        RECT 2904.070 1026.320 2904.350 1026.600 ;
        RECT 2186.930 647.560 2187.210 647.840 ;
      LAYER met3 ;
        RECT 2904.045 1026.610 2904.375 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2904.045 1026.310 2924.800 1026.610 ;
        RECT 2904.045 1026.295 2904.375 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2186.905 647.850 2187.235 647.865 ;
        RECT 2169.670 647.550 2187.235 647.850 ;
        RECT 2169.670 646.880 2169.970 647.550 ;
        RECT 2186.905 647.535 2187.235 647.550 ;
        RECT 2166.000 646.280 2170.000 646.880 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 662.220 2187.230 662.280 ;
        RECT 2903.590 662.220 2903.910 662.280 ;
        RECT 2186.910 662.080 2903.910 662.220 ;
        RECT 2186.910 662.020 2187.230 662.080 ;
        RECT 2903.590 662.020 2903.910 662.080 ;
      LAYER via ;
        RECT 2186.940 662.020 2187.200 662.280 ;
        RECT 2903.620 662.020 2903.880 662.280 ;
      LAYER met2 ;
        RECT 2903.610 1260.875 2903.890 1261.245 ;
        RECT 2903.680 662.310 2903.820 1260.875 ;
        RECT 2186.940 661.990 2187.200 662.310 ;
        RECT 2903.620 661.990 2903.880 662.310 ;
        RECT 2187.000 660.125 2187.140 661.990 ;
        RECT 2186.930 659.755 2187.210 660.125 ;
      LAYER via2 ;
        RECT 2903.610 1260.920 2903.890 1261.200 ;
        RECT 2186.930 659.800 2187.210 660.080 ;
      LAYER met3 ;
        RECT 2903.585 1261.210 2903.915 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2903.585 1260.910 2924.800 1261.210 ;
        RECT 2903.585 1260.895 2903.915 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2186.905 660.090 2187.235 660.105 ;
        RECT 2169.670 659.790 2187.235 660.090 ;
        RECT 2169.670 657.760 2169.970 659.790 ;
        RECT 2186.905 659.775 2187.235 659.790 ;
        RECT 2166.000 657.160 2170.000 657.760 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 669.360 2187.230 669.420 ;
        RECT 2903.130 669.360 2903.450 669.420 ;
        RECT 2186.910 669.220 2903.450 669.360 ;
        RECT 2186.910 669.160 2187.230 669.220 ;
        RECT 2903.130 669.160 2903.450 669.220 ;
      LAYER via ;
        RECT 2186.940 669.160 2187.200 669.420 ;
        RECT 2903.160 669.160 2903.420 669.420 ;
      LAYER met2 ;
        RECT 2903.150 1495.475 2903.430 1495.845 ;
        RECT 2903.220 669.450 2903.360 1495.475 ;
        RECT 2186.940 669.130 2187.200 669.450 ;
        RECT 2903.160 669.130 2903.420 669.450 ;
        RECT 2187.000 668.285 2187.140 669.130 ;
        RECT 2186.930 667.915 2187.210 668.285 ;
      LAYER via2 ;
        RECT 2903.150 1495.520 2903.430 1495.800 ;
        RECT 2186.930 667.960 2187.210 668.240 ;
      LAYER met3 ;
        RECT 2903.125 1495.810 2903.455 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2903.125 1495.510 2924.800 1495.810 ;
        RECT 2903.125 1495.495 2903.455 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2186.905 668.250 2187.235 668.265 ;
        RECT 2169.670 667.960 2187.235 668.250 ;
        RECT 2166.000 667.950 2187.235 667.960 ;
        RECT 2166.000 667.360 2170.000 667.950 ;
        RECT 2186.905 667.935 2187.235 667.950 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2524.090 1725.400 2524.410 1725.460 ;
        RECT 2899.910 1725.400 2900.230 1725.460 ;
        RECT 2524.090 1725.260 2900.230 1725.400 ;
        RECT 2524.090 1725.200 2524.410 1725.260 ;
        RECT 2899.910 1725.200 2900.230 1725.260 ;
        RECT 2521.790 1593.820 2522.110 1593.880 ;
        RECT 2522.250 1593.820 2522.570 1593.880 ;
        RECT 2521.790 1593.680 2522.570 1593.820 ;
        RECT 2521.790 1593.620 2522.110 1593.680 ;
        RECT 2522.250 1593.620 2522.570 1593.680 ;
        RECT 2521.790 1546.220 2522.110 1546.280 ;
        RECT 2522.250 1546.220 2522.570 1546.280 ;
        RECT 2521.790 1546.080 2522.570 1546.220 ;
        RECT 2521.790 1546.020 2522.110 1546.080 ;
        RECT 2522.250 1546.020 2522.570 1546.080 ;
        RECT 2520.870 1545.540 2521.190 1545.600 ;
        RECT 2521.790 1545.540 2522.110 1545.600 ;
        RECT 2520.870 1545.400 2522.110 1545.540 ;
        RECT 2520.870 1545.340 2521.190 1545.400 ;
        RECT 2521.790 1545.340 2522.110 1545.400 ;
        RECT 2520.870 1497.600 2521.190 1497.660 ;
        RECT 2522.250 1497.600 2522.570 1497.660 ;
        RECT 2520.870 1497.460 2522.570 1497.600 ;
        RECT 2520.870 1497.400 2521.190 1497.460 ;
        RECT 2522.250 1497.400 2522.570 1497.460 ;
        RECT 2522.250 1490.460 2522.570 1490.520 ;
        RECT 2523.630 1490.460 2523.950 1490.520 ;
        RECT 2522.250 1490.320 2523.950 1490.460 ;
        RECT 2522.250 1490.260 2522.570 1490.320 ;
        RECT 2523.630 1490.260 2523.950 1490.320 ;
        RECT 2522.710 1442.180 2523.030 1442.240 ;
        RECT 2523.630 1442.180 2523.950 1442.240 ;
        RECT 2522.710 1442.040 2523.950 1442.180 ;
        RECT 2522.710 1441.980 2523.030 1442.040 ;
        RECT 2523.630 1441.980 2523.950 1442.040 ;
        RECT 2522.250 1393.560 2522.570 1393.620 ;
        RECT 2522.710 1393.560 2523.030 1393.620 ;
        RECT 2522.250 1393.420 2523.030 1393.560 ;
        RECT 2522.250 1393.360 2522.570 1393.420 ;
        RECT 2522.710 1393.360 2523.030 1393.420 ;
        RECT 2521.330 1304.140 2521.650 1304.200 ;
        RECT 2522.710 1304.140 2523.030 1304.200 ;
        RECT 2521.330 1304.000 2523.030 1304.140 ;
        RECT 2521.330 1303.940 2521.650 1304.000 ;
        RECT 2522.710 1303.940 2523.030 1304.000 ;
        RECT 2521.330 1269.120 2521.650 1269.180 ;
        RECT 2522.710 1269.120 2523.030 1269.180 ;
        RECT 2521.330 1268.980 2523.030 1269.120 ;
        RECT 2521.330 1268.920 2521.650 1268.980 ;
        RECT 2522.710 1268.920 2523.030 1268.980 ;
        RECT 2520.410 1255.860 2520.730 1255.920 ;
        RECT 2521.330 1255.860 2521.650 1255.920 ;
        RECT 2520.410 1255.720 2521.650 1255.860 ;
        RECT 2520.410 1255.660 2520.730 1255.720 ;
        RECT 2521.330 1255.660 2521.650 1255.720 ;
        RECT 2520.410 1207.580 2520.730 1207.640 ;
        RECT 2522.250 1207.580 2522.570 1207.640 ;
        RECT 2520.410 1207.440 2522.570 1207.580 ;
        RECT 2520.410 1207.380 2520.730 1207.440 ;
        RECT 2522.250 1207.380 2522.570 1207.440 ;
        RECT 2522.250 1173.580 2522.570 1173.640 ;
        RECT 2521.880 1173.440 2522.570 1173.580 ;
        RECT 2521.880 1172.960 2522.020 1173.440 ;
        RECT 2522.250 1173.380 2522.570 1173.440 ;
        RECT 2521.790 1172.700 2522.110 1172.960 ;
        RECT 2520.870 1158.960 2521.190 1159.020 ;
        RECT 2521.790 1158.960 2522.110 1159.020 ;
        RECT 2520.870 1158.820 2522.110 1158.960 ;
        RECT 2520.870 1158.760 2521.190 1158.820 ;
        RECT 2521.790 1158.760 2522.110 1158.820 ;
        RECT 2520.870 1111.020 2521.190 1111.080 ;
        RECT 2522.250 1111.020 2522.570 1111.080 ;
        RECT 2520.870 1110.880 2522.570 1111.020 ;
        RECT 2520.870 1110.820 2521.190 1110.880 ;
        RECT 2522.250 1110.820 2522.570 1110.880 ;
        RECT 2522.250 1077.020 2522.570 1077.080 ;
        RECT 2521.420 1076.880 2522.570 1077.020 ;
        RECT 2521.420 1076.400 2521.560 1076.880 ;
        RECT 2522.250 1076.820 2522.570 1076.880 ;
        RECT 2521.330 1076.140 2521.650 1076.400 ;
        RECT 2520.870 1028.400 2521.190 1028.460 ;
        RECT 2520.870 1028.260 2521.560 1028.400 ;
        RECT 2520.870 1028.200 2521.190 1028.260 ;
        RECT 2521.420 1028.120 2521.560 1028.260 ;
        RECT 2521.330 1027.860 2521.650 1028.120 ;
        RECT 2520.870 1014.460 2521.190 1014.520 ;
        RECT 2521.330 1014.460 2521.650 1014.520 ;
        RECT 2520.870 1014.320 2521.650 1014.460 ;
        RECT 2520.870 1014.260 2521.190 1014.320 ;
        RECT 2521.330 1014.260 2521.650 1014.320 ;
        RECT 2520.870 1013.780 2521.190 1013.840 ;
        RECT 2522.250 1013.780 2522.570 1013.840 ;
        RECT 2520.870 1013.640 2522.570 1013.780 ;
        RECT 2520.870 1013.580 2521.190 1013.640 ;
        RECT 2522.250 1013.580 2522.570 1013.640 ;
        RECT 2522.250 869.620 2522.570 869.680 ;
        RECT 2523.170 869.620 2523.490 869.680 ;
        RECT 2522.250 869.480 2523.490 869.620 ;
        RECT 2522.250 869.420 2522.570 869.480 ;
        RECT 2523.170 869.420 2523.490 869.480 ;
        RECT 2520.870 821.000 2521.190 821.060 ;
        RECT 2521.790 821.000 2522.110 821.060 ;
        RECT 2520.870 820.860 2522.110 821.000 ;
        RECT 2520.870 820.800 2521.190 820.860 ;
        RECT 2521.790 820.800 2522.110 820.860 ;
        RECT 2185.070 682.960 2185.390 683.020 ;
        RECT 2522.250 682.960 2522.570 683.020 ;
        RECT 2185.070 682.820 2522.570 682.960 ;
        RECT 2185.070 682.760 2185.390 682.820 ;
        RECT 2522.250 682.760 2522.570 682.820 ;
      LAYER via ;
        RECT 2524.120 1725.200 2524.380 1725.460 ;
        RECT 2899.940 1725.200 2900.200 1725.460 ;
        RECT 2521.820 1593.620 2522.080 1593.880 ;
        RECT 2522.280 1593.620 2522.540 1593.880 ;
        RECT 2521.820 1546.020 2522.080 1546.280 ;
        RECT 2522.280 1546.020 2522.540 1546.280 ;
        RECT 2520.900 1545.340 2521.160 1545.600 ;
        RECT 2521.820 1545.340 2522.080 1545.600 ;
        RECT 2520.900 1497.400 2521.160 1497.660 ;
        RECT 2522.280 1497.400 2522.540 1497.660 ;
        RECT 2522.280 1490.260 2522.540 1490.520 ;
        RECT 2523.660 1490.260 2523.920 1490.520 ;
        RECT 2522.740 1441.980 2523.000 1442.240 ;
        RECT 2523.660 1441.980 2523.920 1442.240 ;
        RECT 2522.280 1393.360 2522.540 1393.620 ;
        RECT 2522.740 1393.360 2523.000 1393.620 ;
        RECT 2521.360 1303.940 2521.620 1304.200 ;
        RECT 2522.740 1303.940 2523.000 1304.200 ;
        RECT 2521.360 1268.920 2521.620 1269.180 ;
        RECT 2522.740 1268.920 2523.000 1269.180 ;
        RECT 2520.440 1255.660 2520.700 1255.920 ;
        RECT 2521.360 1255.660 2521.620 1255.920 ;
        RECT 2520.440 1207.380 2520.700 1207.640 ;
        RECT 2522.280 1207.380 2522.540 1207.640 ;
        RECT 2522.280 1173.380 2522.540 1173.640 ;
        RECT 2521.820 1172.700 2522.080 1172.960 ;
        RECT 2520.900 1158.760 2521.160 1159.020 ;
        RECT 2521.820 1158.760 2522.080 1159.020 ;
        RECT 2520.900 1110.820 2521.160 1111.080 ;
        RECT 2522.280 1110.820 2522.540 1111.080 ;
        RECT 2522.280 1076.820 2522.540 1077.080 ;
        RECT 2521.360 1076.140 2521.620 1076.400 ;
        RECT 2520.900 1028.200 2521.160 1028.460 ;
        RECT 2521.360 1027.860 2521.620 1028.120 ;
        RECT 2520.900 1014.260 2521.160 1014.520 ;
        RECT 2521.360 1014.260 2521.620 1014.520 ;
        RECT 2520.900 1013.580 2521.160 1013.840 ;
        RECT 2522.280 1013.580 2522.540 1013.840 ;
        RECT 2522.280 869.420 2522.540 869.680 ;
        RECT 2523.200 869.420 2523.460 869.680 ;
        RECT 2520.900 820.800 2521.160 821.060 ;
        RECT 2521.820 820.800 2522.080 821.060 ;
        RECT 2185.100 682.760 2185.360 683.020 ;
        RECT 2522.280 682.760 2522.540 683.020 ;
      LAYER met2 ;
        RECT 2899.930 1730.075 2900.210 1730.445 ;
        RECT 2900.000 1725.490 2900.140 1730.075 ;
        RECT 2524.120 1725.170 2524.380 1725.490 ;
        RECT 2899.940 1725.170 2900.200 1725.490 ;
        RECT 2524.180 1663.010 2524.320 1725.170 ;
        RECT 2522.340 1662.870 2524.320 1663.010 ;
        RECT 2522.340 1656.210 2522.480 1662.870 ;
        RECT 2521.880 1656.070 2522.480 1656.210 ;
        RECT 2521.880 1593.910 2522.020 1656.070 ;
        RECT 2521.820 1593.590 2522.080 1593.910 ;
        RECT 2522.280 1593.590 2522.540 1593.910 ;
        RECT 2522.340 1546.310 2522.480 1593.590 ;
        RECT 2521.820 1545.990 2522.080 1546.310 ;
        RECT 2522.280 1545.990 2522.540 1546.310 ;
        RECT 2521.880 1545.630 2522.020 1545.990 ;
        RECT 2520.900 1545.310 2521.160 1545.630 ;
        RECT 2521.820 1545.310 2522.080 1545.630 ;
        RECT 2520.960 1497.690 2521.100 1545.310 ;
        RECT 2520.900 1497.370 2521.160 1497.690 ;
        RECT 2522.280 1497.370 2522.540 1497.690 ;
        RECT 2522.340 1490.550 2522.480 1497.370 ;
        RECT 2522.280 1490.230 2522.540 1490.550 ;
        RECT 2523.660 1490.230 2523.920 1490.550 ;
        RECT 2523.720 1442.270 2523.860 1490.230 ;
        RECT 2522.740 1441.950 2523.000 1442.270 ;
        RECT 2523.660 1441.950 2523.920 1442.270 ;
        RECT 2522.800 1401.210 2522.940 1441.950 ;
        RECT 2522.340 1401.070 2522.940 1401.210 ;
        RECT 2522.340 1393.650 2522.480 1401.070 ;
        RECT 2522.280 1393.330 2522.540 1393.650 ;
        RECT 2522.740 1393.330 2523.000 1393.650 ;
        RECT 2522.800 1304.765 2522.940 1393.330 ;
        RECT 2521.350 1304.395 2521.630 1304.765 ;
        RECT 2522.730 1304.395 2523.010 1304.765 ;
        RECT 2521.420 1304.230 2521.560 1304.395 ;
        RECT 2521.360 1303.910 2521.620 1304.230 ;
        RECT 2522.740 1303.910 2523.000 1304.230 ;
        RECT 2522.800 1269.210 2522.940 1303.910 ;
        RECT 2521.360 1268.890 2521.620 1269.210 ;
        RECT 2522.740 1268.890 2523.000 1269.210 ;
        RECT 2521.420 1255.950 2521.560 1268.890 ;
        RECT 2520.440 1255.630 2520.700 1255.950 ;
        RECT 2521.360 1255.630 2521.620 1255.950 ;
        RECT 2520.500 1207.670 2520.640 1255.630 ;
        RECT 2520.440 1207.350 2520.700 1207.670 ;
        RECT 2522.280 1207.350 2522.540 1207.670 ;
        RECT 2522.340 1173.670 2522.480 1207.350 ;
        RECT 2522.280 1173.350 2522.540 1173.670 ;
        RECT 2521.820 1172.670 2522.080 1172.990 ;
        RECT 2521.880 1159.050 2522.020 1172.670 ;
        RECT 2520.900 1158.730 2521.160 1159.050 ;
        RECT 2521.820 1158.730 2522.080 1159.050 ;
        RECT 2520.960 1111.110 2521.100 1158.730 ;
        RECT 2520.900 1110.790 2521.160 1111.110 ;
        RECT 2522.280 1110.790 2522.540 1111.110 ;
        RECT 2522.340 1077.110 2522.480 1110.790 ;
        RECT 2522.280 1076.790 2522.540 1077.110 ;
        RECT 2521.360 1076.110 2521.620 1076.430 ;
        RECT 2521.420 1062.570 2521.560 1076.110 ;
        RECT 2520.960 1062.430 2521.560 1062.570 ;
        RECT 2520.960 1028.490 2521.100 1062.430 ;
        RECT 2520.900 1028.170 2521.160 1028.490 ;
        RECT 2521.360 1027.830 2521.620 1028.150 ;
        RECT 2521.420 1014.550 2521.560 1027.830 ;
        RECT 2520.900 1014.230 2521.160 1014.550 ;
        RECT 2521.360 1014.230 2521.620 1014.550 ;
        RECT 2520.960 1013.870 2521.100 1014.230 ;
        RECT 2520.900 1013.550 2521.160 1013.870 ;
        RECT 2522.280 1013.550 2522.540 1013.870 ;
        RECT 2522.340 931.330 2522.480 1013.550 ;
        RECT 2521.880 931.190 2522.480 931.330 ;
        RECT 2521.880 917.845 2522.020 931.190 ;
        RECT 2521.810 917.475 2522.090 917.845 ;
        RECT 2523.190 917.475 2523.470 917.845 ;
        RECT 2523.260 869.710 2523.400 917.475 ;
        RECT 2522.280 869.390 2522.540 869.710 ;
        RECT 2523.200 869.390 2523.460 869.710 ;
        RECT 2522.340 834.770 2522.480 869.390 ;
        RECT 2521.880 834.630 2522.480 834.770 ;
        RECT 2521.880 821.090 2522.020 834.630 ;
        RECT 2520.900 820.770 2521.160 821.090 ;
        RECT 2521.820 820.770 2522.080 821.090 ;
        RECT 2520.960 773.005 2521.100 820.770 ;
        RECT 2520.890 772.635 2521.170 773.005 ;
        RECT 2522.270 772.635 2522.550 773.005 ;
        RECT 2522.340 683.050 2522.480 772.635 ;
        RECT 2185.100 682.730 2185.360 683.050 ;
        RECT 2522.280 682.730 2522.540 683.050 ;
        RECT 2185.160 680.525 2185.300 682.730 ;
        RECT 2185.090 680.155 2185.370 680.525 ;
      LAYER via2 ;
        RECT 2899.930 1730.120 2900.210 1730.400 ;
        RECT 2521.350 1304.440 2521.630 1304.720 ;
        RECT 2522.730 1304.440 2523.010 1304.720 ;
        RECT 2521.810 917.520 2522.090 917.800 ;
        RECT 2523.190 917.520 2523.470 917.800 ;
        RECT 2520.890 772.680 2521.170 772.960 ;
        RECT 2522.270 772.680 2522.550 772.960 ;
        RECT 2185.090 680.200 2185.370 680.480 ;
      LAYER met3 ;
        RECT 2899.905 1730.410 2900.235 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2899.905 1730.110 2924.800 1730.410 ;
        RECT 2899.905 1730.095 2900.235 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2521.325 1304.730 2521.655 1304.745 ;
        RECT 2522.705 1304.730 2523.035 1304.745 ;
        RECT 2521.325 1304.430 2523.035 1304.730 ;
        RECT 2521.325 1304.415 2521.655 1304.430 ;
        RECT 2522.705 1304.415 2523.035 1304.430 ;
        RECT 2521.785 917.810 2522.115 917.825 ;
        RECT 2523.165 917.810 2523.495 917.825 ;
        RECT 2521.785 917.510 2523.495 917.810 ;
        RECT 2521.785 917.495 2522.115 917.510 ;
        RECT 2523.165 917.495 2523.495 917.510 ;
        RECT 2520.865 772.970 2521.195 772.985 ;
        RECT 2522.245 772.970 2522.575 772.985 ;
        RECT 2520.865 772.670 2522.575 772.970 ;
        RECT 2520.865 772.655 2521.195 772.670 ;
        RECT 2522.245 772.655 2522.575 772.670 ;
        RECT 2185.065 680.490 2185.395 680.505 ;
        RECT 2169.670 680.190 2185.395 680.490 ;
        RECT 2169.670 678.840 2169.970 680.190 ;
        RECT 2185.065 680.175 2185.395 680.190 ;
        RECT 2166.000 678.240 2170.000 678.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 689.760 2187.230 689.820 ;
        RECT 2902.670 689.760 2902.990 689.820 ;
        RECT 2186.910 689.620 2902.990 689.760 ;
        RECT 2186.910 689.560 2187.230 689.620 ;
        RECT 2902.670 689.560 2902.990 689.620 ;
      LAYER via ;
        RECT 2186.940 689.560 2187.200 689.820 ;
        RECT 2902.700 689.560 2902.960 689.820 ;
      LAYER met2 ;
        RECT 2902.690 1964.675 2902.970 1965.045 ;
        RECT 2902.760 689.850 2902.900 1964.675 ;
        RECT 2186.940 689.530 2187.200 689.850 ;
        RECT 2902.700 689.530 2902.960 689.850 ;
        RECT 2187.000 689.365 2187.140 689.530 ;
        RECT 2186.930 688.995 2187.210 689.365 ;
      LAYER via2 ;
        RECT 2902.690 1964.720 2902.970 1965.000 ;
        RECT 2186.930 689.040 2187.210 689.320 ;
      LAYER met3 ;
        RECT 2902.665 1965.010 2902.995 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2902.665 1964.710 2924.800 1965.010 ;
        RECT 2902.665 1964.695 2902.995 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2186.905 689.330 2187.235 689.345 ;
        RECT 2169.670 689.040 2187.235 689.330 ;
        RECT 2166.000 689.030 2187.235 689.040 ;
        RECT 2166.000 688.440 2170.000 689.030 ;
        RECT 2186.905 689.015 2187.235 689.030 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2183.690 2194.600 2184.010 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2183.690 2194.460 2901.150 2194.600 ;
        RECT 2183.690 2194.400 2184.010 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
      LAYER via ;
        RECT 2183.720 2194.400 2183.980 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2183.720 2194.370 2183.980 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2183.780 702.285 2183.920 2194.370 ;
        RECT 2183.710 701.915 2183.990 702.285 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2183.710 701.960 2183.990 702.240 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2183.685 702.250 2184.015 702.265 ;
        RECT 2169.670 701.950 2184.015 702.250 ;
        RECT 2169.670 699.920 2169.970 701.950 ;
        RECT 2183.685 701.935 2184.015 701.950 ;
        RECT 2166.000 699.320 2170.000 699.920 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 869.560 207.160 897.760 207.300 ;
        RECT 667.990 206.960 668.310 207.020 ;
        RECT 869.560 206.960 869.700 207.160 ;
        RECT 667.990 206.820 869.700 206.960 ;
        RECT 897.620 206.960 897.760 207.160 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 897.620 206.820 2901.150 206.960 ;
        RECT 667.990 206.760 668.310 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 668.020 206.760 668.280 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 668.010 801.875 668.290 802.245 ;
        RECT 668.080 207.050 668.220 801.875 ;
        RECT 668.020 206.730 668.280 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 668.010 801.920 668.290 802.200 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 667.985 802.210 668.315 802.225 ;
        RECT 670.000 802.210 674.000 802.600 ;
        RECT 667.985 802.000 674.000 802.210 ;
        RECT 667.985 801.910 670.220 802.000 ;
        RECT 667.985 801.895 668.315 801.910 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 661.090 1004.260 661.410 1004.320 ;
        RECT 2902.210 1004.260 2902.530 1004.320 ;
        RECT 661.090 1004.120 2902.530 1004.260 ;
        RECT 661.090 1004.060 661.410 1004.120 ;
        RECT 2902.210 1004.060 2902.530 1004.120 ;
      LAYER via ;
        RECT 661.120 1004.060 661.380 1004.320 ;
        RECT 2902.240 1004.060 2902.500 1004.320 ;
      LAYER met2 ;
        RECT 2902.230 2551.515 2902.510 2551.885 ;
        RECT 2902.300 1004.350 2902.440 2551.515 ;
        RECT 661.120 1004.030 661.380 1004.350 ;
        RECT 2902.240 1004.030 2902.500 1004.350 ;
        RECT 661.180 854.605 661.320 1004.030 ;
        RECT 661.110 854.235 661.390 854.605 ;
      LAYER via2 ;
        RECT 2902.230 2551.560 2902.510 2551.840 ;
        RECT 661.110 854.280 661.390 854.560 ;
      LAYER met3 ;
        RECT 2902.205 2551.850 2902.535 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2902.205 2551.550 2924.800 2551.850 ;
        RECT 2902.205 2551.535 2902.535 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 661.085 854.570 661.415 854.585 ;
        RECT 670.000 854.570 674.000 854.960 ;
        RECT 661.085 854.360 674.000 854.570 ;
        RECT 661.085 854.270 670.220 854.360 ;
        RECT 661.085 854.255 661.415 854.270 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 1004.600 662.330 1004.660 ;
        RECT 2901.290 1004.600 2901.610 1004.660 ;
        RECT 662.010 1004.460 2901.610 1004.600 ;
        RECT 662.010 1004.400 662.330 1004.460 ;
        RECT 2901.290 1004.400 2901.610 1004.460 ;
      LAYER via ;
        RECT 662.040 1004.400 662.300 1004.660 ;
        RECT 2901.320 1004.400 2901.580 1004.660 ;
      LAYER met2 ;
        RECT 2901.310 2786.115 2901.590 2786.485 ;
        RECT 2901.380 1004.690 2901.520 2786.115 ;
        RECT 662.040 1004.370 662.300 1004.690 ;
        RECT 2901.320 1004.370 2901.580 1004.690 ;
        RECT 662.100 860.045 662.240 1004.370 ;
        RECT 662.030 859.675 662.310 860.045 ;
      LAYER via2 ;
        RECT 2901.310 2786.160 2901.590 2786.440 ;
        RECT 662.030 859.720 662.310 860.000 ;
      LAYER met3 ;
        RECT 2901.285 2786.450 2901.615 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2901.285 2786.150 2924.800 2786.450 ;
        RECT 2901.285 2786.135 2901.615 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 662.005 860.010 662.335 860.025 ;
        RECT 670.000 860.010 674.000 860.400 ;
        RECT 662.005 859.800 674.000 860.010 ;
        RECT 662.005 859.710 670.220 859.800 ;
        RECT 662.005 859.695 662.335 859.710 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 785.310 3016.890 785.590 3017.005 ;
        RECT 786.230 3016.890 786.510 3017.005 ;
        RECT 785.310 3016.750 786.510 3016.890 ;
        RECT 785.310 3016.635 785.590 3016.750 ;
        RECT 786.230 3016.635 786.510 3016.750 ;
        RECT 855.230 3016.635 855.510 3017.005 ;
        RECT 855.300 3014.965 855.440 3016.635 ;
        RECT 855.230 3014.595 855.510 3014.965 ;
      LAYER via2 ;
        RECT 785.310 3016.680 785.590 3016.960 ;
        RECT 786.230 3016.680 786.510 3016.960 ;
        RECT 855.230 3016.680 855.510 3016.960 ;
        RECT 855.230 3014.640 855.510 3014.920 ;
      LAYER met3 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2916.710 3020.750 2924.800 3021.050 ;
        RECT 665.430 3016.970 665.810 3016.980 ;
        RECT 785.285 3016.970 785.615 3016.985 ;
        RECT 665.430 3016.670 785.615 3016.970 ;
        RECT 665.430 3016.660 665.810 3016.670 ;
        RECT 785.285 3016.655 785.615 3016.670 ;
        RECT 786.205 3016.970 786.535 3016.985 ;
        RECT 855.205 3016.970 855.535 3016.985 ;
        RECT 786.205 3016.670 797.330 3016.970 ;
        RECT 786.205 3016.655 786.535 3016.670 ;
        RECT 797.030 3016.290 797.330 3016.670 ;
        RECT 855.205 3016.670 904.050 3016.970 ;
        RECT 855.205 3016.655 855.535 3016.670 ;
        RECT 820.910 3016.290 821.290 3016.300 ;
        RECT 797.030 3015.990 821.290 3016.290 ;
        RECT 903.750 3016.290 904.050 3016.670 ;
        RECT 952.510 3016.670 1000.650 3016.970 ;
        RECT 903.750 3015.990 951.890 3016.290 ;
        RECT 820.910 3015.980 821.290 3015.990 ;
        RECT 951.590 3015.610 951.890 3015.990 ;
        RECT 952.510 3015.610 952.810 3016.670 ;
        RECT 1000.350 3016.290 1000.650 3016.670 ;
        RECT 1049.110 3016.670 1097.250 3016.970 ;
        RECT 1000.350 3015.990 1048.490 3016.290 ;
        RECT 951.590 3015.310 952.810 3015.610 ;
        RECT 1048.190 3015.610 1048.490 3015.990 ;
        RECT 1049.110 3015.610 1049.410 3016.670 ;
        RECT 1096.950 3016.290 1097.250 3016.670 ;
        RECT 1145.710 3016.670 1193.850 3016.970 ;
        RECT 1096.950 3015.990 1145.090 3016.290 ;
        RECT 1048.190 3015.310 1049.410 3015.610 ;
        RECT 1144.790 3015.610 1145.090 3015.990 ;
        RECT 1145.710 3015.610 1146.010 3016.670 ;
        RECT 1193.550 3016.290 1193.850 3016.670 ;
        RECT 1242.310 3016.670 1290.450 3016.970 ;
        RECT 1193.550 3015.990 1241.690 3016.290 ;
        RECT 1144.790 3015.310 1146.010 3015.610 ;
        RECT 1241.390 3015.610 1241.690 3015.990 ;
        RECT 1242.310 3015.610 1242.610 3016.670 ;
        RECT 1290.150 3016.290 1290.450 3016.670 ;
        RECT 1338.910 3016.670 1387.050 3016.970 ;
        RECT 1290.150 3015.990 1338.290 3016.290 ;
        RECT 1241.390 3015.310 1242.610 3015.610 ;
        RECT 1337.990 3015.610 1338.290 3015.990 ;
        RECT 1338.910 3015.610 1339.210 3016.670 ;
        RECT 1386.750 3016.290 1387.050 3016.670 ;
        RECT 1435.510 3016.670 1483.650 3016.970 ;
        RECT 1386.750 3015.990 1434.890 3016.290 ;
        RECT 1337.990 3015.310 1339.210 3015.610 ;
        RECT 1434.590 3015.610 1434.890 3015.990 ;
        RECT 1435.510 3015.610 1435.810 3016.670 ;
        RECT 1483.350 3016.290 1483.650 3016.670 ;
        RECT 1532.110 3016.670 1580.250 3016.970 ;
        RECT 1483.350 3015.990 1531.490 3016.290 ;
        RECT 1434.590 3015.310 1435.810 3015.610 ;
        RECT 1531.190 3015.610 1531.490 3015.990 ;
        RECT 1532.110 3015.610 1532.410 3016.670 ;
        RECT 1579.950 3016.290 1580.250 3016.670 ;
        RECT 1628.710 3016.670 1676.850 3016.970 ;
        RECT 1579.950 3015.990 1628.090 3016.290 ;
        RECT 1531.190 3015.310 1532.410 3015.610 ;
        RECT 1627.790 3015.610 1628.090 3015.990 ;
        RECT 1628.710 3015.610 1629.010 3016.670 ;
        RECT 1676.550 3016.290 1676.850 3016.670 ;
        RECT 1725.310 3016.670 1773.450 3016.970 ;
        RECT 1676.550 3015.990 1724.690 3016.290 ;
        RECT 1627.790 3015.310 1629.010 3015.610 ;
        RECT 1724.390 3015.610 1724.690 3015.990 ;
        RECT 1725.310 3015.610 1725.610 3016.670 ;
        RECT 1773.150 3016.290 1773.450 3016.670 ;
        RECT 1821.910 3016.670 1870.050 3016.970 ;
        RECT 1773.150 3015.990 1821.290 3016.290 ;
        RECT 1724.390 3015.310 1725.610 3015.610 ;
        RECT 1820.990 3015.610 1821.290 3015.990 ;
        RECT 1821.910 3015.610 1822.210 3016.670 ;
        RECT 1869.750 3016.290 1870.050 3016.670 ;
        RECT 1918.510 3016.670 1966.650 3016.970 ;
        RECT 1869.750 3015.990 1917.890 3016.290 ;
        RECT 1820.990 3015.310 1822.210 3015.610 ;
        RECT 1917.590 3015.610 1917.890 3015.990 ;
        RECT 1918.510 3015.610 1918.810 3016.670 ;
        RECT 1966.350 3016.290 1966.650 3016.670 ;
        RECT 2015.110 3016.670 2063.250 3016.970 ;
        RECT 1966.350 3015.990 2014.490 3016.290 ;
        RECT 1917.590 3015.310 1918.810 3015.610 ;
        RECT 2014.190 3015.610 2014.490 3015.990 ;
        RECT 2015.110 3015.610 2015.410 3016.670 ;
        RECT 2062.950 3016.290 2063.250 3016.670 ;
        RECT 2111.710 3016.670 2159.850 3016.970 ;
        RECT 2062.950 3015.990 2111.090 3016.290 ;
        RECT 2014.190 3015.310 2015.410 3015.610 ;
        RECT 2110.790 3015.610 2111.090 3015.990 ;
        RECT 2111.710 3015.610 2112.010 3016.670 ;
        RECT 2159.550 3016.290 2159.850 3016.670 ;
        RECT 2208.310 3016.670 2256.450 3016.970 ;
        RECT 2159.550 3015.990 2207.690 3016.290 ;
        RECT 2110.790 3015.310 2112.010 3015.610 ;
        RECT 2207.390 3015.610 2207.690 3015.990 ;
        RECT 2208.310 3015.610 2208.610 3016.670 ;
        RECT 2256.150 3016.290 2256.450 3016.670 ;
        RECT 2304.910 3016.670 2353.050 3016.970 ;
        RECT 2256.150 3015.990 2304.290 3016.290 ;
        RECT 2207.390 3015.310 2208.610 3015.610 ;
        RECT 2303.990 3015.610 2304.290 3015.990 ;
        RECT 2304.910 3015.610 2305.210 3016.670 ;
        RECT 2352.750 3016.290 2353.050 3016.670 ;
        RECT 2401.510 3016.670 2449.650 3016.970 ;
        RECT 2352.750 3015.990 2400.890 3016.290 ;
        RECT 2303.990 3015.310 2305.210 3015.610 ;
        RECT 2400.590 3015.610 2400.890 3015.990 ;
        RECT 2401.510 3015.610 2401.810 3016.670 ;
        RECT 2449.350 3016.290 2449.650 3016.670 ;
        RECT 2498.110 3016.670 2546.250 3016.970 ;
        RECT 2449.350 3015.990 2497.490 3016.290 ;
        RECT 2400.590 3015.310 2401.810 3015.610 ;
        RECT 2497.190 3015.610 2497.490 3015.990 ;
        RECT 2498.110 3015.610 2498.410 3016.670 ;
        RECT 2545.950 3016.290 2546.250 3016.670 ;
        RECT 2594.710 3016.670 2642.850 3016.970 ;
        RECT 2545.950 3015.990 2594.090 3016.290 ;
        RECT 2497.190 3015.310 2498.410 3015.610 ;
        RECT 2593.790 3015.610 2594.090 3015.990 ;
        RECT 2594.710 3015.610 2595.010 3016.670 ;
        RECT 2642.550 3016.290 2642.850 3016.670 ;
        RECT 2691.310 3016.670 2739.450 3016.970 ;
        RECT 2642.550 3015.990 2690.690 3016.290 ;
        RECT 2593.790 3015.310 2595.010 3015.610 ;
        RECT 2690.390 3015.610 2690.690 3015.990 ;
        RECT 2691.310 3015.610 2691.610 3016.670 ;
        RECT 2739.150 3016.290 2739.450 3016.670 ;
        RECT 2787.910 3016.670 2836.050 3016.970 ;
        RECT 2739.150 3015.990 2787.290 3016.290 ;
        RECT 2690.390 3015.310 2691.610 3015.610 ;
        RECT 2786.990 3015.610 2787.290 3015.990 ;
        RECT 2787.910 3015.610 2788.210 3016.670 ;
        RECT 2835.750 3016.290 2836.050 3016.670 ;
        RECT 2916.710 3016.290 2917.010 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2835.750 3015.990 2883.890 3016.290 ;
        RECT 2786.990 3015.310 2788.210 3015.610 ;
        RECT 2883.590 3015.610 2883.890 3015.990 ;
        RECT 2884.510 3015.990 2917.010 3016.290 ;
        RECT 2884.510 3015.610 2884.810 3015.990 ;
        RECT 2883.590 3015.310 2884.810 3015.610 ;
        RECT 820.910 3014.930 821.290 3014.940 ;
        RECT 855.205 3014.930 855.535 3014.945 ;
        RECT 820.910 3014.630 855.535 3014.930 ;
        RECT 820.910 3014.620 821.290 3014.630 ;
        RECT 855.205 3014.615 855.535 3014.630 ;
        RECT 665.430 864.770 665.810 864.780 ;
        RECT 670.000 864.770 674.000 865.160 ;
        RECT 665.430 864.560 674.000 864.770 ;
        RECT 665.430 864.470 670.220 864.560 ;
        RECT 665.430 864.460 665.810 864.470 ;
      LAYER via3 ;
        RECT 665.460 3016.660 665.780 3016.980 ;
        RECT 820.940 3015.980 821.260 3016.300 ;
        RECT 820.940 3014.620 821.260 3014.940 ;
        RECT 665.460 864.460 665.780 864.780 ;
      LAYER met4 ;
        RECT 665.455 3016.655 665.785 3016.985 ;
        RECT 665.470 864.785 665.770 3016.655 ;
        RECT 820.935 3015.975 821.265 3016.305 ;
        RECT 820.950 3014.945 821.250 3015.975 ;
        RECT 820.935 3014.615 821.265 3014.945 ;
        RECT 665.455 864.455 665.785 864.785 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 772.870 3252.000 773.190 3252.060 ;
        RECT 797.250 3252.000 797.570 3252.060 ;
        RECT 772.870 3251.860 797.570 3252.000 ;
        RECT 772.870 3251.800 773.190 3251.860 ;
        RECT 797.250 3251.800 797.570 3251.860 ;
        RECT 676.270 3251.320 676.590 3251.380 ;
        RECT 714.450 3251.320 714.770 3251.380 ;
        RECT 676.270 3251.180 714.770 3251.320 ;
        RECT 676.270 3251.120 676.590 3251.180 ;
        RECT 714.450 3251.120 714.770 3251.180 ;
      LAYER via ;
        RECT 772.900 3251.800 773.160 3252.060 ;
        RECT 797.280 3251.800 797.540 3252.060 ;
        RECT 676.300 3251.120 676.560 3251.380 ;
        RECT 714.480 3251.120 714.740 3251.380 ;
      LAYER met2 ;
        RECT 845.110 3252.595 845.390 3252.965 ;
        RECT 738.850 3252.170 739.130 3252.285 ;
        RECT 738.000 3252.030 739.130 3252.170 ;
        RECT 676.290 3251.235 676.570 3251.605 ;
        RECT 676.300 3251.090 676.560 3251.235 ;
        RECT 714.480 3251.090 714.740 3251.410 ;
        RECT 714.540 3250.245 714.680 3251.090 ;
        RECT 738.000 3250.925 738.140 3252.030 ;
        RECT 738.850 3251.915 739.130 3252.030 ;
        RECT 772.890 3251.915 773.170 3252.285 ;
        RECT 772.900 3251.770 773.160 3251.915 ;
        RECT 797.280 3251.770 797.540 3252.090 ;
        RECT 797.340 3251.605 797.480 3251.770 ;
        RECT 845.180 3251.605 845.320 3252.595 ;
        RECT 797.270 3251.235 797.550 3251.605 ;
        RECT 845.110 3251.235 845.390 3251.605 ;
        RECT 737.930 3250.555 738.210 3250.925 ;
        RECT 714.470 3249.875 714.750 3250.245 ;
      LAYER via2 ;
        RECT 845.110 3252.640 845.390 3252.920 ;
        RECT 676.290 3251.280 676.570 3251.560 ;
        RECT 738.850 3251.960 739.130 3252.240 ;
        RECT 772.890 3251.960 773.170 3252.240 ;
        RECT 797.270 3251.280 797.550 3251.560 ;
        RECT 845.110 3251.280 845.390 3251.560 ;
        RECT 737.930 3250.600 738.210 3250.880 ;
        RECT 714.470 3249.920 714.750 3250.200 ;
      LAYER met3 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2916.710 3255.350 2924.800 3255.650 ;
        RECT 820.910 3252.930 821.290 3252.940 ;
        RECT 845.085 3252.930 845.415 3252.945 ;
        RECT 820.910 3252.630 845.415 3252.930 ;
        RECT 820.910 3252.620 821.290 3252.630 ;
        RECT 845.085 3252.615 845.415 3252.630 ;
        RECT 738.825 3252.250 739.155 3252.265 ;
        RECT 772.865 3252.250 773.195 3252.265 ;
        RECT 738.825 3251.950 773.195 3252.250 ;
        RECT 738.825 3251.935 739.155 3251.950 ;
        RECT 772.865 3251.935 773.195 3251.950 ;
        RECT 667.270 3251.570 667.650 3251.580 ;
        RECT 676.265 3251.570 676.595 3251.585 ;
        RECT 667.270 3251.270 676.595 3251.570 ;
        RECT 667.270 3251.260 667.650 3251.270 ;
        RECT 676.265 3251.255 676.595 3251.270 ;
        RECT 797.245 3251.570 797.575 3251.585 ;
        RECT 820.910 3251.570 821.290 3251.580 ;
        RECT 797.245 3251.270 821.290 3251.570 ;
        RECT 797.245 3251.255 797.575 3251.270 ;
        RECT 820.910 3251.260 821.290 3251.270 ;
        RECT 845.085 3251.570 845.415 3251.585 ;
        RECT 845.085 3251.270 904.050 3251.570 ;
        RECT 845.085 3251.255 845.415 3251.270 ;
        RECT 737.905 3250.890 738.235 3250.905 ;
        RECT 724.350 3250.590 738.235 3250.890 ;
        RECT 903.750 3250.890 904.050 3251.270 ;
        RECT 952.510 3251.270 1000.650 3251.570 ;
        RECT 903.750 3250.590 951.890 3250.890 ;
        RECT 714.445 3250.210 714.775 3250.225 ;
        RECT 724.350 3250.210 724.650 3250.590 ;
        RECT 737.905 3250.575 738.235 3250.590 ;
        RECT 714.445 3249.910 724.650 3250.210 ;
        RECT 951.590 3250.210 951.890 3250.590 ;
        RECT 952.510 3250.210 952.810 3251.270 ;
        RECT 1000.350 3250.890 1000.650 3251.270 ;
        RECT 1049.110 3251.270 1097.250 3251.570 ;
        RECT 1000.350 3250.590 1048.490 3250.890 ;
        RECT 951.590 3249.910 952.810 3250.210 ;
        RECT 1048.190 3250.210 1048.490 3250.590 ;
        RECT 1049.110 3250.210 1049.410 3251.270 ;
        RECT 1096.950 3250.890 1097.250 3251.270 ;
        RECT 1145.710 3251.270 1193.850 3251.570 ;
        RECT 1096.950 3250.590 1145.090 3250.890 ;
        RECT 1048.190 3249.910 1049.410 3250.210 ;
        RECT 1144.790 3250.210 1145.090 3250.590 ;
        RECT 1145.710 3250.210 1146.010 3251.270 ;
        RECT 1193.550 3250.890 1193.850 3251.270 ;
        RECT 1242.310 3251.270 1290.450 3251.570 ;
        RECT 1193.550 3250.590 1241.690 3250.890 ;
        RECT 1144.790 3249.910 1146.010 3250.210 ;
        RECT 1241.390 3250.210 1241.690 3250.590 ;
        RECT 1242.310 3250.210 1242.610 3251.270 ;
        RECT 1290.150 3250.890 1290.450 3251.270 ;
        RECT 1338.910 3251.270 1387.050 3251.570 ;
        RECT 1290.150 3250.590 1338.290 3250.890 ;
        RECT 1241.390 3249.910 1242.610 3250.210 ;
        RECT 1337.990 3250.210 1338.290 3250.590 ;
        RECT 1338.910 3250.210 1339.210 3251.270 ;
        RECT 1386.750 3250.890 1387.050 3251.270 ;
        RECT 1435.510 3251.270 1483.650 3251.570 ;
        RECT 1386.750 3250.590 1434.890 3250.890 ;
        RECT 1337.990 3249.910 1339.210 3250.210 ;
        RECT 1434.590 3250.210 1434.890 3250.590 ;
        RECT 1435.510 3250.210 1435.810 3251.270 ;
        RECT 1483.350 3250.890 1483.650 3251.270 ;
        RECT 1532.110 3251.270 1580.250 3251.570 ;
        RECT 1483.350 3250.590 1531.490 3250.890 ;
        RECT 1434.590 3249.910 1435.810 3250.210 ;
        RECT 1531.190 3250.210 1531.490 3250.590 ;
        RECT 1532.110 3250.210 1532.410 3251.270 ;
        RECT 1579.950 3250.890 1580.250 3251.270 ;
        RECT 1628.710 3251.270 1676.850 3251.570 ;
        RECT 1579.950 3250.590 1628.090 3250.890 ;
        RECT 1531.190 3249.910 1532.410 3250.210 ;
        RECT 1627.790 3250.210 1628.090 3250.590 ;
        RECT 1628.710 3250.210 1629.010 3251.270 ;
        RECT 1676.550 3250.890 1676.850 3251.270 ;
        RECT 1725.310 3251.270 1773.450 3251.570 ;
        RECT 1676.550 3250.590 1724.690 3250.890 ;
        RECT 1627.790 3249.910 1629.010 3250.210 ;
        RECT 1724.390 3250.210 1724.690 3250.590 ;
        RECT 1725.310 3250.210 1725.610 3251.270 ;
        RECT 1773.150 3250.890 1773.450 3251.270 ;
        RECT 1821.910 3251.270 1870.050 3251.570 ;
        RECT 1773.150 3250.590 1821.290 3250.890 ;
        RECT 1724.390 3249.910 1725.610 3250.210 ;
        RECT 1820.990 3250.210 1821.290 3250.590 ;
        RECT 1821.910 3250.210 1822.210 3251.270 ;
        RECT 1869.750 3250.890 1870.050 3251.270 ;
        RECT 1918.510 3251.270 1966.650 3251.570 ;
        RECT 1869.750 3250.590 1917.890 3250.890 ;
        RECT 1820.990 3249.910 1822.210 3250.210 ;
        RECT 1917.590 3250.210 1917.890 3250.590 ;
        RECT 1918.510 3250.210 1918.810 3251.270 ;
        RECT 1966.350 3250.890 1966.650 3251.270 ;
        RECT 2015.110 3251.270 2063.250 3251.570 ;
        RECT 1966.350 3250.590 2014.490 3250.890 ;
        RECT 1917.590 3249.910 1918.810 3250.210 ;
        RECT 2014.190 3250.210 2014.490 3250.590 ;
        RECT 2015.110 3250.210 2015.410 3251.270 ;
        RECT 2062.950 3250.890 2063.250 3251.270 ;
        RECT 2111.710 3251.270 2159.850 3251.570 ;
        RECT 2062.950 3250.590 2111.090 3250.890 ;
        RECT 2014.190 3249.910 2015.410 3250.210 ;
        RECT 2110.790 3250.210 2111.090 3250.590 ;
        RECT 2111.710 3250.210 2112.010 3251.270 ;
        RECT 2159.550 3250.890 2159.850 3251.270 ;
        RECT 2208.310 3251.270 2256.450 3251.570 ;
        RECT 2159.550 3250.590 2207.690 3250.890 ;
        RECT 2110.790 3249.910 2112.010 3250.210 ;
        RECT 2207.390 3250.210 2207.690 3250.590 ;
        RECT 2208.310 3250.210 2208.610 3251.270 ;
        RECT 2256.150 3250.890 2256.450 3251.270 ;
        RECT 2304.910 3251.270 2353.050 3251.570 ;
        RECT 2256.150 3250.590 2304.290 3250.890 ;
        RECT 2207.390 3249.910 2208.610 3250.210 ;
        RECT 2303.990 3250.210 2304.290 3250.590 ;
        RECT 2304.910 3250.210 2305.210 3251.270 ;
        RECT 2352.750 3250.890 2353.050 3251.270 ;
        RECT 2401.510 3251.270 2449.650 3251.570 ;
        RECT 2352.750 3250.590 2400.890 3250.890 ;
        RECT 2303.990 3249.910 2305.210 3250.210 ;
        RECT 2400.590 3250.210 2400.890 3250.590 ;
        RECT 2401.510 3250.210 2401.810 3251.270 ;
        RECT 2449.350 3250.890 2449.650 3251.270 ;
        RECT 2498.110 3251.270 2546.250 3251.570 ;
        RECT 2449.350 3250.590 2497.490 3250.890 ;
        RECT 2400.590 3249.910 2401.810 3250.210 ;
        RECT 2497.190 3250.210 2497.490 3250.590 ;
        RECT 2498.110 3250.210 2498.410 3251.270 ;
        RECT 2545.950 3250.890 2546.250 3251.270 ;
        RECT 2594.710 3251.270 2642.850 3251.570 ;
        RECT 2545.950 3250.590 2594.090 3250.890 ;
        RECT 2497.190 3249.910 2498.410 3250.210 ;
        RECT 2593.790 3250.210 2594.090 3250.590 ;
        RECT 2594.710 3250.210 2595.010 3251.270 ;
        RECT 2642.550 3250.890 2642.850 3251.270 ;
        RECT 2691.310 3251.270 2739.450 3251.570 ;
        RECT 2642.550 3250.590 2690.690 3250.890 ;
        RECT 2593.790 3249.910 2595.010 3250.210 ;
        RECT 2690.390 3250.210 2690.690 3250.590 ;
        RECT 2691.310 3250.210 2691.610 3251.270 ;
        RECT 2739.150 3250.890 2739.450 3251.270 ;
        RECT 2787.910 3251.270 2836.050 3251.570 ;
        RECT 2739.150 3250.590 2787.290 3250.890 ;
        RECT 2690.390 3249.910 2691.610 3250.210 ;
        RECT 2786.990 3250.210 2787.290 3250.590 ;
        RECT 2787.910 3250.210 2788.210 3251.270 ;
        RECT 2835.750 3250.890 2836.050 3251.270 ;
        RECT 2916.710 3250.890 2917.010 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2835.750 3250.590 2883.890 3250.890 ;
        RECT 2786.990 3249.910 2788.210 3250.210 ;
        RECT 2883.590 3250.210 2883.890 3250.590 ;
        RECT 2884.510 3250.590 2917.010 3250.890 ;
        RECT 2884.510 3250.210 2884.810 3250.590 ;
        RECT 2883.590 3249.910 2884.810 3250.210 ;
        RECT 714.445 3249.895 714.775 3249.910 ;
        RECT 667.270 870.210 667.650 870.220 ;
        RECT 670.000 870.210 674.000 870.600 ;
        RECT 667.270 870.000 674.000 870.210 ;
        RECT 667.270 869.910 670.220 870.000 ;
        RECT 667.270 869.900 667.650 869.910 ;
      LAYER via3 ;
        RECT 820.940 3252.620 821.260 3252.940 ;
        RECT 667.300 3251.260 667.620 3251.580 ;
        RECT 820.940 3251.260 821.260 3251.580 ;
        RECT 667.300 869.900 667.620 870.220 ;
      LAYER met4 ;
        RECT 820.935 3252.615 821.265 3252.945 ;
        RECT 820.950 3251.585 821.250 3252.615 ;
        RECT 667.295 3251.255 667.625 3251.585 ;
        RECT 820.935 3251.255 821.265 3251.585 ;
        RECT 667.310 870.225 667.610 3251.255 ;
        RECT 667.295 869.895 667.625 870.225 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 737.910 3485.580 738.230 3485.640 ;
        RECT 772.410 3485.580 772.730 3485.640 ;
        RECT 737.910 3485.440 772.730 3485.580 ;
        RECT 737.910 3485.380 738.230 3485.440 ;
        RECT 772.410 3485.380 772.730 3485.440 ;
        RECT 834.510 3485.580 834.830 3485.640 ;
        RECT 869.010 3485.580 869.330 3485.640 ;
        RECT 834.510 3485.440 869.330 3485.580 ;
        RECT 834.510 3485.380 834.830 3485.440 ;
        RECT 869.010 3485.380 869.330 3485.440 ;
        RECT 931.110 3485.580 931.430 3485.640 ;
        RECT 965.610 3485.580 965.930 3485.640 ;
        RECT 931.110 3485.440 965.930 3485.580 ;
        RECT 931.110 3485.380 931.430 3485.440 ;
        RECT 965.610 3485.380 965.930 3485.440 ;
        RECT 1027.710 3485.580 1028.030 3485.640 ;
        RECT 1062.210 3485.580 1062.530 3485.640 ;
        RECT 1027.710 3485.440 1062.530 3485.580 ;
        RECT 1027.710 3485.380 1028.030 3485.440 ;
        RECT 1062.210 3485.380 1062.530 3485.440 ;
        RECT 1124.310 3485.580 1124.630 3485.640 ;
        RECT 1158.810 3485.580 1159.130 3485.640 ;
        RECT 1124.310 3485.440 1159.130 3485.580 ;
        RECT 1124.310 3485.380 1124.630 3485.440 ;
        RECT 1158.810 3485.380 1159.130 3485.440 ;
        RECT 1220.910 3485.580 1221.230 3485.640 ;
        RECT 1255.410 3485.580 1255.730 3485.640 ;
        RECT 1220.910 3485.440 1255.730 3485.580 ;
        RECT 1220.910 3485.380 1221.230 3485.440 ;
        RECT 1255.410 3485.380 1255.730 3485.440 ;
        RECT 1317.510 3485.580 1317.830 3485.640 ;
        RECT 1352.010 3485.580 1352.330 3485.640 ;
        RECT 1317.510 3485.440 1352.330 3485.580 ;
        RECT 1317.510 3485.380 1317.830 3485.440 ;
        RECT 1352.010 3485.380 1352.330 3485.440 ;
        RECT 1414.110 3485.580 1414.430 3485.640 ;
        RECT 1448.610 3485.580 1448.930 3485.640 ;
        RECT 1414.110 3485.440 1448.930 3485.580 ;
        RECT 1414.110 3485.380 1414.430 3485.440 ;
        RECT 1448.610 3485.380 1448.930 3485.440 ;
        RECT 1510.710 3485.580 1511.030 3485.640 ;
        RECT 1545.210 3485.580 1545.530 3485.640 ;
        RECT 1510.710 3485.440 1545.530 3485.580 ;
        RECT 1510.710 3485.380 1511.030 3485.440 ;
        RECT 1545.210 3485.380 1545.530 3485.440 ;
        RECT 1607.310 3485.580 1607.630 3485.640 ;
        RECT 1641.810 3485.580 1642.130 3485.640 ;
        RECT 1607.310 3485.440 1642.130 3485.580 ;
        RECT 1607.310 3485.380 1607.630 3485.440 ;
        RECT 1641.810 3485.380 1642.130 3485.440 ;
      LAYER via ;
        RECT 737.940 3485.380 738.200 3485.640 ;
        RECT 772.440 3485.380 772.700 3485.640 ;
        RECT 834.540 3485.380 834.800 3485.640 ;
        RECT 869.040 3485.380 869.300 3485.640 ;
        RECT 931.140 3485.380 931.400 3485.640 ;
        RECT 965.640 3485.380 965.900 3485.640 ;
        RECT 1027.740 3485.380 1028.000 3485.640 ;
        RECT 1062.240 3485.380 1062.500 3485.640 ;
        RECT 1124.340 3485.380 1124.600 3485.640 ;
        RECT 1158.840 3485.380 1159.100 3485.640 ;
        RECT 1220.940 3485.380 1221.200 3485.640 ;
        RECT 1255.440 3485.380 1255.700 3485.640 ;
        RECT 1317.540 3485.380 1317.800 3485.640 ;
        RECT 1352.040 3485.380 1352.300 3485.640 ;
        RECT 1414.140 3485.380 1414.400 3485.640 ;
        RECT 1448.640 3485.380 1448.900 3485.640 ;
        RECT 1510.740 3485.380 1511.000 3485.640 ;
        RECT 1545.240 3485.380 1545.500 3485.640 ;
        RECT 1607.340 3485.380 1607.600 3485.640 ;
        RECT 1641.840 3485.380 1642.100 3485.640 ;
      LAYER met2 ;
        RECT 772.430 3485.835 772.710 3486.205 ;
        RECT 869.030 3485.835 869.310 3486.205 ;
        RECT 965.630 3485.835 965.910 3486.205 ;
        RECT 1062.230 3485.835 1062.510 3486.205 ;
        RECT 1158.830 3485.835 1159.110 3486.205 ;
        RECT 1255.430 3485.835 1255.710 3486.205 ;
        RECT 1352.030 3485.835 1352.310 3486.205 ;
        RECT 1448.630 3485.835 1448.910 3486.205 ;
        RECT 1545.230 3485.835 1545.510 3486.205 ;
        RECT 1641.830 3485.835 1642.110 3486.205 ;
        RECT 772.500 3485.670 772.640 3485.835 ;
        RECT 869.100 3485.670 869.240 3485.835 ;
        RECT 965.700 3485.670 965.840 3485.835 ;
        RECT 1062.300 3485.670 1062.440 3485.835 ;
        RECT 1158.900 3485.670 1159.040 3485.835 ;
        RECT 1255.500 3485.670 1255.640 3485.835 ;
        RECT 1352.100 3485.670 1352.240 3485.835 ;
        RECT 1448.700 3485.670 1448.840 3485.835 ;
        RECT 1545.300 3485.670 1545.440 3485.835 ;
        RECT 1641.900 3485.670 1642.040 3485.835 ;
        RECT 737.940 3485.525 738.200 3485.670 ;
        RECT 737.930 3485.155 738.210 3485.525 ;
        RECT 772.440 3485.350 772.700 3485.670 ;
        RECT 834.540 3485.525 834.800 3485.670 ;
        RECT 834.530 3485.155 834.810 3485.525 ;
        RECT 869.040 3485.350 869.300 3485.670 ;
        RECT 931.140 3485.525 931.400 3485.670 ;
        RECT 931.130 3485.155 931.410 3485.525 ;
        RECT 965.640 3485.350 965.900 3485.670 ;
        RECT 1027.740 3485.525 1028.000 3485.670 ;
        RECT 1027.730 3485.155 1028.010 3485.525 ;
        RECT 1062.240 3485.350 1062.500 3485.670 ;
        RECT 1124.340 3485.525 1124.600 3485.670 ;
        RECT 1124.330 3485.155 1124.610 3485.525 ;
        RECT 1158.840 3485.350 1159.100 3485.670 ;
        RECT 1220.940 3485.525 1221.200 3485.670 ;
        RECT 1220.930 3485.155 1221.210 3485.525 ;
        RECT 1255.440 3485.350 1255.700 3485.670 ;
        RECT 1317.540 3485.525 1317.800 3485.670 ;
        RECT 1317.530 3485.155 1317.810 3485.525 ;
        RECT 1352.040 3485.350 1352.300 3485.670 ;
        RECT 1414.140 3485.525 1414.400 3485.670 ;
        RECT 1414.130 3485.155 1414.410 3485.525 ;
        RECT 1448.640 3485.350 1448.900 3485.670 ;
        RECT 1510.740 3485.525 1511.000 3485.670 ;
        RECT 1510.730 3485.155 1511.010 3485.525 ;
        RECT 1545.240 3485.350 1545.500 3485.670 ;
        RECT 1607.340 3485.525 1607.600 3485.670 ;
        RECT 1607.330 3485.155 1607.610 3485.525 ;
        RECT 1641.840 3485.350 1642.100 3485.670 ;
      LAYER via2 ;
        RECT 772.430 3485.880 772.710 3486.160 ;
        RECT 869.030 3485.880 869.310 3486.160 ;
        RECT 965.630 3485.880 965.910 3486.160 ;
        RECT 1062.230 3485.880 1062.510 3486.160 ;
        RECT 1158.830 3485.880 1159.110 3486.160 ;
        RECT 1255.430 3485.880 1255.710 3486.160 ;
        RECT 1352.030 3485.880 1352.310 3486.160 ;
        RECT 1448.630 3485.880 1448.910 3486.160 ;
        RECT 1545.230 3485.880 1545.510 3486.160 ;
        RECT 1641.830 3485.880 1642.110 3486.160 ;
        RECT 737.930 3485.200 738.210 3485.480 ;
        RECT 834.530 3485.200 834.810 3485.480 ;
        RECT 931.130 3485.200 931.410 3485.480 ;
        RECT 1027.730 3485.200 1028.010 3485.480 ;
        RECT 1124.330 3485.200 1124.610 3485.480 ;
        RECT 1220.930 3485.200 1221.210 3485.480 ;
        RECT 1317.530 3485.200 1317.810 3485.480 ;
        RECT 1414.130 3485.200 1414.410 3485.480 ;
        RECT 1510.730 3485.200 1511.010 3485.480 ;
        RECT 1607.330 3485.200 1607.610 3485.480 ;
      LAYER met3 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2916.710 3489.950 2924.800 3490.250 ;
        RECT 668.190 3486.170 668.570 3486.180 ;
        RECT 772.405 3486.170 772.735 3486.185 ;
        RECT 869.005 3486.170 869.335 3486.185 ;
        RECT 965.605 3486.170 965.935 3486.185 ;
        RECT 1062.205 3486.170 1062.535 3486.185 ;
        RECT 1158.805 3486.170 1159.135 3486.185 ;
        RECT 1255.405 3486.170 1255.735 3486.185 ;
        RECT 1352.005 3486.170 1352.335 3486.185 ;
        RECT 1448.605 3486.170 1448.935 3486.185 ;
        RECT 1545.205 3486.170 1545.535 3486.185 ;
        RECT 1641.805 3486.170 1642.135 3486.185 ;
        RECT 668.190 3485.870 690.610 3486.170 ;
        RECT 668.190 3485.860 668.570 3485.870 ;
        RECT 690.310 3485.490 690.610 3485.870 ;
        RECT 772.405 3485.870 787.210 3486.170 ;
        RECT 772.405 3485.855 772.735 3485.870 ;
        RECT 737.905 3485.490 738.235 3485.505 ;
        RECT 690.310 3485.190 738.235 3485.490 ;
        RECT 786.910 3485.490 787.210 3485.870 ;
        RECT 869.005 3485.870 883.810 3486.170 ;
        RECT 869.005 3485.855 869.335 3485.870 ;
        RECT 834.505 3485.490 834.835 3485.505 ;
        RECT 786.910 3485.190 834.835 3485.490 ;
        RECT 883.510 3485.490 883.810 3485.870 ;
        RECT 965.605 3485.870 980.410 3486.170 ;
        RECT 965.605 3485.855 965.935 3485.870 ;
        RECT 931.105 3485.490 931.435 3485.505 ;
        RECT 883.510 3485.190 931.435 3485.490 ;
        RECT 980.110 3485.490 980.410 3485.870 ;
        RECT 1062.205 3485.870 1077.010 3486.170 ;
        RECT 1062.205 3485.855 1062.535 3485.870 ;
        RECT 1027.705 3485.490 1028.035 3485.505 ;
        RECT 980.110 3485.190 1028.035 3485.490 ;
        RECT 1076.710 3485.490 1077.010 3485.870 ;
        RECT 1158.805 3485.870 1173.610 3486.170 ;
        RECT 1158.805 3485.855 1159.135 3485.870 ;
        RECT 1124.305 3485.490 1124.635 3485.505 ;
        RECT 1076.710 3485.190 1124.635 3485.490 ;
        RECT 1173.310 3485.490 1173.610 3485.870 ;
        RECT 1255.405 3485.870 1270.210 3486.170 ;
        RECT 1255.405 3485.855 1255.735 3485.870 ;
        RECT 1220.905 3485.490 1221.235 3485.505 ;
        RECT 1173.310 3485.190 1221.235 3485.490 ;
        RECT 1269.910 3485.490 1270.210 3485.870 ;
        RECT 1352.005 3485.870 1366.810 3486.170 ;
        RECT 1352.005 3485.855 1352.335 3485.870 ;
        RECT 1317.505 3485.490 1317.835 3485.505 ;
        RECT 1269.910 3485.190 1317.835 3485.490 ;
        RECT 1366.510 3485.490 1366.810 3485.870 ;
        RECT 1448.605 3485.870 1463.410 3486.170 ;
        RECT 1448.605 3485.855 1448.935 3485.870 ;
        RECT 1414.105 3485.490 1414.435 3485.505 ;
        RECT 1366.510 3485.190 1414.435 3485.490 ;
        RECT 1463.110 3485.490 1463.410 3485.870 ;
        RECT 1545.205 3485.870 1560.010 3486.170 ;
        RECT 1545.205 3485.855 1545.535 3485.870 ;
        RECT 1510.705 3485.490 1511.035 3485.505 ;
        RECT 1463.110 3485.190 1511.035 3485.490 ;
        RECT 1559.710 3485.490 1560.010 3485.870 ;
        RECT 1641.805 3485.870 1704.450 3486.170 ;
        RECT 1641.805 3485.855 1642.135 3485.870 ;
        RECT 1607.305 3485.490 1607.635 3485.505 ;
        RECT 1559.710 3485.190 1607.635 3485.490 ;
        RECT 1704.150 3485.490 1704.450 3485.870 ;
        RECT 1773.150 3485.870 1801.050 3486.170 ;
        RECT 1704.150 3485.190 1752.290 3485.490 ;
        RECT 737.905 3485.175 738.235 3485.190 ;
        RECT 834.505 3485.175 834.835 3485.190 ;
        RECT 931.105 3485.175 931.435 3485.190 ;
        RECT 1027.705 3485.175 1028.035 3485.190 ;
        RECT 1124.305 3485.175 1124.635 3485.190 ;
        RECT 1220.905 3485.175 1221.235 3485.190 ;
        RECT 1317.505 3485.175 1317.835 3485.190 ;
        RECT 1414.105 3485.175 1414.435 3485.190 ;
        RECT 1510.705 3485.175 1511.035 3485.190 ;
        RECT 1607.305 3485.175 1607.635 3485.190 ;
        RECT 1751.990 3484.810 1752.290 3485.190 ;
        RECT 1773.150 3484.810 1773.450 3485.870 ;
        RECT 1800.750 3485.490 1801.050 3485.870 ;
        RECT 1869.750 3485.870 1917.890 3486.170 ;
        RECT 1800.750 3485.190 1848.890 3485.490 ;
        RECT 1751.990 3484.510 1773.450 3484.810 ;
        RECT 1848.590 3484.810 1848.890 3485.190 ;
        RECT 1869.750 3484.810 1870.050 3485.870 ;
        RECT 1848.590 3484.510 1870.050 3484.810 ;
        RECT 1917.590 3484.810 1917.890 3485.870 ;
        RECT 1918.510 3485.870 1966.650 3486.170 ;
        RECT 1918.510 3484.810 1918.810 3485.870 ;
        RECT 1966.350 3485.490 1966.650 3485.870 ;
        RECT 2015.110 3485.870 2063.250 3486.170 ;
        RECT 1966.350 3485.190 2014.490 3485.490 ;
        RECT 1917.590 3484.510 1918.810 3484.810 ;
        RECT 2014.190 3484.810 2014.490 3485.190 ;
        RECT 2015.110 3484.810 2015.410 3485.870 ;
        RECT 2062.950 3485.490 2063.250 3485.870 ;
        RECT 2111.710 3485.870 2159.850 3486.170 ;
        RECT 2062.950 3485.190 2111.090 3485.490 ;
        RECT 2014.190 3484.510 2015.410 3484.810 ;
        RECT 2110.790 3484.810 2111.090 3485.190 ;
        RECT 2111.710 3484.810 2112.010 3485.870 ;
        RECT 2159.550 3485.490 2159.850 3485.870 ;
        RECT 2208.310 3485.870 2256.450 3486.170 ;
        RECT 2159.550 3485.190 2160.770 3485.490 ;
        RECT 2110.790 3484.510 2112.010 3484.810 ;
        RECT 2160.470 3484.810 2160.770 3485.190 ;
        RECT 2208.310 3484.810 2208.610 3485.870 ;
        RECT 2256.150 3485.490 2256.450 3485.870 ;
        RECT 2304.910 3485.870 2353.050 3486.170 ;
        RECT 2256.150 3485.190 2304.290 3485.490 ;
        RECT 2160.470 3484.510 2208.610 3484.810 ;
        RECT 2303.990 3484.810 2304.290 3485.190 ;
        RECT 2304.910 3484.810 2305.210 3485.870 ;
        RECT 2352.750 3485.490 2353.050 3485.870 ;
        RECT 2401.510 3485.870 2449.650 3486.170 ;
        RECT 2352.750 3485.190 2400.890 3485.490 ;
        RECT 2303.990 3484.510 2305.210 3484.810 ;
        RECT 2400.590 3484.810 2400.890 3485.190 ;
        RECT 2401.510 3484.810 2401.810 3485.870 ;
        RECT 2449.350 3485.490 2449.650 3485.870 ;
        RECT 2498.110 3485.870 2546.250 3486.170 ;
        RECT 2449.350 3485.190 2497.490 3485.490 ;
        RECT 2400.590 3484.510 2401.810 3484.810 ;
        RECT 2497.190 3484.810 2497.490 3485.190 ;
        RECT 2498.110 3484.810 2498.410 3485.870 ;
        RECT 2545.950 3485.490 2546.250 3485.870 ;
        RECT 2594.710 3485.870 2642.850 3486.170 ;
        RECT 2545.950 3485.190 2594.090 3485.490 ;
        RECT 2497.190 3484.510 2498.410 3484.810 ;
        RECT 2593.790 3484.810 2594.090 3485.190 ;
        RECT 2594.710 3484.810 2595.010 3485.870 ;
        RECT 2642.550 3485.490 2642.850 3485.870 ;
        RECT 2691.310 3485.870 2739.450 3486.170 ;
        RECT 2642.550 3485.190 2690.690 3485.490 ;
        RECT 2593.790 3484.510 2595.010 3484.810 ;
        RECT 2690.390 3484.810 2690.690 3485.190 ;
        RECT 2691.310 3484.810 2691.610 3485.870 ;
        RECT 2739.150 3485.490 2739.450 3485.870 ;
        RECT 2787.910 3485.870 2836.050 3486.170 ;
        RECT 2739.150 3485.190 2787.290 3485.490 ;
        RECT 2690.390 3484.510 2691.610 3484.810 ;
        RECT 2786.990 3484.810 2787.290 3485.190 ;
        RECT 2787.910 3484.810 2788.210 3485.870 ;
        RECT 2835.750 3485.490 2836.050 3485.870 ;
        RECT 2916.710 3485.490 2917.010 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2835.750 3485.190 2883.890 3485.490 ;
        RECT 2786.990 3484.510 2788.210 3484.810 ;
        RECT 2883.590 3484.810 2883.890 3485.190 ;
        RECT 2884.510 3485.190 2917.010 3485.490 ;
        RECT 2884.510 3484.810 2884.810 3485.190 ;
        RECT 2883.590 3484.510 2884.810 3484.810 ;
        RECT 668.190 875.650 668.570 875.660 ;
        RECT 670.000 875.650 674.000 876.040 ;
        RECT 668.190 875.440 674.000 875.650 ;
        RECT 668.190 875.350 670.220 875.440 ;
        RECT 668.190 875.340 668.570 875.350 ;
      LAYER via3 ;
        RECT 668.220 3485.860 668.540 3486.180 ;
        RECT 668.220 875.340 668.540 875.660 ;
      LAYER met4 ;
        RECT 668.215 3485.855 668.545 3486.185 ;
        RECT 668.230 875.665 668.530 3485.855 ;
        RECT 668.215 875.335 668.545 875.665 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 1003.525 2636.100 3517.600 ;
        RECT 2635.890 1003.155 2636.170 1003.525 ;
      LAYER via2 ;
        RECT 2635.890 1003.200 2636.170 1003.480 ;
      LAYER met3 ;
        RECT 664.510 1003.490 664.890 1003.500 ;
        RECT 2635.865 1003.490 2636.195 1003.505 ;
        RECT 664.510 1003.190 2636.195 1003.490 ;
        RECT 664.510 1003.180 664.890 1003.190 ;
        RECT 2635.865 1003.175 2636.195 1003.190 ;
        RECT 664.510 881.090 664.890 881.100 ;
        RECT 670.000 881.090 674.000 881.480 ;
        RECT 664.510 880.880 674.000 881.090 ;
        RECT 664.510 880.790 670.220 880.880 ;
        RECT 664.510 880.780 664.890 880.790 ;
      LAYER via3 ;
        RECT 664.540 1003.180 664.860 1003.500 ;
        RECT 664.540 880.780 664.860 881.100 ;
      LAYER met4 ;
        RECT 664.535 1003.175 664.865 1003.505 ;
        RECT 664.550 881.105 664.850 1003.175 ;
        RECT 664.535 880.775 664.865 881.105 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.930 3501.900 663.250 3501.960 ;
        RECT 2311.570 3501.900 2311.890 3501.960 ;
        RECT 662.930 3501.760 2311.890 3501.900 ;
        RECT 662.930 3501.700 663.250 3501.760 ;
        RECT 2311.570 3501.700 2311.890 3501.760 ;
      LAYER via ;
        RECT 662.960 3501.700 663.220 3501.960 ;
        RECT 2311.600 3501.700 2311.860 3501.960 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3501.990 2311.800 3517.600 ;
        RECT 662.960 3501.670 663.220 3501.990 ;
        RECT 2311.600 3501.670 2311.860 3501.990 ;
        RECT 663.020 885.885 663.160 3501.670 ;
        RECT 662.950 885.515 663.230 885.885 ;
      LAYER via2 ;
        RECT 662.950 885.560 663.230 885.840 ;
      LAYER met3 ;
        RECT 662.925 885.850 663.255 885.865 ;
        RECT 670.000 885.850 674.000 886.240 ;
        RECT 662.925 885.640 674.000 885.850 ;
        RECT 662.925 885.550 670.220 885.640 ;
        RECT 662.925 885.535 663.255 885.550 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.030 3502.920 656.350 3502.980 ;
        RECT 1987.270 3502.920 1987.590 3502.980 ;
        RECT 656.030 3502.780 1987.590 3502.920 ;
        RECT 656.030 3502.720 656.350 3502.780 ;
        RECT 1987.270 3502.720 1987.590 3502.780 ;
        RECT 656.030 925.040 656.350 925.100 ;
        RECT 656.030 924.900 656.720 925.040 ;
        RECT 656.030 924.840 656.350 924.900 ;
        RECT 656.030 921.980 656.350 922.040 ;
        RECT 656.580 921.980 656.720 924.900 ;
        RECT 656.030 921.840 656.720 921.980 ;
        RECT 656.030 921.780 656.350 921.840 ;
      LAYER via ;
        RECT 656.060 3502.720 656.320 3502.980 ;
        RECT 1987.300 3502.720 1987.560 3502.980 ;
        RECT 656.060 924.840 656.320 925.100 ;
        RECT 656.060 921.780 656.320 922.040 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3503.010 1987.500 3517.600 ;
        RECT 656.060 3502.690 656.320 3503.010 ;
        RECT 1987.300 3502.690 1987.560 3503.010 ;
        RECT 656.120 925.130 656.260 3502.690 ;
        RECT 656.060 924.810 656.320 925.130 ;
        RECT 656.060 921.750 656.320 922.070 ;
        RECT 656.120 891.325 656.260 921.750 ;
        RECT 656.050 890.955 656.330 891.325 ;
      LAYER via2 ;
        RECT 656.050 891.000 656.330 891.280 ;
      LAYER met3 ;
        RECT 656.025 891.290 656.355 891.305 ;
        RECT 670.000 891.290 674.000 891.680 ;
        RECT 656.025 891.080 674.000 891.290 ;
        RECT 656.025 890.990 670.220 891.080 ;
        RECT 656.025 890.975 656.355 890.990 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.470 3504.280 662.790 3504.340 ;
        RECT 1662.510 3504.280 1662.830 3504.340 ;
        RECT 662.470 3504.140 1662.830 3504.280 ;
        RECT 662.470 3504.080 662.790 3504.140 ;
        RECT 1662.510 3504.080 1662.830 3504.140 ;
      LAYER via ;
        RECT 662.500 3504.080 662.760 3504.340 ;
        RECT 1662.540 3504.080 1662.800 3504.340 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3504.370 1662.740 3517.600 ;
        RECT 662.500 3504.050 662.760 3504.370 ;
        RECT 1662.540 3504.050 1662.800 3504.370 ;
        RECT 662.560 896.765 662.700 3504.050 ;
        RECT 662.490 896.395 662.770 896.765 ;
      LAYER via2 ;
        RECT 662.490 896.440 662.770 896.720 ;
      LAYER met3 ;
        RECT 662.465 896.730 662.795 896.745 ;
        RECT 670.000 896.730 674.000 897.120 ;
        RECT 662.465 896.520 674.000 896.730 ;
        RECT 662.465 896.430 670.220 896.520 ;
        RECT 662.465 896.415 662.795 896.430 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 669.830 3504.960 670.150 3505.020 ;
        RECT 1338.210 3504.960 1338.530 3505.020 ;
        RECT 669.830 3504.820 1338.530 3504.960 ;
        RECT 669.830 3504.760 670.150 3504.820 ;
        RECT 1338.210 3504.760 1338.530 3504.820 ;
      LAYER via ;
        RECT 669.860 3504.760 670.120 3505.020 ;
        RECT 1338.240 3504.760 1338.500 3505.020 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3505.050 1338.440 3517.600 ;
        RECT 669.860 3504.730 670.120 3505.050 ;
        RECT 1338.240 3504.730 1338.500 3505.050 ;
        RECT 669.920 903.565 670.060 3504.730 ;
        RECT 669.850 903.195 670.130 903.565 ;
      LAYER via2 ;
        RECT 669.850 903.240 670.130 903.520 ;
      LAYER met3 ;
        RECT 669.825 903.530 670.155 903.545 ;
        RECT 669.825 903.215 670.370 903.530 ;
        RECT 670.070 902.560 670.370 903.215 ;
        RECT 670.000 901.960 674.000 902.560 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 651.890 759.800 652.210 759.860 ;
        RECT 656.030 759.800 656.350 759.860 ;
        RECT 651.890 759.660 656.350 759.800 ;
        RECT 651.890 759.600 652.210 759.660 ;
        RECT 656.030 759.600 656.350 759.660 ;
        RECT 651.890 737.020 652.210 737.080 ;
        RECT 654.190 737.020 654.510 737.080 ;
        RECT 651.890 736.880 654.510 737.020 ;
        RECT 651.890 736.820 652.210 736.880 ;
        RECT 654.190 736.820 654.510 736.880 ;
        RECT 655.570 669.360 655.890 669.420 ;
        RECT 656.030 669.360 656.350 669.420 ;
        RECT 655.570 669.220 656.350 669.360 ;
        RECT 655.570 669.160 655.890 669.220 ;
        RECT 656.030 669.160 656.350 669.220 ;
        RECT 656.030 621.080 656.350 621.140 ;
        RECT 656.490 621.080 656.810 621.140 ;
        RECT 656.030 620.940 656.810 621.080 ;
        RECT 656.030 620.880 656.350 620.940 ;
        RECT 656.490 620.880 656.810 620.940 ;
        RECT 656.490 579.600 656.810 579.660 ;
        RECT 657.410 579.600 657.730 579.660 ;
        RECT 656.490 579.460 657.730 579.600 ;
        RECT 656.490 579.400 656.810 579.460 ;
        RECT 657.410 579.400 657.730 579.460 ;
        RECT 656.030 572.460 656.350 572.520 ;
        RECT 657.410 572.460 657.730 572.520 ;
        RECT 656.030 572.320 657.730 572.460 ;
        RECT 656.030 572.260 656.350 572.320 ;
        RECT 657.410 572.260 657.730 572.320 ;
        RECT 656.030 524.520 656.350 524.580 ;
        RECT 656.950 524.520 657.270 524.580 ;
        RECT 656.030 524.380 657.270 524.520 ;
        RECT 656.030 524.320 656.350 524.380 ;
        RECT 656.950 524.320 657.270 524.380 ;
        RECT 656.030 476.240 656.350 476.300 ;
        RECT 656.950 476.240 657.270 476.300 ;
        RECT 656.030 476.100 657.270 476.240 ;
        RECT 656.030 476.040 656.350 476.100 ;
        RECT 656.950 476.040 657.270 476.100 ;
        RECT 656.030 441.560 656.350 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 656.030 441.420 2901.150 441.560 ;
        RECT 656.030 441.360 656.350 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 651.920 759.600 652.180 759.860 ;
        RECT 656.060 759.600 656.320 759.860 ;
        RECT 651.920 736.820 652.180 737.080 ;
        RECT 654.220 736.820 654.480 737.080 ;
        RECT 655.600 669.160 655.860 669.420 ;
        RECT 656.060 669.160 656.320 669.420 ;
        RECT 656.060 620.880 656.320 621.140 ;
        RECT 656.520 620.880 656.780 621.140 ;
        RECT 656.520 579.400 656.780 579.660 ;
        RECT 657.440 579.400 657.700 579.660 ;
        RECT 656.060 572.260 656.320 572.520 ;
        RECT 657.440 572.260 657.700 572.520 ;
        RECT 656.060 524.320 656.320 524.580 ;
        RECT 656.980 524.320 657.240 524.580 ;
        RECT 656.060 476.040 656.320 476.300 ;
        RECT 656.980 476.040 657.240 476.300 ;
        RECT 656.060 441.360 656.320 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 656.050 806.635 656.330 807.005 ;
        RECT 656.120 759.890 656.260 806.635 ;
        RECT 651.920 759.570 652.180 759.890 ;
        RECT 656.060 759.570 656.320 759.890 ;
        RECT 651.980 737.110 652.120 759.570 ;
        RECT 651.920 736.790 652.180 737.110 ;
        RECT 654.220 736.790 654.480 737.110 ;
        RECT 654.280 677.125 654.420 736.790 ;
        RECT 654.210 676.755 654.490 677.125 ;
        RECT 655.590 676.075 655.870 676.445 ;
        RECT 655.660 669.450 655.800 676.075 ;
        RECT 655.600 669.130 655.860 669.450 ;
        RECT 656.060 669.130 656.320 669.450 ;
        RECT 656.120 621.170 656.260 669.130 ;
        RECT 656.060 620.850 656.320 621.170 ;
        RECT 656.520 620.850 656.780 621.170 ;
        RECT 656.580 579.690 656.720 620.850 ;
        RECT 656.520 579.370 656.780 579.690 ;
        RECT 657.440 579.370 657.700 579.690 ;
        RECT 657.500 572.550 657.640 579.370 ;
        RECT 656.060 572.230 656.320 572.550 ;
        RECT 657.440 572.230 657.700 572.550 ;
        RECT 656.120 524.610 656.260 572.230 ;
        RECT 656.060 524.290 656.320 524.610 ;
        RECT 656.980 524.290 657.240 524.610 ;
        RECT 657.040 476.330 657.180 524.290 ;
        RECT 656.060 476.010 656.320 476.330 ;
        RECT 656.980 476.010 657.240 476.330 ;
        RECT 656.120 441.650 656.260 476.010 ;
        RECT 656.060 441.330 656.320 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 656.050 806.680 656.330 806.960 ;
        RECT 654.210 676.800 654.490 677.080 ;
        RECT 655.590 676.120 655.870 676.400 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 656.025 806.970 656.355 806.985 ;
        RECT 670.000 806.970 674.000 807.360 ;
        RECT 656.025 806.760 674.000 806.970 ;
        RECT 656.025 806.670 670.220 806.760 ;
        RECT 656.025 806.655 656.355 806.670 ;
        RECT 654.185 677.090 654.515 677.105 ;
        RECT 654.185 676.790 655.880 677.090 ;
        RECT 654.185 676.775 654.515 676.790 ;
        RECT 655.580 676.425 655.880 676.790 ;
        RECT 655.565 676.095 655.895 676.425 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.070 3501.220 667.390 3501.280 ;
        RECT 1013.910 3501.220 1014.230 3501.280 ;
        RECT 667.070 3501.080 1014.230 3501.220 ;
        RECT 667.070 3501.020 667.390 3501.080 ;
        RECT 1013.910 3501.020 1014.230 3501.080 ;
      LAYER via ;
        RECT 667.100 3501.020 667.360 3501.280 ;
        RECT 1013.940 3501.020 1014.200 3501.280 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3501.310 1014.140 3517.600 ;
        RECT 667.100 3500.990 667.360 3501.310 ;
        RECT 1013.940 3500.990 1014.200 3501.310 ;
        RECT 667.160 906.965 667.300 3500.990 ;
        RECT 667.090 906.595 667.370 906.965 ;
      LAYER via2 ;
        RECT 667.090 906.640 667.370 906.920 ;
      LAYER met3 ;
        RECT 667.065 906.930 667.395 906.945 ;
        RECT 670.000 906.930 674.000 907.320 ;
        RECT 667.065 906.720 674.000 906.930 ;
        RECT 667.065 906.630 670.220 906.720 ;
        RECT 667.065 906.615 667.395 906.630 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 666.610 3498.500 666.930 3498.560 ;
        RECT 689.150 3498.500 689.470 3498.560 ;
        RECT 666.610 3498.360 689.470 3498.500 ;
        RECT 666.610 3498.300 666.930 3498.360 ;
        RECT 689.150 3498.300 689.470 3498.360 ;
      LAYER via ;
        RECT 666.640 3498.300 666.900 3498.560 ;
        RECT 689.180 3498.300 689.440 3498.560 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3498.590 689.380 3517.600 ;
        RECT 666.640 3498.270 666.900 3498.590 ;
        RECT 689.180 3498.270 689.440 3498.590 ;
        RECT 666.700 912.405 666.840 3498.270 ;
        RECT 666.630 912.035 666.910 912.405 ;
      LAYER via2 ;
        RECT 666.630 912.080 666.910 912.360 ;
      LAYER met3 ;
        RECT 666.605 912.370 666.935 912.385 ;
        RECT 670.000 912.370 674.000 912.760 ;
        RECT 666.605 912.160 674.000 912.370 ;
        RECT 666.605 912.070 670.220 912.160 ;
        RECT 666.605 912.055 666.935 912.070 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 362.090 3498.500 362.410 3498.560 ;
        RECT 364.850 3498.500 365.170 3498.560 ;
        RECT 362.090 3498.360 365.170 3498.500 ;
        RECT 362.090 3498.300 362.410 3498.360 ;
        RECT 364.850 3498.300 365.170 3498.360 ;
        RECT 362.090 917.560 362.410 917.620 ;
        RECT 652.350 917.560 652.670 917.620 ;
        RECT 362.090 917.420 652.670 917.560 ;
        RECT 362.090 917.360 362.410 917.420 ;
        RECT 652.350 917.360 652.670 917.420 ;
      LAYER via ;
        RECT 362.120 3498.300 362.380 3498.560 ;
        RECT 364.880 3498.300 365.140 3498.560 ;
        RECT 362.120 917.360 362.380 917.620 ;
        RECT 652.380 917.360 652.640 917.620 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3498.590 365.080 3517.600 ;
        RECT 362.120 3498.270 362.380 3498.590 ;
        RECT 364.880 3498.270 365.140 3498.590 ;
        RECT 362.180 917.650 362.320 3498.270 ;
        RECT 362.120 917.330 362.380 917.650 ;
        RECT 652.370 917.475 652.650 917.845 ;
        RECT 652.380 917.330 652.640 917.475 ;
      LAYER via2 ;
        RECT 652.370 917.520 652.650 917.800 ;
      LAYER met3 ;
        RECT 652.345 917.810 652.675 917.825 ;
        RECT 670.000 917.810 674.000 918.200 ;
        RECT 652.345 917.600 674.000 917.810 ;
        RECT 652.345 917.510 670.220 917.600 ;
        RECT 652.345 917.495 652.675 917.510 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3501.900 40.870 3501.960 ;
        RECT 65.390 3501.900 65.710 3501.960 ;
        RECT 40.550 3501.760 65.710 3501.900 ;
        RECT 40.550 3501.700 40.870 3501.760 ;
        RECT 65.390 3501.700 65.710 3501.760 ;
        RECT 65.390 924.360 65.710 924.420 ;
        RECT 656.030 924.360 656.350 924.420 ;
        RECT 65.390 924.220 656.350 924.360 ;
        RECT 65.390 924.160 65.710 924.220 ;
        RECT 656.030 924.160 656.350 924.220 ;
      LAYER via ;
        RECT 40.580 3501.700 40.840 3501.960 ;
        RECT 65.420 3501.700 65.680 3501.960 ;
        RECT 65.420 924.160 65.680 924.420 ;
        RECT 656.060 924.160 656.320 924.420 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.990 40.780 3517.600 ;
        RECT 40.580 3501.670 40.840 3501.990 ;
        RECT 65.420 3501.670 65.680 3501.990 ;
        RECT 65.480 924.450 65.620 3501.670 ;
        RECT 65.420 924.130 65.680 924.450 ;
        RECT 656.060 924.130 656.320 924.450 ;
        RECT 656.120 922.605 656.260 924.130 ;
        RECT 656.050 922.235 656.330 922.605 ;
      LAYER via2 ;
        RECT 656.050 922.280 656.330 922.560 ;
      LAYER met3 ;
        RECT 656.025 922.570 656.355 922.585 ;
        RECT 670.000 922.570 674.000 922.960 ;
        RECT 656.025 922.360 674.000 922.570 ;
        RECT 656.025 922.270 670.220 922.360 ;
        RECT 656.025 922.255 656.355 922.270 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 23.990 931.500 24.310 931.560 ;
        RECT 652.350 931.500 652.670 931.560 ;
        RECT 23.990 931.360 652.670 931.500 ;
        RECT 23.990 931.300 24.310 931.360 ;
        RECT 652.350 931.300 652.670 931.360 ;
      LAYER via ;
        RECT 24.020 931.300 24.280 931.560 ;
        RECT 652.380 931.300 652.640 931.560 ;
      LAYER met2 ;
        RECT 24.010 3267.555 24.290 3267.925 ;
        RECT 24.080 931.590 24.220 3267.555 ;
        RECT 24.020 931.270 24.280 931.590 ;
        RECT 652.380 931.270 652.640 931.590 ;
        RECT 652.440 930.765 652.580 931.270 ;
        RECT 652.370 930.395 652.650 930.765 ;
      LAYER via2 ;
        RECT 24.010 3267.600 24.290 3267.880 ;
        RECT 652.370 930.440 652.650 930.720 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 23.985 3267.890 24.315 3267.905 ;
        RECT -4.800 3267.590 24.315 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 23.985 3267.575 24.315 3267.590 ;
        RECT 652.345 930.730 652.675 930.745 ;
        RECT 652.345 930.430 670.370 930.730 ;
        RECT 652.345 930.415 652.675 930.430 ;
        RECT 670.070 928.400 670.370 930.430 ;
        RECT 670.000 927.800 674.000 928.400 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2974.220 20.630 2974.280 ;
        RECT 24.450 2974.220 24.770 2974.280 ;
        RECT 20.310 2974.080 24.770 2974.220 ;
        RECT 20.310 2974.020 20.630 2974.080 ;
        RECT 24.450 2974.020 24.770 2974.080 ;
        RECT 24.450 938.300 24.770 938.360 ;
        RECT 658.790 938.300 659.110 938.360 ;
        RECT 24.450 938.160 659.110 938.300 ;
        RECT 24.450 938.100 24.770 938.160 ;
        RECT 658.790 938.100 659.110 938.160 ;
      LAYER via ;
        RECT 20.340 2974.020 20.600 2974.280 ;
        RECT 24.480 2974.020 24.740 2974.280 ;
        RECT 24.480 938.100 24.740 938.360 ;
        RECT 658.820 938.100 659.080 938.360 ;
      LAYER met2 ;
        RECT 20.330 2979.915 20.610 2980.285 ;
        RECT 20.400 2974.310 20.540 2979.915 ;
        RECT 20.340 2973.990 20.600 2974.310 ;
        RECT 24.480 2973.990 24.740 2974.310 ;
        RECT 24.540 938.390 24.680 2973.990 ;
        RECT 24.480 938.070 24.740 938.390 ;
        RECT 658.820 938.070 659.080 938.390 ;
        RECT 658.880 933.485 659.020 938.070 ;
        RECT 658.810 933.115 659.090 933.485 ;
      LAYER via2 ;
        RECT 20.330 2979.960 20.610 2980.240 ;
        RECT 658.810 933.160 659.090 933.440 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 20.305 2980.250 20.635 2980.265 ;
        RECT -4.800 2979.950 20.635 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 20.305 2979.935 20.635 2979.950 ;
        RECT 658.785 933.450 659.115 933.465 ;
        RECT 670.000 933.450 674.000 933.840 ;
        RECT 658.785 933.240 674.000 933.450 ;
        RECT 658.785 933.150 670.220 933.240 ;
        RECT 658.785 933.135 659.115 933.150 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 945.100 17.870 945.160 ;
        RECT 17.550 944.960 659.480 945.100 ;
        RECT 17.550 944.900 17.870 944.960 ;
        RECT 658.790 943.060 659.110 943.120 ;
        RECT 659.340 943.060 659.480 944.960 ;
        RECT 658.790 942.920 659.480 943.060 ;
        RECT 658.790 942.860 659.110 942.920 ;
      LAYER via ;
        RECT 17.580 944.900 17.840 945.160 ;
        RECT 658.820 942.860 659.080 943.120 ;
      LAYER met2 ;
        RECT 17.570 2692.955 17.850 2693.325 ;
        RECT 17.640 945.190 17.780 2692.955 ;
        RECT 17.580 944.870 17.840 945.190 ;
        RECT 658.820 942.830 659.080 943.150 ;
        RECT 658.880 938.925 659.020 942.830 ;
        RECT 658.810 938.555 659.090 938.925 ;
      LAYER via2 ;
        RECT 17.570 2693.000 17.850 2693.280 ;
        RECT 658.810 938.600 659.090 938.880 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 17.545 2693.290 17.875 2693.305 ;
        RECT -4.800 2692.990 17.875 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 17.545 2692.975 17.875 2692.990 ;
        RECT 658.785 938.890 659.115 938.905 ;
        RECT 670.000 938.890 674.000 939.280 ;
        RECT 658.785 938.680 674.000 938.890 ;
        RECT 658.785 938.590 670.220 938.680 ;
        RECT 658.785 938.575 659.115 938.590 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2403.360 20.630 2403.420 ;
        RECT 24.910 2403.360 25.230 2403.420 ;
        RECT 20.310 2403.220 25.230 2403.360 ;
        RECT 20.310 2403.160 20.630 2403.220 ;
        RECT 24.910 2403.160 25.230 2403.220 ;
        RECT 24.910 944.760 25.230 944.820 ;
        RECT 658.790 944.760 659.110 944.820 ;
        RECT 24.910 944.620 659.110 944.760 ;
        RECT 24.910 944.560 25.230 944.620 ;
        RECT 658.790 944.560 659.110 944.620 ;
      LAYER via ;
        RECT 20.340 2403.160 20.600 2403.420 ;
        RECT 24.940 2403.160 25.200 2403.420 ;
        RECT 24.940 944.560 25.200 944.820 ;
        RECT 658.820 944.560 659.080 944.820 ;
      LAYER met2 ;
        RECT 20.330 2405.315 20.610 2405.685 ;
        RECT 20.400 2403.450 20.540 2405.315 ;
        RECT 20.340 2403.130 20.600 2403.450 ;
        RECT 24.940 2403.130 25.200 2403.450 ;
        RECT 25.000 944.850 25.140 2403.130 ;
        RECT 24.940 944.530 25.200 944.850 ;
        RECT 658.820 944.530 659.080 944.850 ;
        RECT 658.880 943.685 659.020 944.530 ;
        RECT 658.810 943.315 659.090 943.685 ;
      LAYER via2 ;
        RECT 20.330 2405.360 20.610 2405.640 ;
        RECT 658.810 943.360 659.090 943.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 20.305 2405.650 20.635 2405.665 ;
        RECT -4.800 2405.350 20.635 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 20.305 2405.335 20.635 2405.350 ;
        RECT 658.785 943.650 659.115 943.665 ;
        RECT 670.000 943.650 674.000 944.040 ;
        RECT 658.785 943.440 674.000 943.650 ;
        RECT 658.785 943.350 670.220 943.440 ;
        RECT 658.785 943.335 659.115 943.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2118.440 20.630 2118.500 ;
        RECT 25.370 2118.440 25.690 2118.500 ;
        RECT 20.310 2118.300 25.690 2118.440 ;
        RECT 20.310 2118.240 20.630 2118.300 ;
        RECT 25.370 2118.240 25.690 2118.300 ;
        RECT 25.370 952.240 25.690 952.300 ;
        RECT 658.790 952.240 659.110 952.300 ;
        RECT 25.370 952.100 659.110 952.240 ;
        RECT 25.370 952.040 25.690 952.100 ;
        RECT 658.790 952.040 659.110 952.100 ;
      LAYER via ;
        RECT 20.340 2118.240 20.600 2118.500 ;
        RECT 25.400 2118.240 25.660 2118.500 ;
        RECT 25.400 952.040 25.660 952.300 ;
        RECT 658.820 952.040 659.080 952.300 ;
      LAYER met2 ;
        RECT 20.330 2118.355 20.610 2118.725 ;
        RECT 20.340 2118.210 20.600 2118.355 ;
        RECT 25.400 2118.210 25.660 2118.530 ;
        RECT 25.460 952.330 25.600 2118.210 ;
        RECT 25.400 952.010 25.660 952.330 ;
        RECT 658.820 952.010 659.080 952.330 ;
        RECT 658.880 949.125 659.020 952.010 ;
        RECT 658.810 948.755 659.090 949.125 ;
      LAYER via2 ;
        RECT 20.330 2118.400 20.610 2118.680 ;
        RECT 658.810 948.800 659.090 949.080 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 20.305 2118.690 20.635 2118.705 ;
        RECT -4.800 2118.390 20.635 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 20.305 2118.375 20.635 2118.390 ;
        RECT 658.785 949.090 659.115 949.105 ;
        RECT 670.000 949.090 674.000 949.480 ;
        RECT 658.785 948.880 674.000 949.090 ;
        RECT 658.785 948.790 670.220 948.880 ;
        RECT 658.785 948.775 659.115 948.790 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 1828.760 14.190 1828.820 ;
        RECT 25.830 1828.760 26.150 1828.820 ;
        RECT 13.870 1828.620 26.150 1828.760 ;
        RECT 13.870 1828.560 14.190 1828.620 ;
        RECT 25.830 1828.560 26.150 1828.620 ;
        RECT 25.830 959.040 26.150 959.100 ;
        RECT 658.790 959.040 659.110 959.100 ;
        RECT 25.830 958.900 659.110 959.040 ;
        RECT 25.830 958.840 26.150 958.900 ;
        RECT 658.790 958.840 659.110 958.900 ;
      LAYER via ;
        RECT 13.900 1828.560 14.160 1828.820 ;
        RECT 25.860 1828.560 26.120 1828.820 ;
        RECT 25.860 958.840 26.120 959.100 ;
        RECT 658.820 958.840 659.080 959.100 ;
      LAYER met2 ;
        RECT 13.890 1830.715 14.170 1831.085 ;
        RECT 13.960 1828.850 14.100 1830.715 ;
        RECT 13.900 1828.530 14.160 1828.850 ;
        RECT 25.860 1828.530 26.120 1828.850 ;
        RECT 25.920 959.130 26.060 1828.530 ;
        RECT 25.860 958.810 26.120 959.130 ;
        RECT 658.820 958.810 659.080 959.130 ;
        RECT 658.880 954.565 659.020 958.810 ;
        RECT 658.810 954.195 659.090 954.565 ;
      LAYER via2 ;
        RECT 13.890 1830.760 14.170 1831.040 ;
        RECT 658.810 954.240 659.090 954.520 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 13.865 1831.050 14.195 1831.065 ;
        RECT -4.800 1830.750 14.195 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 13.865 1830.735 14.195 1830.750 ;
        RECT 658.785 954.530 659.115 954.545 ;
        RECT 670.000 954.530 674.000 954.920 ;
        RECT 658.785 954.320 674.000 954.530 ;
        RECT 658.785 954.230 670.220 954.320 ;
        RECT 658.785 954.215 659.115 954.230 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 603.740 662.330 603.800 ;
        RECT 2901.750 603.740 2902.070 603.800 ;
        RECT 662.010 603.600 2902.070 603.740 ;
        RECT 662.010 603.540 662.330 603.600 ;
        RECT 2901.750 603.540 2902.070 603.600 ;
      LAYER via ;
        RECT 662.040 603.540 662.300 603.800 ;
        RECT 2901.780 603.540 2902.040 603.800 ;
      LAYER met2 ;
        RECT 662.030 812.075 662.310 812.445 ;
        RECT 662.100 603.830 662.240 812.075 ;
        RECT 2901.770 674.035 2902.050 674.405 ;
        RECT 2901.840 603.830 2901.980 674.035 ;
        RECT 662.040 603.510 662.300 603.830 ;
        RECT 2901.780 603.510 2902.040 603.830 ;
      LAYER via2 ;
        RECT 662.030 812.120 662.310 812.400 ;
        RECT 2901.770 674.080 2902.050 674.360 ;
      LAYER met3 ;
        RECT 662.005 812.410 662.335 812.425 ;
        RECT 670.000 812.410 674.000 812.800 ;
        RECT 662.005 812.200 674.000 812.410 ;
        RECT 662.005 812.110 670.220 812.200 ;
        RECT 662.005 812.095 662.335 812.110 ;
        RECT 2901.745 674.370 2902.075 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2901.745 674.070 2924.800 674.370 ;
        RECT 2901.745 674.055 2902.075 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 1539.080 20.630 1539.140 ;
        RECT 26.290 1539.080 26.610 1539.140 ;
        RECT 20.310 1538.940 26.610 1539.080 ;
        RECT 20.310 1538.880 20.630 1538.940 ;
        RECT 26.290 1538.880 26.610 1538.940 ;
        RECT 26.290 965.840 26.610 965.900 ;
        RECT 26.290 965.700 659.480 965.840 ;
        RECT 26.290 965.640 26.610 965.700 ;
        RECT 658.790 964.140 659.110 964.200 ;
        RECT 659.340 964.140 659.480 965.700 ;
        RECT 658.790 964.000 659.480 964.140 ;
        RECT 658.790 963.940 659.110 964.000 ;
      LAYER via ;
        RECT 20.340 1538.880 20.600 1539.140 ;
        RECT 26.320 1538.880 26.580 1539.140 ;
        RECT 26.320 965.640 26.580 965.900 ;
        RECT 658.820 963.940 659.080 964.200 ;
      LAYER met2 ;
        RECT 20.330 1543.755 20.610 1544.125 ;
        RECT 20.400 1539.170 20.540 1543.755 ;
        RECT 20.340 1538.850 20.600 1539.170 ;
        RECT 26.320 1538.850 26.580 1539.170 ;
        RECT 26.380 965.930 26.520 1538.850 ;
        RECT 26.320 965.610 26.580 965.930 ;
        RECT 658.820 963.910 659.080 964.230 ;
        RECT 658.880 960.005 659.020 963.910 ;
        RECT 658.810 959.635 659.090 960.005 ;
      LAYER via2 ;
        RECT 20.330 1543.800 20.610 1544.080 ;
        RECT 658.810 959.680 659.090 959.960 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 20.305 1544.090 20.635 1544.105 ;
        RECT -4.800 1543.790 20.635 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 20.305 1543.775 20.635 1543.790 ;
        RECT 658.785 959.970 659.115 959.985 ;
        RECT 670.000 959.970 674.000 960.360 ;
        RECT 658.785 959.760 674.000 959.970 ;
        RECT 658.785 959.670 670.220 959.760 ;
        RECT 658.785 959.655 659.115 959.670 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 1324.880 14.190 1324.940 ;
        RECT 27.210 1324.880 27.530 1324.940 ;
        RECT 13.870 1324.740 27.530 1324.880 ;
        RECT 13.870 1324.680 14.190 1324.740 ;
        RECT 27.210 1324.680 27.530 1324.740 ;
        RECT 27.210 965.500 27.530 965.560 ;
        RECT 658.790 965.500 659.110 965.560 ;
        RECT 27.210 965.360 659.110 965.500 ;
        RECT 27.210 965.300 27.530 965.360 ;
        RECT 658.790 965.300 659.110 965.360 ;
      LAYER via ;
        RECT 13.900 1324.680 14.160 1324.940 ;
        RECT 27.240 1324.680 27.500 1324.940 ;
        RECT 27.240 965.300 27.500 965.560 ;
        RECT 658.820 965.300 659.080 965.560 ;
      LAYER met2 ;
        RECT 13.890 1328.195 14.170 1328.565 ;
        RECT 13.960 1324.970 14.100 1328.195 ;
        RECT 13.900 1324.650 14.160 1324.970 ;
        RECT 27.240 1324.650 27.500 1324.970 ;
        RECT 27.300 965.590 27.440 1324.650 ;
        RECT 27.240 965.270 27.500 965.590 ;
        RECT 658.820 965.270 659.080 965.590 ;
        RECT 658.880 964.765 659.020 965.270 ;
        RECT 658.810 964.395 659.090 964.765 ;
      LAYER via2 ;
        RECT 13.890 1328.240 14.170 1328.520 ;
        RECT 658.810 964.440 659.090 964.720 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 13.865 1328.530 14.195 1328.545 ;
        RECT -4.800 1328.230 14.195 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 13.865 1328.215 14.195 1328.230 ;
        RECT 658.785 964.730 659.115 964.745 ;
        RECT 670.000 964.730 674.000 965.120 ;
        RECT 658.785 964.520 674.000 964.730 ;
        RECT 658.785 964.430 670.220 964.520 ;
        RECT 658.785 964.415 659.115 964.430 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 1111.020 15.110 1111.080 ;
        RECT 72.290 1111.020 72.610 1111.080 ;
        RECT 14.790 1110.880 72.610 1111.020 ;
        RECT 14.790 1110.820 15.110 1110.880 ;
        RECT 72.290 1110.820 72.610 1110.880 ;
        RECT 72.290 972.300 72.610 972.360 ;
        RECT 658.790 972.300 659.110 972.360 ;
        RECT 72.290 972.160 659.110 972.300 ;
        RECT 72.290 972.100 72.610 972.160 ;
        RECT 658.790 972.100 659.110 972.160 ;
      LAYER via ;
        RECT 14.820 1110.820 15.080 1111.080 ;
        RECT 72.320 1110.820 72.580 1111.080 ;
        RECT 72.320 972.100 72.580 972.360 ;
        RECT 658.820 972.100 659.080 972.360 ;
      LAYER met2 ;
        RECT 14.810 1112.635 15.090 1113.005 ;
        RECT 14.880 1111.110 15.020 1112.635 ;
        RECT 14.820 1110.790 15.080 1111.110 ;
        RECT 72.320 1110.790 72.580 1111.110 ;
        RECT 72.380 972.390 72.520 1110.790 ;
        RECT 72.320 972.070 72.580 972.390 ;
        RECT 658.820 972.070 659.080 972.390 ;
        RECT 658.880 970.205 659.020 972.070 ;
        RECT 658.810 969.835 659.090 970.205 ;
      LAYER via2 ;
        RECT 14.810 1112.680 15.090 1112.960 ;
        RECT 658.810 969.880 659.090 970.160 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 14.785 1112.970 15.115 1112.985 ;
        RECT -4.800 1112.670 15.115 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 14.785 1112.655 15.115 1112.670 ;
        RECT 658.785 970.170 659.115 970.185 ;
        RECT 670.000 970.170 674.000 970.560 ;
        RECT 658.785 969.960 674.000 970.170 ;
        RECT 658.785 969.870 670.220 969.960 ;
        RECT 658.785 969.855 659.115 969.870 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 79.190 972.980 79.510 973.040 ;
        RECT 658.790 972.980 659.110 973.040 ;
        RECT 79.190 972.840 659.110 972.980 ;
        RECT 79.190 972.780 79.510 972.840 ;
        RECT 658.790 972.780 659.110 972.840 ;
        RECT 14.330 903.960 14.650 904.020 ;
        RECT 79.190 903.960 79.510 904.020 ;
        RECT 14.330 903.820 79.510 903.960 ;
        RECT 14.330 903.760 14.650 903.820 ;
        RECT 79.190 903.760 79.510 903.820 ;
      LAYER via ;
        RECT 79.220 972.780 79.480 973.040 ;
        RECT 658.820 972.780 659.080 973.040 ;
        RECT 14.360 903.760 14.620 904.020 ;
        RECT 79.220 903.760 79.480 904.020 ;
      LAYER met2 ;
        RECT 658.810 975.275 659.090 975.645 ;
        RECT 658.880 973.070 659.020 975.275 ;
        RECT 79.220 972.750 79.480 973.070 ;
        RECT 658.820 972.750 659.080 973.070 ;
        RECT 79.280 904.050 79.420 972.750 ;
        RECT 14.360 903.730 14.620 904.050 ;
        RECT 79.220 903.730 79.480 904.050 ;
        RECT 14.420 897.445 14.560 903.730 ;
        RECT 14.350 897.075 14.630 897.445 ;
      LAYER via2 ;
        RECT 658.810 975.320 659.090 975.600 ;
        RECT 14.350 897.120 14.630 897.400 ;
      LAYER met3 ;
        RECT 658.785 975.610 659.115 975.625 ;
        RECT 670.000 975.610 674.000 976.000 ;
        RECT 658.785 975.400 674.000 975.610 ;
        RECT 658.785 975.310 670.220 975.400 ;
        RECT 658.785 975.295 659.115 975.310 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 14.325 897.410 14.655 897.425 ;
        RECT -4.800 897.110 14.655 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 14.325 897.095 14.655 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 654.190 980.600 654.510 980.860 ;
        RECT 86.090 980.460 86.410 980.520 ;
        RECT 654.280 980.460 654.420 980.600 ;
        RECT 86.090 980.320 654.420 980.460 ;
        RECT 86.090 980.260 86.410 980.320 ;
        RECT 16.630 682.960 16.950 683.020 ;
        RECT 86.090 682.960 86.410 683.020 ;
        RECT 16.630 682.820 86.410 682.960 ;
        RECT 16.630 682.760 16.950 682.820 ;
        RECT 86.090 682.760 86.410 682.820 ;
      LAYER via ;
        RECT 654.220 980.600 654.480 980.860 ;
        RECT 86.120 980.260 86.380 980.520 ;
        RECT 16.660 682.760 16.920 683.020 ;
        RECT 86.120 682.760 86.380 683.020 ;
      LAYER met2 ;
        RECT 654.210 980.715 654.490 981.085 ;
        RECT 654.220 980.570 654.480 980.715 ;
        RECT 86.120 980.230 86.380 980.550 ;
        RECT 86.180 683.050 86.320 980.230 ;
        RECT 16.660 682.730 16.920 683.050 ;
        RECT 86.120 682.730 86.380 683.050 ;
        RECT 16.720 681.885 16.860 682.730 ;
        RECT 16.650 681.515 16.930 681.885 ;
      LAYER via2 ;
        RECT 654.210 980.760 654.490 981.040 ;
        RECT 16.650 681.560 16.930 681.840 ;
      LAYER met3 ;
        RECT 654.185 981.050 654.515 981.065 ;
        RECT 670.000 981.050 674.000 981.440 ;
        RECT 654.185 980.840 674.000 981.050 ;
        RECT 654.185 980.750 670.220 980.840 ;
        RECT 654.185 980.735 654.515 980.750 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.625 681.850 16.955 681.865 ;
        RECT -4.800 681.550 16.955 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.625 681.535 16.955 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.750 981.480 27.070 981.540 ;
        RECT 656.950 981.480 657.270 981.540 ;
        RECT 26.750 981.340 657.270 981.480 ;
        RECT 26.750 981.280 27.070 981.340 ;
        RECT 656.950 981.280 657.270 981.340 ;
        RECT 13.870 466.720 14.190 466.780 ;
        RECT 26.750 466.720 27.070 466.780 ;
        RECT 13.870 466.580 27.070 466.720 ;
        RECT 13.870 466.520 14.190 466.580 ;
        RECT 26.750 466.520 27.070 466.580 ;
      LAYER via ;
        RECT 26.780 981.280 27.040 981.540 ;
        RECT 656.980 981.280 657.240 981.540 ;
        RECT 13.900 466.520 14.160 466.780 ;
        RECT 26.780 466.520 27.040 466.780 ;
      LAYER met2 ;
        RECT 656.970 985.475 657.250 985.845 ;
        RECT 657.040 981.570 657.180 985.475 ;
        RECT 26.780 981.250 27.040 981.570 ;
        RECT 656.980 981.250 657.240 981.570 ;
        RECT 26.840 466.810 26.980 981.250 ;
        RECT 13.900 466.490 14.160 466.810 ;
        RECT 26.780 466.490 27.040 466.810 ;
        RECT 13.960 466.325 14.100 466.490 ;
        RECT 13.890 465.955 14.170 466.325 ;
      LAYER via2 ;
        RECT 656.970 985.520 657.250 985.800 ;
        RECT 13.890 466.000 14.170 466.280 ;
      LAYER met3 ;
        RECT 656.945 985.810 657.275 985.825 ;
        RECT 670.000 985.810 674.000 986.200 ;
        RECT 656.945 985.600 674.000 985.810 ;
        RECT 656.945 985.510 670.220 985.600 ;
        RECT 656.945 985.495 657.275 985.510 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 13.865 466.290 14.195 466.305 ;
        RECT -4.800 465.990 14.195 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 13.865 465.975 14.195 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 986.920 17.410 986.980 ;
        RECT 656.950 986.920 657.270 986.980 ;
        RECT 17.090 986.780 657.270 986.920 ;
        RECT 17.090 986.720 17.410 986.780 ;
        RECT 656.950 986.720 657.270 986.780 ;
      LAYER via ;
        RECT 17.120 986.720 17.380 986.980 ;
        RECT 656.980 986.720 657.240 986.980 ;
      LAYER met2 ;
        RECT 656.970 990.915 657.250 991.285 ;
        RECT 657.040 987.010 657.180 990.915 ;
        RECT 17.120 986.690 17.380 987.010 ;
        RECT 656.980 986.690 657.240 987.010 ;
        RECT 17.180 250.765 17.320 986.690 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 656.970 990.960 657.250 991.240 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 656.945 991.250 657.275 991.265 ;
        RECT 670.000 991.250 674.000 991.640 ;
        RECT 656.945 991.040 674.000 991.250 ;
        RECT 656.945 990.950 670.220 991.040 ;
        RECT 656.945 990.935 657.275 990.950 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 658.790 41.380 659.110 41.440 ;
        RECT 17.090 41.240 659.110 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 658.790 41.180 659.110 41.240 ;
      LAYER via ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 658.820 41.180 659.080 41.440 ;
      LAYER met2 ;
        RECT 658.810 996.355 659.090 996.725 ;
        RECT 658.880 980.405 659.020 996.355 ;
        RECT 658.810 980.035 659.090 980.405 ;
        RECT 658.810 932.435 659.090 932.805 ;
        RECT 658.880 41.470 659.020 932.435 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 658.820 41.150 659.080 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 658.810 996.400 659.090 996.680 ;
        RECT 658.810 980.080 659.090 980.360 ;
        RECT 658.810 932.480 659.090 932.760 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 658.785 996.690 659.115 996.705 ;
        RECT 670.000 996.690 674.000 997.080 ;
        RECT 658.785 996.480 674.000 996.690 ;
        RECT 658.785 996.390 670.220 996.480 ;
        RECT 658.785 996.375 659.115 996.390 ;
        RECT 658.070 980.370 658.450 980.380 ;
        RECT 658.785 980.370 659.115 980.385 ;
        RECT 658.070 980.070 659.115 980.370 ;
        RECT 658.070 980.060 658.450 980.070 ;
        RECT 658.785 980.055 659.115 980.070 ;
        RECT 658.070 932.770 658.450 932.780 ;
        RECT 658.785 932.770 659.115 932.785 ;
        RECT 658.070 932.470 659.115 932.770 ;
        RECT 658.070 932.460 658.450 932.470 ;
        RECT 658.785 932.455 659.115 932.470 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
      LAYER via3 ;
        RECT 658.100 980.060 658.420 980.380 ;
        RECT 658.100 932.460 658.420 932.780 ;
      LAYER met4 ;
        RECT 658.095 980.055 658.425 980.385 ;
        RECT 658.110 932.785 658.410 980.055 ;
        RECT 658.095 932.455 658.425 932.785 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.990 999.160 668.310 999.220 ;
        RECT 2901.290 999.160 2901.610 999.220 ;
        RECT 667.990 999.020 2901.610 999.160 ;
        RECT 667.990 998.960 668.310 999.020 ;
        RECT 2901.290 998.960 2901.610 999.020 ;
      LAYER via ;
        RECT 668.020 998.960 668.280 999.220 ;
        RECT 2901.320 998.960 2901.580 999.220 ;
      LAYER met2 ;
        RECT 668.020 998.930 668.280 999.250 ;
        RECT 2901.320 998.930 2901.580 999.250 ;
        RECT 668.080 817.885 668.220 998.930 ;
        RECT 2901.380 909.685 2901.520 998.930 ;
        RECT 2901.310 909.315 2901.590 909.685 ;
        RECT 668.010 817.515 668.290 817.885 ;
      LAYER via2 ;
        RECT 2901.310 909.360 2901.590 909.640 ;
        RECT 668.010 817.560 668.290 817.840 ;
      LAYER met3 ;
        RECT 2901.285 909.650 2901.615 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2901.285 909.350 2924.800 909.650 ;
        RECT 2901.285 909.335 2901.615 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT 667.985 817.850 668.315 817.865 ;
        RECT 670.000 817.850 674.000 818.240 ;
        RECT 667.985 817.640 674.000 817.850 ;
        RECT 667.985 817.550 670.220 817.640 ;
        RECT 667.985 817.535 668.315 817.550 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.490 1138.900 656.810 1138.960 ;
        RECT 2900.830 1138.900 2901.150 1138.960 ;
        RECT 656.490 1138.760 2901.150 1138.900 ;
        RECT 656.490 1138.700 656.810 1138.760 ;
        RECT 2900.830 1138.700 2901.150 1138.760 ;
      LAYER via ;
        RECT 656.520 1138.700 656.780 1138.960 ;
        RECT 2900.860 1138.700 2901.120 1138.960 ;
      LAYER met2 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
        RECT 2900.920 1138.990 2901.060 1143.915 ;
        RECT 656.520 1138.670 656.780 1138.990 ;
        RECT 2900.860 1138.670 2901.120 1138.990 ;
        RECT 656.580 822.645 656.720 1138.670 ;
        RECT 656.510 822.275 656.790 822.645 ;
      LAYER via2 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
        RECT 656.510 822.320 656.790 822.600 ;
      LAYER met3 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 656.485 822.610 656.815 822.625 ;
        RECT 670.000 822.610 674.000 823.000 ;
        RECT 656.485 822.400 674.000 822.610 ;
        RECT 656.485 822.310 670.220 822.400 ;
        RECT 656.485 822.295 656.815 822.310 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 663.390 1373.500 663.710 1373.560 ;
        RECT 2898.070 1373.500 2898.390 1373.560 ;
        RECT 663.390 1373.360 2898.390 1373.500 ;
        RECT 663.390 1373.300 663.710 1373.360 ;
        RECT 2898.070 1373.300 2898.390 1373.360 ;
      LAYER via ;
        RECT 663.420 1373.300 663.680 1373.560 ;
        RECT 2898.100 1373.300 2898.360 1373.560 ;
      LAYER met2 ;
        RECT 2898.090 1378.515 2898.370 1378.885 ;
        RECT 2898.160 1373.590 2898.300 1378.515 ;
        RECT 663.420 1373.270 663.680 1373.590 ;
        RECT 2898.100 1373.270 2898.360 1373.590 ;
        RECT 663.480 828.085 663.620 1373.270 ;
        RECT 663.410 827.715 663.690 828.085 ;
      LAYER via2 ;
        RECT 2898.090 1378.560 2898.370 1378.840 ;
        RECT 663.410 827.760 663.690 828.040 ;
      LAYER met3 ;
        RECT 2898.065 1378.850 2898.395 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2898.065 1378.550 2924.800 1378.850 ;
        RECT 2898.065 1378.535 2898.395 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 663.385 828.050 663.715 828.065 ;
        RECT 670.000 828.050 674.000 828.440 ;
        RECT 663.385 827.840 674.000 828.050 ;
        RECT 663.385 827.750 670.220 827.840 ;
        RECT 663.385 827.735 663.715 827.750 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 663.850 1608.100 664.170 1608.160 ;
        RECT 2898.070 1608.100 2898.390 1608.160 ;
        RECT 663.850 1607.960 2898.390 1608.100 ;
        RECT 663.850 1607.900 664.170 1607.960 ;
        RECT 2898.070 1607.900 2898.390 1607.960 ;
      LAYER via ;
        RECT 663.880 1607.900 664.140 1608.160 ;
        RECT 2898.100 1607.900 2898.360 1608.160 ;
      LAYER met2 ;
        RECT 2898.090 1613.115 2898.370 1613.485 ;
        RECT 2898.160 1608.190 2898.300 1613.115 ;
        RECT 663.880 1607.870 664.140 1608.190 ;
        RECT 2898.100 1607.870 2898.360 1608.190 ;
        RECT 663.940 833.525 664.080 1607.870 ;
        RECT 663.870 833.155 664.150 833.525 ;
      LAYER via2 ;
        RECT 2898.090 1613.160 2898.370 1613.440 ;
        RECT 663.870 833.200 664.150 833.480 ;
      LAYER met3 ;
        RECT 2898.065 1613.450 2898.395 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2898.065 1613.150 2924.800 1613.450 ;
        RECT 2898.065 1613.135 2898.395 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 663.845 833.490 664.175 833.505 ;
        RECT 670.000 833.490 674.000 833.880 ;
        RECT 663.845 833.280 674.000 833.490 ;
        RECT 663.845 833.190 670.220 833.280 ;
        RECT 663.845 833.175 664.175 833.190 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 658.330 1707.720 658.650 1707.780 ;
        RECT 2903.590 1707.720 2903.910 1707.780 ;
        RECT 658.330 1707.580 2903.910 1707.720 ;
        RECT 658.330 1707.520 658.650 1707.580 ;
        RECT 2903.590 1707.520 2903.910 1707.580 ;
      LAYER via ;
        RECT 658.360 1707.520 658.620 1707.780 ;
        RECT 2903.620 1707.520 2903.880 1707.780 ;
      LAYER met2 ;
        RECT 2903.610 1847.715 2903.890 1848.085 ;
        RECT 2903.680 1707.810 2903.820 1847.715 ;
        RECT 658.360 1707.490 658.620 1707.810 ;
        RECT 2903.620 1707.490 2903.880 1707.810 ;
        RECT 658.420 838.965 658.560 1707.490 ;
        RECT 658.350 838.595 658.630 838.965 ;
      LAYER via2 ;
        RECT 2903.610 1847.760 2903.890 1848.040 ;
        RECT 658.350 838.640 658.630 838.920 ;
      LAYER met3 ;
        RECT 2903.585 1848.050 2903.915 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2903.585 1847.750 2924.800 1848.050 ;
        RECT 2903.585 1847.735 2903.915 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 658.325 838.930 658.655 838.945 ;
        RECT 670.000 838.930 674.000 839.320 ;
        RECT 658.325 838.720 674.000 838.930 ;
        RECT 658.325 838.630 670.220 838.720 ;
        RECT 658.325 838.615 658.655 838.630 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 664.770 2077.300 665.090 2077.360 ;
        RECT 2898.990 2077.300 2899.310 2077.360 ;
        RECT 664.770 2077.160 2899.310 2077.300 ;
        RECT 664.770 2077.100 665.090 2077.160 ;
        RECT 2898.990 2077.100 2899.310 2077.160 ;
      LAYER via ;
        RECT 664.800 2077.100 665.060 2077.360 ;
        RECT 2899.020 2077.100 2899.280 2077.360 ;
      LAYER met2 ;
        RECT 2899.010 2082.315 2899.290 2082.685 ;
        RECT 2899.080 2077.390 2899.220 2082.315 ;
        RECT 664.800 2077.070 665.060 2077.390 ;
        RECT 2899.020 2077.070 2899.280 2077.390 ;
        RECT 664.860 843.725 665.000 2077.070 ;
        RECT 664.790 843.355 665.070 843.725 ;
      LAYER via2 ;
        RECT 2899.010 2082.360 2899.290 2082.640 ;
        RECT 664.790 843.400 665.070 843.680 ;
      LAYER met3 ;
        RECT 2898.985 2082.650 2899.315 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2898.985 2082.350 2924.800 2082.650 ;
        RECT 2898.985 2082.335 2899.315 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 664.765 843.690 665.095 843.705 ;
        RECT 670.000 843.690 674.000 844.080 ;
        RECT 664.765 843.480 674.000 843.690 ;
        RECT 664.765 843.390 670.220 843.480 ;
        RECT 664.765 843.375 665.095 843.390 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 665.690 2311.900 666.010 2311.960 ;
        RECT 2898.990 2311.900 2899.310 2311.960 ;
        RECT 665.690 2311.760 2899.310 2311.900 ;
        RECT 665.690 2311.700 666.010 2311.760 ;
        RECT 2898.990 2311.700 2899.310 2311.760 ;
      LAYER via ;
        RECT 665.720 2311.700 665.980 2311.960 ;
        RECT 2899.020 2311.700 2899.280 2311.960 ;
      LAYER met2 ;
        RECT 2899.010 2316.915 2899.290 2317.285 ;
        RECT 2899.080 2311.990 2899.220 2316.915 ;
        RECT 665.720 2311.670 665.980 2311.990 ;
        RECT 2899.020 2311.670 2899.280 2311.990 ;
        RECT 665.780 849.165 665.920 2311.670 ;
        RECT 665.710 848.795 665.990 849.165 ;
      LAYER via2 ;
        RECT 2899.010 2316.960 2899.290 2317.240 ;
        RECT 665.710 848.840 665.990 849.120 ;
      LAYER met3 ;
        RECT 2898.985 2317.250 2899.315 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2898.985 2316.950 2924.800 2317.250 ;
        RECT 2898.985 2316.935 2899.315 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 665.685 849.130 666.015 849.145 ;
        RECT 670.000 849.130 674.000 849.520 ;
        RECT 665.685 848.920 674.000 849.130 ;
        RECT 665.685 848.830 670.220 848.920 ;
        RECT 665.685 848.815 666.015 848.830 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 151.540 662.330 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 662.010 151.400 2901.150 151.540 ;
        RECT 662.010 151.340 662.330 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 662.040 151.340 662.300 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 662.030 601.955 662.310 602.325 ;
        RECT 662.100 151.630 662.240 601.955 ;
        RECT 662.040 151.310 662.300 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 662.030 602.000 662.310 602.280 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 662.005 602.290 662.335 602.305 ;
        RECT 670.000 602.290 674.000 602.680 ;
        RECT 662.005 602.080 674.000 602.290 ;
        RECT 662.005 601.990 670.220 602.080 ;
        RECT 662.005 601.975 662.335 601.990 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 660.630 2491.080 660.950 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 660.630 2490.940 2901.150 2491.080 ;
        RECT 660.630 2490.880 660.950 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
      LAYER via ;
        RECT 660.660 2490.880 660.920 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 660.660 2490.850 660.920 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 660.720 654.685 660.860 2490.850 ;
        RECT 660.650 654.315 660.930 654.685 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
        RECT 660.650 654.360 660.930 654.640 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 660.625 654.650 660.955 654.665 ;
        RECT 670.000 654.650 674.000 655.040 ;
        RECT 660.625 654.440 674.000 654.650 ;
        RECT 660.625 654.350 670.220 654.440 ;
        RECT 660.625 654.335 660.955 654.350 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 1003.920 657.270 1003.980 ;
        RECT 2901.750 1003.920 2902.070 1003.980 ;
        RECT 656.950 1003.780 2902.070 1003.920 ;
        RECT 656.950 1003.720 657.270 1003.780 ;
        RECT 2901.750 1003.720 2902.070 1003.780 ;
        RECT 656.950 991.680 657.270 991.740 ;
        RECT 656.950 991.540 657.640 991.680 ;
        RECT 656.950 991.480 657.270 991.540 ;
        RECT 656.950 980.120 657.270 980.180 ;
        RECT 657.500 980.120 657.640 991.540 ;
        RECT 656.950 979.980 657.640 980.120 ;
        RECT 656.950 979.920 657.270 979.980 ;
      LAYER via ;
        RECT 656.980 1003.720 657.240 1003.980 ;
        RECT 2901.780 1003.720 2902.040 1003.980 ;
        RECT 656.980 991.480 657.240 991.740 ;
        RECT 656.980 979.920 657.240 980.180 ;
      LAYER met2 ;
        RECT 2901.770 2727.635 2902.050 2728.005 ;
        RECT 2901.840 1004.010 2901.980 2727.635 ;
        RECT 656.980 1003.690 657.240 1004.010 ;
        RECT 2901.780 1003.690 2902.040 1004.010 ;
        RECT 657.040 991.770 657.180 1003.690 ;
        RECT 656.980 991.450 657.240 991.770 ;
        RECT 656.980 979.890 657.240 980.210 ;
        RECT 657.040 660.125 657.180 979.890 ;
        RECT 656.970 659.755 657.250 660.125 ;
      LAYER via2 ;
        RECT 2901.770 2727.680 2902.050 2727.960 ;
        RECT 656.970 659.800 657.250 660.080 ;
      LAYER met3 ;
        RECT 2901.745 2727.970 2902.075 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2901.745 2727.670 2924.800 2727.970 ;
        RECT 2901.745 2727.655 2902.075 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 656.945 660.090 657.275 660.105 ;
        RECT 670.000 660.090 674.000 660.480 ;
        RECT 656.945 659.880 674.000 660.090 ;
        RECT 656.945 659.790 670.220 659.880 ;
        RECT 656.945 659.775 657.275 659.790 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 785.310 2961.810 785.590 2961.925 ;
        RECT 786.230 2961.810 786.510 2961.925 ;
        RECT 785.310 2961.670 786.510 2961.810 ;
        RECT 785.310 2961.555 785.590 2961.670 ;
        RECT 786.230 2961.555 786.510 2961.670 ;
        RECT 855.230 2961.555 855.510 2961.925 ;
        RECT 855.300 2959.885 855.440 2961.555 ;
        RECT 855.230 2959.515 855.510 2959.885 ;
      LAYER via2 ;
        RECT 785.310 2961.600 785.590 2961.880 ;
        RECT 786.230 2961.600 786.510 2961.880 ;
        RECT 855.230 2961.600 855.510 2961.880 ;
        RECT 855.230 2959.560 855.510 2959.840 ;
      LAYER met3 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2916.710 2962.270 2924.800 2962.570 ;
        RECT 666.350 2961.890 666.730 2961.900 ;
        RECT 785.285 2961.890 785.615 2961.905 ;
        RECT 666.350 2961.590 785.615 2961.890 ;
        RECT 666.350 2961.580 666.730 2961.590 ;
        RECT 785.285 2961.575 785.615 2961.590 ;
        RECT 786.205 2961.890 786.535 2961.905 ;
        RECT 855.205 2961.890 855.535 2961.905 ;
        RECT 786.205 2961.590 796.410 2961.890 ;
        RECT 786.205 2961.575 786.535 2961.590 ;
        RECT 796.110 2961.210 796.410 2961.590 ;
        RECT 855.205 2961.590 904.050 2961.890 ;
        RECT 855.205 2961.575 855.535 2961.590 ;
        RECT 820.910 2961.210 821.290 2961.220 ;
        RECT 796.110 2960.910 821.290 2961.210 ;
        RECT 903.750 2961.210 904.050 2961.590 ;
        RECT 952.510 2961.590 1000.650 2961.890 ;
        RECT 903.750 2960.910 951.890 2961.210 ;
        RECT 820.910 2960.900 821.290 2960.910 ;
        RECT 951.590 2960.530 951.890 2960.910 ;
        RECT 952.510 2960.530 952.810 2961.590 ;
        RECT 1000.350 2961.210 1000.650 2961.590 ;
        RECT 1049.110 2961.590 1097.250 2961.890 ;
        RECT 1000.350 2960.910 1048.490 2961.210 ;
        RECT 951.590 2960.230 952.810 2960.530 ;
        RECT 1048.190 2960.530 1048.490 2960.910 ;
        RECT 1049.110 2960.530 1049.410 2961.590 ;
        RECT 1096.950 2961.210 1097.250 2961.590 ;
        RECT 1145.710 2961.590 1193.850 2961.890 ;
        RECT 1096.950 2960.910 1145.090 2961.210 ;
        RECT 1048.190 2960.230 1049.410 2960.530 ;
        RECT 1144.790 2960.530 1145.090 2960.910 ;
        RECT 1145.710 2960.530 1146.010 2961.590 ;
        RECT 1193.550 2961.210 1193.850 2961.590 ;
        RECT 1242.310 2961.590 1290.450 2961.890 ;
        RECT 1193.550 2960.910 1241.690 2961.210 ;
        RECT 1144.790 2960.230 1146.010 2960.530 ;
        RECT 1241.390 2960.530 1241.690 2960.910 ;
        RECT 1242.310 2960.530 1242.610 2961.590 ;
        RECT 1290.150 2961.210 1290.450 2961.590 ;
        RECT 1338.910 2961.590 1387.050 2961.890 ;
        RECT 1290.150 2960.910 1338.290 2961.210 ;
        RECT 1241.390 2960.230 1242.610 2960.530 ;
        RECT 1337.990 2960.530 1338.290 2960.910 ;
        RECT 1338.910 2960.530 1339.210 2961.590 ;
        RECT 1386.750 2961.210 1387.050 2961.590 ;
        RECT 1435.510 2961.590 1483.650 2961.890 ;
        RECT 1386.750 2960.910 1434.890 2961.210 ;
        RECT 1337.990 2960.230 1339.210 2960.530 ;
        RECT 1434.590 2960.530 1434.890 2960.910 ;
        RECT 1435.510 2960.530 1435.810 2961.590 ;
        RECT 1483.350 2961.210 1483.650 2961.590 ;
        RECT 1532.110 2961.590 1580.250 2961.890 ;
        RECT 1483.350 2960.910 1531.490 2961.210 ;
        RECT 1434.590 2960.230 1435.810 2960.530 ;
        RECT 1531.190 2960.530 1531.490 2960.910 ;
        RECT 1532.110 2960.530 1532.410 2961.590 ;
        RECT 1579.950 2961.210 1580.250 2961.590 ;
        RECT 1628.710 2961.590 1676.850 2961.890 ;
        RECT 1579.950 2960.910 1628.090 2961.210 ;
        RECT 1531.190 2960.230 1532.410 2960.530 ;
        RECT 1627.790 2960.530 1628.090 2960.910 ;
        RECT 1628.710 2960.530 1629.010 2961.590 ;
        RECT 1676.550 2961.210 1676.850 2961.590 ;
        RECT 1725.310 2961.590 1773.450 2961.890 ;
        RECT 1676.550 2960.910 1724.690 2961.210 ;
        RECT 1627.790 2960.230 1629.010 2960.530 ;
        RECT 1724.390 2960.530 1724.690 2960.910 ;
        RECT 1725.310 2960.530 1725.610 2961.590 ;
        RECT 1773.150 2961.210 1773.450 2961.590 ;
        RECT 1821.910 2961.590 1870.050 2961.890 ;
        RECT 1773.150 2960.910 1821.290 2961.210 ;
        RECT 1724.390 2960.230 1725.610 2960.530 ;
        RECT 1820.990 2960.530 1821.290 2960.910 ;
        RECT 1821.910 2960.530 1822.210 2961.590 ;
        RECT 1869.750 2961.210 1870.050 2961.590 ;
        RECT 1918.510 2961.590 1966.650 2961.890 ;
        RECT 1869.750 2960.910 1917.890 2961.210 ;
        RECT 1820.990 2960.230 1822.210 2960.530 ;
        RECT 1917.590 2960.530 1917.890 2960.910 ;
        RECT 1918.510 2960.530 1918.810 2961.590 ;
        RECT 1966.350 2961.210 1966.650 2961.590 ;
        RECT 2015.110 2961.590 2063.250 2961.890 ;
        RECT 1966.350 2960.910 2014.490 2961.210 ;
        RECT 1917.590 2960.230 1918.810 2960.530 ;
        RECT 2014.190 2960.530 2014.490 2960.910 ;
        RECT 2015.110 2960.530 2015.410 2961.590 ;
        RECT 2062.950 2961.210 2063.250 2961.590 ;
        RECT 2111.710 2961.590 2159.850 2961.890 ;
        RECT 2062.950 2960.910 2111.090 2961.210 ;
        RECT 2014.190 2960.230 2015.410 2960.530 ;
        RECT 2110.790 2960.530 2111.090 2960.910 ;
        RECT 2111.710 2960.530 2112.010 2961.590 ;
        RECT 2159.550 2961.210 2159.850 2961.590 ;
        RECT 2208.310 2961.590 2256.450 2961.890 ;
        RECT 2159.550 2960.910 2207.690 2961.210 ;
        RECT 2110.790 2960.230 2112.010 2960.530 ;
        RECT 2207.390 2960.530 2207.690 2960.910 ;
        RECT 2208.310 2960.530 2208.610 2961.590 ;
        RECT 2256.150 2961.210 2256.450 2961.590 ;
        RECT 2304.910 2961.590 2353.050 2961.890 ;
        RECT 2256.150 2960.910 2304.290 2961.210 ;
        RECT 2207.390 2960.230 2208.610 2960.530 ;
        RECT 2303.990 2960.530 2304.290 2960.910 ;
        RECT 2304.910 2960.530 2305.210 2961.590 ;
        RECT 2352.750 2961.210 2353.050 2961.590 ;
        RECT 2401.510 2961.590 2449.650 2961.890 ;
        RECT 2352.750 2960.910 2400.890 2961.210 ;
        RECT 2303.990 2960.230 2305.210 2960.530 ;
        RECT 2400.590 2960.530 2400.890 2960.910 ;
        RECT 2401.510 2960.530 2401.810 2961.590 ;
        RECT 2449.350 2961.210 2449.650 2961.590 ;
        RECT 2498.110 2961.590 2546.250 2961.890 ;
        RECT 2449.350 2960.910 2497.490 2961.210 ;
        RECT 2400.590 2960.230 2401.810 2960.530 ;
        RECT 2497.190 2960.530 2497.490 2960.910 ;
        RECT 2498.110 2960.530 2498.410 2961.590 ;
        RECT 2545.950 2961.210 2546.250 2961.590 ;
        RECT 2594.710 2961.590 2642.850 2961.890 ;
        RECT 2545.950 2960.910 2594.090 2961.210 ;
        RECT 2497.190 2960.230 2498.410 2960.530 ;
        RECT 2593.790 2960.530 2594.090 2960.910 ;
        RECT 2594.710 2960.530 2595.010 2961.590 ;
        RECT 2642.550 2961.210 2642.850 2961.590 ;
        RECT 2691.310 2961.590 2739.450 2961.890 ;
        RECT 2642.550 2960.910 2690.690 2961.210 ;
        RECT 2593.790 2960.230 2595.010 2960.530 ;
        RECT 2690.390 2960.530 2690.690 2960.910 ;
        RECT 2691.310 2960.530 2691.610 2961.590 ;
        RECT 2739.150 2961.210 2739.450 2961.590 ;
        RECT 2787.910 2961.590 2836.050 2961.890 ;
        RECT 2739.150 2960.910 2787.290 2961.210 ;
        RECT 2690.390 2960.230 2691.610 2960.530 ;
        RECT 2786.990 2960.530 2787.290 2960.910 ;
        RECT 2787.910 2960.530 2788.210 2961.590 ;
        RECT 2835.750 2961.210 2836.050 2961.590 ;
        RECT 2916.710 2961.210 2917.010 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 2835.750 2960.910 2883.890 2961.210 ;
        RECT 2786.990 2960.230 2788.210 2960.530 ;
        RECT 2883.590 2960.530 2883.890 2960.910 ;
        RECT 2884.510 2960.910 2917.010 2961.210 ;
        RECT 2884.510 2960.530 2884.810 2960.910 ;
        RECT 2883.590 2960.230 2884.810 2960.530 ;
        RECT 820.910 2959.850 821.290 2959.860 ;
        RECT 855.205 2959.850 855.535 2959.865 ;
        RECT 820.910 2959.550 855.535 2959.850 ;
        RECT 820.910 2959.540 821.290 2959.550 ;
        RECT 855.205 2959.535 855.535 2959.550 ;
        RECT 666.350 664.850 666.730 664.860 ;
        RECT 670.000 664.850 674.000 665.240 ;
        RECT 666.350 664.640 674.000 664.850 ;
        RECT 666.350 664.550 670.220 664.640 ;
        RECT 666.350 664.540 666.730 664.550 ;
      LAYER via3 ;
        RECT 666.380 2961.580 666.700 2961.900 ;
        RECT 820.940 2960.900 821.260 2961.220 ;
        RECT 820.940 2959.540 821.260 2959.860 ;
        RECT 666.380 664.540 666.700 664.860 ;
      LAYER met4 ;
        RECT 666.375 2961.575 666.705 2961.905 ;
        RECT 666.390 664.865 666.690 2961.575 ;
        RECT 820.935 2960.895 821.265 2961.225 ;
        RECT 820.950 2959.865 821.250 2960.895 ;
        RECT 820.935 2959.535 821.265 2959.865 ;
        RECT 666.375 664.535 666.705 664.865 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 785.310 3196.410 785.590 3196.525 ;
        RECT 786.230 3196.410 786.510 3196.525 ;
        RECT 785.310 3196.270 786.510 3196.410 ;
        RECT 785.310 3196.155 785.590 3196.270 ;
        RECT 786.230 3196.155 786.510 3196.270 ;
        RECT 855.230 3196.155 855.510 3196.525 ;
        RECT 855.300 3194.485 855.440 3196.155 ;
        RECT 855.230 3194.115 855.510 3194.485 ;
      LAYER via2 ;
        RECT 785.310 3196.200 785.590 3196.480 ;
        RECT 786.230 3196.200 786.510 3196.480 ;
        RECT 855.230 3196.200 855.510 3196.480 ;
        RECT 855.230 3194.160 855.510 3194.440 ;
      LAYER met3 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2916.710 3196.870 2924.800 3197.170 ;
        RECT 785.285 3196.490 785.615 3196.505 ;
        RECT 662.710 3196.190 785.615 3196.490 ;
        RECT 658.990 3195.130 659.370 3195.140 ;
        RECT 662.710 3195.130 663.010 3196.190 ;
        RECT 785.285 3196.175 785.615 3196.190 ;
        RECT 786.205 3196.490 786.535 3196.505 ;
        RECT 855.205 3196.490 855.535 3196.505 ;
        RECT 786.205 3196.190 796.410 3196.490 ;
        RECT 786.205 3196.175 786.535 3196.190 ;
        RECT 796.110 3195.810 796.410 3196.190 ;
        RECT 855.205 3196.190 904.050 3196.490 ;
        RECT 855.205 3196.175 855.535 3196.190 ;
        RECT 820.910 3195.810 821.290 3195.820 ;
        RECT 796.110 3195.510 821.290 3195.810 ;
        RECT 903.750 3195.810 904.050 3196.190 ;
        RECT 952.510 3196.190 1000.650 3196.490 ;
        RECT 903.750 3195.510 951.890 3195.810 ;
        RECT 820.910 3195.500 821.290 3195.510 ;
        RECT 658.990 3194.830 663.010 3195.130 ;
        RECT 951.590 3195.130 951.890 3195.510 ;
        RECT 952.510 3195.130 952.810 3196.190 ;
        RECT 1000.350 3195.810 1000.650 3196.190 ;
        RECT 1049.110 3196.190 1097.250 3196.490 ;
        RECT 1000.350 3195.510 1048.490 3195.810 ;
        RECT 951.590 3194.830 952.810 3195.130 ;
        RECT 1048.190 3195.130 1048.490 3195.510 ;
        RECT 1049.110 3195.130 1049.410 3196.190 ;
        RECT 1096.950 3195.810 1097.250 3196.190 ;
        RECT 1145.710 3196.190 1193.850 3196.490 ;
        RECT 1096.950 3195.510 1145.090 3195.810 ;
        RECT 1048.190 3194.830 1049.410 3195.130 ;
        RECT 1144.790 3195.130 1145.090 3195.510 ;
        RECT 1145.710 3195.130 1146.010 3196.190 ;
        RECT 1193.550 3195.810 1193.850 3196.190 ;
        RECT 1242.310 3196.190 1290.450 3196.490 ;
        RECT 1193.550 3195.510 1241.690 3195.810 ;
        RECT 1144.790 3194.830 1146.010 3195.130 ;
        RECT 1241.390 3195.130 1241.690 3195.510 ;
        RECT 1242.310 3195.130 1242.610 3196.190 ;
        RECT 1290.150 3195.810 1290.450 3196.190 ;
        RECT 1338.910 3196.190 1387.050 3196.490 ;
        RECT 1290.150 3195.510 1338.290 3195.810 ;
        RECT 1241.390 3194.830 1242.610 3195.130 ;
        RECT 1337.990 3195.130 1338.290 3195.510 ;
        RECT 1338.910 3195.130 1339.210 3196.190 ;
        RECT 1386.750 3195.810 1387.050 3196.190 ;
        RECT 1435.510 3196.190 1483.650 3196.490 ;
        RECT 1386.750 3195.510 1434.890 3195.810 ;
        RECT 1337.990 3194.830 1339.210 3195.130 ;
        RECT 1434.590 3195.130 1434.890 3195.510 ;
        RECT 1435.510 3195.130 1435.810 3196.190 ;
        RECT 1483.350 3195.810 1483.650 3196.190 ;
        RECT 1532.110 3196.190 1580.250 3196.490 ;
        RECT 1483.350 3195.510 1531.490 3195.810 ;
        RECT 1434.590 3194.830 1435.810 3195.130 ;
        RECT 1531.190 3195.130 1531.490 3195.510 ;
        RECT 1532.110 3195.130 1532.410 3196.190 ;
        RECT 1579.950 3195.810 1580.250 3196.190 ;
        RECT 1628.710 3196.190 1676.850 3196.490 ;
        RECT 1579.950 3195.510 1628.090 3195.810 ;
        RECT 1531.190 3194.830 1532.410 3195.130 ;
        RECT 1627.790 3195.130 1628.090 3195.510 ;
        RECT 1628.710 3195.130 1629.010 3196.190 ;
        RECT 1676.550 3195.810 1676.850 3196.190 ;
        RECT 1725.310 3196.190 1773.450 3196.490 ;
        RECT 1676.550 3195.510 1724.690 3195.810 ;
        RECT 1627.790 3194.830 1629.010 3195.130 ;
        RECT 1724.390 3195.130 1724.690 3195.510 ;
        RECT 1725.310 3195.130 1725.610 3196.190 ;
        RECT 1773.150 3195.810 1773.450 3196.190 ;
        RECT 1821.910 3196.190 1870.050 3196.490 ;
        RECT 1773.150 3195.510 1821.290 3195.810 ;
        RECT 1724.390 3194.830 1725.610 3195.130 ;
        RECT 1820.990 3195.130 1821.290 3195.510 ;
        RECT 1821.910 3195.130 1822.210 3196.190 ;
        RECT 1869.750 3195.810 1870.050 3196.190 ;
        RECT 1918.510 3196.190 1966.650 3196.490 ;
        RECT 1869.750 3195.510 1917.890 3195.810 ;
        RECT 1820.990 3194.830 1822.210 3195.130 ;
        RECT 1917.590 3195.130 1917.890 3195.510 ;
        RECT 1918.510 3195.130 1918.810 3196.190 ;
        RECT 1966.350 3195.810 1966.650 3196.190 ;
        RECT 2015.110 3196.190 2063.250 3196.490 ;
        RECT 1966.350 3195.510 2014.490 3195.810 ;
        RECT 1917.590 3194.830 1918.810 3195.130 ;
        RECT 2014.190 3195.130 2014.490 3195.510 ;
        RECT 2015.110 3195.130 2015.410 3196.190 ;
        RECT 2062.950 3195.810 2063.250 3196.190 ;
        RECT 2111.710 3196.190 2159.850 3196.490 ;
        RECT 2062.950 3195.510 2111.090 3195.810 ;
        RECT 2014.190 3194.830 2015.410 3195.130 ;
        RECT 2110.790 3195.130 2111.090 3195.510 ;
        RECT 2111.710 3195.130 2112.010 3196.190 ;
        RECT 2159.550 3195.810 2159.850 3196.190 ;
        RECT 2208.310 3196.190 2256.450 3196.490 ;
        RECT 2159.550 3195.510 2207.690 3195.810 ;
        RECT 2110.790 3194.830 2112.010 3195.130 ;
        RECT 2207.390 3195.130 2207.690 3195.510 ;
        RECT 2208.310 3195.130 2208.610 3196.190 ;
        RECT 2256.150 3195.810 2256.450 3196.190 ;
        RECT 2304.910 3196.190 2353.050 3196.490 ;
        RECT 2256.150 3195.510 2304.290 3195.810 ;
        RECT 2207.390 3194.830 2208.610 3195.130 ;
        RECT 2303.990 3195.130 2304.290 3195.510 ;
        RECT 2304.910 3195.130 2305.210 3196.190 ;
        RECT 2352.750 3195.810 2353.050 3196.190 ;
        RECT 2401.510 3196.190 2449.650 3196.490 ;
        RECT 2352.750 3195.510 2400.890 3195.810 ;
        RECT 2303.990 3194.830 2305.210 3195.130 ;
        RECT 2400.590 3195.130 2400.890 3195.510 ;
        RECT 2401.510 3195.130 2401.810 3196.190 ;
        RECT 2449.350 3195.810 2449.650 3196.190 ;
        RECT 2498.110 3196.190 2546.250 3196.490 ;
        RECT 2449.350 3195.510 2497.490 3195.810 ;
        RECT 2400.590 3194.830 2401.810 3195.130 ;
        RECT 2497.190 3195.130 2497.490 3195.510 ;
        RECT 2498.110 3195.130 2498.410 3196.190 ;
        RECT 2545.950 3195.810 2546.250 3196.190 ;
        RECT 2594.710 3196.190 2642.850 3196.490 ;
        RECT 2545.950 3195.510 2594.090 3195.810 ;
        RECT 2497.190 3194.830 2498.410 3195.130 ;
        RECT 2593.790 3195.130 2594.090 3195.510 ;
        RECT 2594.710 3195.130 2595.010 3196.190 ;
        RECT 2642.550 3195.810 2642.850 3196.190 ;
        RECT 2691.310 3196.190 2739.450 3196.490 ;
        RECT 2642.550 3195.510 2690.690 3195.810 ;
        RECT 2593.790 3194.830 2595.010 3195.130 ;
        RECT 2690.390 3195.130 2690.690 3195.510 ;
        RECT 2691.310 3195.130 2691.610 3196.190 ;
        RECT 2739.150 3195.810 2739.450 3196.190 ;
        RECT 2787.910 3196.190 2836.050 3196.490 ;
        RECT 2739.150 3195.510 2787.290 3195.810 ;
        RECT 2690.390 3194.830 2691.610 3195.130 ;
        RECT 2786.990 3195.130 2787.290 3195.510 ;
        RECT 2787.910 3195.130 2788.210 3196.190 ;
        RECT 2835.750 3195.810 2836.050 3196.190 ;
        RECT 2916.710 3195.810 2917.010 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 2835.750 3195.510 2883.890 3195.810 ;
        RECT 2786.990 3194.830 2788.210 3195.130 ;
        RECT 2883.590 3195.130 2883.890 3195.510 ;
        RECT 2884.510 3195.510 2917.010 3195.810 ;
        RECT 2884.510 3195.130 2884.810 3195.510 ;
        RECT 2883.590 3194.830 2884.810 3195.130 ;
        RECT 658.990 3194.820 659.370 3194.830 ;
        RECT 820.910 3194.450 821.290 3194.460 ;
        RECT 855.205 3194.450 855.535 3194.465 ;
        RECT 820.910 3194.150 855.535 3194.450 ;
        RECT 820.910 3194.140 821.290 3194.150 ;
        RECT 855.205 3194.135 855.535 3194.150 ;
        RECT 658.990 670.290 659.370 670.300 ;
        RECT 670.000 670.290 674.000 670.680 ;
        RECT 658.990 670.080 674.000 670.290 ;
        RECT 658.990 669.990 670.220 670.080 ;
        RECT 658.990 669.980 659.370 669.990 ;
      LAYER via3 ;
        RECT 659.020 3194.820 659.340 3195.140 ;
        RECT 820.940 3195.500 821.260 3195.820 ;
        RECT 820.940 3194.140 821.260 3194.460 ;
        RECT 659.020 669.980 659.340 670.300 ;
      LAYER met4 ;
        RECT 820.935 3195.495 821.265 3195.825 ;
        RECT 659.015 3194.815 659.345 3195.145 ;
        RECT 659.030 670.305 659.330 3194.815 ;
        RECT 820.950 3194.465 821.250 3195.495 ;
        RECT 820.935 3194.135 821.265 3194.465 ;
        RECT 659.015 669.975 659.345 670.305 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 772.870 3431.520 773.190 3431.580 ;
        RECT 797.250 3431.520 797.570 3431.580 ;
        RECT 772.870 3431.380 797.570 3431.520 ;
        RECT 772.870 3431.320 773.190 3431.380 ;
        RECT 797.250 3431.320 797.570 3431.380 ;
        RECT 676.270 3430.840 676.590 3430.900 ;
        RECT 714.450 3430.840 714.770 3430.900 ;
        RECT 676.270 3430.700 714.770 3430.840 ;
        RECT 676.270 3430.640 676.590 3430.700 ;
        RECT 714.450 3430.640 714.770 3430.700 ;
      LAYER via ;
        RECT 772.900 3431.320 773.160 3431.580 ;
        RECT 797.280 3431.320 797.540 3431.580 ;
        RECT 676.300 3430.640 676.560 3430.900 ;
        RECT 714.480 3430.640 714.740 3430.900 ;
      LAYER met2 ;
        RECT 845.110 3432.115 845.390 3432.485 ;
        RECT 738.850 3431.690 739.130 3431.805 ;
        RECT 738.000 3431.550 739.130 3431.690 ;
        RECT 676.290 3430.755 676.570 3431.125 ;
        RECT 676.300 3430.610 676.560 3430.755 ;
        RECT 714.480 3430.610 714.740 3430.930 ;
        RECT 714.540 3429.765 714.680 3430.610 ;
        RECT 738.000 3430.445 738.140 3431.550 ;
        RECT 738.850 3431.435 739.130 3431.550 ;
        RECT 772.890 3431.435 773.170 3431.805 ;
        RECT 772.900 3431.290 773.160 3431.435 ;
        RECT 797.280 3431.290 797.540 3431.610 ;
        RECT 797.340 3431.125 797.480 3431.290 ;
        RECT 845.180 3431.125 845.320 3432.115 ;
        RECT 797.270 3430.755 797.550 3431.125 ;
        RECT 845.110 3430.755 845.390 3431.125 ;
        RECT 737.930 3430.075 738.210 3430.445 ;
        RECT 714.470 3429.395 714.750 3429.765 ;
      LAYER via2 ;
        RECT 845.110 3432.160 845.390 3432.440 ;
        RECT 676.290 3430.800 676.570 3431.080 ;
        RECT 738.850 3431.480 739.130 3431.760 ;
        RECT 772.890 3431.480 773.170 3431.760 ;
        RECT 797.270 3430.800 797.550 3431.080 ;
        RECT 845.110 3430.800 845.390 3431.080 ;
        RECT 737.930 3430.120 738.210 3430.400 ;
        RECT 714.470 3429.440 714.750 3429.720 ;
      LAYER met3 ;
        RECT 820.910 3432.450 821.290 3432.460 ;
        RECT 845.085 3432.450 845.415 3432.465 ;
        RECT 820.910 3432.150 845.415 3432.450 ;
        RECT 820.910 3432.140 821.290 3432.150 ;
        RECT 845.085 3432.135 845.415 3432.150 ;
        RECT 738.825 3431.770 739.155 3431.785 ;
        RECT 772.865 3431.770 773.195 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 738.825 3431.470 773.195 3431.770 ;
        RECT 738.825 3431.455 739.155 3431.470 ;
        RECT 772.865 3431.455 773.195 3431.470 ;
        RECT 2916.710 3431.470 2924.800 3431.770 ;
        RECT 676.265 3431.090 676.595 3431.105 ;
        RECT 662.710 3430.790 676.595 3431.090 ;
        RECT 659.910 3429.730 660.290 3429.740 ;
        RECT 662.710 3429.730 663.010 3430.790 ;
        RECT 676.265 3430.775 676.595 3430.790 ;
        RECT 797.245 3431.090 797.575 3431.105 ;
        RECT 820.910 3431.090 821.290 3431.100 ;
        RECT 797.245 3430.790 821.290 3431.090 ;
        RECT 797.245 3430.775 797.575 3430.790 ;
        RECT 820.910 3430.780 821.290 3430.790 ;
        RECT 845.085 3431.090 845.415 3431.105 ;
        RECT 845.085 3430.790 904.050 3431.090 ;
        RECT 845.085 3430.775 845.415 3430.790 ;
        RECT 737.905 3430.410 738.235 3430.425 ;
        RECT 724.350 3430.110 738.235 3430.410 ;
        RECT 903.750 3430.410 904.050 3430.790 ;
        RECT 952.510 3430.790 1000.650 3431.090 ;
        RECT 903.750 3430.110 951.890 3430.410 ;
        RECT 659.910 3429.430 663.010 3429.730 ;
        RECT 714.445 3429.730 714.775 3429.745 ;
        RECT 724.350 3429.730 724.650 3430.110 ;
        RECT 737.905 3430.095 738.235 3430.110 ;
        RECT 714.445 3429.430 724.650 3429.730 ;
        RECT 951.590 3429.730 951.890 3430.110 ;
        RECT 952.510 3429.730 952.810 3430.790 ;
        RECT 1000.350 3430.410 1000.650 3430.790 ;
        RECT 1049.110 3430.790 1097.250 3431.090 ;
        RECT 1000.350 3430.110 1048.490 3430.410 ;
        RECT 951.590 3429.430 952.810 3429.730 ;
        RECT 1048.190 3429.730 1048.490 3430.110 ;
        RECT 1049.110 3429.730 1049.410 3430.790 ;
        RECT 1096.950 3430.410 1097.250 3430.790 ;
        RECT 1145.710 3430.790 1193.850 3431.090 ;
        RECT 1096.950 3430.110 1145.090 3430.410 ;
        RECT 1048.190 3429.430 1049.410 3429.730 ;
        RECT 1144.790 3429.730 1145.090 3430.110 ;
        RECT 1145.710 3429.730 1146.010 3430.790 ;
        RECT 1193.550 3430.410 1193.850 3430.790 ;
        RECT 1242.310 3430.790 1290.450 3431.090 ;
        RECT 1193.550 3430.110 1241.690 3430.410 ;
        RECT 1144.790 3429.430 1146.010 3429.730 ;
        RECT 1241.390 3429.730 1241.690 3430.110 ;
        RECT 1242.310 3429.730 1242.610 3430.790 ;
        RECT 1290.150 3430.410 1290.450 3430.790 ;
        RECT 1338.910 3430.790 1387.050 3431.090 ;
        RECT 1290.150 3430.110 1338.290 3430.410 ;
        RECT 1241.390 3429.430 1242.610 3429.730 ;
        RECT 1337.990 3429.730 1338.290 3430.110 ;
        RECT 1338.910 3429.730 1339.210 3430.790 ;
        RECT 1386.750 3430.410 1387.050 3430.790 ;
        RECT 1435.510 3430.790 1483.650 3431.090 ;
        RECT 1386.750 3430.110 1434.890 3430.410 ;
        RECT 1337.990 3429.430 1339.210 3429.730 ;
        RECT 1434.590 3429.730 1434.890 3430.110 ;
        RECT 1435.510 3429.730 1435.810 3430.790 ;
        RECT 1483.350 3430.410 1483.650 3430.790 ;
        RECT 1532.110 3430.790 1580.250 3431.090 ;
        RECT 1483.350 3430.110 1531.490 3430.410 ;
        RECT 1434.590 3429.430 1435.810 3429.730 ;
        RECT 1531.190 3429.730 1531.490 3430.110 ;
        RECT 1532.110 3429.730 1532.410 3430.790 ;
        RECT 1579.950 3430.410 1580.250 3430.790 ;
        RECT 1628.710 3430.790 1676.850 3431.090 ;
        RECT 1579.950 3430.110 1628.090 3430.410 ;
        RECT 1531.190 3429.430 1532.410 3429.730 ;
        RECT 1627.790 3429.730 1628.090 3430.110 ;
        RECT 1628.710 3429.730 1629.010 3430.790 ;
        RECT 1676.550 3430.410 1676.850 3430.790 ;
        RECT 1725.310 3430.790 1773.450 3431.090 ;
        RECT 1676.550 3430.110 1724.690 3430.410 ;
        RECT 1627.790 3429.430 1629.010 3429.730 ;
        RECT 1724.390 3429.730 1724.690 3430.110 ;
        RECT 1725.310 3429.730 1725.610 3430.790 ;
        RECT 1773.150 3430.410 1773.450 3430.790 ;
        RECT 1821.910 3430.790 1870.050 3431.090 ;
        RECT 1773.150 3430.110 1821.290 3430.410 ;
        RECT 1724.390 3429.430 1725.610 3429.730 ;
        RECT 1820.990 3429.730 1821.290 3430.110 ;
        RECT 1821.910 3429.730 1822.210 3430.790 ;
        RECT 1869.750 3430.410 1870.050 3430.790 ;
        RECT 1918.510 3430.790 1966.650 3431.090 ;
        RECT 1869.750 3430.110 1917.890 3430.410 ;
        RECT 1820.990 3429.430 1822.210 3429.730 ;
        RECT 1917.590 3429.730 1917.890 3430.110 ;
        RECT 1918.510 3429.730 1918.810 3430.790 ;
        RECT 1966.350 3430.410 1966.650 3430.790 ;
        RECT 2015.110 3430.790 2063.250 3431.090 ;
        RECT 1966.350 3430.110 2014.490 3430.410 ;
        RECT 1917.590 3429.430 1918.810 3429.730 ;
        RECT 2014.190 3429.730 2014.490 3430.110 ;
        RECT 2015.110 3429.730 2015.410 3430.790 ;
        RECT 2062.950 3430.410 2063.250 3430.790 ;
        RECT 2111.710 3430.790 2159.850 3431.090 ;
        RECT 2062.950 3430.110 2111.090 3430.410 ;
        RECT 2014.190 3429.430 2015.410 3429.730 ;
        RECT 2110.790 3429.730 2111.090 3430.110 ;
        RECT 2111.710 3429.730 2112.010 3430.790 ;
        RECT 2159.550 3430.410 2159.850 3430.790 ;
        RECT 2208.310 3430.790 2256.450 3431.090 ;
        RECT 2159.550 3430.110 2207.690 3430.410 ;
        RECT 2110.790 3429.430 2112.010 3429.730 ;
        RECT 2207.390 3429.730 2207.690 3430.110 ;
        RECT 2208.310 3429.730 2208.610 3430.790 ;
        RECT 2256.150 3430.410 2256.450 3430.790 ;
        RECT 2304.910 3430.790 2353.050 3431.090 ;
        RECT 2256.150 3430.110 2304.290 3430.410 ;
        RECT 2207.390 3429.430 2208.610 3429.730 ;
        RECT 2303.990 3429.730 2304.290 3430.110 ;
        RECT 2304.910 3429.730 2305.210 3430.790 ;
        RECT 2352.750 3430.410 2353.050 3430.790 ;
        RECT 2401.510 3430.790 2449.650 3431.090 ;
        RECT 2352.750 3430.110 2400.890 3430.410 ;
        RECT 2303.990 3429.430 2305.210 3429.730 ;
        RECT 2400.590 3429.730 2400.890 3430.110 ;
        RECT 2401.510 3429.730 2401.810 3430.790 ;
        RECT 2449.350 3430.410 2449.650 3430.790 ;
        RECT 2498.110 3430.790 2546.250 3431.090 ;
        RECT 2449.350 3430.110 2497.490 3430.410 ;
        RECT 2400.590 3429.430 2401.810 3429.730 ;
        RECT 2497.190 3429.730 2497.490 3430.110 ;
        RECT 2498.110 3429.730 2498.410 3430.790 ;
        RECT 2545.950 3430.410 2546.250 3430.790 ;
        RECT 2594.710 3430.790 2642.850 3431.090 ;
        RECT 2545.950 3430.110 2594.090 3430.410 ;
        RECT 2497.190 3429.430 2498.410 3429.730 ;
        RECT 2593.790 3429.730 2594.090 3430.110 ;
        RECT 2594.710 3429.730 2595.010 3430.790 ;
        RECT 2642.550 3430.410 2642.850 3430.790 ;
        RECT 2691.310 3430.790 2739.450 3431.090 ;
        RECT 2642.550 3430.110 2690.690 3430.410 ;
        RECT 2593.790 3429.430 2595.010 3429.730 ;
        RECT 2690.390 3429.730 2690.690 3430.110 ;
        RECT 2691.310 3429.730 2691.610 3430.790 ;
        RECT 2739.150 3430.410 2739.450 3430.790 ;
        RECT 2787.910 3430.790 2836.050 3431.090 ;
        RECT 2739.150 3430.110 2787.290 3430.410 ;
        RECT 2690.390 3429.430 2691.610 3429.730 ;
        RECT 2786.990 3429.730 2787.290 3430.110 ;
        RECT 2787.910 3429.730 2788.210 3430.790 ;
        RECT 2835.750 3430.410 2836.050 3430.790 ;
        RECT 2916.710 3430.410 2917.010 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2835.750 3430.110 2883.890 3430.410 ;
        RECT 2786.990 3429.430 2788.210 3429.730 ;
        RECT 2883.590 3429.730 2883.890 3430.110 ;
        RECT 2884.510 3430.110 2917.010 3430.410 ;
        RECT 2884.510 3429.730 2884.810 3430.110 ;
        RECT 2883.590 3429.430 2884.810 3429.730 ;
        RECT 659.910 3429.420 660.290 3429.430 ;
        RECT 714.445 3429.415 714.775 3429.430 ;
        RECT 659.910 675.730 660.290 675.740 ;
        RECT 670.000 675.730 674.000 676.120 ;
        RECT 659.910 675.520 674.000 675.730 ;
        RECT 659.910 675.430 670.220 675.520 ;
        RECT 659.910 675.420 660.290 675.430 ;
      LAYER via3 ;
        RECT 820.940 3432.140 821.260 3432.460 ;
        RECT 659.940 3429.420 660.260 3429.740 ;
        RECT 820.940 3430.780 821.260 3431.100 ;
        RECT 659.940 675.420 660.260 675.740 ;
      LAYER met4 ;
        RECT 820.935 3432.135 821.265 3432.465 ;
        RECT 820.950 3431.105 821.250 3432.135 ;
        RECT 820.935 3430.775 821.265 3431.105 ;
        RECT 659.935 3429.415 660.265 3429.745 ;
        RECT 659.950 675.745 660.250 3429.415 ;
        RECT 659.935 675.415 660.265 675.745 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.845 2717.520 3517.600 ;
        RECT 2717.310 3501.475 2717.590 3501.845 ;
      LAYER via2 ;
        RECT 2717.310 3501.520 2717.590 3501.800 ;
      LAYER met3 ;
        RECT 661.750 3501.810 662.130 3501.820 ;
        RECT 2717.285 3501.810 2717.615 3501.825 ;
        RECT 661.750 3501.510 2717.615 3501.810 ;
        RECT 661.750 3501.500 662.130 3501.510 ;
        RECT 2717.285 3501.495 2717.615 3501.510 ;
        RECT 661.750 681.170 662.130 681.180 ;
        RECT 670.000 681.170 674.000 681.560 ;
        RECT 661.750 680.960 674.000 681.170 ;
        RECT 661.750 680.870 670.220 680.960 ;
        RECT 661.750 680.860 662.130 680.870 ;
      LAYER via3 ;
        RECT 661.780 3501.500 662.100 3501.820 ;
        RECT 661.780 680.860 662.100 681.180 ;
      LAYER met4 ;
        RECT 661.775 3501.495 662.105 3501.825 ;
        RECT 661.790 681.185 662.090 3501.495 ;
        RECT 661.775 680.855 662.105 681.185 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3502.525 2392.760 3517.600 ;
        RECT 2392.550 3502.155 2392.830 3502.525 ;
      LAYER via2 ;
        RECT 2392.550 3502.200 2392.830 3502.480 ;
      LAYER met3 ;
        RECT 660.830 3502.490 661.210 3502.500 ;
        RECT 2392.525 3502.490 2392.855 3502.505 ;
        RECT 660.830 3502.190 2392.855 3502.490 ;
        RECT 660.830 3502.180 661.210 3502.190 ;
        RECT 2392.525 3502.175 2392.855 3502.190 ;
        RECT 660.830 685.930 661.210 685.940 ;
        RECT 670.000 685.930 674.000 686.320 ;
        RECT 660.830 685.720 674.000 685.930 ;
        RECT 660.830 685.630 670.220 685.720 ;
        RECT 660.830 685.620 661.210 685.630 ;
      LAYER via3 ;
        RECT 660.860 3502.180 661.180 3502.500 ;
        RECT 660.860 685.620 661.180 685.940 ;
      LAYER met4 ;
        RECT 660.855 3502.175 661.185 3502.505 ;
        RECT 660.870 685.945 661.170 3502.175 ;
        RECT 660.855 685.615 661.185 685.945 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 661.550 3502.580 661.870 3502.640 ;
        RECT 2068.230 3502.580 2068.550 3502.640 ;
        RECT 661.550 3502.440 2068.550 3502.580 ;
        RECT 661.550 3502.380 661.870 3502.440 ;
        RECT 2068.230 3502.380 2068.550 3502.440 ;
      LAYER via ;
        RECT 661.580 3502.380 661.840 3502.640 ;
        RECT 2068.260 3502.380 2068.520 3502.640 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3502.670 2068.460 3517.600 ;
        RECT 661.580 3502.350 661.840 3502.670 ;
        RECT 2068.260 3502.350 2068.520 3502.670 ;
        RECT 661.640 691.405 661.780 3502.350 ;
        RECT 661.570 691.035 661.850 691.405 ;
      LAYER via2 ;
        RECT 661.570 691.080 661.850 691.360 ;
      LAYER met3 ;
        RECT 661.545 691.370 661.875 691.385 ;
        RECT 670.000 691.370 674.000 691.760 ;
        RECT 661.545 691.160 674.000 691.370 ;
        RECT 661.545 691.070 670.220 691.160 ;
        RECT 661.545 691.055 661.875 691.070 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 655.570 3503.600 655.890 3503.660 ;
        RECT 1743.930 3503.600 1744.250 3503.660 ;
        RECT 655.570 3503.460 1744.250 3503.600 ;
        RECT 655.570 3503.400 655.890 3503.460 ;
        RECT 1743.930 3503.400 1744.250 3503.460 ;
        RECT 655.570 781.560 655.890 781.620 ;
        RECT 655.570 781.420 657.180 781.560 ;
        RECT 655.570 781.360 655.890 781.420 ;
        RECT 656.490 779.860 656.810 779.920 ;
        RECT 657.040 779.860 657.180 781.420 ;
        RECT 656.490 779.720 657.180 779.860 ;
        RECT 656.490 779.660 656.810 779.720 ;
        RECT 656.490 765.580 656.810 765.640 ;
        RECT 656.490 765.440 657.180 765.580 ;
        RECT 656.490 765.380 656.810 765.440 ;
        RECT 655.570 764.220 655.890 764.280 ;
        RECT 657.040 764.220 657.180 765.440 ;
        RECT 655.570 764.080 657.180 764.220 ;
        RECT 655.570 764.020 655.890 764.080 ;
      LAYER via ;
        RECT 655.600 3503.400 655.860 3503.660 ;
        RECT 1743.960 3503.400 1744.220 3503.660 ;
        RECT 655.600 781.360 655.860 781.620 ;
        RECT 656.520 779.660 656.780 779.920 ;
        RECT 656.520 765.380 656.780 765.640 ;
        RECT 655.600 764.020 655.860 764.280 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3503.690 1744.160 3517.600 ;
        RECT 655.600 3503.370 655.860 3503.690 ;
        RECT 1743.960 3503.370 1744.220 3503.690 ;
        RECT 655.660 781.650 655.800 3503.370 ;
        RECT 655.600 781.330 655.860 781.650 ;
        RECT 656.520 779.630 656.780 779.950 ;
        RECT 656.580 765.670 656.720 779.630 ;
        RECT 656.520 765.350 656.780 765.670 ;
        RECT 655.600 763.990 655.860 764.310 ;
        RECT 655.660 759.290 655.800 763.990 ;
        RECT 655.660 759.150 656.720 759.290 ;
        RECT 656.580 696.845 656.720 759.150 ;
        RECT 656.510 696.475 656.790 696.845 ;
      LAYER via2 ;
        RECT 656.510 696.520 656.790 696.800 ;
      LAYER met3 ;
        RECT 656.485 696.810 656.815 696.825 ;
        RECT 670.000 696.810 674.000 697.200 ;
        RECT 656.485 696.600 674.000 696.810 ;
        RECT 656.485 696.510 670.220 696.600 ;
        RECT 656.485 696.495 656.815 696.510 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 668.910 3504.620 669.230 3504.680 ;
        RECT 1419.170 3504.620 1419.490 3504.680 ;
        RECT 668.910 3504.480 1419.490 3504.620 ;
        RECT 668.910 3504.420 669.230 3504.480 ;
        RECT 1419.170 3504.420 1419.490 3504.480 ;
      LAYER via ;
        RECT 668.940 3504.420 669.200 3504.680 ;
        RECT 1419.200 3504.420 1419.460 3504.680 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3504.710 1419.400 3517.600 ;
        RECT 668.940 3504.390 669.200 3504.710 ;
        RECT 1419.200 3504.390 1419.460 3504.710 ;
        RECT 669.000 702.285 669.140 3504.390 ;
        RECT 668.930 701.915 669.210 702.285 ;
      LAYER via2 ;
        RECT 668.930 701.960 669.210 702.240 ;
      LAYER met3 ;
        RECT 668.905 702.250 669.235 702.265 ;
        RECT 670.000 702.250 674.000 702.640 ;
        RECT 668.905 702.040 674.000 702.250 ;
        RECT 668.905 701.950 670.220 702.040 ;
        RECT 668.905 701.935 669.235 701.950 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 660.630 386.140 660.950 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 660.630 386.000 2901.150 386.140 ;
        RECT 660.630 385.940 660.950 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 660.660 385.940 660.920 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 660.650 606.715 660.930 607.085 ;
        RECT 660.720 386.230 660.860 606.715 ;
        RECT 660.660 385.910 660.920 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 660.650 606.760 660.930 607.040 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 660.625 607.050 660.955 607.065 ;
        RECT 670.000 607.050 674.000 607.440 ;
        RECT 660.625 606.840 674.000 607.050 ;
        RECT 660.625 606.750 670.220 606.840 ;
        RECT 660.625 606.735 660.955 606.750 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 668.450 3503.940 668.770 3504.000 ;
        RECT 1094.870 3503.940 1095.190 3504.000 ;
        RECT 668.450 3503.800 1095.190 3503.940 ;
        RECT 668.450 3503.740 668.770 3503.800 ;
        RECT 1094.870 3503.740 1095.190 3503.800 ;
      LAYER via ;
        RECT 668.480 3503.740 668.740 3504.000 ;
        RECT 1094.900 3503.740 1095.160 3504.000 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3504.030 1095.100 3517.600 ;
        RECT 668.480 3503.710 668.740 3504.030 ;
        RECT 1094.900 3503.710 1095.160 3504.030 ;
        RECT 668.540 707.045 668.680 3503.710 ;
        RECT 668.470 706.675 668.750 707.045 ;
      LAYER via2 ;
        RECT 668.470 706.720 668.750 707.000 ;
      LAYER met3 ;
        RECT 668.445 707.010 668.775 707.025 ;
        RECT 670.000 707.010 674.000 707.400 ;
        RECT 668.445 706.800 674.000 707.010 ;
        RECT 668.445 706.710 670.220 706.800 ;
        RECT 668.445 706.695 668.775 706.710 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 767.810 3491.360 768.130 3491.420 ;
        RECT 771.030 3491.360 771.350 3491.420 ;
        RECT 767.810 3491.220 771.350 3491.360 ;
        RECT 767.810 3491.160 768.130 3491.220 ;
        RECT 771.030 3491.160 771.350 3491.220 ;
        RECT 766.430 3429.820 766.750 3429.880 ;
        RECT 768.270 3429.820 768.590 3429.880 ;
        RECT 766.430 3429.680 768.590 3429.820 ;
        RECT 766.430 3429.620 766.750 3429.680 ;
        RECT 768.270 3429.620 768.590 3429.680 ;
        RECT 766.430 3422.340 766.750 3422.400 ;
        RECT 767.350 3422.340 767.670 3422.400 ;
        RECT 766.430 3422.200 767.670 3422.340 ;
        RECT 766.430 3422.140 766.750 3422.200 ;
        RECT 767.350 3422.140 767.670 3422.200 ;
        RECT 766.430 3284.300 766.750 3284.360 ;
        RECT 767.350 3284.300 767.670 3284.360 ;
        RECT 766.430 3284.160 767.670 3284.300 ;
        RECT 766.430 3284.100 766.750 3284.160 ;
        RECT 767.350 3284.100 767.670 3284.160 ;
        RECT 766.430 3236.360 766.750 3236.420 ;
        RECT 767.810 3236.360 768.130 3236.420 ;
        RECT 766.430 3236.220 768.130 3236.360 ;
        RECT 766.430 3236.160 766.750 3236.220 ;
        RECT 767.810 3236.160 768.130 3236.220 ;
        RECT 766.430 3188.420 766.750 3188.480 ;
        RECT 767.810 3188.420 768.130 3188.480 ;
        RECT 766.430 3188.280 768.130 3188.420 ;
        RECT 766.430 3188.220 766.750 3188.280 ;
        RECT 767.810 3188.220 768.130 3188.280 ;
        RECT 766.890 3153.540 767.210 3153.800 ;
        RECT 766.980 3152.720 767.120 3153.540 ;
        RECT 767.810 3152.720 768.130 3152.780 ;
        RECT 766.980 3152.580 768.130 3152.720 ;
        RECT 767.810 3152.520 768.130 3152.580 ;
        RECT 765.970 3132.660 766.290 3132.720 ;
        RECT 767.810 3132.660 768.130 3132.720 ;
        RECT 765.970 3132.520 768.130 3132.660 ;
        RECT 765.970 3132.460 766.290 3132.520 ;
        RECT 767.810 3132.460 768.130 3132.520 ;
        RECT 765.970 3084.380 766.290 3084.440 ;
        RECT 766.430 3084.380 766.750 3084.440 ;
        RECT 765.970 3084.240 766.750 3084.380 ;
        RECT 765.970 3084.180 766.290 3084.240 ;
        RECT 766.430 3084.180 766.750 3084.240 ;
        RECT 766.430 3056.160 766.750 3056.220 ;
        RECT 767.810 3056.160 768.130 3056.220 ;
        RECT 766.430 3056.020 768.130 3056.160 ;
        RECT 766.430 3055.960 766.750 3056.020 ;
        RECT 767.810 3055.960 768.130 3056.020 ;
        RECT 766.890 2994.960 767.210 2995.020 ;
        RECT 767.810 2994.960 768.130 2995.020 ;
        RECT 766.890 2994.820 768.130 2994.960 ;
        RECT 766.890 2994.760 767.210 2994.820 ;
        RECT 767.810 2994.760 768.130 2994.820 ;
        RECT 765.510 2970.820 765.830 2970.880 ;
        RECT 766.890 2970.820 767.210 2970.880 ;
        RECT 765.510 2970.680 767.210 2970.820 ;
        RECT 765.510 2970.620 765.830 2970.680 ;
        RECT 766.890 2970.620 767.210 2970.680 ;
        RECT 765.510 2912.340 765.830 2912.400 ;
        RECT 766.890 2912.340 767.210 2912.400 ;
        RECT 765.510 2912.200 767.210 2912.340 ;
        RECT 765.510 2912.140 765.830 2912.200 ;
        RECT 766.890 2912.140 767.210 2912.200 ;
        RECT 765.510 2884.800 765.830 2884.860 ;
        RECT 766.430 2884.800 766.750 2884.860 ;
        RECT 765.510 2884.660 766.750 2884.800 ;
        RECT 765.510 2884.600 765.830 2884.660 ;
        RECT 766.430 2884.600 766.750 2884.660 ;
        RECT 765.050 2884.120 765.370 2884.180 ;
        RECT 766.430 2884.120 766.750 2884.180 ;
        RECT 765.050 2883.980 766.750 2884.120 ;
        RECT 765.050 2883.920 765.370 2883.980 ;
        RECT 766.430 2883.920 766.750 2883.980 ;
        RECT 766.430 2670.260 766.750 2670.320 ;
        RECT 767.350 2670.260 767.670 2670.320 ;
        RECT 766.430 2670.120 767.670 2670.260 ;
        RECT 766.430 2670.060 766.750 2670.120 ;
        RECT 767.350 2670.060 767.670 2670.120 ;
        RECT 767.810 2608.380 768.130 2608.440 ;
        RECT 768.730 2608.380 769.050 2608.440 ;
        RECT 767.810 2608.240 769.050 2608.380 ;
        RECT 767.810 2608.180 768.130 2608.240 ;
        RECT 768.730 2608.180 769.050 2608.240 ;
        RECT 766.890 2525.560 767.210 2525.820 ;
        RECT 766.980 2525.420 767.120 2525.560 ;
        RECT 767.350 2525.420 767.670 2525.480 ;
        RECT 766.980 2525.280 767.670 2525.420 ;
        RECT 767.350 2525.220 767.670 2525.280 ;
        RECT 766.890 2511.820 767.210 2511.880 ;
        RECT 767.350 2511.820 767.670 2511.880 ;
        RECT 766.890 2511.680 767.670 2511.820 ;
        RECT 766.890 2511.620 767.210 2511.680 ;
        RECT 767.350 2511.620 767.670 2511.680 ;
        RECT 766.890 2477.140 767.210 2477.200 ;
        RECT 767.810 2477.140 768.130 2477.200 ;
        RECT 766.890 2477.000 768.130 2477.140 ;
        RECT 766.890 2476.940 767.210 2477.000 ;
        RECT 767.810 2476.940 768.130 2477.000 ;
        RECT 766.430 2463.200 766.750 2463.260 ;
        RECT 767.810 2463.200 768.130 2463.260 ;
        RECT 766.430 2463.060 768.130 2463.200 ;
        RECT 766.430 2463.000 766.750 2463.060 ;
        RECT 767.810 2463.000 768.130 2463.060 ;
        RECT 766.430 2380.580 766.750 2380.640 ;
        RECT 767.350 2380.580 767.670 2380.640 ;
        RECT 766.430 2380.440 767.670 2380.580 ;
        RECT 766.430 2380.380 766.750 2380.440 ;
        RECT 767.350 2380.380 767.670 2380.440 ;
        RECT 766.890 2332.100 767.210 2332.360 ;
        RECT 766.980 2331.960 767.120 2332.100 ;
        RECT 767.350 2331.960 767.670 2332.020 ;
        RECT 766.980 2331.820 767.670 2331.960 ;
        RECT 767.350 2331.760 767.670 2331.820 ;
        RECT 767.350 2318.360 767.670 2318.420 ;
        RECT 767.810 2318.360 768.130 2318.420 ;
        RECT 767.350 2318.220 768.130 2318.360 ;
        RECT 767.350 2318.160 767.670 2318.220 ;
        RECT 767.810 2318.160 768.130 2318.220 ;
        RECT 767.810 2284.020 768.130 2284.080 ;
        RECT 767.440 2283.880 768.130 2284.020 ;
        RECT 767.440 2283.740 767.580 2283.880 ;
        RECT 767.810 2283.820 768.130 2283.880 ;
        RECT 767.350 2283.480 767.670 2283.740 ;
        RECT 766.890 2235.740 767.210 2235.800 ;
        RECT 767.810 2235.740 768.130 2235.800 ;
        RECT 766.890 2235.600 768.130 2235.740 ;
        RECT 766.890 2235.540 767.210 2235.600 ;
        RECT 767.810 2235.540 768.130 2235.600 ;
        RECT 766.890 2221.800 767.210 2221.860 ;
        RECT 767.350 2221.800 767.670 2221.860 ;
        RECT 766.890 2221.660 767.670 2221.800 ;
        RECT 766.890 2221.600 767.210 2221.660 ;
        RECT 767.350 2221.600 767.670 2221.660 ;
        RECT 767.350 2187.460 767.670 2187.520 ;
        RECT 766.980 2187.320 767.670 2187.460 ;
        RECT 766.980 2187.180 767.120 2187.320 ;
        RECT 767.350 2187.260 767.670 2187.320 ;
        RECT 766.890 2186.920 767.210 2187.180 ;
        RECT 766.430 2149.380 766.750 2149.440 ;
        RECT 767.350 2149.380 767.670 2149.440 ;
        RECT 766.430 2149.240 767.670 2149.380 ;
        RECT 766.430 2149.180 766.750 2149.240 ;
        RECT 767.350 2149.180 767.670 2149.240 ;
        RECT 765.050 2125.240 765.370 2125.300 ;
        RECT 766.430 2125.240 766.750 2125.300 ;
        RECT 765.050 2125.100 766.750 2125.240 ;
        RECT 765.050 2125.040 765.370 2125.100 ;
        RECT 766.430 2125.040 766.750 2125.100 ;
        RECT 765.970 2042.420 766.290 2042.680 ;
        RECT 766.060 2042.280 766.200 2042.420 ;
        RECT 766.890 2042.280 767.210 2042.340 ;
        RECT 766.060 2042.140 767.210 2042.280 ;
        RECT 766.890 2042.080 767.210 2042.140 ;
        RECT 766.890 1994.480 767.210 1994.740 ;
        RECT 766.980 1994.060 767.120 1994.480 ;
        RECT 766.890 1993.800 767.210 1994.060 ;
        RECT 765.970 1931.780 766.290 1931.840 ;
        RECT 766.430 1931.780 766.750 1931.840 ;
        RECT 765.970 1931.640 766.750 1931.780 ;
        RECT 765.970 1931.580 766.290 1931.640 ;
        RECT 766.430 1931.580 766.750 1931.640 ;
        RECT 765.970 1883.840 766.290 1883.900 ;
        RECT 767.350 1883.840 767.670 1883.900 ;
        RECT 765.970 1883.700 767.670 1883.840 ;
        RECT 765.970 1883.640 766.290 1883.700 ;
        RECT 767.350 1883.640 767.670 1883.700 ;
        RECT 766.430 1835.220 766.750 1835.280 ;
        RECT 767.810 1835.220 768.130 1835.280 ;
        RECT 766.430 1835.080 768.130 1835.220 ;
        RECT 766.430 1835.020 766.750 1835.080 ;
        RECT 767.810 1835.020 768.130 1835.080 ;
        RECT 766.430 1787.280 766.750 1787.340 ;
        RECT 767.350 1787.280 767.670 1787.340 ;
        RECT 766.430 1787.140 767.670 1787.280 ;
        RECT 766.430 1787.080 766.750 1787.140 ;
        RECT 767.350 1787.080 767.670 1787.140 ;
        RECT 767.350 1752.940 767.670 1753.000 ;
        RECT 766.980 1752.800 767.670 1752.940 ;
        RECT 766.980 1752.660 767.120 1752.800 ;
        RECT 767.350 1752.740 767.670 1752.800 ;
        RECT 766.890 1752.400 767.210 1752.660 ;
        RECT 766.890 1594.160 767.210 1594.220 ;
        RECT 767.350 1594.160 767.670 1594.220 ;
        RECT 766.890 1594.020 767.670 1594.160 ;
        RECT 766.890 1593.960 767.210 1594.020 ;
        RECT 767.350 1593.960 767.670 1594.020 ;
        RECT 766.890 1559.820 767.210 1559.880 ;
        RECT 767.350 1559.820 767.670 1559.880 ;
        RECT 766.890 1559.680 767.670 1559.820 ;
        RECT 766.890 1559.620 767.210 1559.680 ;
        RECT 767.350 1559.620 767.670 1559.680 ;
        RECT 766.430 1511.200 766.750 1511.260 ;
        RECT 767.350 1511.200 767.670 1511.260 ;
        RECT 766.430 1511.060 767.670 1511.200 ;
        RECT 766.430 1511.000 766.750 1511.060 ;
        RECT 767.350 1511.000 767.670 1511.060 ;
        RECT 766.430 1414.640 766.750 1414.700 ;
        RECT 767.350 1414.640 767.670 1414.700 ;
        RECT 766.430 1414.500 767.670 1414.640 ;
        RECT 766.430 1414.440 766.750 1414.500 ;
        RECT 767.350 1414.440 767.670 1414.500 ;
        RECT 766.430 1400.700 766.750 1400.760 ;
        RECT 766.890 1400.700 767.210 1400.760 ;
        RECT 766.430 1400.560 767.210 1400.700 ;
        RECT 766.430 1400.500 766.750 1400.560 ;
        RECT 766.890 1400.500 767.210 1400.560 ;
        RECT 766.430 1366.360 766.750 1366.420 ;
        RECT 767.810 1366.360 768.130 1366.420 ;
        RECT 766.430 1366.220 768.130 1366.360 ;
        RECT 766.430 1366.160 766.750 1366.220 ;
        RECT 767.810 1366.160 768.130 1366.220 ;
        RECT 766.890 1352.420 767.210 1352.480 ;
        RECT 767.810 1352.420 768.130 1352.480 ;
        RECT 766.890 1352.280 768.130 1352.420 ;
        RECT 766.890 1352.220 767.210 1352.280 ;
        RECT 767.810 1352.220 768.130 1352.280 ;
        RECT 766.890 1304.480 767.210 1304.540 ;
        RECT 768.270 1304.480 768.590 1304.540 ;
        RECT 766.890 1304.340 768.590 1304.480 ;
        RECT 766.890 1304.280 767.210 1304.340 ;
        RECT 768.270 1304.280 768.590 1304.340 ;
        RECT 768.270 1270.140 768.590 1270.200 ;
        RECT 767.900 1270.000 768.590 1270.140 ;
        RECT 767.900 1269.520 768.040 1270.000 ;
        RECT 768.270 1269.940 768.590 1270.000 ;
        RECT 767.810 1269.260 768.130 1269.520 ;
        RECT 766.430 1173.380 766.750 1173.640 ;
        RECT 766.520 1172.960 766.660 1173.380 ;
        RECT 766.430 1172.700 766.750 1172.960 ;
        RECT 765.970 1124.960 766.290 1125.020 ;
        RECT 765.970 1124.820 766.660 1124.960 ;
        RECT 765.970 1124.760 766.290 1124.820 ;
        RECT 766.520 1124.680 766.660 1124.820 ;
        RECT 766.430 1124.420 766.750 1124.680 ;
        RECT 765.970 1111.020 766.290 1111.080 ;
        RECT 766.430 1111.020 766.750 1111.080 ;
        RECT 765.970 1110.880 766.750 1111.020 ;
        RECT 765.970 1110.820 766.290 1110.880 ;
        RECT 766.430 1110.820 766.750 1110.880 ;
        RECT 765.970 1076.480 766.290 1076.740 ;
        RECT 766.060 1076.000 766.200 1076.480 ;
        RECT 766.430 1076.000 766.750 1076.060 ;
        RECT 766.060 1075.860 766.750 1076.000 ;
        RECT 766.430 1075.800 766.750 1075.860 ;
        RECT 765.970 1062.400 766.290 1062.460 ;
        RECT 766.430 1062.400 766.750 1062.460 ;
        RECT 765.970 1062.260 766.750 1062.400 ;
        RECT 765.970 1062.200 766.290 1062.260 ;
        RECT 766.430 1062.200 766.750 1062.260 ;
        RECT 765.970 1014.460 766.290 1014.520 ;
        RECT 766.890 1014.460 767.210 1014.520 ;
        RECT 765.970 1014.320 767.210 1014.460 ;
        RECT 765.970 1014.260 766.290 1014.320 ;
        RECT 766.890 1014.260 767.210 1014.320 ;
        RECT 667.530 1005.960 667.850 1006.020 ;
        RECT 766.890 1005.960 767.210 1006.020 ;
        RECT 667.530 1005.820 767.210 1005.960 ;
        RECT 667.530 1005.760 667.850 1005.820 ;
        RECT 766.890 1005.760 767.210 1005.820 ;
      LAYER via ;
        RECT 767.840 3491.160 768.100 3491.420 ;
        RECT 771.060 3491.160 771.320 3491.420 ;
        RECT 766.460 3429.620 766.720 3429.880 ;
        RECT 768.300 3429.620 768.560 3429.880 ;
        RECT 766.460 3422.140 766.720 3422.400 ;
        RECT 767.380 3422.140 767.640 3422.400 ;
        RECT 766.460 3284.100 766.720 3284.360 ;
        RECT 767.380 3284.100 767.640 3284.360 ;
        RECT 766.460 3236.160 766.720 3236.420 ;
        RECT 767.840 3236.160 768.100 3236.420 ;
        RECT 766.460 3188.220 766.720 3188.480 ;
        RECT 767.840 3188.220 768.100 3188.480 ;
        RECT 766.920 3153.540 767.180 3153.800 ;
        RECT 767.840 3152.520 768.100 3152.780 ;
        RECT 766.000 3132.460 766.260 3132.720 ;
        RECT 767.840 3132.460 768.100 3132.720 ;
        RECT 766.000 3084.180 766.260 3084.440 ;
        RECT 766.460 3084.180 766.720 3084.440 ;
        RECT 766.460 3055.960 766.720 3056.220 ;
        RECT 767.840 3055.960 768.100 3056.220 ;
        RECT 766.920 2994.760 767.180 2995.020 ;
        RECT 767.840 2994.760 768.100 2995.020 ;
        RECT 765.540 2970.620 765.800 2970.880 ;
        RECT 766.920 2970.620 767.180 2970.880 ;
        RECT 765.540 2912.140 765.800 2912.400 ;
        RECT 766.920 2912.140 767.180 2912.400 ;
        RECT 765.540 2884.600 765.800 2884.860 ;
        RECT 766.460 2884.600 766.720 2884.860 ;
        RECT 765.080 2883.920 765.340 2884.180 ;
        RECT 766.460 2883.920 766.720 2884.180 ;
        RECT 766.460 2670.060 766.720 2670.320 ;
        RECT 767.380 2670.060 767.640 2670.320 ;
        RECT 767.840 2608.180 768.100 2608.440 ;
        RECT 768.760 2608.180 769.020 2608.440 ;
        RECT 766.920 2525.560 767.180 2525.820 ;
        RECT 767.380 2525.220 767.640 2525.480 ;
        RECT 766.920 2511.620 767.180 2511.880 ;
        RECT 767.380 2511.620 767.640 2511.880 ;
        RECT 766.920 2476.940 767.180 2477.200 ;
        RECT 767.840 2476.940 768.100 2477.200 ;
        RECT 766.460 2463.000 766.720 2463.260 ;
        RECT 767.840 2463.000 768.100 2463.260 ;
        RECT 766.460 2380.380 766.720 2380.640 ;
        RECT 767.380 2380.380 767.640 2380.640 ;
        RECT 766.920 2332.100 767.180 2332.360 ;
        RECT 767.380 2331.760 767.640 2332.020 ;
        RECT 767.380 2318.160 767.640 2318.420 ;
        RECT 767.840 2318.160 768.100 2318.420 ;
        RECT 767.840 2283.820 768.100 2284.080 ;
        RECT 767.380 2283.480 767.640 2283.740 ;
        RECT 766.920 2235.540 767.180 2235.800 ;
        RECT 767.840 2235.540 768.100 2235.800 ;
        RECT 766.920 2221.600 767.180 2221.860 ;
        RECT 767.380 2221.600 767.640 2221.860 ;
        RECT 767.380 2187.260 767.640 2187.520 ;
        RECT 766.920 2186.920 767.180 2187.180 ;
        RECT 766.460 2149.180 766.720 2149.440 ;
        RECT 767.380 2149.180 767.640 2149.440 ;
        RECT 765.080 2125.040 765.340 2125.300 ;
        RECT 766.460 2125.040 766.720 2125.300 ;
        RECT 766.000 2042.420 766.260 2042.680 ;
        RECT 766.920 2042.080 767.180 2042.340 ;
        RECT 766.920 1994.480 767.180 1994.740 ;
        RECT 766.920 1993.800 767.180 1994.060 ;
        RECT 766.000 1931.580 766.260 1931.840 ;
        RECT 766.460 1931.580 766.720 1931.840 ;
        RECT 766.000 1883.640 766.260 1883.900 ;
        RECT 767.380 1883.640 767.640 1883.900 ;
        RECT 766.460 1835.020 766.720 1835.280 ;
        RECT 767.840 1835.020 768.100 1835.280 ;
        RECT 766.460 1787.080 766.720 1787.340 ;
        RECT 767.380 1787.080 767.640 1787.340 ;
        RECT 767.380 1752.740 767.640 1753.000 ;
        RECT 766.920 1752.400 767.180 1752.660 ;
        RECT 766.920 1593.960 767.180 1594.220 ;
        RECT 767.380 1593.960 767.640 1594.220 ;
        RECT 766.920 1559.620 767.180 1559.880 ;
        RECT 767.380 1559.620 767.640 1559.880 ;
        RECT 766.460 1511.000 766.720 1511.260 ;
        RECT 767.380 1511.000 767.640 1511.260 ;
        RECT 766.460 1414.440 766.720 1414.700 ;
        RECT 767.380 1414.440 767.640 1414.700 ;
        RECT 766.460 1400.500 766.720 1400.760 ;
        RECT 766.920 1400.500 767.180 1400.760 ;
        RECT 766.460 1366.160 766.720 1366.420 ;
        RECT 767.840 1366.160 768.100 1366.420 ;
        RECT 766.920 1352.220 767.180 1352.480 ;
        RECT 767.840 1352.220 768.100 1352.480 ;
        RECT 766.920 1304.280 767.180 1304.540 ;
        RECT 768.300 1304.280 768.560 1304.540 ;
        RECT 768.300 1269.940 768.560 1270.200 ;
        RECT 767.840 1269.260 768.100 1269.520 ;
        RECT 766.460 1173.380 766.720 1173.640 ;
        RECT 766.460 1172.700 766.720 1172.960 ;
        RECT 766.000 1124.760 766.260 1125.020 ;
        RECT 766.460 1124.420 766.720 1124.680 ;
        RECT 766.000 1110.820 766.260 1111.080 ;
        RECT 766.460 1110.820 766.720 1111.080 ;
        RECT 766.000 1076.480 766.260 1076.740 ;
        RECT 766.460 1075.800 766.720 1076.060 ;
        RECT 766.000 1062.200 766.260 1062.460 ;
        RECT 766.460 1062.200 766.720 1062.460 ;
        RECT 766.000 1014.260 766.260 1014.520 ;
        RECT 766.920 1014.260 767.180 1014.520 ;
        RECT 667.560 1005.760 667.820 1006.020 ;
        RECT 766.920 1005.760 767.180 1006.020 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3517.370 770.800 3517.600 ;
        RECT 770.660 3517.230 771.260 3517.370 ;
        RECT 771.120 3491.450 771.260 3517.230 ;
        RECT 767.840 3491.130 768.100 3491.450 ;
        RECT 771.060 3491.130 771.320 3491.450 ;
        RECT 767.900 3443.930 768.040 3491.130 ;
        RECT 767.900 3443.790 768.500 3443.930 ;
        RECT 768.360 3429.910 768.500 3443.790 ;
        RECT 766.460 3429.590 766.720 3429.910 ;
        RECT 768.300 3429.590 768.560 3429.910 ;
        RECT 766.520 3422.430 766.660 3429.590 ;
        RECT 766.460 3422.110 766.720 3422.430 ;
        RECT 767.380 3422.110 767.640 3422.430 ;
        RECT 767.440 3346.010 767.580 3422.110 ;
        RECT 767.440 3345.870 768.500 3346.010 ;
        RECT 768.360 3298.410 768.500 3345.870 ;
        RECT 767.440 3298.270 768.500 3298.410 ;
        RECT 767.440 3284.390 767.580 3298.270 ;
        RECT 766.460 3284.070 766.720 3284.390 ;
        RECT 767.380 3284.070 767.640 3284.390 ;
        RECT 766.520 3236.450 766.660 3284.070 ;
        RECT 766.460 3236.130 766.720 3236.450 ;
        RECT 767.840 3236.130 768.100 3236.450 ;
        RECT 767.900 3188.510 768.040 3236.130 ;
        RECT 766.460 3188.250 766.720 3188.510 ;
        RECT 766.460 3188.190 767.120 3188.250 ;
        RECT 767.840 3188.190 768.100 3188.510 ;
        RECT 766.520 3188.110 767.120 3188.190 ;
        RECT 766.980 3153.830 767.120 3188.110 ;
        RECT 766.920 3153.510 767.180 3153.830 ;
        RECT 767.840 3152.490 768.100 3152.810 ;
        RECT 767.900 3132.750 768.040 3152.490 ;
        RECT 766.000 3132.430 766.260 3132.750 ;
        RECT 767.840 3132.430 768.100 3132.750 ;
        RECT 766.060 3084.470 766.200 3132.430 ;
        RECT 766.000 3084.150 766.260 3084.470 ;
        RECT 766.460 3084.150 766.720 3084.470 ;
        RECT 766.520 3056.250 766.660 3084.150 ;
        RECT 766.460 3055.930 766.720 3056.250 ;
        RECT 767.840 3055.930 768.100 3056.250 ;
        RECT 767.900 2995.050 768.040 3055.930 ;
        RECT 766.920 2994.730 767.180 2995.050 ;
        RECT 767.840 2994.730 768.100 2995.050 ;
        RECT 766.980 2970.910 767.120 2994.730 ;
        RECT 765.540 2970.590 765.800 2970.910 ;
        RECT 766.920 2970.590 767.180 2970.910 ;
        RECT 765.600 2946.965 765.740 2970.590 ;
        RECT 765.530 2946.595 765.810 2946.965 ;
        RECT 766.450 2946.850 766.730 2946.965 ;
        RECT 766.450 2946.710 767.120 2946.850 ;
        RECT 766.450 2946.595 766.730 2946.710 ;
        RECT 766.980 2912.430 767.120 2946.710 ;
        RECT 765.540 2912.110 765.800 2912.430 ;
        RECT 766.920 2912.110 767.180 2912.430 ;
        RECT 765.600 2884.890 765.740 2912.110 ;
        RECT 765.540 2884.570 765.800 2884.890 ;
        RECT 766.460 2884.570 766.720 2884.890 ;
        RECT 766.520 2884.210 766.660 2884.570 ;
        RECT 765.080 2883.890 765.340 2884.210 ;
        RECT 766.460 2883.890 766.720 2884.210 ;
        RECT 765.140 2836.125 765.280 2883.890 ;
        RECT 765.070 2835.755 765.350 2836.125 ;
        RECT 765.990 2835.755 766.270 2836.125 ;
        RECT 766.060 2691.170 766.200 2835.755 ;
        RECT 766.060 2691.030 766.660 2691.170 ;
        RECT 766.520 2670.350 766.660 2691.030 ;
        RECT 766.460 2670.030 766.720 2670.350 ;
        RECT 767.380 2670.030 767.640 2670.350 ;
        RECT 767.440 2656.605 767.580 2670.030 ;
        RECT 767.370 2656.235 767.650 2656.605 ;
        RECT 768.750 2656.235 769.030 2656.605 ;
        RECT 768.820 2608.470 768.960 2656.235 ;
        RECT 767.840 2608.150 768.100 2608.470 ;
        RECT 768.760 2608.150 769.020 2608.470 ;
        RECT 767.900 2573.530 768.040 2608.150 ;
        RECT 767.440 2573.390 768.040 2573.530 ;
        RECT 767.440 2559.930 767.580 2573.390 ;
        RECT 766.980 2559.790 767.580 2559.930 ;
        RECT 766.980 2525.850 767.120 2559.790 ;
        RECT 766.920 2525.530 767.180 2525.850 ;
        RECT 767.380 2525.190 767.640 2525.510 ;
        RECT 767.440 2511.910 767.580 2525.190 ;
        RECT 766.920 2511.590 767.180 2511.910 ;
        RECT 767.380 2511.590 767.640 2511.910 ;
        RECT 766.980 2477.230 767.120 2511.590 ;
        RECT 766.920 2476.910 767.180 2477.230 ;
        RECT 767.840 2476.910 768.100 2477.230 ;
        RECT 767.900 2463.290 768.040 2476.910 ;
        RECT 766.460 2462.970 766.720 2463.290 ;
        RECT 767.840 2462.970 768.100 2463.290 ;
        RECT 766.520 2415.205 766.660 2462.970 ;
        RECT 766.450 2414.835 766.730 2415.205 ;
        RECT 767.370 2414.835 767.650 2415.205 ;
        RECT 767.440 2380.670 767.580 2414.835 ;
        RECT 766.460 2380.410 766.720 2380.670 ;
        RECT 766.460 2380.350 767.120 2380.410 ;
        RECT 767.380 2380.350 767.640 2380.670 ;
        RECT 766.520 2380.270 767.120 2380.350 ;
        RECT 766.980 2332.390 767.120 2380.270 ;
        RECT 766.920 2332.070 767.180 2332.390 ;
        RECT 767.380 2331.730 767.640 2332.050 ;
        RECT 767.440 2318.450 767.580 2331.730 ;
        RECT 767.380 2318.130 767.640 2318.450 ;
        RECT 767.840 2318.130 768.100 2318.450 ;
        RECT 767.900 2284.110 768.040 2318.130 ;
        RECT 767.840 2283.790 768.100 2284.110 ;
        RECT 767.380 2283.450 767.640 2283.770 ;
        RECT 767.440 2270.250 767.580 2283.450 ;
        RECT 767.440 2270.110 768.040 2270.250 ;
        RECT 767.900 2235.830 768.040 2270.110 ;
        RECT 766.920 2235.510 767.180 2235.830 ;
        RECT 767.840 2235.510 768.100 2235.830 ;
        RECT 766.980 2221.890 767.120 2235.510 ;
        RECT 766.920 2221.570 767.180 2221.890 ;
        RECT 767.380 2221.570 767.640 2221.890 ;
        RECT 767.440 2187.550 767.580 2221.570 ;
        RECT 767.380 2187.230 767.640 2187.550 ;
        RECT 766.920 2186.890 767.180 2187.210 ;
        RECT 766.980 2173.690 767.120 2186.890 ;
        RECT 766.980 2173.550 767.580 2173.690 ;
        RECT 767.440 2149.470 767.580 2173.550 ;
        RECT 766.460 2149.150 766.720 2149.470 ;
        RECT 767.380 2149.150 767.640 2149.470 ;
        RECT 766.520 2125.330 766.660 2149.150 ;
        RECT 765.080 2125.010 765.340 2125.330 ;
        RECT 766.460 2125.010 766.720 2125.330 ;
        RECT 765.140 2077.245 765.280 2125.010 ;
        RECT 765.070 2076.875 765.350 2077.245 ;
        RECT 765.990 2076.875 766.270 2077.245 ;
        RECT 766.060 2042.710 766.200 2076.875 ;
        RECT 766.000 2042.390 766.260 2042.710 ;
        RECT 766.920 2042.050 767.180 2042.370 ;
        RECT 766.980 1994.770 767.120 2042.050 ;
        RECT 766.920 1994.450 767.180 1994.770 ;
        RECT 766.920 1993.770 767.180 1994.090 ;
        RECT 766.980 1945.890 767.120 1993.770 ;
        RECT 766.520 1945.750 767.120 1945.890 ;
        RECT 766.520 1931.870 766.660 1945.750 ;
        RECT 766.000 1931.550 766.260 1931.870 ;
        RECT 766.460 1931.550 766.720 1931.870 ;
        RECT 766.060 1883.930 766.200 1931.550 ;
        RECT 766.000 1883.610 766.260 1883.930 ;
        RECT 767.380 1883.610 767.640 1883.930 ;
        RECT 767.440 1859.530 767.580 1883.610 ;
        RECT 767.440 1859.390 768.040 1859.530 ;
        RECT 767.900 1835.310 768.040 1859.390 ;
        RECT 766.460 1834.990 766.720 1835.310 ;
        RECT 767.840 1834.990 768.100 1835.310 ;
        RECT 766.520 1787.370 766.660 1834.990 ;
        RECT 766.460 1787.050 766.720 1787.370 ;
        RECT 767.380 1787.050 767.640 1787.370 ;
        RECT 767.440 1753.030 767.580 1787.050 ;
        RECT 767.380 1752.710 767.640 1753.030 ;
        RECT 766.920 1752.370 767.180 1752.690 ;
        RECT 766.980 1705.285 767.120 1752.370 ;
        RECT 766.910 1704.915 767.190 1705.285 ;
        RECT 766.910 1703.555 767.190 1703.925 ;
        RECT 766.980 1656.210 767.120 1703.555 ;
        RECT 766.980 1656.070 767.580 1656.210 ;
        RECT 767.440 1594.250 767.580 1656.070 ;
        RECT 766.920 1593.930 767.180 1594.250 ;
        RECT 767.380 1593.930 767.640 1594.250 ;
        RECT 766.980 1559.910 767.120 1593.930 ;
        RECT 766.920 1559.590 767.180 1559.910 ;
        RECT 767.380 1559.590 767.640 1559.910 ;
        RECT 767.440 1511.290 767.580 1559.590 ;
        RECT 766.460 1510.970 766.720 1511.290 ;
        RECT 767.380 1510.970 767.640 1511.290 ;
        RECT 766.520 1510.690 766.660 1510.970 ;
        RECT 766.520 1510.550 767.120 1510.690 ;
        RECT 766.980 1463.090 767.120 1510.550 ;
        RECT 766.980 1462.950 767.580 1463.090 ;
        RECT 767.440 1414.730 767.580 1462.950 ;
        RECT 766.460 1414.410 766.720 1414.730 ;
        RECT 767.380 1414.410 767.640 1414.730 ;
        RECT 766.520 1414.130 766.660 1414.410 ;
        RECT 766.520 1413.990 767.120 1414.130 ;
        RECT 766.980 1400.790 767.120 1413.990 ;
        RECT 766.460 1400.470 766.720 1400.790 ;
        RECT 766.920 1400.470 767.180 1400.790 ;
        RECT 766.520 1366.450 766.660 1400.470 ;
        RECT 766.460 1366.130 766.720 1366.450 ;
        RECT 767.840 1366.130 768.100 1366.450 ;
        RECT 767.900 1352.510 768.040 1366.130 ;
        RECT 766.920 1352.190 767.180 1352.510 ;
        RECT 767.840 1352.190 768.100 1352.510 ;
        RECT 766.980 1304.570 767.120 1352.190 ;
        RECT 766.920 1304.250 767.180 1304.570 ;
        RECT 768.300 1304.250 768.560 1304.570 ;
        RECT 768.360 1270.230 768.500 1304.250 ;
        RECT 768.300 1269.910 768.560 1270.230 ;
        RECT 767.840 1269.230 768.100 1269.550 ;
        RECT 767.900 1221.010 768.040 1269.230 ;
        RECT 766.980 1220.870 768.040 1221.010 ;
        RECT 766.980 1207.410 767.120 1220.870 ;
        RECT 766.520 1207.270 767.120 1207.410 ;
        RECT 766.520 1173.670 766.660 1207.270 ;
        RECT 766.460 1173.350 766.720 1173.670 ;
        RECT 766.460 1172.670 766.720 1172.990 ;
        RECT 766.520 1159.130 766.660 1172.670 ;
        RECT 766.060 1158.990 766.660 1159.130 ;
        RECT 766.060 1125.050 766.200 1158.990 ;
        RECT 766.000 1124.730 766.260 1125.050 ;
        RECT 766.460 1124.390 766.720 1124.710 ;
        RECT 766.520 1111.110 766.660 1124.390 ;
        RECT 766.000 1110.790 766.260 1111.110 ;
        RECT 766.460 1110.790 766.720 1111.110 ;
        RECT 766.060 1076.770 766.200 1110.790 ;
        RECT 766.000 1076.450 766.260 1076.770 ;
        RECT 766.460 1075.770 766.720 1076.090 ;
        RECT 766.520 1062.490 766.660 1075.770 ;
        RECT 766.000 1062.170 766.260 1062.490 ;
        RECT 766.460 1062.170 766.720 1062.490 ;
        RECT 766.060 1014.550 766.200 1062.170 ;
        RECT 766.000 1014.230 766.260 1014.550 ;
        RECT 766.920 1014.230 767.180 1014.550 ;
        RECT 766.980 1006.050 767.120 1014.230 ;
        RECT 667.560 1005.730 667.820 1006.050 ;
        RECT 766.920 1005.730 767.180 1006.050 ;
        RECT 667.620 712.485 667.760 1005.730 ;
        RECT 667.550 712.115 667.830 712.485 ;
      LAYER via2 ;
        RECT 765.530 2946.640 765.810 2946.920 ;
        RECT 766.450 2946.640 766.730 2946.920 ;
        RECT 765.070 2835.800 765.350 2836.080 ;
        RECT 765.990 2835.800 766.270 2836.080 ;
        RECT 767.370 2656.280 767.650 2656.560 ;
        RECT 768.750 2656.280 769.030 2656.560 ;
        RECT 766.450 2414.880 766.730 2415.160 ;
        RECT 767.370 2414.880 767.650 2415.160 ;
        RECT 765.070 2076.920 765.350 2077.200 ;
        RECT 765.990 2076.920 766.270 2077.200 ;
        RECT 766.910 1704.960 767.190 1705.240 ;
        RECT 766.910 1703.600 767.190 1703.880 ;
        RECT 667.550 712.160 667.830 712.440 ;
      LAYER met3 ;
        RECT 765.505 2946.930 765.835 2946.945 ;
        RECT 766.425 2946.930 766.755 2946.945 ;
        RECT 765.505 2946.630 766.755 2946.930 ;
        RECT 765.505 2946.615 765.835 2946.630 ;
        RECT 766.425 2946.615 766.755 2946.630 ;
        RECT 765.045 2836.090 765.375 2836.105 ;
        RECT 765.965 2836.090 766.295 2836.105 ;
        RECT 765.045 2835.790 766.295 2836.090 ;
        RECT 765.045 2835.775 765.375 2835.790 ;
        RECT 765.965 2835.775 766.295 2835.790 ;
        RECT 767.345 2656.570 767.675 2656.585 ;
        RECT 768.725 2656.570 769.055 2656.585 ;
        RECT 767.345 2656.270 769.055 2656.570 ;
        RECT 767.345 2656.255 767.675 2656.270 ;
        RECT 768.725 2656.255 769.055 2656.270 ;
        RECT 766.425 2415.170 766.755 2415.185 ;
        RECT 767.345 2415.170 767.675 2415.185 ;
        RECT 766.425 2414.870 767.675 2415.170 ;
        RECT 766.425 2414.855 766.755 2414.870 ;
        RECT 767.345 2414.855 767.675 2414.870 ;
        RECT 765.045 2077.210 765.375 2077.225 ;
        RECT 765.965 2077.210 766.295 2077.225 ;
        RECT 765.045 2076.910 766.295 2077.210 ;
        RECT 765.045 2076.895 765.375 2076.910 ;
        RECT 765.965 2076.895 766.295 2076.910 ;
        RECT 766.885 1705.250 767.215 1705.265 ;
        RECT 766.670 1704.935 767.215 1705.250 ;
        RECT 766.670 1703.905 766.970 1704.935 ;
        RECT 766.670 1703.590 767.215 1703.905 ;
        RECT 766.885 1703.575 767.215 1703.590 ;
        RECT 667.525 712.450 667.855 712.465 ;
        RECT 670.000 712.450 674.000 712.840 ;
        RECT 667.525 712.240 674.000 712.450 ;
        RECT 667.525 712.150 670.220 712.240 ;
        RECT 667.525 712.135 667.855 712.150 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3501.900 446.130 3501.960 ;
        RECT 631.190 3501.900 631.510 3501.960 ;
        RECT 445.810 3501.760 631.510 3501.900 ;
        RECT 445.810 3501.700 446.130 3501.760 ;
        RECT 631.190 3501.700 631.510 3501.760 ;
        RECT 631.190 1657.200 631.510 1657.460 ;
        RECT 631.280 1656.780 631.420 1657.200 ;
        RECT 631.190 1656.520 631.510 1656.780 ;
        RECT 631.190 722.060 631.510 722.120 ;
        RECT 655.570 722.060 655.890 722.120 ;
        RECT 631.190 721.920 655.890 722.060 ;
        RECT 631.190 721.860 631.510 721.920 ;
        RECT 655.570 721.860 655.890 721.920 ;
      LAYER via ;
        RECT 445.840 3501.700 446.100 3501.960 ;
        RECT 631.220 3501.700 631.480 3501.960 ;
        RECT 631.220 1657.200 631.480 1657.460 ;
        RECT 631.220 1656.520 631.480 1656.780 ;
        RECT 631.220 721.860 631.480 722.120 ;
        RECT 655.600 721.860 655.860 722.120 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3501.990 446.040 3517.600 ;
        RECT 445.840 3501.670 446.100 3501.990 ;
        RECT 631.220 3501.670 631.480 3501.990 ;
        RECT 631.280 1657.490 631.420 3501.670 ;
        RECT 631.220 1657.170 631.480 1657.490 ;
        RECT 631.220 1656.490 631.480 1656.810 ;
        RECT 631.280 722.150 631.420 1656.490 ;
        RECT 631.220 721.830 631.480 722.150 ;
        RECT 655.600 721.830 655.860 722.150 ;
        RECT 655.660 717.925 655.800 721.830 ;
        RECT 655.590 717.555 655.870 717.925 ;
      LAYER via2 ;
        RECT 655.590 717.600 655.870 717.880 ;
      LAYER met3 ;
        RECT 655.565 717.890 655.895 717.905 ;
        RECT 670.000 717.890 674.000 718.280 ;
        RECT 655.565 717.680 674.000 717.890 ;
        RECT 655.565 717.590 670.220 717.680 ;
        RECT 655.565 717.575 655.895 717.590 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 448.200 724.300 483.300 724.440 ;
        RECT 304.130 724.100 304.450 724.160 ;
        RECT 338.170 724.100 338.490 724.160 ;
        RECT 304.130 723.960 338.490 724.100 ;
        RECT 304.130 723.900 304.450 723.960 ;
        RECT 338.170 723.900 338.490 723.960 ;
        RECT 192.810 723.760 193.130 723.820 ;
        RECT 206.610 723.760 206.930 723.820 ;
        RECT 192.810 723.620 206.930 723.760 ;
        RECT 192.810 723.560 193.130 723.620 ;
        RECT 206.610 723.560 206.930 723.620 ;
        RECT 207.070 723.760 207.390 723.820 ;
        RECT 289.410 723.760 289.730 723.820 ;
        RECT 303.210 723.760 303.530 723.820 ;
        RECT 448.200 723.760 448.340 724.300 ;
        RECT 483.160 724.160 483.300 724.300 ;
        RECT 483.070 723.900 483.390 724.160 ;
        RECT 655.570 724.100 655.890 724.160 ;
        RECT 531.000 723.960 544.940 724.100 ;
        RECT 207.070 723.620 213.280 723.760 ;
        RECT 207.070 723.560 207.390 723.620 ;
        RECT 123.810 723.420 124.130 723.480 ;
        RECT 144.970 723.420 145.290 723.480 ;
        RECT 123.810 723.280 145.290 723.420 ;
        RECT 213.140 723.420 213.280 723.620 ;
        RECT 289.410 723.620 303.530 723.760 ;
        RECT 289.410 723.560 289.730 723.620 ;
        RECT 303.210 723.560 303.530 723.620 ;
        RECT 406.340 723.620 448.340 723.760 ;
        RECT 241.570 723.420 241.890 723.480 ;
        RECT 213.140 723.280 241.890 723.420 ;
        RECT 123.810 723.220 124.130 723.280 ;
        RECT 144.970 723.220 145.290 723.280 ;
        RECT 241.570 723.220 241.890 723.280 ;
        RECT 386.010 723.420 386.330 723.480 ;
        RECT 399.810 723.420 400.130 723.480 ;
        RECT 386.010 723.280 400.130 723.420 ;
        RECT 386.010 723.220 386.330 723.280 ;
        RECT 399.810 723.220 400.130 723.280 ;
        RECT 400.270 723.420 400.590 723.480 ;
        RECT 406.340 723.420 406.480 723.620 ;
        RECT 400.270 723.280 406.480 723.420 ;
        RECT 507.450 723.420 507.770 723.480 ;
        RECT 531.000 723.420 531.140 723.960 ;
        RECT 507.450 723.280 531.140 723.420 ;
        RECT 544.800 723.420 544.940 723.960 ;
        RECT 641.400 723.960 655.890 724.100 ;
        RECT 627.510 723.760 627.830 723.820 ;
        RECT 641.400 723.760 641.540 723.960 ;
        RECT 655.570 723.900 655.890 723.960 ;
        RECT 627.510 723.620 641.540 723.760 ;
        RECT 627.510 723.560 627.830 723.620 ;
        RECT 579.670 723.420 579.990 723.480 ;
        RECT 544.800 723.280 579.990 723.420 ;
        RECT 400.270 723.220 400.590 723.280 ;
        RECT 507.450 723.220 507.770 723.280 ;
        RECT 579.670 723.220 579.990 723.280 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 304.160 723.900 304.420 724.160 ;
        RECT 338.200 723.900 338.460 724.160 ;
        RECT 192.840 723.560 193.100 723.820 ;
        RECT 206.640 723.560 206.900 723.820 ;
        RECT 207.100 723.560 207.360 723.820 ;
        RECT 123.840 723.220 124.100 723.480 ;
        RECT 145.000 723.220 145.260 723.480 ;
        RECT 289.440 723.560 289.700 723.820 ;
        RECT 303.240 723.560 303.500 723.820 ;
        RECT 483.100 723.900 483.360 724.160 ;
        RECT 241.600 723.220 241.860 723.480 ;
        RECT 386.040 723.220 386.300 723.480 ;
        RECT 399.840 723.220 400.100 723.480 ;
        RECT 400.300 723.220 400.560 723.480 ;
        RECT 507.480 723.220 507.740 723.480 ;
        RECT 627.540 723.560 627.800 723.820 ;
        RECT 655.600 723.900 655.860 724.160 ;
        RECT 579.700 723.220 579.960 723.480 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 723.510 124.040 3498.270 ;
        RECT 304.160 723.930 304.420 724.190 ;
        RECT 338.200 724.045 338.460 724.190 ;
        RECT 206.700 723.850 207.300 723.930 ;
        RECT 303.300 723.870 304.420 723.930 ;
        RECT 303.300 723.850 304.360 723.870 ;
        RECT 192.840 723.530 193.100 723.850 ;
        RECT 206.640 723.790 207.360 723.850 ;
        RECT 206.640 723.530 206.900 723.790 ;
        RECT 207.100 723.530 207.360 723.790 ;
        RECT 289.440 723.530 289.700 723.850 ;
        RECT 303.240 723.790 304.360 723.850 ;
        RECT 303.240 723.530 303.500 723.790 ;
        RECT 338.190 723.675 338.470 724.045 ;
        RECT 386.030 723.675 386.310 724.045 ;
        RECT 483.100 723.930 483.360 724.190 ;
        RECT 483.550 723.930 483.830 724.045 ;
        RECT 483.100 723.870 483.830 723.930 ;
        RECT 483.160 723.790 483.830 723.870 ;
        RECT 483.550 723.675 483.830 723.790 ;
        RECT 507.470 723.675 507.750 724.045 ;
        RECT 655.600 723.870 655.860 724.190 ;
        RECT 123.840 723.190 124.100 723.510 ;
        RECT 145.000 723.365 145.260 723.510 ;
        RECT 192.900 723.365 193.040 723.530 ;
        RECT 241.600 723.365 241.860 723.510 ;
        RECT 289.500 723.365 289.640 723.530 ;
        RECT 386.100 723.510 386.240 723.675 ;
        RECT 507.540 723.510 507.680 723.675 ;
        RECT 627.540 723.530 627.800 723.850 ;
        RECT 144.990 722.995 145.270 723.365 ;
        RECT 192.830 722.995 193.110 723.365 ;
        RECT 241.590 722.995 241.870 723.365 ;
        RECT 289.430 722.995 289.710 723.365 ;
        RECT 386.040 723.190 386.300 723.510 ;
        RECT 399.840 723.250 400.100 723.510 ;
        RECT 400.300 723.250 400.560 723.510 ;
        RECT 399.840 723.190 400.560 723.250 ;
        RECT 507.480 723.190 507.740 723.510 ;
        RECT 579.700 723.365 579.960 723.510 ;
        RECT 627.600 723.365 627.740 723.530 ;
        RECT 399.900 723.110 400.500 723.190 ;
        RECT 579.690 722.995 579.970 723.365 ;
        RECT 627.530 722.995 627.810 723.365 ;
        RECT 655.660 722.685 655.800 723.870 ;
        RECT 655.590 722.315 655.870 722.685 ;
      LAYER via2 ;
        RECT 338.190 723.720 338.470 724.000 ;
        RECT 386.030 723.720 386.310 724.000 ;
        RECT 483.550 723.720 483.830 724.000 ;
        RECT 507.470 723.720 507.750 724.000 ;
        RECT 144.990 723.040 145.270 723.320 ;
        RECT 192.830 723.040 193.110 723.320 ;
        RECT 241.590 723.040 241.870 723.320 ;
        RECT 289.430 723.040 289.710 723.320 ;
        RECT 579.690 723.040 579.970 723.320 ;
        RECT 627.530 723.040 627.810 723.320 ;
        RECT 655.590 722.360 655.870 722.640 ;
      LAYER met3 ;
        RECT 338.165 724.010 338.495 724.025 ;
        RECT 386.005 724.010 386.335 724.025 ;
        RECT 338.165 723.710 386.335 724.010 ;
        RECT 338.165 723.695 338.495 723.710 ;
        RECT 386.005 723.695 386.335 723.710 ;
        RECT 483.525 724.010 483.855 724.025 ;
        RECT 507.445 724.010 507.775 724.025 ;
        RECT 483.525 723.710 507.775 724.010 ;
        RECT 483.525 723.695 483.855 723.710 ;
        RECT 507.445 723.695 507.775 723.710 ;
        RECT 144.965 723.330 145.295 723.345 ;
        RECT 192.805 723.330 193.135 723.345 ;
        RECT 144.965 723.030 193.135 723.330 ;
        RECT 144.965 723.015 145.295 723.030 ;
        RECT 192.805 723.015 193.135 723.030 ;
        RECT 241.565 723.330 241.895 723.345 ;
        RECT 289.405 723.330 289.735 723.345 ;
        RECT 241.565 723.030 289.735 723.330 ;
        RECT 241.565 723.015 241.895 723.030 ;
        RECT 289.405 723.015 289.735 723.030 ;
        RECT 579.665 723.330 579.995 723.345 ;
        RECT 627.505 723.330 627.835 723.345 ;
        RECT 579.665 723.030 627.835 723.330 ;
        RECT 579.665 723.015 579.995 723.030 ;
        RECT 627.505 723.015 627.835 723.030 ;
        RECT 655.565 722.650 655.895 722.665 ;
        RECT 670.000 722.650 674.000 723.040 ;
        RECT 655.565 722.440 674.000 722.650 ;
        RECT 655.565 722.350 670.220 722.440 ;
        RECT 655.565 722.335 655.895 722.350 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 99.890 3339.720 100.210 3339.780 ;
        RECT 17.090 3339.580 100.210 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 99.890 3339.520 100.210 3339.580 ;
        RECT 99.890 731.240 100.210 731.300 ;
        RECT 655.570 731.240 655.890 731.300 ;
        RECT 99.890 731.100 655.890 731.240 ;
        RECT 99.890 731.040 100.210 731.100 ;
        RECT 655.570 731.040 655.890 731.100 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 99.920 3339.520 100.180 3339.780 ;
        RECT 99.920 731.040 100.180 731.300 ;
        RECT 655.600 731.040 655.860 731.300 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 99.920 3339.490 100.180 3339.810 ;
        RECT 99.980 731.330 100.120 3339.490 ;
        RECT 99.920 731.010 100.180 731.330 ;
        RECT 655.600 731.010 655.860 731.330 ;
        RECT 655.660 728.125 655.800 731.010 ;
        RECT 655.590 727.755 655.870 728.125 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 655.590 727.800 655.870 728.080 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 655.565 728.090 655.895 728.105 ;
        RECT 670.000 728.090 674.000 728.480 ;
        RECT 655.565 727.880 674.000 728.090 ;
        RECT 655.565 727.790 670.220 727.880 ;
        RECT 655.565 727.775 655.895 727.790 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 106.790 3050.040 107.110 3050.100 ;
        RECT 17.090 3049.900 107.110 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 106.790 3049.840 107.110 3049.900 ;
        RECT 106.790 738.040 107.110 738.100 ;
        RECT 655.570 738.040 655.890 738.100 ;
        RECT 106.790 737.900 655.890 738.040 ;
        RECT 106.790 737.840 107.110 737.900 ;
        RECT 655.570 737.840 655.890 737.900 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 106.820 3049.840 107.080 3050.100 ;
        RECT 106.820 737.840 107.080 738.100 ;
        RECT 655.600 737.840 655.860 738.100 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 106.820 3049.810 107.080 3050.130 ;
        RECT 106.880 738.130 107.020 3049.810 ;
        RECT 106.820 737.810 107.080 738.130 ;
        RECT 655.600 737.810 655.860 738.130 ;
        RECT 655.660 733.565 655.800 737.810 ;
        RECT 655.590 733.195 655.870 733.565 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 655.590 733.240 655.870 733.520 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 655.565 733.530 655.895 733.545 ;
        RECT 670.000 733.530 674.000 733.920 ;
        RECT 655.565 733.320 674.000 733.530 ;
        RECT 655.565 733.230 670.220 733.320 ;
        RECT 655.565 733.215 655.895 733.230 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2760.360 16.030 2760.420 ;
        RECT 141.290 2760.360 141.610 2760.420 ;
        RECT 15.710 2760.220 141.610 2760.360 ;
        RECT 15.710 2760.160 16.030 2760.220 ;
        RECT 141.290 2760.160 141.610 2760.220 ;
        RECT 141.290 745.180 141.610 745.240 ;
        RECT 141.290 745.040 656.260 745.180 ;
        RECT 141.290 744.980 141.610 745.040 ;
        RECT 656.120 744.500 656.260 745.040 ;
        RECT 655.660 744.360 656.260 744.500 ;
        RECT 655.660 743.200 655.800 744.360 ;
        RECT 655.570 742.940 655.890 743.200 ;
      LAYER via ;
        RECT 15.740 2760.160 16.000 2760.420 ;
        RECT 141.320 2760.160 141.580 2760.420 ;
        RECT 141.320 744.980 141.580 745.240 ;
        RECT 655.600 742.940 655.860 743.200 ;
      LAYER met2 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
        RECT 15.800 2760.450 15.940 2765.035 ;
        RECT 15.740 2760.130 16.000 2760.450 ;
        RECT 141.320 2760.130 141.580 2760.450 ;
        RECT 141.380 745.270 141.520 2760.130 ;
        RECT 141.320 744.950 141.580 745.270 ;
        RECT 655.600 742.910 655.860 743.230 ;
        RECT 655.660 739.005 655.800 742.910 ;
        RECT 655.590 738.635 655.870 739.005 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
        RECT 655.590 738.680 655.870 738.960 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.800 2765.070 16.035 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
        RECT 655.565 738.970 655.895 738.985 ;
        RECT 670.000 738.970 674.000 739.360 ;
        RECT 655.565 738.760 674.000 738.970 ;
        RECT 655.565 738.670 670.220 738.760 ;
        RECT 655.565 738.655 655.895 738.670 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2477.480 16.950 2477.540 ;
        RECT 155.090 2477.480 155.410 2477.540 ;
        RECT 16.630 2477.340 155.410 2477.480 ;
        RECT 16.630 2477.280 16.950 2477.340 ;
        RECT 155.090 2477.280 155.410 2477.340 ;
        RECT 155.090 744.840 155.410 744.900 ;
        RECT 655.570 744.840 655.890 744.900 ;
        RECT 155.090 744.700 655.890 744.840 ;
        RECT 155.090 744.640 155.410 744.700 ;
        RECT 655.570 744.640 655.890 744.700 ;
      LAYER via ;
        RECT 16.660 2477.280 16.920 2477.540 ;
        RECT 155.120 2477.280 155.380 2477.540 ;
        RECT 155.120 744.640 155.380 744.900 ;
        RECT 655.600 744.640 655.860 744.900 ;
      LAYER met2 ;
        RECT 16.650 2477.395 16.930 2477.765 ;
        RECT 16.660 2477.250 16.920 2477.395 ;
        RECT 155.120 2477.250 155.380 2477.570 ;
        RECT 155.180 744.930 155.320 2477.250 ;
        RECT 155.120 744.610 155.380 744.930 ;
        RECT 655.600 744.610 655.860 744.930 ;
        RECT 655.660 743.765 655.800 744.610 ;
        RECT 655.590 743.395 655.870 743.765 ;
      LAYER via2 ;
        RECT 16.650 2477.440 16.930 2477.720 ;
        RECT 655.590 743.440 655.870 743.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 16.625 2477.730 16.955 2477.745 ;
        RECT -4.800 2477.430 16.955 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 16.625 2477.415 16.955 2477.430 ;
        RECT 655.565 743.730 655.895 743.745 ;
        RECT 670.000 743.730 674.000 744.120 ;
        RECT 655.565 743.520 674.000 743.730 ;
        RECT 655.565 743.430 670.220 743.520 ;
        RECT 655.565 743.415 655.895 743.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 751.980 18.790 752.040 ;
        RECT 655.570 751.980 655.890 752.040 ;
        RECT 18.470 751.840 655.890 751.980 ;
        RECT 18.470 751.780 18.790 751.840 ;
        RECT 655.570 751.780 655.890 751.840 ;
      LAYER via ;
        RECT 18.500 751.780 18.760 752.040 ;
        RECT 655.600 751.780 655.860 752.040 ;
      LAYER met2 ;
        RECT 18.490 2189.755 18.770 2190.125 ;
        RECT 18.560 752.070 18.700 2189.755 ;
        RECT 18.500 751.750 18.760 752.070 ;
        RECT 655.600 751.750 655.860 752.070 ;
        RECT 655.660 749.205 655.800 751.750 ;
        RECT 655.590 748.835 655.870 749.205 ;
      LAYER via2 ;
        RECT 18.490 2189.800 18.770 2190.080 ;
        RECT 655.590 748.880 655.870 749.160 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 18.465 2190.090 18.795 2190.105 ;
        RECT -4.800 2189.790 18.795 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 18.465 2189.775 18.795 2189.790 ;
        RECT 655.565 749.170 655.895 749.185 ;
        RECT 670.000 749.170 674.000 749.560 ;
        RECT 655.565 748.960 674.000 749.170 ;
        RECT 655.565 748.870 670.220 748.960 ;
        RECT 655.565 748.855 655.895 748.870 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 758.780 19.250 758.840 ;
        RECT 655.570 758.780 655.890 758.840 ;
        RECT 18.930 758.640 655.890 758.780 ;
        RECT 18.930 758.580 19.250 758.640 ;
        RECT 655.570 758.580 655.890 758.640 ;
      LAYER via ;
        RECT 18.960 758.580 19.220 758.840 ;
        RECT 655.600 758.580 655.860 758.840 ;
      LAYER met2 ;
        RECT 18.950 1902.795 19.230 1903.165 ;
        RECT 19.020 758.870 19.160 1902.795 ;
        RECT 18.960 758.550 19.220 758.870 ;
        RECT 655.600 758.550 655.860 758.870 ;
        RECT 655.660 754.645 655.800 758.550 ;
        RECT 655.590 754.275 655.870 754.645 ;
      LAYER via2 ;
        RECT 18.950 1902.840 19.230 1903.120 ;
        RECT 655.590 754.320 655.870 754.600 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 18.925 1903.130 19.255 1903.145 ;
        RECT -4.800 1902.830 19.255 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 18.925 1902.815 19.255 1902.830 ;
        RECT 655.565 754.610 655.895 754.625 ;
        RECT 670.000 754.610 674.000 755.000 ;
        RECT 655.565 754.400 674.000 754.610 ;
        RECT 655.565 754.310 670.220 754.400 ;
        RECT 655.565 754.295 655.895 754.310 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 670.290 604.080 670.610 604.140 ;
        RECT 2904.510 604.080 2904.830 604.140 ;
        RECT 670.290 603.940 2904.830 604.080 ;
        RECT 670.290 603.880 670.610 603.940 ;
        RECT 2904.510 603.880 2904.830 603.940 ;
      LAYER via ;
        RECT 670.320 603.880 670.580 604.140 ;
        RECT 2904.540 603.880 2904.800 604.140 ;
      LAYER met2 ;
        RECT 2904.530 615.555 2904.810 615.925 ;
        RECT 670.310 609.435 670.590 609.805 ;
        RECT 670.380 604.170 670.520 609.435 ;
        RECT 2904.600 604.170 2904.740 615.555 ;
        RECT 670.320 603.850 670.580 604.170 ;
        RECT 2904.540 603.850 2904.800 604.170 ;
      LAYER via2 ;
        RECT 2904.530 615.600 2904.810 615.880 ;
        RECT 670.310 609.480 670.590 609.760 ;
      LAYER met3 ;
        RECT 2904.505 615.890 2904.835 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2904.505 615.590 2924.800 615.890 ;
        RECT 2904.505 615.575 2904.835 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
        RECT 670.000 612.280 674.000 612.880 ;
        RECT 670.070 609.785 670.370 612.280 ;
        RECT 670.070 609.470 670.615 609.785 ;
        RECT 670.285 609.455 670.615 609.470 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.770 765.580 435.090 765.640 ;
        RECT 186.000 765.440 303.900 765.580 ;
        RECT 96.210 765.240 96.530 765.300 ;
        RECT 61.800 765.100 96.530 765.240 ;
        RECT 48.000 764.760 48.600 764.900 ;
        RECT 19.850 764.560 20.170 764.620 ;
        RECT 48.000 764.560 48.140 764.760 ;
        RECT 19.850 764.420 48.140 764.560 ;
        RECT 48.460 764.560 48.600 764.760 ;
        RECT 61.800 764.560 61.940 765.100 ;
        RECT 96.210 765.040 96.530 765.100 ;
        RECT 111.390 765.240 111.710 765.300 ;
        RECT 138.070 765.240 138.390 765.300 ;
        RECT 111.390 765.100 138.390 765.240 ;
        RECT 111.390 765.040 111.710 765.100 ;
        RECT 138.070 765.040 138.390 765.100 ;
        RECT 169.350 765.240 169.670 765.300 ;
        RECT 186.000 765.240 186.140 765.440 ;
        RECT 169.350 765.100 186.140 765.240 ;
        RECT 303.760 765.240 303.900 765.440 ;
        RECT 427.500 765.440 435.090 765.580 ;
        RECT 427.500 765.300 427.640 765.440 ;
        RECT 434.770 765.380 435.090 765.440 ;
        RECT 303.760 765.100 362.320 765.240 ;
        RECT 169.350 765.040 169.670 765.100 ;
        RECT 362.180 764.900 362.320 765.100 ;
        RECT 427.410 765.040 427.730 765.300 ;
        RECT 579.300 765.100 596.460 765.240 ;
        RECT 379.570 764.900 379.890 764.960 ;
        RECT 362.180 764.760 379.890 764.900 ;
        RECT 379.570 764.700 379.890 764.760 ;
        RECT 524.010 764.900 524.330 764.960 ;
        RECT 544.710 764.900 545.030 764.960 ;
        RECT 524.010 764.760 545.030 764.900 ;
        RECT 524.010 764.700 524.330 764.760 ;
        RECT 544.710 764.700 545.030 764.760 ;
        RECT 545.170 764.900 545.490 764.960 ;
        RECT 579.300 764.900 579.440 765.100 ;
        RECT 545.170 764.760 579.440 764.900 ;
        RECT 545.170 764.700 545.490 764.760 ;
        RECT 48.460 764.420 61.940 764.560 ;
        RECT 596.320 764.560 596.460 765.100 ;
        RECT 656.490 764.560 656.810 764.620 ;
        RECT 596.320 764.420 656.810 764.560 ;
        RECT 19.850 764.360 20.170 764.420 ;
        RECT 656.490 764.360 656.810 764.420 ;
      LAYER via ;
        RECT 19.880 764.360 20.140 764.620 ;
        RECT 96.240 765.040 96.500 765.300 ;
        RECT 111.420 765.040 111.680 765.300 ;
        RECT 138.100 765.040 138.360 765.300 ;
        RECT 169.380 765.040 169.640 765.300 ;
        RECT 434.800 765.380 435.060 765.640 ;
        RECT 427.440 765.040 427.700 765.300 ;
        RECT 379.600 764.700 379.860 764.960 ;
        RECT 524.040 764.700 524.300 764.960 ;
        RECT 544.740 764.700 545.000 764.960 ;
        RECT 545.200 764.700 545.460 764.960 ;
        RECT 656.520 764.360 656.780 764.620 ;
      LAYER met2 ;
        RECT 19.870 1615.155 20.150 1615.525 ;
        RECT 19.940 764.650 20.080 1615.155 ;
        RECT 434.800 765.525 435.060 765.670 ;
        RECT 96.230 765.155 96.510 765.525 ;
        RECT 111.410 765.155 111.690 765.525 ;
        RECT 138.090 765.155 138.370 765.525 ;
        RECT 169.370 765.155 169.650 765.525 ;
        RECT 96.240 765.010 96.500 765.155 ;
        RECT 111.420 765.010 111.680 765.155 ;
        RECT 138.100 765.010 138.360 765.155 ;
        RECT 169.380 765.010 169.640 765.155 ;
        RECT 427.440 765.010 427.700 765.330 ;
        RECT 434.790 765.155 435.070 765.525 ;
        RECT 523.570 765.155 523.850 765.525 ;
        RECT 379.600 764.845 379.860 764.990 ;
        RECT 427.500 764.845 427.640 765.010 ;
        RECT 19.880 764.330 20.140 764.650 ;
        RECT 379.590 764.475 379.870 764.845 ;
        RECT 427.430 764.475 427.710 764.845 ;
        RECT 523.640 764.730 523.780 765.155 ;
        RECT 524.040 764.730 524.300 764.990 ;
        RECT 523.640 764.670 524.300 764.730 ;
        RECT 544.740 764.730 545.000 764.990 ;
        RECT 545.200 764.730 545.460 764.990 ;
        RECT 544.740 764.670 545.460 764.730 ;
        RECT 523.640 764.590 524.240 764.670 ;
        RECT 544.800 764.590 545.400 764.670 ;
        RECT 656.520 764.330 656.780 764.650 ;
        RECT 656.580 760.085 656.720 764.330 ;
        RECT 656.510 759.715 656.790 760.085 ;
      LAYER via2 ;
        RECT 19.870 1615.200 20.150 1615.480 ;
        RECT 96.230 765.200 96.510 765.480 ;
        RECT 111.410 765.200 111.690 765.480 ;
        RECT 138.090 765.200 138.370 765.480 ;
        RECT 169.370 765.200 169.650 765.480 ;
        RECT 434.790 765.200 435.070 765.480 ;
        RECT 523.570 765.200 523.850 765.480 ;
        RECT 379.590 764.520 379.870 764.800 ;
        RECT 427.430 764.520 427.710 764.800 ;
        RECT 656.510 759.760 656.790 760.040 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 19.845 1615.490 20.175 1615.505 ;
        RECT -4.800 1615.190 20.175 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 19.845 1615.175 20.175 1615.190 ;
        RECT 96.205 765.490 96.535 765.505 ;
        RECT 111.385 765.490 111.715 765.505 ;
        RECT 96.205 765.190 111.715 765.490 ;
        RECT 96.205 765.175 96.535 765.190 ;
        RECT 111.385 765.175 111.715 765.190 ;
        RECT 138.065 765.490 138.395 765.505 ;
        RECT 169.345 765.490 169.675 765.505 ;
        RECT 138.065 765.190 169.675 765.490 ;
        RECT 138.065 765.175 138.395 765.190 ;
        RECT 169.345 765.175 169.675 765.190 ;
        RECT 434.765 765.490 435.095 765.505 ;
        RECT 523.545 765.490 523.875 765.505 ;
        RECT 434.765 765.190 523.875 765.490 ;
        RECT 434.765 765.175 435.095 765.190 ;
        RECT 523.545 765.175 523.875 765.190 ;
        RECT 379.565 764.810 379.895 764.825 ;
        RECT 427.405 764.810 427.735 764.825 ;
        RECT 379.565 764.510 427.735 764.810 ;
        RECT 379.565 764.495 379.895 764.510 ;
        RECT 427.405 764.495 427.735 764.510 ;
        RECT 656.485 760.050 656.815 760.065 ;
        RECT 670.000 760.050 674.000 760.440 ;
        RECT 656.485 759.840 674.000 760.050 ;
        RECT 656.485 759.750 670.220 759.840 ;
        RECT 656.485 759.735 656.815 759.750 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 765.920 20.630 765.980 ;
        RECT 655.570 765.920 655.890 765.980 ;
        RECT 20.310 765.780 655.890 765.920 ;
        RECT 20.310 765.720 20.630 765.780 ;
        RECT 655.570 765.720 655.890 765.780 ;
      LAYER via ;
        RECT 20.340 765.720 20.600 765.980 ;
        RECT 655.600 765.720 655.860 765.980 ;
      LAYER met2 ;
        RECT 20.330 1400.275 20.610 1400.645 ;
        RECT 20.400 766.010 20.540 1400.275 ;
        RECT 20.340 765.690 20.600 766.010 ;
        RECT 655.600 765.690 655.860 766.010 ;
        RECT 655.660 764.845 655.800 765.690 ;
        RECT 655.590 764.475 655.870 764.845 ;
      LAYER via2 ;
        RECT 20.330 1400.320 20.610 1400.600 ;
        RECT 655.590 764.520 655.870 764.800 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 20.305 1400.610 20.635 1400.625 ;
        RECT -4.800 1400.310 20.635 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 20.305 1400.295 20.635 1400.310 ;
        RECT 655.565 764.810 655.895 764.825 ;
        RECT 670.000 764.810 674.000 765.200 ;
        RECT 655.565 764.600 674.000 764.810 ;
        RECT 655.565 764.510 670.220 764.600 ;
        RECT 655.565 764.495 655.895 764.510 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 303.210 772.720 303.530 772.780 ;
        RECT 158.400 772.580 303.530 772.720 ;
        RECT 158.400 772.380 158.540 772.580 ;
        RECT 303.210 772.520 303.530 772.580 ;
        RECT 448.570 772.380 448.890 772.440 ;
        RECT 655.570 772.380 655.890 772.440 ;
        RECT 110.560 772.240 158.540 772.380 ;
        RECT 304.220 772.240 351.740 772.380 ;
        RECT 62.170 772.040 62.490 772.100 ;
        RECT 110.560 772.040 110.700 772.240 ;
        RECT 62.170 771.900 110.700 772.040 ;
        RECT 303.210 772.040 303.530 772.100 ;
        RECT 304.220 772.040 304.360 772.240 ;
        RECT 303.210 771.900 304.360 772.040 ;
        RECT 351.600 772.040 351.740 772.240 ;
        RECT 448.570 772.240 497.100 772.380 ;
        RECT 448.570 772.180 448.890 772.240 ;
        RECT 496.960 772.040 497.100 772.240 ;
        RECT 579.760 772.240 655.890 772.380 ;
        RECT 351.600 771.900 410.620 772.040 ;
        RECT 496.960 771.900 544.940 772.040 ;
        RECT 62.170 771.840 62.490 771.900 ;
        RECT 303.210 771.840 303.530 771.900 ;
        RECT 16.630 771.700 16.950 771.760 ;
        RECT 61.710 771.700 62.030 771.760 ;
        RECT 16.630 771.560 62.030 771.700 ;
        RECT 410.480 771.700 410.620 771.900 ;
        RECT 448.110 771.700 448.430 771.760 ;
        RECT 410.480 771.560 448.430 771.700 ;
        RECT 544.800 771.700 544.940 771.900 ;
        RECT 579.760 771.700 579.900 772.240 ;
        RECT 655.570 772.180 655.890 772.240 ;
        RECT 544.800 771.560 579.900 771.700 ;
        RECT 16.630 771.500 16.950 771.560 ;
        RECT 61.710 771.500 62.030 771.560 ;
        RECT 448.110 771.500 448.430 771.560 ;
      LAYER via ;
        RECT 303.240 772.520 303.500 772.780 ;
        RECT 62.200 771.840 62.460 772.100 ;
        RECT 303.240 771.840 303.500 772.100 ;
        RECT 448.600 772.180 448.860 772.440 ;
        RECT 16.660 771.500 16.920 771.760 ;
        RECT 61.740 771.500 62.000 771.760 ;
        RECT 448.140 771.500 448.400 771.760 ;
        RECT 655.600 772.180 655.860 772.440 ;
      LAYER met2 ;
        RECT 16.650 1184.715 16.930 1185.085 ;
        RECT 16.720 771.790 16.860 1184.715 ;
        RECT 303.240 772.490 303.500 772.810 ;
        RECT 303.300 772.130 303.440 772.490 ;
        RECT 448.600 772.210 448.860 772.470 ;
        RECT 448.200 772.150 448.860 772.210 ;
        RECT 655.600 772.150 655.860 772.470 ;
        RECT 62.200 771.810 62.460 772.130 ;
        RECT 303.240 771.810 303.500 772.130 ;
        RECT 448.200 772.070 448.800 772.150 ;
        RECT 16.660 771.470 16.920 771.790 ;
        RECT 61.740 771.530 62.000 771.790 ;
        RECT 62.260 771.530 62.400 771.810 ;
        RECT 448.200 771.790 448.340 772.070 ;
        RECT 61.740 771.470 62.400 771.530 ;
        RECT 448.140 771.470 448.400 771.790 ;
        RECT 61.800 771.390 62.400 771.470 ;
        RECT 655.660 770.285 655.800 772.150 ;
        RECT 655.590 769.915 655.870 770.285 ;
      LAYER via2 ;
        RECT 16.650 1184.760 16.930 1185.040 ;
        RECT 655.590 769.960 655.870 770.240 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 16.625 1185.050 16.955 1185.065 ;
        RECT -4.800 1184.750 16.955 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 16.625 1184.735 16.955 1184.750 ;
        RECT 655.565 770.250 655.895 770.265 ;
        RECT 670.000 770.250 674.000 770.640 ;
        RECT 655.565 770.040 674.000 770.250 ;
        RECT 655.565 769.950 670.220 770.040 ;
        RECT 655.565 769.935 655.895 769.950 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 779.520 18.330 779.580 ;
        RECT 655.570 779.520 655.890 779.580 ;
        RECT 18.010 779.380 655.890 779.520 ;
        RECT 18.010 779.320 18.330 779.380 ;
        RECT 655.570 779.320 655.890 779.380 ;
      LAYER via ;
        RECT 18.040 779.320 18.300 779.580 ;
        RECT 655.600 779.320 655.860 779.580 ;
      LAYER met2 ;
        RECT 18.030 969.155 18.310 969.525 ;
        RECT 18.100 779.610 18.240 969.155 ;
        RECT 18.040 779.290 18.300 779.610 ;
        RECT 655.600 779.290 655.860 779.610 ;
        RECT 655.660 775.725 655.800 779.290 ;
        RECT 655.590 775.355 655.870 775.725 ;
      LAYER via2 ;
        RECT 18.030 969.200 18.310 969.480 ;
        RECT 655.590 775.400 655.870 775.680 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 18.005 969.490 18.335 969.505 ;
        RECT -4.800 969.190 18.335 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 18.005 969.175 18.335 969.190 ;
        RECT 655.565 775.690 655.895 775.705 ;
        RECT 670.000 775.690 674.000 776.080 ;
        RECT 655.565 775.480 674.000 775.690 ;
        RECT 655.565 775.390 670.220 775.480 ;
        RECT 655.565 775.375 655.895 775.390 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 780.200 16.490 780.260 ;
        RECT 655.570 780.200 655.890 780.260 ;
        RECT 16.170 780.060 655.890 780.200 ;
        RECT 16.170 780.000 16.490 780.060 ;
        RECT 655.570 780.000 655.890 780.060 ;
      LAYER via ;
        RECT 16.200 780.000 16.460 780.260 ;
        RECT 655.600 780.000 655.860 780.260 ;
      LAYER met2 ;
        RECT 655.590 780.795 655.870 781.165 ;
        RECT 655.660 780.290 655.800 780.795 ;
        RECT 16.200 779.970 16.460 780.290 ;
        RECT 655.600 779.970 655.860 780.290 ;
        RECT 16.260 753.965 16.400 779.970 ;
        RECT 16.190 753.595 16.470 753.965 ;
      LAYER via2 ;
        RECT 655.590 780.840 655.870 781.120 ;
        RECT 16.190 753.640 16.470 753.920 ;
      LAYER met3 ;
        RECT 655.565 781.130 655.895 781.145 ;
        RECT 670.000 781.130 674.000 781.520 ;
        RECT 655.565 780.920 674.000 781.130 ;
        RECT 655.565 780.830 670.220 780.920 ;
        RECT 655.565 780.815 655.895 780.830 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 16.165 753.930 16.495 753.945 ;
        RECT -4.800 753.630 16.495 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 16.165 753.615 16.495 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 780.540 17.870 780.600 ;
        RECT 656.490 780.540 656.810 780.600 ;
        RECT 17.550 780.400 656.810 780.540 ;
        RECT 17.550 780.340 17.870 780.400 ;
        RECT 656.490 780.340 656.810 780.400 ;
      LAYER via ;
        RECT 17.580 780.340 17.840 780.600 ;
        RECT 656.520 780.340 656.780 780.600 ;
      LAYER met2 ;
        RECT 656.510 785.555 656.790 785.925 ;
        RECT 656.580 780.630 656.720 785.555 ;
        RECT 17.580 780.310 17.840 780.630 ;
        RECT 656.520 780.310 656.780 780.630 ;
        RECT 17.640 538.405 17.780 780.310 ;
        RECT 17.570 538.035 17.850 538.405 ;
      LAYER via2 ;
        RECT 656.510 785.600 656.790 785.880 ;
        RECT 17.570 538.080 17.850 538.360 ;
      LAYER met3 ;
        RECT 656.485 785.890 656.815 785.905 ;
        RECT 670.000 785.890 674.000 786.280 ;
        RECT 656.485 785.680 674.000 785.890 ;
        RECT 656.485 785.590 670.220 785.680 ;
        RECT 656.485 785.575 656.815 785.590 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 17.545 538.370 17.875 538.385 ;
        RECT -4.800 538.070 17.875 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 17.545 538.055 17.875 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 658.330 324.260 658.650 324.320 ;
        RECT 16.630 324.120 658.650 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 658.330 324.060 658.650 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 658.360 324.060 658.620 324.320 ;
      LAYER met2 ;
        RECT 658.350 790.995 658.630 791.365 ;
        RECT 658.420 324.350 658.560 790.995 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 658.360 324.030 658.620 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 658.350 791.040 658.630 791.320 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 658.325 791.330 658.655 791.345 ;
        RECT 670.000 791.330 674.000 791.720 ;
        RECT 658.325 791.120 674.000 791.330 ;
        RECT 658.325 791.030 670.220 791.120 ;
        RECT 658.325 791.015 658.655 791.030 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 661.090 110.400 661.410 110.460 ;
        RECT 15.710 110.260 661.410 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 661.090 110.200 661.410 110.260 ;
      LAYER via ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 661.120 110.200 661.380 110.460 ;
      LAYER met2 ;
        RECT 661.110 796.435 661.390 796.805 ;
        RECT 661.180 110.490 661.320 796.435 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 661.120 110.170 661.380 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 661.110 796.480 661.390 796.760 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 661.085 796.770 661.415 796.785 ;
        RECT 670.000 796.770 674.000 797.160 ;
        RECT 661.085 796.560 674.000 796.770 ;
        RECT 661.085 796.470 670.220 796.560 ;
        RECT 661.085 796.455 661.415 796.470 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 669.830 603.400 670.150 603.460 ;
        RECT 2901.290 603.400 2901.610 603.460 ;
        RECT 669.830 603.260 2901.610 603.400 ;
        RECT 669.830 603.200 670.150 603.260 ;
        RECT 2901.290 603.200 2901.610 603.260 ;
      LAYER via ;
        RECT 669.860 603.200 670.120 603.460 ;
        RECT 2901.320 603.200 2901.580 603.460 ;
      LAYER met2 ;
        RECT 2901.310 850.155 2901.590 850.525 ;
        RECT 669.850 614.875 670.130 615.245 ;
        RECT 669.920 603.490 670.060 614.875 ;
        RECT 2901.380 603.490 2901.520 850.155 ;
        RECT 669.860 603.170 670.120 603.490 ;
        RECT 2901.320 603.170 2901.580 603.490 ;
      LAYER via2 ;
        RECT 2901.310 850.200 2901.590 850.480 ;
        RECT 669.850 614.920 670.130 615.200 ;
      LAYER met3 ;
        RECT 2901.285 850.490 2901.615 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2901.285 850.190 2924.800 850.490 ;
        RECT 2901.285 850.175 2901.615 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT 670.000 617.720 674.000 618.320 ;
        RECT 670.070 615.225 670.370 617.720 ;
        RECT 669.825 614.910 670.370 615.225 ;
        RECT 669.825 614.895 670.155 614.910 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 657.410 1083.480 657.730 1083.540 ;
        RECT 2898.070 1083.480 2898.390 1083.540 ;
        RECT 657.410 1083.340 2898.390 1083.480 ;
        RECT 657.410 1083.280 657.730 1083.340 ;
        RECT 2898.070 1083.280 2898.390 1083.340 ;
      LAYER via ;
        RECT 657.440 1083.280 657.700 1083.540 ;
        RECT 2898.100 1083.280 2898.360 1083.540 ;
      LAYER met2 ;
        RECT 2898.090 1084.755 2898.370 1085.125 ;
        RECT 2898.160 1083.570 2898.300 1084.755 ;
        RECT 657.440 1083.250 657.700 1083.570 ;
        RECT 2898.100 1083.250 2898.360 1083.570 ;
        RECT 657.500 622.725 657.640 1083.250 ;
        RECT 657.430 622.355 657.710 622.725 ;
      LAYER via2 ;
        RECT 2898.090 1084.800 2898.370 1085.080 ;
        RECT 657.430 622.400 657.710 622.680 ;
      LAYER met3 ;
        RECT 2898.065 1085.090 2898.395 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2898.065 1084.790 2924.800 1085.090 ;
        RECT 2898.065 1084.775 2898.395 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
        RECT 657.405 622.690 657.735 622.705 ;
        RECT 670.000 622.690 674.000 623.080 ;
        RECT 657.405 622.480 674.000 622.690 ;
        RECT 657.405 622.390 670.220 622.480 ;
        RECT 657.405 622.375 657.735 622.390 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 657.870 1318.080 658.190 1318.140 ;
        RECT 2900.830 1318.080 2901.150 1318.140 ;
        RECT 657.870 1317.940 2901.150 1318.080 ;
        RECT 657.870 1317.880 658.190 1317.940 ;
        RECT 2900.830 1317.880 2901.150 1317.940 ;
      LAYER via ;
        RECT 657.900 1317.880 658.160 1318.140 ;
        RECT 2900.860 1317.880 2901.120 1318.140 ;
      LAYER met2 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
        RECT 2900.920 1318.170 2901.060 1319.355 ;
        RECT 657.900 1317.850 658.160 1318.170 ;
        RECT 2900.860 1317.850 2901.120 1318.170 ;
        RECT 657.960 628.165 658.100 1317.850 ;
        RECT 657.890 627.795 658.170 628.165 ;
      LAYER via2 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
        RECT 657.890 627.840 658.170 628.120 ;
      LAYER met3 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 657.865 628.130 658.195 628.145 ;
        RECT 670.000 628.130 674.000 628.520 ;
        RECT 657.865 627.920 674.000 628.130 ;
        RECT 657.865 627.830 670.220 627.920 ;
        RECT 657.865 627.815 658.195 627.830 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 659.250 1552.680 659.570 1552.740 ;
        RECT 2898.530 1552.680 2898.850 1552.740 ;
        RECT 659.250 1552.540 2898.850 1552.680 ;
        RECT 659.250 1552.480 659.570 1552.540 ;
        RECT 2898.530 1552.480 2898.850 1552.540 ;
      LAYER via ;
        RECT 659.280 1552.480 659.540 1552.740 ;
        RECT 2898.560 1552.480 2898.820 1552.740 ;
      LAYER met2 ;
        RECT 2898.550 1553.955 2898.830 1554.325 ;
        RECT 2898.620 1552.770 2898.760 1553.955 ;
        RECT 659.280 1552.450 659.540 1552.770 ;
        RECT 2898.560 1552.450 2898.820 1552.770 ;
        RECT 659.340 633.605 659.480 1552.450 ;
        RECT 659.270 633.235 659.550 633.605 ;
      LAYER via2 ;
        RECT 2898.550 1554.000 2898.830 1554.280 ;
        RECT 659.270 633.280 659.550 633.560 ;
      LAYER met3 ;
        RECT 2898.525 1554.290 2898.855 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2898.525 1553.990 2924.800 1554.290 ;
        RECT 2898.525 1553.975 2898.855 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 659.245 633.570 659.575 633.585 ;
        RECT 670.000 633.570 674.000 633.960 ;
        RECT 659.245 633.360 674.000 633.570 ;
        RECT 659.245 633.270 670.220 633.360 ;
        RECT 659.245 633.255 659.575 633.270 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 660.170 1708.060 660.490 1708.120 ;
        RECT 2904.050 1708.060 2904.370 1708.120 ;
        RECT 660.170 1707.920 2904.370 1708.060 ;
        RECT 660.170 1707.860 660.490 1707.920 ;
        RECT 2904.050 1707.860 2904.370 1707.920 ;
      LAYER via ;
        RECT 660.200 1707.860 660.460 1708.120 ;
        RECT 2904.080 1707.860 2904.340 1708.120 ;
      LAYER met2 ;
        RECT 2904.070 1789.235 2904.350 1789.605 ;
        RECT 2904.140 1708.150 2904.280 1789.235 ;
        RECT 660.200 1707.830 660.460 1708.150 ;
        RECT 2904.080 1707.830 2904.340 1708.150 ;
        RECT 660.260 639.045 660.400 1707.830 ;
        RECT 660.190 638.675 660.470 639.045 ;
      LAYER via2 ;
        RECT 2904.070 1789.280 2904.350 1789.560 ;
        RECT 660.190 638.720 660.470 639.000 ;
      LAYER met3 ;
        RECT 2904.045 1789.570 2904.375 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2904.045 1789.270 2924.800 1789.570 ;
        RECT 2904.045 1789.255 2904.375 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 660.165 639.010 660.495 639.025 ;
        RECT 670.000 639.010 674.000 639.400 ;
        RECT 660.165 638.800 674.000 639.010 ;
        RECT 660.165 638.710 670.220 638.800 ;
        RECT 660.165 638.695 660.495 638.710 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 659.710 1708.400 660.030 1708.460 ;
        RECT 2903.130 1708.400 2903.450 1708.460 ;
        RECT 659.710 1708.260 2903.450 1708.400 ;
        RECT 659.710 1708.200 660.030 1708.260 ;
        RECT 2903.130 1708.200 2903.450 1708.260 ;
      LAYER via ;
        RECT 659.740 1708.200 660.000 1708.460 ;
        RECT 2903.160 1708.200 2903.420 1708.460 ;
      LAYER met2 ;
        RECT 2903.150 2023.835 2903.430 2024.205 ;
        RECT 2903.220 1708.490 2903.360 2023.835 ;
        RECT 659.740 1708.170 660.000 1708.490 ;
        RECT 2903.160 1708.170 2903.420 1708.490 ;
        RECT 659.800 643.805 659.940 1708.170 ;
        RECT 659.730 643.435 660.010 643.805 ;
      LAYER via2 ;
        RECT 2903.150 2023.880 2903.430 2024.160 ;
        RECT 659.730 643.480 660.010 643.760 ;
      LAYER met3 ;
        RECT 2903.125 2024.170 2903.455 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2903.125 2023.870 2924.800 2024.170 ;
        RECT 2903.125 2023.855 2903.455 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 659.705 643.770 660.035 643.785 ;
        RECT 670.000 643.770 674.000 644.160 ;
        RECT 659.705 643.560 674.000 643.770 ;
        RECT 659.705 643.470 670.220 643.560 ;
        RECT 659.705 643.455 660.035 643.470 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 666.150 2256.480 666.470 2256.540 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 666.150 2256.340 2901.150 2256.480 ;
        RECT 666.150 2256.280 666.470 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
      LAYER via ;
        RECT 666.180 2256.280 666.440 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 666.180 2256.250 666.440 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 666.240 649.245 666.380 2256.250 ;
        RECT 666.170 648.875 666.450 649.245 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
        RECT 666.170 648.920 666.450 649.200 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 666.145 649.210 666.475 649.225 ;
        RECT 670.000 649.210 674.000 649.600 ;
        RECT 666.145 649.000 674.000 649.210 ;
        RECT 666.145 648.910 670.220 649.000 ;
        RECT 666.145 648.895 666.475 648.910 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 37.300 633.350 37.360 ;
        RECT 994.130 37.300 994.450 37.360 ;
        RECT 633.030 37.160 994.450 37.300 ;
        RECT 633.030 37.100 633.350 37.160 ;
        RECT 994.130 37.100 994.450 37.160 ;
      LAYER via ;
        RECT 633.060 37.100 633.320 37.360 ;
        RECT 994.160 37.100 994.420 37.360 ;
      LAYER met2 ;
        RECT 995.770 600.170 996.050 604.000 ;
        RECT 994.220 600.030 996.050 600.170 ;
        RECT 994.220 37.390 994.360 600.030 ;
        RECT 995.770 600.000 996.050 600.030 ;
        RECT 633.060 37.070 633.320 37.390 ;
        RECT 994.160 37.070 994.420 37.390 ;
        RECT 633.120 2.400 633.260 37.070 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1914.590 579.940 1914.910 580.000 ;
        RECT 1915.510 579.940 1915.830 580.000 ;
        RECT 1914.590 579.800 1915.830 579.940 ;
        RECT 1914.590 579.740 1914.910 579.800 ;
        RECT 1915.510 579.740 1915.830 579.800 ;
        RECT 1916.430 497.320 1916.750 497.380 ;
        RECT 1916.060 497.180 1916.750 497.320 ;
        RECT 1916.060 496.700 1916.200 497.180 ;
        RECT 1916.430 497.120 1916.750 497.180 ;
        RECT 1915.970 496.440 1916.290 496.700 ;
        RECT 1914.590 483.040 1914.910 483.100 ;
        RECT 1915.970 483.040 1916.290 483.100 ;
        RECT 1914.590 482.900 1916.290 483.040 ;
        RECT 1914.590 482.840 1914.910 482.900 ;
        RECT 1915.970 482.840 1916.290 482.900 ;
        RECT 1914.590 435.100 1914.910 435.160 ;
        RECT 1915.510 435.100 1915.830 435.160 ;
        RECT 1914.590 434.960 1915.830 435.100 ;
        RECT 1914.590 434.900 1914.910 434.960 ;
        RECT 1915.510 434.900 1915.830 434.960 ;
        RECT 1916.430 338.200 1916.750 338.260 ;
        RECT 1918.270 338.200 1918.590 338.260 ;
        RECT 1916.430 338.060 1918.590 338.200 ;
        RECT 1916.430 338.000 1916.750 338.060 ;
        RECT 1918.270 338.000 1918.590 338.060 ;
        RECT 1916.430 304.200 1916.750 304.260 ;
        RECT 1916.060 304.060 1916.750 304.200 ;
        RECT 1916.060 303.580 1916.200 304.060 ;
        RECT 1916.430 304.000 1916.750 304.060 ;
        RECT 1915.970 303.320 1916.290 303.580 ;
        RECT 1915.050 289.580 1915.370 289.640 ;
        RECT 1915.970 289.580 1916.290 289.640 ;
        RECT 1915.050 289.440 1916.290 289.580 ;
        RECT 1915.050 289.380 1915.370 289.440 ;
        RECT 1915.970 289.380 1916.290 289.440 ;
        RECT 1915.050 241.640 1915.370 241.700 ;
        RECT 1916.430 241.640 1916.750 241.700 ;
        RECT 1915.050 241.500 1916.750 241.640 ;
        RECT 1915.050 241.440 1915.370 241.500 ;
        RECT 1916.430 241.440 1916.750 241.500 ;
        RECT 1915.050 193.020 1915.370 193.080 ;
        RECT 1915.970 193.020 1916.290 193.080 ;
        RECT 1915.050 192.880 1916.290 193.020 ;
        RECT 1915.050 192.820 1915.370 192.880 ;
        RECT 1915.970 192.820 1916.290 192.880 ;
        RECT 1915.050 145.080 1915.370 145.140 ;
        RECT 1916.430 145.080 1916.750 145.140 ;
        RECT 1915.050 144.940 1916.750 145.080 ;
        RECT 1915.050 144.880 1915.370 144.940 ;
        RECT 1916.430 144.880 1916.750 144.940 ;
        RECT 1915.050 144.400 1915.370 144.460 ;
        RECT 1916.430 144.400 1916.750 144.460 ;
        RECT 1915.050 144.260 1916.750 144.400 ;
        RECT 1915.050 144.200 1915.370 144.260 ;
        RECT 1916.430 144.200 1916.750 144.260 ;
        RECT 1915.050 96.800 1915.370 96.860 ;
        RECT 1916.890 96.800 1917.210 96.860 ;
        RECT 1915.050 96.660 1917.210 96.800 ;
        RECT 1915.050 96.600 1915.370 96.660 ;
        RECT 1916.890 96.600 1917.210 96.660 ;
        RECT 1916.890 62.460 1917.210 62.520 ;
        RECT 1916.520 62.320 1917.210 62.460 ;
        RECT 1916.520 62.180 1916.660 62.320 ;
        RECT 1916.890 62.260 1917.210 62.320 ;
        RECT 1916.430 61.920 1916.750 62.180 ;
        RECT 1916.430 37.640 1916.750 37.700 ;
        RECT 1916.430 37.500 2387.240 37.640 ;
        RECT 1916.430 37.440 1916.750 37.500 ;
        RECT 2387.100 37.300 2387.240 37.500 ;
        RECT 2417.370 37.300 2417.690 37.360 ;
        RECT 2387.100 37.160 2417.690 37.300 ;
        RECT 2417.370 37.100 2417.690 37.160 ;
      LAYER via ;
        RECT 1914.620 579.740 1914.880 580.000 ;
        RECT 1915.540 579.740 1915.800 580.000 ;
        RECT 1916.460 497.120 1916.720 497.380 ;
        RECT 1916.000 496.440 1916.260 496.700 ;
        RECT 1914.620 482.840 1914.880 483.100 ;
        RECT 1916.000 482.840 1916.260 483.100 ;
        RECT 1914.620 434.900 1914.880 435.160 ;
        RECT 1915.540 434.900 1915.800 435.160 ;
        RECT 1916.460 338.000 1916.720 338.260 ;
        RECT 1918.300 338.000 1918.560 338.260 ;
        RECT 1916.460 304.000 1916.720 304.260 ;
        RECT 1916.000 303.320 1916.260 303.580 ;
        RECT 1915.080 289.380 1915.340 289.640 ;
        RECT 1916.000 289.380 1916.260 289.640 ;
        RECT 1915.080 241.440 1915.340 241.700 ;
        RECT 1916.460 241.440 1916.720 241.700 ;
        RECT 1915.080 192.820 1915.340 193.080 ;
        RECT 1916.000 192.820 1916.260 193.080 ;
        RECT 1915.080 144.880 1915.340 145.140 ;
        RECT 1916.460 144.880 1916.720 145.140 ;
        RECT 1915.080 144.200 1915.340 144.460 ;
        RECT 1916.460 144.200 1916.720 144.460 ;
        RECT 1915.080 96.600 1915.340 96.860 ;
        RECT 1916.920 96.600 1917.180 96.860 ;
        RECT 1916.920 62.260 1917.180 62.520 ;
        RECT 1916.460 61.920 1916.720 62.180 ;
        RECT 1916.460 37.440 1916.720 37.700 ;
        RECT 2417.400 37.100 2417.660 37.360 ;
      LAYER met2 ;
        RECT 1913.930 600.170 1914.210 604.000 ;
        RECT 1913.930 600.030 1914.820 600.170 ;
        RECT 1913.930 600.000 1914.210 600.030 ;
        RECT 1914.680 580.030 1914.820 600.030 ;
        RECT 1914.620 579.710 1914.880 580.030 ;
        RECT 1915.540 579.710 1915.800 580.030 ;
        RECT 1915.600 545.090 1915.740 579.710 ;
        RECT 1915.600 544.950 1916.660 545.090 ;
        RECT 1916.520 497.410 1916.660 544.950 ;
        RECT 1916.460 497.090 1916.720 497.410 ;
        RECT 1916.000 496.410 1916.260 496.730 ;
        RECT 1916.060 483.130 1916.200 496.410 ;
        RECT 1914.620 482.810 1914.880 483.130 ;
        RECT 1916.000 482.810 1916.260 483.130 ;
        RECT 1914.680 435.190 1914.820 482.810 ;
        RECT 1914.620 434.870 1914.880 435.190 ;
        RECT 1915.540 434.870 1915.800 435.190 ;
        RECT 1915.600 399.570 1915.740 434.870 ;
        RECT 1915.600 399.430 1916.200 399.570 ;
        RECT 1916.060 386.085 1916.200 399.430 ;
        RECT 1915.990 385.715 1916.270 386.085 ;
        RECT 1918.290 385.715 1918.570 386.085 ;
        RECT 1918.360 338.290 1918.500 385.715 ;
        RECT 1916.460 337.970 1916.720 338.290 ;
        RECT 1918.300 337.970 1918.560 338.290 ;
        RECT 1916.520 304.290 1916.660 337.970 ;
        RECT 1916.460 303.970 1916.720 304.290 ;
        RECT 1916.000 303.290 1916.260 303.610 ;
        RECT 1916.060 289.670 1916.200 303.290 ;
        RECT 1915.080 289.350 1915.340 289.670 ;
        RECT 1916.000 289.350 1916.260 289.670 ;
        RECT 1915.140 241.730 1915.280 289.350 ;
        RECT 1915.080 241.410 1915.340 241.730 ;
        RECT 1916.460 241.410 1916.720 241.730 ;
        RECT 1916.520 217.330 1916.660 241.410 ;
        RECT 1916.060 217.190 1916.660 217.330 ;
        RECT 1916.060 193.110 1916.200 217.190 ;
        RECT 1915.080 192.790 1915.340 193.110 ;
        RECT 1916.000 192.790 1916.260 193.110 ;
        RECT 1915.140 145.170 1915.280 192.790 ;
        RECT 1915.080 144.850 1915.340 145.170 ;
        RECT 1916.460 144.850 1916.720 145.170 ;
        RECT 1916.520 144.490 1916.660 144.850 ;
        RECT 1915.080 144.170 1915.340 144.490 ;
        RECT 1916.460 144.170 1916.720 144.490 ;
        RECT 1915.140 96.890 1915.280 144.170 ;
        RECT 1915.080 96.570 1915.340 96.890 ;
        RECT 1916.920 96.570 1917.180 96.890 ;
        RECT 1916.980 62.550 1917.120 96.570 ;
        RECT 1916.920 62.230 1917.180 62.550 ;
        RECT 1916.460 61.890 1916.720 62.210 ;
        RECT 1916.520 37.730 1916.660 61.890 ;
        RECT 1916.460 37.410 1916.720 37.730 ;
        RECT 2417.400 37.070 2417.660 37.390 ;
        RECT 2417.460 2.400 2417.600 37.070 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
      LAYER via2 ;
        RECT 1915.990 385.760 1916.270 386.040 ;
        RECT 1918.290 385.760 1918.570 386.040 ;
      LAYER met3 ;
        RECT 1915.965 386.050 1916.295 386.065 ;
        RECT 1918.265 386.050 1918.595 386.065 ;
        RECT 1915.965 385.750 1918.595 386.050 ;
        RECT 1915.965 385.735 1916.295 385.750 ;
        RECT 1918.265 385.735 1918.595 385.750 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1924.710 41.380 1925.030 41.440 ;
        RECT 2434.850 41.380 2435.170 41.440 ;
        RECT 1924.710 41.240 2435.170 41.380 ;
        RECT 1924.710 41.180 1925.030 41.240 ;
        RECT 2434.850 41.180 2435.170 41.240 ;
      LAYER via ;
        RECT 1924.740 41.180 1925.000 41.440 ;
        RECT 2434.880 41.180 2435.140 41.440 ;
      LAYER met2 ;
        RECT 1923.130 600.170 1923.410 604.000 ;
        RECT 1923.130 600.030 1924.940 600.170 ;
        RECT 1923.130 600.000 1923.410 600.030 ;
        RECT 1924.800 41.470 1924.940 600.030 ;
        RECT 1924.740 41.150 1925.000 41.470 ;
        RECT 2434.880 41.150 2435.140 41.470 ;
        RECT 2434.940 2.400 2435.080 41.150 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1933.910 586.740 1934.230 586.800 ;
        RECT 1938.050 586.740 1938.370 586.800 ;
        RECT 1933.910 586.600 1938.370 586.740 ;
        RECT 1933.910 586.540 1934.230 586.600 ;
        RECT 1938.050 586.540 1938.370 586.600 ;
        RECT 1938.050 41.040 1938.370 41.100 ;
        RECT 2452.790 41.040 2453.110 41.100 ;
        RECT 1938.050 40.900 2453.110 41.040 ;
        RECT 1938.050 40.840 1938.370 40.900 ;
        RECT 2452.790 40.840 2453.110 40.900 ;
      LAYER via ;
        RECT 1933.940 586.540 1934.200 586.800 ;
        RECT 1938.080 586.540 1938.340 586.800 ;
        RECT 1938.080 40.840 1938.340 41.100 ;
        RECT 2452.820 40.840 2453.080 41.100 ;
      LAYER met2 ;
        RECT 1932.330 600.170 1932.610 604.000 ;
        RECT 1932.330 600.030 1934.140 600.170 ;
        RECT 1932.330 600.000 1932.610 600.030 ;
        RECT 1934.000 586.830 1934.140 600.030 ;
        RECT 1933.940 586.510 1934.200 586.830 ;
        RECT 1938.080 586.510 1938.340 586.830 ;
        RECT 1938.140 41.130 1938.280 586.510 ;
        RECT 1938.080 40.810 1938.340 41.130 ;
        RECT 2452.820 40.810 2453.080 41.130 ;
        RECT 2452.880 2.400 2453.020 40.810 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1943.570 579.600 1943.890 579.660 ;
        RECT 1944.490 579.600 1944.810 579.660 ;
        RECT 1943.570 579.460 1944.810 579.600 ;
        RECT 1943.570 579.400 1943.890 579.460 ;
        RECT 1944.490 579.400 1944.810 579.460 ;
        RECT 1943.570 531.320 1943.890 531.380 ;
        RECT 1944.030 531.320 1944.350 531.380 ;
        RECT 1943.570 531.180 1944.350 531.320 ;
        RECT 1943.570 531.120 1943.890 531.180 ;
        RECT 1944.030 531.120 1944.350 531.180 ;
        RECT 1943.570 483.040 1943.890 483.100 ;
        RECT 1944.490 483.040 1944.810 483.100 ;
        RECT 1943.570 482.900 1944.810 483.040 ;
        RECT 1943.570 482.840 1943.890 482.900 ;
        RECT 1944.490 482.840 1944.810 482.900 ;
        RECT 1943.570 434.760 1943.890 434.820 ;
        RECT 1944.030 434.760 1944.350 434.820 ;
        RECT 1943.570 434.620 1944.350 434.760 ;
        RECT 1943.570 434.560 1943.890 434.620 ;
        RECT 1944.030 434.560 1944.350 434.620 ;
        RECT 1944.030 338.200 1944.350 338.260 ;
        RECT 1945.870 338.200 1946.190 338.260 ;
        RECT 1944.030 338.060 1946.190 338.200 ;
        RECT 1944.030 338.000 1944.350 338.060 ;
        RECT 1945.870 338.000 1946.190 338.060 ;
        RECT 1944.030 304.200 1944.350 304.260 ;
        RECT 1943.660 304.060 1944.350 304.200 ;
        RECT 1943.660 303.580 1943.800 304.060 ;
        RECT 1944.030 304.000 1944.350 304.060 ;
        RECT 1943.570 303.320 1943.890 303.580 ;
        RECT 1942.650 289.580 1942.970 289.640 ;
        RECT 1943.570 289.580 1943.890 289.640 ;
        RECT 1942.650 289.440 1943.890 289.580 ;
        RECT 1942.650 289.380 1942.970 289.440 ;
        RECT 1943.570 289.380 1943.890 289.440 ;
        RECT 1942.650 241.640 1942.970 241.700 ;
        RECT 1944.030 241.640 1944.350 241.700 ;
        RECT 1942.650 241.500 1944.350 241.640 ;
        RECT 1942.650 241.440 1942.970 241.500 ;
        RECT 1944.030 241.440 1944.350 241.500 ;
        RECT 1943.570 158.680 1943.890 158.740 ;
        RECT 1944.490 158.680 1944.810 158.740 ;
        RECT 1943.570 158.540 1944.810 158.680 ;
        RECT 1943.570 158.480 1943.890 158.540 ;
        RECT 1944.490 158.480 1944.810 158.540 ;
        RECT 1943.570 120.940 1943.890 121.000 ;
        RECT 1944.490 120.940 1944.810 121.000 ;
        RECT 1943.570 120.800 1944.810 120.940 ;
        RECT 1943.570 120.740 1943.890 120.800 ;
        RECT 1944.490 120.740 1944.810 120.800 ;
        RECT 1944.490 40.700 1944.810 40.760 ;
        RECT 2470.730 40.700 2471.050 40.760 ;
        RECT 1944.490 40.560 2471.050 40.700 ;
        RECT 1944.490 40.500 1944.810 40.560 ;
        RECT 2470.730 40.500 2471.050 40.560 ;
      LAYER via ;
        RECT 1943.600 579.400 1943.860 579.660 ;
        RECT 1944.520 579.400 1944.780 579.660 ;
        RECT 1943.600 531.120 1943.860 531.380 ;
        RECT 1944.060 531.120 1944.320 531.380 ;
        RECT 1943.600 482.840 1943.860 483.100 ;
        RECT 1944.520 482.840 1944.780 483.100 ;
        RECT 1943.600 434.560 1943.860 434.820 ;
        RECT 1944.060 434.560 1944.320 434.820 ;
        RECT 1944.060 338.000 1944.320 338.260 ;
        RECT 1945.900 338.000 1946.160 338.260 ;
        RECT 1944.060 304.000 1944.320 304.260 ;
        RECT 1943.600 303.320 1943.860 303.580 ;
        RECT 1942.680 289.380 1942.940 289.640 ;
        RECT 1943.600 289.380 1943.860 289.640 ;
        RECT 1942.680 241.440 1942.940 241.700 ;
        RECT 1944.060 241.440 1944.320 241.700 ;
        RECT 1943.600 158.480 1943.860 158.740 ;
        RECT 1944.520 158.480 1944.780 158.740 ;
        RECT 1943.600 120.740 1943.860 121.000 ;
        RECT 1944.520 120.740 1944.780 121.000 ;
        RECT 1944.520 40.500 1944.780 40.760 ;
        RECT 2470.760 40.500 2471.020 40.760 ;
      LAYER met2 ;
        RECT 1941.530 600.850 1941.810 604.000 ;
        RECT 1941.530 600.710 1942.420 600.850 ;
        RECT 1941.530 600.000 1941.810 600.710 ;
        RECT 1942.280 580.565 1942.420 600.710 ;
        RECT 1942.210 580.195 1942.490 580.565 ;
        RECT 1943.590 579.515 1943.870 579.885 ;
        RECT 1943.600 579.370 1943.860 579.515 ;
        RECT 1944.520 579.370 1944.780 579.690 ;
        RECT 1944.580 531.605 1944.720 579.370 ;
        RECT 1943.590 531.235 1943.870 531.605 ;
        RECT 1943.600 531.090 1943.860 531.235 ;
        RECT 1944.060 531.090 1944.320 531.410 ;
        RECT 1944.510 531.235 1944.790 531.605 ;
        RECT 1944.120 483.210 1944.260 531.090 ;
        RECT 1943.660 483.130 1944.260 483.210 ;
        RECT 1943.600 483.070 1944.260 483.130 ;
        RECT 1943.600 482.810 1943.860 483.070 ;
        RECT 1944.520 482.810 1944.780 483.130 ;
        RECT 1943.660 482.655 1943.800 482.810 ;
        RECT 1944.580 447.850 1944.720 482.810 ;
        RECT 1943.660 447.710 1944.720 447.850 ;
        RECT 1943.660 434.850 1943.800 447.710 ;
        RECT 1943.600 434.530 1943.860 434.850 ;
        RECT 1944.060 434.530 1944.320 434.850 ;
        RECT 1944.120 399.570 1944.260 434.530 ;
        RECT 1943.660 399.430 1944.260 399.570 ;
        RECT 1943.660 386.085 1943.800 399.430 ;
        RECT 1943.590 385.715 1943.870 386.085 ;
        RECT 1945.890 385.715 1946.170 386.085 ;
        RECT 1945.960 338.290 1946.100 385.715 ;
        RECT 1944.060 337.970 1944.320 338.290 ;
        RECT 1945.900 337.970 1946.160 338.290 ;
        RECT 1944.120 304.290 1944.260 337.970 ;
        RECT 1944.060 303.970 1944.320 304.290 ;
        RECT 1943.600 303.290 1943.860 303.610 ;
        RECT 1943.660 289.670 1943.800 303.290 ;
        RECT 1942.680 289.350 1942.940 289.670 ;
        RECT 1943.600 289.350 1943.860 289.670 ;
        RECT 1942.740 241.730 1942.880 289.350 ;
        RECT 1942.680 241.410 1942.940 241.730 ;
        RECT 1944.060 241.410 1944.320 241.730 ;
        RECT 1944.120 217.330 1944.260 241.410 ;
        RECT 1943.660 217.190 1944.260 217.330 ;
        RECT 1943.660 158.770 1943.800 217.190 ;
        RECT 1943.600 158.450 1943.860 158.770 ;
        RECT 1944.520 158.450 1944.780 158.770 ;
        RECT 1944.580 121.030 1944.720 158.450 ;
        RECT 1943.600 120.710 1943.860 121.030 ;
        RECT 1944.520 120.710 1944.780 121.030 ;
        RECT 1943.660 62.290 1943.800 120.710 ;
        RECT 1943.660 62.150 1944.720 62.290 ;
        RECT 1944.580 40.790 1944.720 62.150 ;
        RECT 1944.520 40.470 1944.780 40.790 ;
        RECT 2470.760 40.470 2471.020 40.790 ;
        RECT 2470.820 2.400 2470.960 40.470 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
      LAYER via2 ;
        RECT 1942.210 580.240 1942.490 580.520 ;
        RECT 1943.590 579.560 1943.870 579.840 ;
        RECT 1943.590 531.280 1943.870 531.560 ;
        RECT 1944.510 531.280 1944.790 531.560 ;
        RECT 1943.590 385.760 1943.870 386.040 ;
        RECT 1945.890 385.760 1946.170 386.040 ;
      LAYER met3 ;
        RECT 1942.185 580.530 1942.515 580.545 ;
        RECT 1942.185 580.230 1944.570 580.530 ;
        RECT 1942.185 580.215 1942.515 580.230 ;
        RECT 1943.565 579.850 1943.895 579.865 ;
        RECT 1944.270 579.850 1944.570 580.230 ;
        RECT 1943.565 579.550 1944.570 579.850 ;
        RECT 1943.565 579.535 1943.895 579.550 ;
        RECT 1943.565 531.570 1943.895 531.585 ;
        RECT 1944.485 531.570 1944.815 531.585 ;
        RECT 1943.565 531.270 1944.815 531.570 ;
        RECT 1943.565 531.255 1943.895 531.270 ;
        RECT 1944.485 531.255 1944.815 531.270 ;
        RECT 1943.565 386.050 1943.895 386.065 ;
        RECT 1945.865 386.050 1946.195 386.065 ;
        RECT 1943.565 385.750 1946.195 386.050 ;
        RECT 1943.565 385.735 1943.895 385.750 ;
        RECT 1945.865 385.735 1946.195 385.750 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1952.310 40.360 1952.630 40.420 ;
        RECT 2488.670 40.360 2488.990 40.420 ;
        RECT 1952.310 40.220 2488.990 40.360 ;
        RECT 1952.310 40.160 1952.630 40.220 ;
        RECT 2488.670 40.160 2488.990 40.220 ;
      LAYER via ;
        RECT 1952.340 40.160 1952.600 40.420 ;
        RECT 2488.700 40.160 2488.960 40.420 ;
      LAYER met2 ;
        RECT 1950.730 600.170 1951.010 604.000 ;
        RECT 1950.730 600.030 1952.540 600.170 ;
        RECT 1950.730 600.000 1951.010 600.030 ;
        RECT 1952.400 40.450 1952.540 600.030 ;
        RECT 1952.340 40.130 1952.600 40.450 ;
        RECT 2488.700 40.130 2488.960 40.450 ;
        RECT 2488.760 2.400 2488.900 40.130 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1961.510 586.740 1961.830 586.800 ;
        RECT 1965.650 586.740 1965.970 586.800 ;
        RECT 1961.510 586.600 1965.970 586.740 ;
        RECT 1961.510 586.540 1961.830 586.600 ;
        RECT 1965.650 586.540 1965.970 586.600 ;
        RECT 1965.650 40.020 1965.970 40.080 ;
        RECT 2506.150 40.020 2506.470 40.080 ;
        RECT 1965.650 39.880 2506.470 40.020 ;
        RECT 1965.650 39.820 1965.970 39.880 ;
        RECT 2506.150 39.820 2506.470 39.880 ;
      LAYER via ;
        RECT 1961.540 586.540 1961.800 586.800 ;
        RECT 1965.680 586.540 1965.940 586.800 ;
        RECT 1965.680 39.820 1965.940 40.080 ;
        RECT 2506.180 39.820 2506.440 40.080 ;
      LAYER met2 ;
        RECT 1959.930 600.170 1960.210 604.000 ;
        RECT 1959.930 600.030 1961.740 600.170 ;
        RECT 1959.930 600.000 1960.210 600.030 ;
        RECT 1961.600 586.830 1961.740 600.030 ;
        RECT 1961.540 586.510 1961.800 586.830 ;
        RECT 1965.680 586.510 1965.940 586.830 ;
        RECT 1965.740 40.110 1965.880 586.510 ;
        RECT 1965.680 39.790 1965.940 40.110 ;
        RECT 2506.180 39.790 2506.440 40.110 ;
        RECT 2506.240 2.400 2506.380 39.790 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1972.090 531.320 1972.410 531.380 ;
        RECT 1972.550 531.320 1972.870 531.380 ;
        RECT 1972.090 531.180 1972.870 531.320 ;
        RECT 1972.090 531.120 1972.410 531.180 ;
        RECT 1972.550 531.120 1972.870 531.180 ;
        RECT 1972.550 496.980 1972.870 497.040 ;
        RECT 1972.180 496.840 1972.870 496.980 ;
        RECT 1972.180 496.700 1972.320 496.840 ;
        RECT 1972.550 496.780 1972.870 496.840 ;
        RECT 1972.090 496.440 1972.410 496.700 ;
        RECT 1971.630 448.700 1971.950 448.760 ;
        RECT 1972.550 448.700 1972.870 448.760 ;
        RECT 1971.630 448.560 1972.870 448.700 ;
        RECT 1971.630 448.500 1971.950 448.560 ;
        RECT 1972.550 448.500 1972.870 448.560 ;
        RECT 1971.170 434.760 1971.490 434.820 ;
        RECT 1972.090 434.760 1972.410 434.820 ;
        RECT 1971.170 434.620 1972.410 434.760 ;
        RECT 1971.170 434.560 1971.490 434.620 ;
        RECT 1972.090 434.560 1972.410 434.620 ;
        RECT 1971.170 386.480 1971.490 386.540 ;
        RECT 1972.550 386.480 1972.870 386.540 ;
        RECT 1971.170 386.340 1972.870 386.480 ;
        RECT 1971.170 386.280 1971.490 386.340 ;
        RECT 1972.550 386.280 1972.870 386.340 ;
        RECT 1972.090 338.200 1972.410 338.260 ;
        RECT 1972.550 338.200 1972.870 338.260 ;
        RECT 1972.090 338.060 1972.870 338.200 ;
        RECT 1972.090 338.000 1972.410 338.060 ;
        RECT 1972.550 338.000 1972.870 338.060 ;
        RECT 1972.090 241.640 1972.410 241.700 ;
        RECT 1972.550 241.640 1972.870 241.700 ;
        RECT 1972.090 241.500 1972.870 241.640 ;
        RECT 1972.090 241.440 1972.410 241.500 ;
        RECT 1972.550 241.440 1972.870 241.500 ;
        RECT 1972.090 145.080 1972.410 145.140 ;
        RECT 1972.550 145.080 1972.870 145.140 ;
        RECT 1972.090 144.940 1972.870 145.080 ;
        RECT 1972.090 144.880 1972.410 144.940 ;
        RECT 1972.550 144.880 1972.870 144.940 ;
        RECT 1971.630 62.260 1971.950 62.520 ;
        RECT 1971.720 61.780 1971.860 62.260 ;
        RECT 1972.090 61.780 1972.410 61.840 ;
        RECT 1971.720 61.640 1972.410 61.780 ;
        RECT 1972.090 61.580 1972.410 61.640 ;
        RECT 1971.630 39.680 1971.950 39.740 ;
        RECT 2524.090 39.680 2524.410 39.740 ;
        RECT 1971.630 39.540 2524.410 39.680 ;
        RECT 1971.630 39.480 1971.950 39.540 ;
        RECT 2524.090 39.480 2524.410 39.540 ;
      LAYER via ;
        RECT 1972.120 531.120 1972.380 531.380 ;
        RECT 1972.580 531.120 1972.840 531.380 ;
        RECT 1972.580 496.780 1972.840 497.040 ;
        RECT 1972.120 496.440 1972.380 496.700 ;
        RECT 1971.660 448.500 1971.920 448.760 ;
        RECT 1972.580 448.500 1972.840 448.760 ;
        RECT 1971.200 434.560 1971.460 434.820 ;
        RECT 1972.120 434.560 1972.380 434.820 ;
        RECT 1971.200 386.280 1971.460 386.540 ;
        RECT 1972.580 386.280 1972.840 386.540 ;
        RECT 1972.120 338.000 1972.380 338.260 ;
        RECT 1972.580 338.000 1972.840 338.260 ;
        RECT 1972.120 241.440 1972.380 241.700 ;
        RECT 1972.580 241.440 1972.840 241.700 ;
        RECT 1972.120 144.880 1972.380 145.140 ;
        RECT 1972.580 144.880 1972.840 145.140 ;
        RECT 1971.660 62.260 1971.920 62.520 ;
        RECT 1972.120 61.580 1972.380 61.840 ;
        RECT 1971.660 39.480 1971.920 39.740 ;
        RECT 2524.120 39.480 2524.380 39.740 ;
      LAYER met2 ;
        RECT 1969.130 601.530 1969.410 604.000 ;
        RECT 1969.130 601.390 1970.940 601.530 ;
        RECT 1969.130 600.000 1969.410 601.390 ;
        RECT 1970.800 545.090 1970.940 601.390 ;
        RECT 1970.800 544.950 1971.860 545.090 ;
        RECT 1971.720 544.410 1971.860 544.950 ;
        RECT 1971.720 544.270 1972.320 544.410 ;
        RECT 1972.180 531.410 1972.320 544.270 ;
        RECT 1972.120 531.090 1972.380 531.410 ;
        RECT 1972.580 531.090 1972.840 531.410 ;
        RECT 1972.640 497.070 1972.780 531.090 ;
        RECT 1972.580 496.750 1972.840 497.070 ;
        RECT 1972.120 496.410 1972.380 496.730 ;
        RECT 1972.180 483.210 1972.320 496.410 ;
        RECT 1972.180 483.070 1972.780 483.210 ;
        RECT 1972.640 448.790 1972.780 483.070 ;
        RECT 1971.660 448.530 1971.920 448.790 ;
        RECT 1971.660 448.470 1972.320 448.530 ;
        RECT 1972.580 448.470 1972.840 448.790 ;
        RECT 1971.720 448.390 1972.320 448.470 ;
        RECT 1972.180 434.850 1972.320 448.390 ;
        RECT 1971.200 434.530 1971.460 434.850 ;
        RECT 1972.120 434.530 1972.380 434.850 ;
        RECT 1971.260 386.570 1971.400 434.530 ;
        RECT 1971.200 386.250 1971.460 386.570 ;
        RECT 1972.580 386.250 1972.840 386.570 ;
        RECT 1972.640 338.290 1972.780 386.250 ;
        RECT 1972.120 337.970 1972.380 338.290 ;
        RECT 1972.580 337.970 1972.840 338.290 ;
        RECT 1972.180 303.690 1972.320 337.970 ;
        RECT 1972.180 303.550 1972.780 303.690 ;
        RECT 1972.640 241.730 1972.780 303.550 ;
        RECT 1972.120 241.410 1972.380 241.730 ;
        RECT 1972.580 241.410 1972.840 241.730 ;
        RECT 1972.180 207.130 1972.320 241.410 ;
        RECT 1972.180 206.990 1972.780 207.130 ;
        RECT 1972.640 145.170 1972.780 206.990 ;
        RECT 1972.120 144.850 1972.380 145.170 ;
        RECT 1972.580 144.850 1972.840 145.170 ;
        RECT 1972.180 96.970 1972.320 144.850 ;
        RECT 1971.720 96.830 1972.320 96.970 ;
        RECT 1971.720 62.550 1971.860 96.830 ;
        RECT 1971.660 62.230 1971.920 62.550 ;
        RECT 1972.120 61.550 1972.380 61.870 ;
        RECT 1972.180 48.010 1972.320 61.550 ;
        RECT 1971.720 47.870 1972.320 48.010 ;
        RECT 1971.720 39.770 1971.860 47.870 ;
        RECT 1971.660 39.450 1971.920 39.770 ;
        RECT 2524.120 39.450 2524.380 39.770 ;
        RECT 2524.180 2.400 2524.320 39.450 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1979.450 39.340 1979.770 39.400 ;
        RECT 2542.030 39.340 2542.350 39.400 ;
        RECT 1979.450 39.200 2542.350 39.340 ;
        RECT 1979.450 39.140 1979.770 39.200 ;
        RECT 2542.030 39.140 2542.350 39.200 ;
      LAYER via ;
        RECT 1979.480 39.140 1979.740 39.400 ;
        RECT 2542.060 39.140 2542.320 39.400 ;
      LAYER met2 ;
        RECT 1978.330 600.170 1978.610 604.000 ;
        RECT 1978.330 600.030 1979.680 600.170 ;
        RECT 1978.330 600.000 1978.610 600.030 ;
        RECT 1979.540 39.430 1979.680 600.030 ;
        RECT 1979.480 39.110 1979.740 39.430 ;
        RECT 2542.060 39.110 2542.320 39.430 ;
        RECT 2542.120 2.400 2542.260 39.110 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1989.110 586.740 1989.430 586.800 ;
        RECT 1993.710 586.740 1994.030 586.800 ;
        RECT 1989.110 586.600 1994.030 586.740 ;
        RECT 1989.110 586.540 1989.430 586.600 ;
        RECT 1993.710 586.540 1994.030 586.600 ;
        RECT 1993.710 20.980 1994.030 21.040 ;
        RECT 2559.970 20.980 2560.290 21.040 ;
        RECT 1993.710 20.840 2560.290 20.980 ;
        RECT 1993.710 20.780 1994.030 20.840 ;
        RECT 2559.970 20.780 2560.290 20.840 ;
      LAYER via ;
        RECT 1989.140 586.540 1989.400 586.800 ;
        RECT 1993.740 586.540 1994.000 586.800 ;
        RECT 1993.740 20.780 1994.000 21.040 ;
        RECT 2560.000 20.780 2560.260 21.040 ;
      LAYER met2 ;
        RECT 1987.530 600.170 1987.810 604.000 ;
        RECT 1987.530 600.030 1989.340 600.170 ;
        RECT 1987.530 600.000 1987.810 600.030 ;
        RECT 1989.200 586.830 1989.340 600.030 ;
        RECT 1989.140 586.510 1989.400 586.830 ;
        RECT 1993.740 586.510 1994.000 586.830 ;
        RECT 1993.800 21.070 1993.940 586.510 ;
        RECT 1993.740 20.750 1994.000 21.070 ;
        RECT 2560.000 20.750 2560.260 21.070 ;
        RECT 2560.060 2.400 2560.200 20.750 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1998.310 587.420 1998.630 587.480 ;
        RECT 2000.150 587.420 2000.470 587.480 ;
        RECT 1998.310 587.280 2000.470 587.420 ;
        RECT 1998.310 587.220 1998.630 587.280 ;
        RECT 2000.150 587.220 2000.470 587.280 ;
        RECT 2000.150 21.320 2000.470 21.380 ;
        RECT 2577.910 21.320 2578.230 21.380 ;
        RECT 2000.150 21.180 2578.230 21.320 ;
        RECT 2000.150 21.120 2000.470 21.180 ;
        RECT 2577.910 21.120 2578.230 21.180 ;
      LAYER via ;
        RECT 1998.340 587.220 1998.600 587.480 ;
        RECT 2000.180 587.220 2000.440 587.480 ;
        RECT 2000.180 21.120 2000.440 21.380 ;
        RECT 2577.940 21.120 2578.200 21.380 ;
      LAYER met2 ;
        RECT 1996.730 600.170 1997.010 604.000 ;
        RECT 1996.730 600.030 1998.540 600.170 ;
        RECT 1996.730 600.000 1997.010 600.030 ;
        RECT 1998.400 587.510 1998.540 600.030 ;
        RECT 1998.340 587.190 1998.600 587.510 ;
        RECT 2000.180 587.190 2000.440 587.510 ;
        RECT 2000.240 21.410 2000.380 587.190 ;
        RECT 2000.180 21.090 2000.440 21.410 ;
        RECT 2577.940 21.090 2578.200 21.410 ;
        RECT 2578.000 2.400 2578.140 21.090 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1084.750 476.380 1085.070 476.640 ;
        RECT 1084.290 476.240 1084.610 476.300 ;
        RECT 1084.840 476.240 1084.980 476.380 ;
        RECT 1084.290 476.100 1084.980 476.240 ;
        RECT 1084.290 476.040 1084.610 476.100 ;
        RECT 1084.290 448.500 1084.610 448.760 ;
        RECT 1083.830 448.360 1084.150 448.420 ;
        RECT 1084.380 448.360 1084.520 448.500 ;
        RECT 1083.830 448.220 1084.520 448.360 ;
        RECT 1083.830 448.160 1084.150 448.220 ;
        RECT 1083.830 427.960 1084.150 428.020 ;
        RECT 1084.290 427.960 1084.610 428.020 ;
        RECT 1083.830 427.820 1084.610 427.960 ;
        RECT 1083.830 427.760 1084.150 427.820 ;
        RECT 1084.290 427.760 1084.610 427.820 ;
        RECT 1084.290 379.680 1084.610 379.740 ;
        RECT 1085.210 379.680 1085.530 379.740 ;
        RECT 1084.290 379.540 1085.530 379.680 ;
        RECT 1084.290 379.480 1084.610 379.540 ;
        RECT 1085.210 379.480 1085.530 379.540 ;
        RECT 1084.290 337.860 1084.610 337.920 ;
        RECT 1085.210 337.860 1085.530 337.920 ;
        RECT 1084.290 337.720 1085.530 337.860 ;
        RECT 1084.290 337.660 1084.610 337.720 ;
        RECT 1085.210 337.660 1085.530 337.720 ;
        RECT 811.510 17.920 811.830 17.980 ;
        RECT 966.070 17.920 966.390 17.980 ;
        RECT 811.510 17.780 966.390 17.920 ;
        RECT 811.510 17.720 811.830 17.780 ;
        RECT 966.070 17.720 966.390 17.780 ;
        RECT 1013.910 17.580 1014.230 17.640 ;
        RECT 1027.710 17.580 1028.030 17.640 ;
        RECT 1013.910 17.440 1028.030 17.580 ;
        RECT 1013.910 17.380 1014.230 17.440 ;
        RECT 1027.710 17.380 1028.030 17.440 ;
        RECT 1028.170 17.580 1028.490 17.640 ;
        RECT 1084.290 17.580 1084.610 17.640 ;
        RECT 1028.170 17.440 1084.610 17.580 ;
        RECT 1028.170 17.380 1028.490 17.440 ;
        RECT 1084.290 17.380 1084.610 17.440 ;
      LAYER via ;
        RECT 1084.780 476.380 1085.040 476.640 ;
        RECT 1084.320 476.040 1084.580 476.300 ;
        RECT 1084.320 448.500 1084.580 448.760 ;
        RECT 1083.860 448.160 1084.120 448.420 ;
        RECT 1083.860 427.760 1084.120 428.020 ;
        RECT 1084.320 427.760 1084.580 428.020 ;
        RECT 1084.320 379.480 1084.580 379.740 ;
        RECT 1085.240 379.480 1085.500 379.740 ;
        RECT 1084.320 337.660 1084.580 337.920 ;
        RECT 1085.240 337.660 1085.500 337.920 ;
        RECT 811.540 17.720 811.800 17.980 ;
        RECT 966.100 17.720 966.360 17.980 ;
        RECT 1013.940 17.380 1014.200 17.640 ;
        RECT 1027.740 17.380 1028.000 17.640 ;
        RECT 1028.200 17.380 1028.460 17.640 ;
        RECT 1084.320 17.380 1084.580 17.640 ;
      LAYER met2 ;
        RECT 1087.770 600.170 1088.050 604.000 ;
        RECT 1086.680 600.030 1088.050 600.170 ;
        RECT 1086.680 579.885 1086.820 600.030 ;
        RECT 1087.770 600.000 1088.050 600.030 ;
        RECT 1084.770 579.515 1085.050 579.885 ;
        RECT 1086.610 579.515 1086.890 579.885 ;
        RECT 1084.840 476.670 1084.980 579.515 ;
        RECT 1084.780 476.350 1085.040 476.670 ;
        RECT 1084.320 476.010 1084.580 476.330 ;
        RECT 1084.380 448.790 1084.520 476.010 ;
        RECT 1084.320 448.470 1084.580 448.790 ;
        RECT 1083.860 448.130 1084.120 448.450 ;
        RECT 1083.920 428.050 1084.060 448.130 ;
        RECT 1083.860 427.730 1084.120 428.050 ;
        RECT 1084.320 427.730 1084.580 428.050 ;
        RECT 1084.380 427.450 1084.520 427.730 ;
        RECT 1084.380 427.310 1085.440 427.450 ;
        RECT 1085.300 379.770 1085.440 427.310 ;
        RECT 1084.320 379.450 1084.580 379.770 ;
        RECT 1085.240 379.450 1085.500 379.770 ;
        RECT 1084.380 337.950 1084.520 379.450 ;
        RECT 1084.320 337.630 1084.580 337.950 ;
        RECT 1085.240 337.630 1085.500 337.950 ;
        RECT 1085.300 313.210 1085.440 337.630 ;
        RECT 1084.380 313.070 1085.440 313.210 ;
        RECT 1084.380 207.130 1084.520 313.070 ;
        RECT 1083.920 206.990 1084.520 207.130 ;
        RECT 1083.920 206.450 1084.060 206.990 ;
        RECT 1083.920 206.310 1084.520 206.450 ;
        RECT 1084.380 110.570 1084.520 206.310 ;
        RECT 1083.920 110.430 1084.520 110.570 ;
        RECT 1083.920 109.890 1084.060 110.430 ;
        RECT 1083.920 109.750 1084.520 109.890 ;
        RECT 811.540 17.690 811.800 18.010 ;
        RECT 966.090 17.835 966.370 18.205 ;
        RECT 1013.930 17.835 1014.210 18.205 ;
        RECT 966.100 17.690 966.360 17.835 ;
        RECT 811.600 2.400 811.740 17.690 ;
        RECT 1014.000 17.670 1014.140 17.835 ;
        RECT 1084.380 17.670 1084.520 109.750 ;
        RECT 1013.940 17.350 1014.200 17.670 ;
        RECT 1027.740 17.580 1028.000 17.670 ;
        RECT 1028.200 17.580 1028.460 17.670 ;
        RECT 1027.740 17.440 1028.460 17.580 ;
        RECT 1027.740 17.350 1028.000 17.440 ;
        RECT 1028.200 17.350 1028.460 17.440 ;
        RECT 1084.320 17.350 1084.580 17.670 ;
        RECT 811.390 -4.800 811.950 2.400 ;
      LAYER via2 ;
        RECT 1084.770 579.560 1085.050 579.840 ;
        RECT 1086.610 579.560 1086.890 579.840 ;
        RECT 966.090 17.880 966.370 18.160 ;
        RECT 1013.930 17.880 1014.210 18.160 ;
      LAYER met3 ;
        RECT 1084.745 579.850 1085.075 579.865 ;
        RECT 1086.585 579.850 1086.915 579.865 ;
        RECT 1084.745 579.550 1086.915 579.850 ;
        RECT 1084.745 579.535 1085.075 579.550 ;
        RECT 1086.585 579.535 1086.915 579.550 ;
        RECT 966.065 18.170 966.395 18.185 ;
        RECT 1013.905 18.170 1014.235 18.185 ;
        RECT 966.065 17.870 1014.235 18.170 ;
        RECT 966.065 17.855 966.395 17.870 ;
        RECT 1013.905 17.855 1014.235 17.870 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.510 22.000 2007.830 22.060 ;
        RECT 2595.390 22.000 2595.710 22.060 ;
        RECT 2007.510 21.860 2595.710 22.000 ;
        RECT 2007.510 21.800 2007.830 21.860 ;
        RECT 2595.390 21.800 2595.710 21.860 ;
      LAYER via ;
        RECT 2007.540 21.800 2007.800 22.060 ;
        RECT 2595.420 21.800 2595.680 22.060 ;
      LAYER met2 ;
        RECT 2005.930 600.170 2006.210 604.000 ;
        RECT 2005.930 600.030 2007.740 600.170 ;
        RECT 2005.930 600.000 2006.210 600.030 ;
        RECT 2007.600 22.090 2007.740 600.030 ;
        RECT 2007.540 21.770 2007.800 22.090 ;
        RECT 2595.420 21.770 2595.680 22.090 ;
        RECT 2595.480 2.400 2595.620 21.770 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2016.710 586.740 2017.030 586.800 ;
        RECT 2021.310 586.740 2021.630 586.800 ;
        RECT 2016.710 586.600 2021.630 586.740 ;
        RECT 2016.710 586.540 2017.030 586.600 ;
        RECT 2021.310 586.540 2021.630 586.600 ;
        RECT 2021.310 21.660 2021.630 21.720 ;
        RECT 2613.330 21.660 2613.650 21.720 ;
        RECT 2021.310 21.520 2613.650 21.660 ;
        RECT 2021.310 21.460 2021.630 21.520 ;
        RECT 2613.330 21.460 2613.650 21.520 ;
      LAYER via ;
        RECT 2016.740 586.540 2017.000 586.800 ;
        RECT 2021.340 586.540 2021.600 586.800 ;
        RECT 2021.340 21.460 2021.600 21.720 ;
        RECT 2613.360 21.460 2613.620 21.720 ;
      LAYER met2 ;
        RECT 2015.130 600.170 2015.410 604.000 ;
        RECT 2015.130 600.030 2016.940 600.170 ;
        RECT 2015.130 600.000 2015.410 600.030 ;
        RECT 2016.800 586.830 2016.940 600.030 ;
        RECT 2016.740 586.510 2017.000 586.830 ;
        RECT 2021.340 586.510 2021.600 586.830 ;
        RECT 2021.400 21.750 2021.540 586.510 ;
        RECT 2021.340 21.430 2021.600 21.750 ;
        RECT 2613.360 21.430 2613.620 21.750 ;
        RECT 2613.420 2.400 2613.560 21.430 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2025.910 587.080 2026.230 587.140 ;
        RECT 2028.210 587.080 2028.530 587.140 ;
        RECT 2025.910 586.940 2028.530 587.080 ;
        RECT 2025.910 586.880 2026.230 586.940 ;
        RECT 2028.210 586.880 2028.530 586.940 ;
        RECT 2028.210 22.340 2028.530 22.400 ;
        RECT 2631.270 22.340 2631.590 22.400 ;
        RECT 2028.210 22.200 2631.590 22.340 ;
        RECT 2028.210 22.140 2028.530 22.200 ;
        RECT 2631.270 22.140 2631.590 22.200 ;
      LAYER via ;
        RECT 2025.940 586.880 2026.200 587.140 ;
        RECT 2028.240 586.880 2028.500 587.140 ;
        RECT 2028.240 22.140 2028.500 22.400 ;
        RECT 2631.300 22.140 2631.560 22.400 ;
      LAYER met2 ;
        RECT 2024.330 600.170 2024.610 604.000 ;
        RECT 2024.330 600.030 2026.140 600.170 ;
        RECT 2024.330 600.000 2024.610 600.030 ;
        RECT 2026.000 587.170 2026.140 600.030 ;
        RECT 2025.940 586.850 2026.200 587.170 ;
        RECT 2028.240 586.850 2028.500 587.170 ;
        RECT 2028.300 22.430 2028.440 586.850 ;
        RECT 2028.240 22.110 2028.500 22.430 ;
        RECT 2631.300 22.110 2631.560 22.430 ;
        RECT 2631.360 2.400 2631.500 22.110 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2034.650 22.680 2034.970 22.740 ;
        RECT 2649.210 22.680 2649.530 22.740 ;
        RECT 2034.650 22.540 2649.530 22.680 ;
        RECT 2034.650 22.480 2034.970 22.540 ;
        RECT 2649.210 22.480 2649.530 22.540 ;
      LAYER via ;
        RECT 2034.680 22.480 2034.940 22.740 ;
        RECT 2649.240 22.480 2649.500 22.740 ;
      LAYER met2 ;
        RECT 2033.530 600.170 2033.810 604.000 ;
        RECT 2033.530 600.030 2034.880 600.170 ;
        RECT 2033.530 600.000 2033.810 600.030 ;
        RECT 2034.740 22.770 2034.880 600.030 ;
        RECT 2034.680 22.450 2034.940 22.770 ;
        RECT 2649.240 22.450 2649.500 22.770 ;
        RECT 2649.300 2.400 2649.440 22.450 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2044.310 586.740 2044.630 586.800 ;
        RECT 2048.450 586.740 2048.770 586.800 ;
        RECT 2044.310 586.600 2048.770 586.740 ;
        RECT 2044.310 586.540 2044.630 586.600 ;
        RECT 2048.450 586.540 2048.770 586.600 ;
        RECT 2048.910 23.020 2049.230 23.080 ;
        RECT 2667.150 23.020 2667.470 23.080 ;
        RECT 2048.910 22.880 2667.470 23.020 ;
        RECT 2048.910 22.820 2049.230 22.880 ;
        RECT 2667.150 22.820 2667.470 22.880 ;
      LAYER via ;
        RECT 2044.340 586.540 2044.600 586.800 ;
        RECT 2048.480 586.540 2048.740 586.800 ;
        RECT 2048.940 22.820 2049.200 23.080 ;
        RECT 2667.180 22.820 2667.440 23.080 ;
      LAYER met2 ;
        RECT 2042.730 600.170 2043.010 604.000 ;
        RECT 2042.730 600.030 2044.540 600.170 ;
        RECT 2042.730 600.000 2043.010 600.030 ;
        RECT 2044.400 586.830 2044.540 600.030 ;
        RECT 2044.340 586.510 2044.600 586.830 ;
        RECT 2048.480 586.510 2048.740 586.830 ;
        RECT 2048.540 42.570 2048.680 586.510 ;
        RECT 2048.540 42.430 2049.140 42.570 ;
        RECT 2049.000 23.110 2049.140 42.430 ;
        RECT 2048.940 22.790 2049.200 23.110 ;
        RECT 2667.180 22.790 2667.440 23.110 ;
        RECT 2667.240 2.400 2667.380 22.790 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2053.510 586.740 2053.830 586.800 ;
        RECT 2055.810 586.740 2056.130 586.800 ;
        RECT 2053.510 586.600 2056.130 586.740 ;
        RECT 2053.510 586.540 2053.830 586.600 ;
        RECT 2055.810 586.540 2056.130 586.600 ;
        RECT 2055.810 23.360 2056.130 23.420 ;
        RECT 2684.630 23.360 2684.950 23.420 ;
        RECT 2055.810 23.220 2684.950 23.360 ;
        RECT 2055.810 23.160 2056.130 23.220 ;
        RECT 2684.630 23.160 2684.950 23.220 ;
      LAYER via ;
        RECT 2053.540 586.540 2053.800 586.800 ;
        RECT 2055.840 586.540 2056.100 586.800 ;
        RECT 2055.840 23.160 2056.100 23.420 ;
        RECT 2684.660 23.160 2684.920 23.420 ;
      LAYER met2 ;
        RECT 2051.930 600.170 2052.210 604.000 ;
        RECT 2051.930 600.030 2053.740 600.170 ;
        RECT 2051.930 600.000 2052.210 600.030 ;
        RECT 2053.600 586.830 2053.740 600.030 ;
        RECT 2053.540 586.510 2053.800 586.830 ;
        RECT 2055.840 586.510 2056.100 586.830 ;
        RECT 2055.900 23.450 2056.040 586.510 ;
        RECT 2055.840 23.130 2056.100 23.450 ;
        RECT 2684.660 23.130 2684.920 23.450 ;
        RECT 2684.720 2.400 2684.860 23.130 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2062.710 23.700 2063.030 23.760 ;
        RECT 2702.570 23.700 2702.890 23.760 ;
        RECT 2062.710 23.560 2702.890 23.700 ;
        RECT 2062.710 23.500 2063.030 23.560 ;
        RECT 2702.570 23.500 2702.890 23.560 ;
      LAYER via ;
        RECT 2062.740 23.500 2063.000 23.760 ;
        RECT 2702.600 23.500 2702.860 23.760 ;
      LAYER met2 ;
        RECT 2061.130 600.170 2061.410 604.000 ;
        RECT 2061.130 600.030 2062.940 600.170 ;
        RECT 2061.130 600.000 2061.410 600.030 ;
        RECT 2062.800 23.790 2062.940 600.030 ;
        RECT 2062.740 23.470 2063.000 23.790 ;
        RECT 2702.600 23.470 2702.860 23.790 ;
        RECT 2702.660 2.400 2702.800 23.470 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2071.910 586.740 2072.230 586.800 ;
        RECT 2076.510 586.740 2076.830 586.800 ;
        RECT 2071.910 586.600 2076.830 586.740 ;
        RECT 2071.910 586.540 2072.230 586.600 ;
        RECT 2076.510 586.540 2076.830 586.600 ;
        RECT 2076.510 27.440 2076.830 27.500 ;
        RECT 2720.510 27.440 2720.830 27.500 ;
        RECT 2076.510 27.300 2720.830 27.440 ;
        RECT 2076.510 27.240 2076.830 27.300 ;
        RECT 2720.510 27.240 2720.830 27.300 ;
      LAYER via ;
        RECT 2071.940 586.540 2072.200 586.800 ;
        RECT 2076.540 586.540 2076.800 586.800 ;
        RECT 2076.540 27.240 2076.800 27.500 ;
        RECT 2720.540 27.240 2720.800 27.500 ;
      LAYER met2 ;
        RECT 2070.330 600.170 2070.610 604.000 ;
        RECT 2070.330 600.030 2072.140 600.170 ;
        RECT 2070.330 600.000 2070.610 600.030 ;
        RECT 2072.000 586.830 2072.140 600.030 ;
        RECT 2071.940 586.510 2072.200 586.830 ;
        RECT 2076.540 586.510 2076.800 586.830 ;
        RECT 2076.600 27.530 2076.740 586.510 ;
        RECT 2076.540 27.210 2076.800 27.530 ;
        RECT 2720.540 27.210 2720.800 27.530 ;
        RECT 2720.600 2.400 2720.740 27.210 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2081.110 586.740 2081.430 586.800 ;
        RECT 2083.410 586.740 2083.730 586.800 ;
        RECT 2081.110 586.600 2083.730 586.740 ;
        RECT 2081.110 586.540 2081.430 586.600 ;
        RECT 2083.410 586.540 2083.730 586.600 ;
        RECT 2083.410 27.100 2083.730 27.160 ;
        RECT 2738.450 27.100 2738.770 27.160 ;
        RECT 2083.410 26.960 2738.770 27.100 ;
        RECT 2083.410 26.900 2083.730 26.960 ;
        RECT 2738.450 26.900 2738.770 26.960 ;
      LAYER via ;
        RECT 2081.140 586.540 2081.400 586.800 ;
        RECT 2083.440 586.540 2083.700 586.800 ;
        RECT 2083.440 26.900 2083.700 27.160 ;
        RECT 2738.480 26.900 2738.740 27.160 ;
      LAYER met2 ;
        RECT 2079.530 600.170 2079.810 604.000 ;
        RECT 2079.530 600.030 2081.340 600.170 ;
        RECT 2079.530 600.000 2079.810 600.030 ;
        RECT 2081.200 586.830 2081.340 600.030 ;
        RECT 2081.140 586.510 2081.400 586.830 ;
        RECT 2083.440 586.510 2083.700 586.830 ;
        RECT 2083.500 27.190 2083.640 586.510 ;
        RECT 2083.440 26.870 2083.700 27.190 ;
        RECT 2738.480 26.870 2738.740 27.190 ;
        RECT 2738.540 2.400 2738.680 26.870 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 26.760 2090.630 26.820 ;
        RECT 2755.930 26.760 2756.250 26.820 ;
        RECT 2090.310 26.620 2756.250 26.760 ;
        RECT 2090.310 26.560 2090.630 26.620 ;
        RECT 2755.930 26.560 2756.250 26.620 ;
      LAYER via ;
        RECT 2090.340 26.560 2090.600 26.820 ;
        RECT 2755.960 26.560 2756.220 26.820 ;
      LAYER met2 ;
        RECT 2088.730 600.170 2089.010 604.000 ;
        RECT 2088.730 600.030 2090.540 600.170 ;
        RECT 2088.730 600.000 2089.010 600.030 ;
        RECT 2090.400 26.850 2090.540 600.030 ;
        RECT 2090.340 26.530 2090.600 26.850 ;
        RECT 2755.960 26.530 2756.220 26.850 ;
        RECT 2756.020 2.400 2756.160 26.530 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 829.450 18.260 829.770 18.320 ;
        RECT 1098.090 18.260 1098.410 18.320 ;
        RECT 829.450 18.120 1098.410 18.260 ;
        RECT 829.450 18.060 829.770 18.120 ;
        RECT 1098.090 18.060 1098.410 18.120 ;
      LAYER via ;
        RECT 829.480 18.060 829.740 18.320 ;
        RECT 1098.120 18.060 1098.380 18.320 ;
      LAYER met2 ;
        RECT 1096.970 600.170 1097.250 604.000 ;
        RECT 1096.970 600.030 1098.320 600.170 ;
        RECT 1096.970 600.000 1097.250 600.030 ;
        RECT 1098.180 18.350 1098.320 600.030 ;
        RECT 829.480 18.030 829.740 18.350 ;
        RECT 1098.120 18.030 1098.380 18.350 ;
        RECT 829.540 2.400 829.680 18.030 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2099.510 587.420 2099.830 587.480 ;
        RECT 2104.110 587.420 2104.430 587.480 ;
        RECT 2099.510 587.280 2104.430 587.420 ;
        RECT 2099.510 587.220 2099.830 587.280 ;
        RECT 2104.110 587.220 2104.430 587.280 ;
        RECT 2104.110 26.420 2104.430 26.480 ;
        RECT 2773.870 26.420 2774.190 26.480 ;
        RECT 2104.110 26.280 2774.190 26.420 ;
        RECT 2104.110 26.220 2104.430 26.280 ;
        RECT 2773.870 26.220 2774.190 26.280 ;
      LAYER via ;
        RECT 2099.540 587.220 2099.800 587.480 ;
        RECT 2104.140 587.220 2104.400 587.480 ;
        RECT 2104.140 26.220 2104.400 26.480 ;
        RECT 2773.900 26.220 2774.160 26.480 ;
      LAYER met2 ;
        RECT 2097.930 600.170 2098.210 604.000 ;
        RECT 2097.930 600.030 2099.740 600.170 ;
        RECT 2097.930 600.000 2098.210 600.030 ;
        RECT 2099.600 587.510 2099.740 600.030 ;
        RECT 2099.540 587.190 2099.800 587.510 ;
        RECT 2104.140 587.190 2104.400 587.510 ;
        RECT 2104.200 26.510 2104.340 587.190 ;
        RECT 2104.140 26.190 2104.400 26.510 ;
        RECT 2773.900 26.190 2774.160 26.510 ;
        RECT 2773.960 2.400 2774.100 26.190 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2108.710 587.420 2109.030 587.480 ;
        RECT 2111.010 587.420 2111.330 587.480 ;
        RECT 2108.710 587.280 2111.330 587.420 ;
        RECT 2108.710 587.220 2109.030 587.280 ;
        RECT 2111.010 587.220 2111.330 587.280 ;
        RECT 2111.010 26.080 2111.330 26.140 ;
        RECT 2791.810 26.080 2792.130 26.140 ;
        RECT 2111.010 25.940 2792.130 26.080 ;
        RECT 2111.010 25.880 2111.330 25.940 ;
        RECT 2791.810 25.880 2792.130 25.940 ;
      LAYER via ;
        RECT 2108.740 587.220 2109.000 587.480 ;
        RECT 2111.040 587.220 2111.300 587.480 ;
        RECT 2111.040 25.880 2111.300 26.140 ;
        RECT 2791.840 25.880 2792.100 26.140 ;
      LAYER met2 ;
        RECT 2107.130 600.170 2107.410 604.000 ;
        RECT 2107.130 600.030 2108.940 600.170 ;
        RECT 2107.130 600.000 2107.410 600.030 ;
        RECT 2108.800 587.510 2108.940 600.030 ;
        RECT 2108.740 587.190 2109.000 587.510 ;
        RECT 2111.040 587.190 2111.300 587.510 ;
        RECT 2111.100 26.170 2111.240 587.190 ;
        RECT 2111.040 25.850 2111.300 26.170 ;
        RECT 2791.840 25.850 2792.100 26.170 ;
        RECT 2791.900 2.400 2792.040 25.850 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2117.910 25.400 2118.230 25.460 ;
        RECT 2809.750 25.400 2810.070 25.460 ;
        RECT 2117.910 25.260 2810.070 25.400 ;
        RECT 2117.910 25.200 2118.230 25.260 ;
        RECT 2809.750 25.200 2810.070 25.260 ;
      LAYER via ;
        RECT 2117.940 25.200 2118.200 25.460 ;
        RECT 2809.780 25.200 2810.040 25.460 ;
      LAYER met2 ;
        RECT 2116.330 600.170 2116.610 604.000 ;
        RECT 2116.330 600.030 2118.140 600.170 ;
        RECT 2116.330 600.000 2116.610 600.030 ;
        RECT 2118.000 25.490 2118.140 600.030 ;
        RECT 2117.940 25.170 2118.200 25.490 ;
        RECT 2809.780 25.170 2810.040 25.490 ;
        RECT 2809.840 2.400 2809.980 25.170 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2127.110 587.420 2127.430 587.480 ;
        RECT 2131.710 587.420 2132.030 587.480 ;
        RECT 2127.110 587.280 2132.030 587.420 ;
        RECT 2127.110 587.220 2127.430 587.280 ;
        RECT 2131.710 587.220 2132.030 587.280 ;
        RECT 2131.710 25.740 2132.030 25.800 ;
        RECT 2827.690 25.740 2828.010 25.800 ;
        RECT 2131.710 25.600 2828.010 25.740 ;
        RECT 2131.710 25.540 2132.030 25.600 ;
        RECT 2827.690 25.540 2828.010 25.600 ;
      LAYER via ;
        RECT 2127.140 587.220 2127.400 587.480 ;
        RECT 2131.740 587.220 2132.000 587.480 ;
        RECT 2131.740 25.540 2132.000 25.800 ;
        RECT 2827.720 25.540 2827.980 25.800 ;
      LAYER met2 ;
        RECT 2125.530 600.170 2125.810 604.000 ;
        RECT 2125.530 600.030 2127.340 600.170 ;
        RECT 2125.530 600.000 2125.810 600.030 ;
        RECT 2127.200 587.510 2127.340 600.030 ;
        RECT 2127.140 587.190 2127.400 587.510 ;
        RECT 2131.740 587.190 2132.000 587.510 ;
        RECT 2131.800 25.830 2131.940 587.190 ;
        RECT 2131.740 25.510 2132.000 25.830 ;
        RECT 2827.720 25.510 2827.980 25.830 ;
        RECT 2827.780 2.400 2827.920 25.510 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2136.310 573.820 2136.630 573.880 ;
        RECT 2138.610 573.820 2138.930 573.880 ;
        RECT 2136.310 573.680 2138.930 573.820 ;
        RECT 2136.310 573.620 2136.630 573.680 ;
        RECT 2138.610 573.620 2138.930 573.680 ;
        RECT 2138.610 25.060 2138.930 25.120 ;
        RECT 2845.170 25.060 2845.490 25.120 ;
        RECT 2138.610 24.920 2845.490 25.060 ;
        RECT 2138.610 24.860 2138.930 24.920 ;
        RECT 2845.170 24.860 2845.490 24.920 ;
      LAYER via ;
        RECT 2136.340 573.620 2136.600 573.880 ;
        RECT 2138.640 573.620 2138.900 573.880 ;
        RECT 2138.640 24.860 2138.900 25.120 ;
        RECT 2845.200 24.860 2845.460 25.120 ;
      LAYER met2 ;
        RECT 2134.730 600.170 2135.010 604.000 ;
        RECT 2134.730 600.030 2136.540 600.170 ;
        RECT 2134.730 600.000 2135.010 600.030 ;
        RECT 2136.400 573.910 2136.540 600.030 ;
        RECT 2136.340 573.590 2136.600 573.910 ;
        RECT 2138.640 573.590 2138.900 573.910 ;
        RECT 2138.700 25.150 2138.840 573.590 ;
        RECT 2138.640 24.830 2138.900 25.150 ;
        RECT 2845.200 24.830 2845.460 25.150 ;
        RECT 2845.260 2.400 2845.400 24.830 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.510 24.720 2145.830 24.780 ;
        RECT 2863.110 24.720 2863.430 24.780 ;
        RECT 2145.510 24.580 2863.430 24.720 ;
        RECT 2145.510 24.520 2145.830 24.580 ;
        RECT 2863.110 24.520 2863.430 24.580 ;
      LAYER via ;
        RECT 2145.540 24.520 2145.800 24.780 ;
        RECT 2863.140 24.520 2863.400 24.780 ;
      LAYER met2 ;
        RECT 2143.930 600.170 2144.210 604.000 ;
        RECT 2143.930 600.030 2145.740 600.170 ;
        RECT 2143.930 600.000 2144.210 600.030 ;
        RECT 2145.600 24.810 2145.740 600.030 ;
        RECT 2145.540 24.490 2145.800 24.810 ;
        RECT 2863.140 24.490 2863.400 24.810 ;
        RECT 2863.200 2.400 2863.340 24.490 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2154.710 588.440 2155.030 588.500 ;
        RECT 2159.310 588.440 2159.630 588.500 ;
        RECT 2154.710 588.300 2159.630 588.440 ;
        RECT 2154.710 588.240 2155.030 588.300 ;
        RECT 2159.310 588.240 2159.630 588.300 ;
        RECT 2159.310 24.380 2159.630 24.440 ;
        RECT 2881.050 24.380 2881.370 24.440 ;
        RECT 2159.310 24.240 2881.370 24.380 ;
        RECT 2159.310 24.180 2159.630 24.240 ;
        RECT 2881.050 24.180 2881.370 24.240 ;
      LAYER via ;
        RECT 2154.740 588.240 2155.000 588.500 ;
        RECT 2159.340 588.240 2159.600 588.500 ;
        RECT 2159.340 24.180 2159.600 24.440 ;
        RECT 2881.080 24.180 2881.340 24.440 ;
      LAYER met2 ;
        RECT 2153.130 600.170 2153.410 604.000 ;
        RECT 2153.130 600.030 2154.940 600.170 ;
        RECT 2153.130 600.000 2153.410 600.030 ;
        RECT 2154.800 588.530 2154.940 600.030 ;
        RECT 2154.740 588.210 2155.000 588.530 ;
        RECT 2159.340 588.210 2159.600 588.530 ;
        RECT 2159.400 24.470 2159.540 588.210 ;
        RECT 2159.340 24.150 2159.600 24.470 ;
        RECT 2881.080 24.150 2881.340 24.470 ;
        RECT 2881.140 2.400 2881.280 24.150 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2163.910 587.420 2164.230 587.480 ;
        RECT 2166.210 587.420 2166.530 587.480 ;
        RECT 2163.910 587.280 2166.530 587.420 ;
        RECT 2163.910 587.220 2164.230 587.280 ;
        RECT 2166.210 587.220 2166.530 587.280 ;
        RECT 2166.210 24.040 2166.530 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 2166.210 23.900 2899.310 24.040 ;
        RECT 2166.210 23.840 2166.530 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 2163.940 587.220 2164.200 587.480 ;
        RECT 2166.240 587.220 2166.500 587.480 ;
        RECT 2166.240 23.840 2166.500 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 2162.330 600.170 2162.610 604.000 ;
        RECT 2162.330 600.030 2164.140 600.170 ;
        RECT 2162.330 600.000 2162.610 600.030 ;
        RECT 2164.000 587.510 2164.140 600.030 ;
        RECT 2163.940 587.190 2164.200 587.510 ;
        RECT 2166.240 587.190 2166.500 587.510 ;
        RECT 2166.300 24.130 2166.440 587.190 ;
        RECT 2166.240 23.810 2166.500 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.400 2899.220 23.810 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 846.930 18.600 847.250 18.660 ;
        RECT 1036.910 18.600 1037.230 18.660 ;
        RECT 846.930 18.460 1037.230 18.600 ;
        RECT 846.930 18.400 847.250 18.460 ;
        RECT 1036.910 18.400 1037.230 18.460 ;
        RECT 1036.910 16.220 1037.230 16.280 ;
        RECT 1102.230 16.220 1102.550 16.280 ;
        RECT 1036.910 16.080 1102.550 16.220 ;
        RECT 1036.910 16.020 1037.230 16.080 ;
        RECT 1102.230 16.020 1102.550 16.080 ;
      LAYER via ;
        RECT 846.960 18.400 847.220 18.660 ;
        RECT 1036.940 18.400 1037.200 18.660 ;
        RECT 1036.940 16.020 1037.200 16.280 ;
        RECT 1102.260 16.020 1102.520 16.280 ;
      LAYER met2 ;
        RECT 1106.170 600.170 1106.450 604.000 ;
        RECT 1104.160 600.030 1106.450 600.170 ;
        RECT 846.960 18.370 847.220 18.690 ;
        RECT 1036.940 18.370 1037.200 18.690 ;
        RECT 847.020 2.400 847.160 18.370 ;
        RECT 1037.000 16.310 1037.140 18.370 ;
        RECT 1104.160 16.730 1104.300 600.030 ;
        RECT 1106.170 600.000 1106.450 600.030 ;
        RECT 1102.320 16.590 1104.300 16.730 ;
        RECT 1102.320 16.310 1102.460 16.590 ;
        RECT 1036.940 15.990 1037.200 16.310 ;
        RECT 1102.260 15.990 1102.520 16.310 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1111.890 545.400 1112.210 545.660 ;
        RECT 1111.980 544.980 1112.120 545.400 ;
        RECT 1111.890 544.720 1112.210 544.980 ;
        RECT 1111.430 524.520 1111.750 524.580 ;
        RECT 1111.890 524.520 1112.210 524.580 ;
        RECT 1111.430 524.380 1112.210 524.520 ;
        RECT 1111.430 524.320 1111.750 524.380 ;
        RECT 1111.890 524.320 1112.210 524.380 ;
        RECT 1111.430 458.900 1111.750 458.960 ;
        RECT 1112.350 458.900 1112.670 458.960 ;
        RECT 1111.430 458.760 1112.670 458.900 ;
        RECT 1111.430 458.700 1111.750 458.760 ;
        RECT 1112.350 458.700 1112.670 458.760 ;
        RECT 1111.430 386.480 1111.750 386.540 ;
        RECT 1111.890 386.480 1112.210 386.540 ;
        RECT 1111.430 386.340 1112.210 386.480 ;
        RECT 1111.430 386.280 1111.750 386.340 ;
        RECT 1111.890 386.280 1112.210 386.340 ;
        RECT 1111.430 110.540 1111.750 110.800 ;
        RECT 1111.520 110.120 1111.660 110.540 ;
        RECT 1111.430 109.860 1111.750 110.120 ;
        RECT 864.870 18.940 865.190 19.000 ;
        RECT 1111.430 18.940 1111.750 19.000 ;
        RECT 864.870 18.800 1111.750 18.940 ;
        RECT 864.870 18.740 865.190 18.800 ;
        RECT 1111.430 18.740 1111.750 18.800 ;
      LAYER via ;
        RECT 1111.920 545.400 1112.180 545.660 ;
        RECT 1111.920 544.720 1112.180 544.980 ;
        RECT 1111.460 524.320 1111.720 524.580 ;
        RECT 1111.920 524.320 1112.180 524.580 ;
        RECT 1111.460 458.700 1111.720 458.960 ;
        RECT 1112.380 458.700 1112.640 458.960 ;
        RECT 1111.460 386.280 1111.720 386.540 ;
        RECT 1111.920 386.280 1112.180 386.540 ;
        RECT 1111.460 110.540 1111.720 110.800 ;
        RECT 1111.460 109.860 1111.720 110.120 ;
        RECT 864.900 18.740 865.160 19.000 ;
        RECT 1111.460 18.740 1111.720 19.000 ;
      LAYER met2 ;
        RECT 1114.910 600.170 1115.190 604.000 ;
        RECT 1113.820 600.030 1115.190 600.170 ;
        RECT 1113.820 596.770 1113.960 600.030 ;
        RECT 1114.910 600.000 1115.190 600.030 ;
        RECT 1111.980 596.630 1113.960 596.770 ;
        RECT 1111.980 545.690 1112.120 596.630 ;
        RECT 1111.920 545.370 1112.180 545.690 ;
        RECT 1111.920 544.690 1112.180 545.010 ;
        RECT 1111.980 524.610 1112.120 544.690 ;
        RECT 1111.460 524.290 1111.720 524.610 ;
        RECT 1111.920 524.290 1112.180 524.610 ;
        RECT 1111.520 524.125 1111.660 524.290 ;
        RECT 1111.450 523.755 1111.730 524.125 ;
        RECT 1112.370 523.075 1112.650 523.445 ;
        RECT 1112.440 458.990 1112.580 523.075 ;
        RECT 1111.460 458.670 1111.720 458.990 ;
        RECT 1112.380 458.670 1112.640 458.990 ;
        RECT 1111.520 386.570 1111.660 458.670 ;
        RECT 1111.460 386.250 1111.720 386.570 ;
        RECT 1111.920 386.250 1112.180 386.570 ;
        RECT 1111.980 303.690 1112.120 386.250 ;
        RECT 1111.520 303.550 1112.120 303.690 ;
        RECT 1111.520 303.010 1111.660 303.550 ;
        RECT 1111.520 302.870 1112.120 303.010 ;
        RECT 1111.980 207.130 1112.120 302.870 ;
        RECT 1111.520 206.990 1112.120 207.130 ;
        RECT 1111.520 206.450 1111.660 206.990 ;
        RECT 1111.520 206.310 1112.120 206.450 ;
        RECT 1111.980 145.250 1112.120 206.310 ;
        RECT 1111.520 145.110 1112.120 145.250 ;
        RECT 1111.520 110.830 1111.660 145.110 ;
        RECT 1111.460 110.510 1111.720 110.830 ;
        RECT 1111.460 109.830 1111.720 110.150 ;
        RECT 1111.520 19.030 1111.660 109.830 ;
        RECT 864.900 18.710 865.160 19.030 ;
        RECT 1111.460 18.710 1111.720 19.030 ;
        RECT 864.960 2.400 865.100 18.710 ;
        RECT 864.750 -4.800 865.310 2.400 ;
      LAYER via2 ;
        RECT 1111.450 523.800 1111.730 524.080 ;
        RECT 1112.370 523.120 1112.650 523.400 ;
      LAYER met3 ;
        RECT 1111.425 524.090 1111.755 524.105 ;
        RECT 1110.750 523.790 1111.755 524.090 ;
        RECT 1110.750 523.410 1111.050 523.790 ;
        RECT 1111.425 523.775 1111.755 523.790 ;
        RECT 1112.345 523.410 1112.675 523.425 ;
        RECT 1110.750 523.110 1112.675 523.410 ;
        RECT 1112.345 523.095 1112.675 523.110 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1118.330 524.180 1118.650 524.240 ;
        RECT 1118.790 524.180 1119.110 524.240 ;
        RECT 1118.330 524.040 1119.110 524.180 ;
        RECT 1118.330 523.980 1118.650 524.040 ;
        RECT 1118.790 523.980 1119.110 524.040 ;
        RECT 1118.330 255.720 1118.650 255.980 ;
        RECT 1118.420 255.300 1118.560 255.720 ;
        RECT 1118.330 255.040 1118.650 255.300 ;
        RECT 1118.330 110.540 1118.650 110.800 ;
        RECT 1118.420 110.120 1118.560 110.540 ;
        RECT 1118.330 109.860 1118.650 110.120 ;
        RECT 1117.870 90.000 1118.190 90.060 ;
        RECT 1118.330 90.000 1118.650 90.060 ;
        RECT 1117.870 89.860 1118.650 90.000 ;
        RECT 1117.870 89.800 1118.190 89.860 ;
        RECT 1118.330 89.800 1118.650 89.860 ;
        RECT 882.810 19.280 883.130 19.340 ;
        RECT 1090.270 19.280 1090.590 19.340 ;
        RECT 882.810 19.140 1090.590 19.280 ;
        RECT 882.810 19.080 883.130 19.140 ;
        RECT 1090.270 19.080 1090.590 19.140 ;
        RECT 1090.270 17.580 1090.590 17.640 ;
        RECT 1118.330 17.580 1118.650 17.640 ;
        RECT 1090.270 17.440 1118.650 17.580 ;
        RECT 1090.270 17.380 1090.590 17.440 ;
        RECT 1118.330 17.380 1118.650 17.440 ;
      LAYER via ;
        RECT 1118.360 523.980 1118.620 524.240 ;
        RECT 1118.820 523.980 1119.080 524.240 ;
        RECT 1118.360 255.720 1118.620 255.980 ;
        RECT 1118.360 255.040 1118.620 255.300 ;
        RECT 1118.360 110.540 1118.620 110.800 ;
        RECT 1118.360 109.860 1118.620 110.120 ;
        RECT 1117.900 89.800 1118.160 90.060 ;
        RECT 1118.360 89.800 1118.620 90.060 ;
        RECT 882.840 19.080 883.100 19.340 ;
        RECT 1090.300 19.080 1090.560 19.340 ;
        RECT 1090.300 17.380 1090.560 17.640 ;
        RECT 1118.360 17.380 1118.620 17.640 ;
      LAYER met2 ;
        RECT 1124.110 600.850 1124.390 604.000 ;
        RECT 1122.100 600.710 1124.390 600.850 ;
        RECT 1122.100 596.770 1122.240 600.710 ;
        RECT 1124.110 600.000 1124.390 600.710 ;
        RECT 1120.260 596.630 1122.240 596.770 ;
        RECT 1120.260 569.570 1120.400 596.630 ;
        RECT 1118.420 569.430 1120.400 569.570 ;
        RECT 1118.420 524.270 1118.560 569.430 ;
        RECT 1118.360 523.950 1118.620 524.270 ;
        RECT 1118.820 523.950 1119.080 524.270 ;
        RECT 1118.880 400.930 1119.020 523.950 ;
        RECT 1118.880 400.790 1119.480 400.930 ;
        RECT 1119.340 400.250 1119.480 400.790 ;
        RECT 1118.420 400.110 1119.480 400.250 ;
        RECT 1118.420 351.970 1118.560 400.110 ;
        RECT 1117.960 351.830 1118.560 351.970 ;
        RECT 1117.960 351.290 1118.100 351.830 ;
        RECT 1117.960 351.150 1118.560 351.290 ;
        RECT 1118.420 256.010 1118.560 351.150 ;
        RECT 1118.360 255.690 1118.620 256.010 ;
        RECT 1118.360 255.010 1118.620 255.330 ;
        RECT 1118.420 110.830 1118.560 255.010 ;
        RECT 1118.360 110.510 1118.620 110.830 ;
        RECT 1118.360 109.830 1118.620 110.150 ;
        RECT 1118.420 90.090 1118.560 109.830 ;
        RECT 1117.900 89.770 1118.160 90.090 ;
        RECT 1118.360 89.770 1118.620 90.090 ;
        RECT 1117.960 41.210 1118.100 89.770 ;
        RECT 1117.960 41.070 1118.560 41.210 ;
        RECT 882.840 19.050 883.100 19.370 ;
        RECT 1090.300 19.050 1090.560 19.370 ;
        RECT 882.900 2.400 883.040 19.050 ;
        RECT 1090.360 17.670 1090.500 19.050 ;
        RECT 1118.420 17.670 1118.560 41.070 ;
        RECT 1090.300 17.350 1090.560 17.670 ;
        RECT 1118.360 17.350 1118.620 17.670 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 900.750 19.620 901.070 19.680 ;
        RECT 1132.130 19.620 1132.450 19.680 ;
        RECT 900.750 19.480 1132.450 19.620 ;
        RECT 900.750 19.420 901.070 19.480 ;
        RECT 1132.130 19.420 1132.450 19.480 ;
      LAYER via ;
        RECT 900.780 19.420 901.040 19.680 ;
        RECT 1132.160 19.420 1132.420 19.680 ;
      LAYER met2 ;
        RECT 1133.310 600.170 1133.590 604.000 ;
        RECT 1132.220 600.030 1133.590 600.170 ;
        RECT 1132.220 19.710 1132.360 600.030 ;
        RECT 1133.310 600.000 1133.590 600.030 ;
        RECT 900.780 19.390 901.040 19.710 ;
        RECT 1132.160 19.390 1132.420 19.710 ;
        RECT 900.840 2.400 900.980 19.390 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1139.490 548.660 1139.810 548.720 ;
        RECT 1140.410 548.660 1140.730 548.720 ;
        RECT 1139.490 548.520 1140.730 548.660 ;
        RECT 1139.490 548.460 1139.810 548.520 ;
        RECT 1140.410 548.460 1140.730 548.520 ;
        RECT 1139.030 524.860 1139.350 524.920 ;
        RECT 1140.410 524.860 1140.730 524.920 ;
        RECT 1139.030 524.720 1140.730 524.860 ;
        RECT 1139.030 524.660 1139.350 524.720 ;
        RECT 1140.410 524.660 1140.730 524.720 ;
        RECT 1137.650 524.180 1137.970 524.240 ;
        RECT 1139.030 524.180 1139.350 524.240 ;
        RECT 1137.650 524.040 1139.350 524.180 ;
        RECT 1137.650 523.980 1137.970 524.040 ;
        RECT 1139.030 523.980 1139.350 524.040 ;
        RECT 1139.030 475.900 1139.350 475.960 ;
        RECT 1140.410 475.900 1140.730 475.960 ;
        RECT 1139.030 475.760 1140.730 475.900 ;
        RECT 1139.030 475.700 1139.350 475.760 ;
        RECT 1140.410 475.700 1140.730 475.760 ;
        RECT 1139.490 338.200 1139.810 338.260 ;
        RECT 1139.950 338.200 1140.270 338.260 ;
        RECT 1139.490 338.060 1140.270 338.200 ;
        RECT 1139.490 338.000 1139.810 338.060 ;
        RECT 1139.950 338.000 1140.270 338.060 ;
        RECT 1139.030 137.940 1139.350 138.000 ;
        RECT 1139.490 137.940 1139.810 138.000 ;
        RECT 1139.030 137.800 1139.810 137.940 ;
        RECT 1139.030 137.740 1139.350 137.800 ;
        RECT 1139.490 137.740 1139.810 137.800 ;
        RECT 1139.490 110.740 1139.810 110.800 ;
        RECT 1139.120 110.600 1139.810 110.740 ;
        RECT 1139.120 110.460 1139.260 110.600 ;
        RECT 1139.490 110.540 1139.810 110.600 ;
        RECT 1139.030 110.200 1139.350 110.460 ;
        RECT 918.690 19.960 919.010 20.020 ;
        RECT 1139.030 19.960 1139.350 20.020 ;
        RECT 918.690 19.820 1139.350 19.960 ;
        RECT 918.690 19.760 919.010 19.820 ;
        RECT 1139.030 19.760 1139.350 19.820 ;
      LAYER via ;
        RECT 1139.520 548.460 1139.780 548.720 ;
        RECT 1140.440 548.460 1140.700 548.720 ;
        RECT 1139.060 524.660 1139.320 524.920 ;
        RECT 1140.440 524.660 1140.700 524.920 ;
        RECT 1137.680 523.980 1137.940 524.240 ;
        RECT 1139.060 523.980 1139.320 524.240 ;
        RECT 1139.060 475.700 1139.320 475.960 ;
        RECT 1140.440 475.700 1140.700 475.960 ;
        RECT 1139.520 338.000 1139.780 338.260 ;
        RECT 1139.980 338.000 1140.240 338.260 ;
        RECT 1139.060 137.740 1139.320 138.000 ;
        RECT 1139.520 137.740 1139.780 138.000 ;
        RECT 1139.520 110.540 1139.780 110.800 ;
        RECT 1139.060 110.200 1139.320 110.460 ;
        RECT 918.720 19.760 918.980 20.020 ;
        RECT 1139.060 19.760 1139.320 20.020 ;
      LAYER met2 ;
        RECT 1142.510 600.170 1142.790 604.000 ;
        RECT 1140.500 600.030 1142.790 600.170 ;
        RECT 1140.500 596.770 1140.640 600.030 ;
        RECT 1142.510 600.000 1142.790 600.030 ;
        RECT 1139.580 596.630 1140.640 596.770 ;
        RECT 1139.580 548.750 1139.720 596.630 ;
        RECT 1139.520 548.430 1139.780 548.750 ;
        RECT 1140.440 548.430 1140.700 548.750 ;
        RECT 1140.500 524.950 1140.640 548.430 ;
        RECT 1139.060 524.630 1139.320 524.950 ;
        RECT 1140.440 524.630 1140.700 524.950 ;
        RECT 1139.120 524.270 1139.260 524.630 ;
        RECT 1137.680 523.950 1137.940 524.270 ;
        RECT 1139.060 523.950 1139.320 524.270 ;
        RECT 1137.740 476.525 1137.880 523.950 ;
        RECT 1137.670 476.155 1137.950 476.525 ;
        RECT 1139.050 476.155 1139.330 476.525 ;
        RECT 1139.120 475.990 1139.260 476.155 ;
        RECT 1139.060 475.670 1139.320 475.990 ;
        RECT 1140.440 475.670 1140.700 475.990 ;
        RECT 1140.500 433.570 1140.640 475.670 ;
        RECT 1139.120 433.430 1140.640 433.570 ;
        RECT 1139.120 400.930 1139.260 433.430 ;
        RECT 1139.120 400.790 1140.180 400.930 ;
        RECT 1140.040 338.290 1140.180 400.790 ;
        RECT 1139.520 337.970 1139.780 338.290 ;
        RECT 1139.980 337.970 1140.240 338.290 ;
        RECT 1139.580 303.690 1139.720 337.970 ;
        RECT 1139.120 303.550 1139.720 303.690 ;
        RECT 1139.120 303.010 1139.260 303.550 ;
        RECT 1139.120 302.870 1139.720 303.010 ;
        RECT 1139.580 207.130 1139.720 302.870 ;
        RECT 1139.120 206.990 1139.720 207.130 ;
        RECT 1139.120 206.450 1139.260 206.990 ;
        RECT 1139.120 206.310 1139.720 206.450 ;
        RECT 1139.580 145.250 1139.720 206.310 ;
        RECT 1139.120 145.110 1139.720 145.250 ;
        RECT 1139.120 138.030 1139.260 145.110 ;
        RECT 1139.060 137.710 1139.320 138.030 ;
        RECT 1139.520 137.710 1139.780 138.030 ;
        RECT 1139.580 110.830 1139.720 137.710 ;
        RECT 1139.520 110.510 1139.780 110.830 ;
        RECT 1139.060 110.170 1139.320 110.490 ;
        RECT 1139.120 20.050 1139.260 110.170 ;
        RECT 918.720 19.730 918.980 20.050 ;
        RECT 1139.060 19.730 1139.320 20.050 ;
        RECT 918.780 2.400 918.920 19.730 ;
        RECT 918.570 -4.800 919.130 2.400 ;
      LAYER via2 ;
        RECT 1137.670 476.200 1137.950 476.480 ;
        RECT 1139.050 476.200 1139.330 476.480 ;
      LAYER met3 ;
        RECT 1137.645 476.490 1137.975 476.505 ;
        RECT 1139.025 476.490 1139.355 476.505 ;
        RECT 1137.645 476.190 1139.355 476.490 ;
        RECT 1137.645 476.175 1137.975 476.190 ;
        RECT 1139.025 476.175 1139.355 476.190 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.930 255.720 1146.250 255.980 ;
        RECT 1146.020 255.300 1146.160 255.720 ;
        RECT 1145.930 255.040 1146.250 255.300 ;
        RECT 936.170 27.100 936.490 27.160 ;
        RECT 1145.470 27.100 1145.790 27.160 ;
        RECT 936.170 26.960 1145.790 27.100 ;
        RECT 936.170 26.900 936.490 26.960 ;
        RECT 1145.470 26.900 1145.790 26.960 ;
      LAYER via ;
        RECT 1145.960 255.720 1146.220 255.980 ;
        RECT 1145.960 255.040 1146.220 255.300 ;
        RECT 936.200 26.900 936.460 27.160 ;
        RECT 1145.500 26.900 1145.760 27.160 ;
      LAYER met2 ;
        RECT 1151.710 600.170 1151.990 604.000 ;
        RECT 1149.700 600.030 1151.990 600.170 ;
        RECT 1149.700 596.770 1149.840 600.030 ;
        RECT 1151.710 600.000 1151.990 600.030 ;
        RECT 1147.860 596.630 1149.840 596.770 ;
        RECT 1147.860 569.570 1148.000 596.630 ;
        RECT 1146.020 569.430 1148.000 569.570 ;
        RECT 1146.020 500.210 1146.160 569.430 ;
        RECT 1146.020 500.070 1146.620 500.210 ;
        RECT 1146.480 458.730 1146.620 500.070 ;
        RECT 1146.480 458.590 1147.080 458.730 ;
        RECT 1146.940 447.170 1147.080 458.590 ;
        RECT 1146.480 447.030 1147.080 447.170 ;
        RECT 1146.480 410.450 1146.620 447.030 ;
        RECT 1146.020 410.310 1146.620 410.450 ;
        RECT 1146.020 351.970 1146.160 410.310 ;
        RECT 1145.560 351.830 1146.160 351.970 ;
        RECT 1145.560 351.290 1145.700 351.830 ;
        RECT 1145.560 351.150 1146.160 351.290 ;
        RECT 1146.020 256.010 1146.160 351.150 ;
        RECT 1145.960 255.690 1146.220 256.010 ;
        RECT 1145.960 255.010 1146.220 255.330 ;
        RECT 1146.020 158.850 1146.160 255.010 ;
        RECT 1145.560 158.710 1146.160 158.850 ;
        RECT 1145.560 158.170 1145.700 158.710 ;
        RECT 1145.560 158.030 1146.160 158.170 ;
        RECT 1146.020 62.290 1146.160 158.030 ;
        RECT 1145.560 62.150 1146.160 62.290 ;
        RECT 1145.560 27.190 1145.700 62.150 ;
        RECT 936.200 26.870 936.460 27.190 ;
        RECT 1145.500 26.870 1145.760 27.190 ;
        RECT 936.260 2.400 936.400 26.870 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 954.110 20.640 954.430 20.700 ;
        RECT 1131.670 20.640 1131.990 20.700 ;
        RECT 954.110 20.500 1131.990 20.640 ;
        RECT 954.110 20.440 954.430 20.500 ;
        RECT 1131.670 20.440 1131.990 20.500 ;
        RECT 1131.670 19.280 1131.990 19.340 ;
        RECT 1159.730 19.280 1160.050 19.340 ;
        RECT 1131.670 19.140 1160.050 19.280 ;
        RECT 1131.670 19.080 1131.990 19.140 ;
        RECT 1159.730 19.080 1160.050 19.140 ;
      LAYER via ;
        RECT 954.140 20.440 954.400 20.700 ;
        RECT 1131.700 20.440 1131.960 20.700 ;
        RECT 1131.700 19.080 1131.960 19.340 ;
        RECT 1159.760 19.080 1160.020 19.340 ;
      LAYER met2 ;
        RECT 1160.910 600.170 1161.190 604.000 ;
        RECT 1159.820 600.030 1161.190 600.170 ;
        RECT 954.140 20.410 954.400 20.730 ;
        RECT 1131.700 20.410 1131.960 20.730 ;
        RECT 954.200 2.400 954.340 20.410 ;
        RECT 1131.760 19.370 1131.900 20.410 ;
        RECT 1159.820 19.370 1159.960 600.030 ;
        RECT 1160.910 600.000 1161.190 600.030 ;
        RECT 1131.700 19.050 1131.960 19.370 ;
        RECT 1159.760 19.050 1160.020 19.370 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1167.090 572.460 1167.410 572.520 ;
        RECT 1168.010 572.460 1168.330 572.520 ;
        RECT 1167.090 572.320 1168.330 572.460 ;
        RECT 1167.090 572.260 1167.410 572.320 ;
        RECT 1168.010 572.260 1168.330 572.320 ;
        RECT 1166.630 524.520 1166.950 524.580 ;
        RECT 1168.010 524.520 1168.330 524.580 ;
        RECT 1166.630 524.380 1168.330 524.520 ;
        RECT 1166.630 524.320 1166.950 524.380 ;
        RECT 1168.010 524.320 1168.330 524.380 ;
        RECT 1166.630 476.240 1166.950 476.300 ;
        RECT 1167.090 476.240 1167.410 476.300 ;
        RECT 1166.630 476.100 1167.410 476.240 ;
        RECT 1166.630 476.040 1166.950 476.100 ;
        RECT 1167.090 476.040 1167.410 476.100 ;
        RECT 1167.090 420.820 1167.410 420.880 ;
        RECT 1168.010 420.820 1168.330 420.880 ;
        RECT 1167.090 420.680 1168.330 420.820 ;
        RECT 1167.090 420.620 1167.410 420.680 ;
        RECT 1168.010 420.620 1168.330 420.680 ;
        RECT 1167.090 396.680 1167.410 396.740 ;
        RECT 1168.010 396.680 1168.330 396.740 ;
        RECT 1167.090 396.540 1168.330 396.680 ;
        RECT 1167.090 396.480 1167.410 396.540 ;
        RECT 1168.010 396.480 1168.330 396.540 ;
        RECT 1126.150 18.940 1126.470 19.000 ;
        RECT 1167.090 18.940 1167.410 19.000 ;
        RECT 1126.150 18.800 1167.410 18.940 ;
        RECT 1126.150 18.740 1126.470 18.800 ;
        RECT 1167.090 18.740 1167.410 18.800 ;
        RECT 972.050 16.900 972.370 16.960 ;
        RECT 1126.150 16.900 1126.470 16.960 ;
        RECT 972.050 16.760 1126.470 16.900 ;
        RECT 972.050 16.700 972.370 16.760 ;
        RECT 1126.150 16.700 1126.470 16.760 ;
      LAYER via ;
        RECT 1167.120 572.260 1167.380 572.520 ;
        RECT 1168.040 572.260 1168.300 572.520 ;
        RECT 1166.660 524.320 1166.920 524.580 ;
        RECT 1168.040 524.320 1168.300 524.580 ;
        RECT 1166.660 476.040 1166.920 476.300 ;
        RECT 1167.120 476.040 1167.380 476.300 ;
        RECT 1167.120 420.620 1167.380 420.880 ;
        RECT 1168.040 420.620 1168.300 420.880 ;
        RECT 1167.120 396.480 1167.380 396.740 ;
        RECT 1168.040 396.480 1168.300 396.740 ;
        RECT 1126.180 18.740 1126.440 19.000 ;
        RECT 1167.120 18.740 1167.380 19.000 ;
        RECT 972.080 16.700 972.340 16.960 ;
        RECT 1126.180 16.700 1126.440 16.960 ;
      LAYER met2 ;
        RECT 1170.110 600.170 1170.390 604.000 ;
        RECT 1168.100 600.030 1170.390 600.170 ;
        RECT 1168.100 596.770 1168.240 600.030 ;
        RECT 1170.110 600.000 1170.390 600.030 ;
        RECT 1167.180 596.630 1168.240 596.770 ;
        RECT 1167.180 572.550 1167.320 596.630 ;
        RECT 1167.120 572.230 1167.380 572.550 ;
        RECT 1168.040 572.230 1168.300 572.550 ;
        RECT 1168.100 524.610 1168.240 572.230 ;
        RECT 1166.660 524.290 1166.920 524.610 ;
        RECT 1168.040 524.290 1168.300 524.610 ;
        RECT 1166.720 476.330 1166.860 524.290 ;
        RECT 1166.660 476.010 1166.920 476.330 ;
        RECT 1167.120 476.010 1167.380 476.330 ;
        RECT 1167.180 420.910 1167.320 476.010 ;
        RECT 1167.120 420.590 1167.380 420.910 ;
        RECT 1168.040 420.590 1168.300 420.910 ;
        RECT 1168.100 396.770 1168.240 420.590 ;
        RECT 1167.120 396.450 1167.380 396.770 ;
        RECT 1168.040 396.450 1168.300 396.770 ;
        RECT 1167.180 303.690 1167.320 396.450 ;
        RECT 1166.720 303.550 1167.320 303.690 ;
        RECT 1166.720 303.010 1166.860 303.550 ;
        RECT 1166.720 302.870 1167.320 303.010 ;
        RECT 1167.180 207.130 1167.320 302.870 ;
        RECT 1166.720 206.990 1167.320 207.130 ;
        RECT 1166.720 206.450 1166.860 206.990 ;
        RECT 1166.720 206.310 1167.320 206.450 ;
        RECT 1167.180 110.570 1167.320 206.310 ;
        RECT 1166.720 110.430 1167.320 110.570 ;
        RECT 1166.720 109.890 1166.860 110.430 ;
        RECT 1166.720 109.750 1167.320 109.890 ;
        RECT 1167.180 19.030 1167.320 109.750 ;
        RECT 1126.180 18.710 1126.440 19.030 ;
        RECT 1167.120 18.710 1167.380 19.030 ;
        RECT 1126.240 16.990 1126.380 18.710 ;
        RECT 972.080 16.670 972.340 16.990 ;
        RECT 1126.180 16.670 1126.440 16.990 ;
        RECT 972.140 2.400 972.280 16.670 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1000.570 583.000 1000.890 583.060 ;
        RECT 1003.330 583.000 1003.650 583.060 ;
        RECT 1000.570 582.860 1003.650 583.000 ;
        RECT 1000.570 582.800 1000.890 582.860 ;
        RECT 1003.330 582.800 1003.650 582.860 ;
        RECT 650.970 35.600 651.290 35.660 ;
        RECT 1000.570 35.600 1000.890 35.660 ;
        RECT 650.970 35.460 1000.890 35.600 ;
        RECT 650.970 35.400 651.290 35.460 ;
        RECT 1000.570 35.400 1000.890 35.460 ;
      LAYER via ;
        RECT 1000.600 582.800 1000.860 583.060 ;
        RECT 1003.360 582.800 1003.620 583.060 ;
        RECT 651.000 35.400 651.260 35.660 ;
        RECT 1000.600 35.400 1000.860 35.660 ;
      LAYER met2 ;
        RECT 1004.970 600.170 1005.250 604.000 ;
        RECT 1003.420 600.030 1005.250 600.170 ;
        RECT 1003.420 583.090 1003.560 600.030 ;
        RECT 1004.970 600.000 1005.250 600.030 ;
        RECT 1000.600 582.770 1000.860 583.090 ;
        RECT 1003.360 582.770 1003.620 583.090 ;
        RECT 1000.660 35.690 1000.800 582.770 ;
        RECT 651.000 35.370 651.260 35.690 ;
        RECT 1000.600 35.370 1000.860 35.690 ;
        RECT 651.060 2.400 651.200 35.370 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1173.990 400.760 1174.310 400.820 ;
        RECT 1173.620 400.620 1174.310 400.760 ;
        RECT 1173.620 400.480 1173.760 400.620 ;
        RECT 1173.990 400.560 1174.310 400.620 ;
        RECT 1173.530 400.220 1173.850 400.480 ;
        RECT 1014.830 23.020 1015.150 23.080 ;
        RECT 1173.070 23.020 1173.390 23.080 ;
        RECT 1014.830 22.880 1173.390 23.020 ;
        RECT 1014.830 22.820 1015.150 22.880 ;
        RECT 1173.070 22.820 1173.390 22.880 ;
        RECT 989.990 14.860 990.310 14.920 ;
        RECT 1014.830 14.860 1015.150 14.920 ;
        RECT 989.990 14.720 1015.150 14.860 ;
        RECT 989.990 14.660 990.310 14.720 ;
        RECT 1014.830 14.660 1015.150 14.720 ;
      LAYER via ;
        RECT 1174.020 400.560 1174.280 400.820 ;
        RECT 1173.560 400.220 1173.820 400.480 ;
        RECT 1014.860 22.820 1015.120 23.080 ;
        RECT 1173.100 22.820 1173.360 23.080 ;
        RECT 990.020 14.660 990.280 14.920 ;
        RECT 1014.860 14.660 1015.120 14.920 ;
      LAYER met2 ;
        RECT 1179.310 600.170 1179.590 604.000 ;
        RECT 1177.300 600.030 1179.590 600.170 ;
        RECT 1177.300 596.770 1177.440 600.030 ;
        RECT 1179.310 600.000 1179.590 600.030 ;
        RECT 1175.460 596.630 1177.440 596.770 ;
        RECT 1175.460 569.570 1175.600 596.630 ;
        RECT 1173.620 569.430 1175.600 569.570 ;
        RECT 1173.620 500.210 1173.760 569.430 ;
        RECT 1173.620 500.070 1174.680 500.210 ;
        RECT 1174.540 496.130 1174.680 500.070 ;
        RECT 1174.080 495.990 1174.680 496.130 ;
        RECT 1174.080 400.850 1174.220 495.990 ;
        RECT 1174.020 400.530 1174.280 400.850 ;
        RECT 1173.560 400.190 1173.820 400.510 ;
        RECT 1173.620 351.970 1173.760 400.190 ;
        RECT 1173.160 351.830 1173.760 351.970 ;
        RECT 1173.160 351.290 1173.300 351.830 ;
        RECT 1173.160 351.150 1173.760 351.290 ;
        RECT 1173.620 255.410 1173.760 351.150 ;
        RECT 1173.160 255.270 1173.760 255.410 ;
        RECT 1173.160 254.730 1173.300 255.270 ;
        RECT 1173.160 254.590 1173.760 254.730 ;
        RECT 1173.620 158.850 1173.760 254.590 ;
        RECT 1173.160 158.710 1173.760 158.850 ;
        RECT 1173.160 158.170 1173.300 158.710 ;
        RECT 1173.160 158.030 1173.760 158.170 ;
        RECT 1173.620 62.290 1173.760 158.030 ;
        RECT 1173.160 62.150 1173.760 62.290 ;
        RECT 1173.160 23.110 1173.300 62.150 ;
        RECT 1014.860 22.790 1015.120 23.110 ;
        RECT 1173.100 22.790 1173.360 23.110 ;
        RECT 1014.920 14.950 1015.060 22.790 ;
        RECT 990.020 14.630 990.280 14.950 ;
        RECT 1014.860 14.630 1015.120 14.950 ;
        RECT 990.080 2.400 990.220 14.630 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1014.370 23.700 1014.690 23.760 ;
        RECT 1187.330 23.700 1187.650 23.760 ;
        RECT 1014.370 23.560 1187.650 23.700 ;
        RECT 1014.370 23.500 1014.690 23.560 ;
        RECT 1187.330 23.500 1187.650 23.560 ;
        RECT 1007.470 15.880 1007.790 15.940 ;
        RECT 1014.370 15.880 1014.690 15.940 ;
        RECT 1007.470 15.740 1014.690 15.880 ;
        RECT 1007.470 15.680 1007.790 15.740 ;
        RECT 1014.370 15.680 1014.690 15.740 ;
      LAYER via ;
        RECT 1014.400 23.500 1014.660 23.760 ;
        RECT 1187.360 23.500 1187.620 23.760 ;
        RECT 1007.500 15.680 1007.760 15.940 ;
        RECT 1014.400 15.680 1014.660 15.940 ;
      LAYER met2 ;
        RECT 1188.510 600.170 1188.790 604.000 ;
        RECT 1187.420 600.030 1188.790 600.170 ;
        RECT 1187.420 23.790 1187.560 600.030 ;
        RECT 1188.510 600.000 1188.790 600.030 ;
        RECT 1014.400 23.470 1014.660 23.790 ;
        RECT 1187.360 23.470 1187.620 23.790 ;
        RECT 1014.460 15.970 1014.600 23.470 ;
        RECT 1007.500 15.650 1007.760 15.970 ;
        RECT 1014.400 15.650 1014.660 15.970 ;
        RECT 1007.560 2.400 1007.700 15.650 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1194.690 572.460 1195.010 572.520 ;
        RECT 1195.610 572.460 1195.930 572.520 ;
        RECT 1194.690 572.320 1195.930 572.460 ;
        RECT 1194.690 572.260 1195.010 572.320 ;
        RECT 1195.610 572.260 1195.930 572.320 ;
        RECT 1194.230 524.520 1194.550 524.580 ;
        RECT 1195.610 524.520 1195.930 524.580 ;
        RECT 1194.230 524.380 1195.930 524.520 ;
        RECT 1194.230 524.320 1194.550 524.380 ;
        RECT 1195.610 524.320 1195.930 524.380 ;
        RECT 1194.690 337.860 1195.010 337.920 ;
        RECT 1195.610 337.860 1195.930 337.920 ;
        RECT 1194.690 337.720 1195.930 337.860 ;
        RECT 1194.690 337.660 1195.010 337.720 ;
        RECT 1195.610 337.660 1195.930 337.720 ;
        RECT 1194.690 289.920 1195.010 289.980 ;
        RECT 1195.610 289.920 1195.930 289.980 ;
        RECT 1194.690 289.780 1195.930 289.920 ;
        RECT 1194.690 289.720 1195.010 289.780 ;
        RECT 1195.610 289.720 1195.930 289.780 ;
        RECT 1194.690 120.940 1195.010 121.000 ;
        RECT 1195.610 120.940 1195.930 121.000 ;
        RECT 1194.690 120.800 1195.930 120.940 ;
        RECT 1194.690 120.740 1195.010 120.800 ;
        RECT 1195.610 120.740 1195.930 120.800 ;
        RECT 1194.690 96.800 1195.010 96.860 ;
        RECT 1195.610 96.800 1195.930 96.860 ;
        RECT 1194.690 96.660 1195.930 96.800 ;
        RECT 1194.690 96.600 1195.010 96.660 ;
        RECT 1195.610 96.600 1195.930 96.660 ;
        RECT 1025.410 23.360 1025.730 23.420 ;
        RECT 1194.690 23.360 1195.010 23.420 ;
        RECT 1025.410 23.220 1195.010 23.360 ;
        RECT 1025.410 23.160 1025.730 23.220 ;
        RECT 1194.690 23.160 1195.010 23.220 ;
      LAYER via ;
        RECT 1194.720 572.260 1194.980 572.520 ;
        RECT 1195.640 572.260 1195.900 572.520 ;
        RECT 1194.260 524.320 1194.520 524.580 ;
        RECT 1195.640 524.320 1195.900 524.580 ;
        RECT 1194.720 337.660 1194.980 337.920 ;
        RECT 1195.640 337.660 1195.900 337.920 ;
        RECT 1194.720 289.720 1194.980 289.980 ;
        RECT 1195.640 289.720 1195.900 289.980 ;
        RECT 1194.720 120.740 1194.980 121.000 ;
        RECT 1195.640 120.740 1195.900 121.000 ;
        RECT 1194.720 96.600 1194.980 96.860 ;
        RECT 1195.640 96.600 1195.900 96.860 ;
        RECT 1025.440 23.160 1025.700 23.420 ;
        RECT 1194.720 23.160 1194.980 23.420 ;
      LAYER met2 ;
        RECT 1197.710 600.170 1197.990 604.000 ;
        RECT 1195.700 600.030 1197.990 600.170 ;
        RECT 1195.700 596.770 1195.840 600.030 ;
        RECT 1197.710 600.000 1197.990 600.030 ;
        RECT 1194.780 596.630 1195.840 596.770 ;
        RECT 1194.780 572.550 1194.920 596.630 ;
        RECT 1194.720 572.230 1194.980 572.550 ;
        RECT 1195.640 572.230 1195.900 572.550 ;
        RECT 1195.700 524.610 1195.840 572.230 ;
        RECT 1194.260 524.290 1194.520 524.610 ;
        RECT 1195.640 524.290 1195.900 524.610 ;
        RECT 1194.320 524.010 1194.460 524.290 ;
        RECT 1194.320 523.870 1194.920 524.010 ;
        RECT 1194.780 400.930 1194.920 523.870 ;
        RECT 1194.320 400.790 1194.920 400.930 ;
        RECT 1194.320 400.250 1194.460 400.790 ;
        RECT 1194.320 400.110 1194.920 400.250 ;
        RECT 1194.780 337.950 1194.920 400.110 ;
        RECT 1194.720 337.630 1194.980 337.950 ;
        RECT 1195.640 337.630 1195.900 337.950 ;
        RECT 1195.700 290.010 1195.840 337.630 ;
        RECT 1194.720 289.690 1194.980 290.010 ;
        RECT 1195.640 289.690 1195.900 290.010 ;
        RECT 1194.780 207.130 1194.920 289.690 ;
        RECT 1194.320 206.990 1194.920 207.130 ;
        RECT 1194.320 206.450 1194.460 206.990 ;
        RECT 1194.320 206.310 1194.920 206.450 ;
        RECT 1194.780 121.030 1194.920 206.310 ;
        RECT 1194.720 120.710 1194.980 121.030 ;
        RECT 1195.640 120.710 1195.900 121.030 ;
        RECT 1195.700 96.890 1195.840 120.710 ;
        RECT 1194.720 96.570 1194.980 96.890 ;
        RECT 1195.640 96.570 1195.900 96.890 ;
        RECT 1194.780 23.450 1194.920 96.570 ;
        RECT 1025.440 23.130 1025.700 23.450 ;
        RECT 1194.720 23.130 1194.980 23.450 ;
        RECT 1025.500 2.400 1025.640 23.130 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1201.130 496.780 1201.450 497.040 ;
        RECT 1200.670 496.640 1200.990 496.700 ;
        RECT 1201.220 496.640 1201.360 496.780 ;
        RECT 1200.670 496.500 1201.360 496.640 ;
        RECT 1200.670 496.440 1200.990 496.500 ;
        RECT 1200.670 476.240 1200.990 476.300 ;
        RECT 1201.590 476.240 1201.910 476.300 ;
        RECT 1200.670 476.100 1201.910 476.240 ;
        RECT 1200.670 476.040 1200.990 476.100 ;
        RECT 1201.590 476.040 1201.910 476.100 ;
        RECT 1201.590 400.760 1201.910 400.820 ;
        RECT 1201.220 400.620 1201.910 400.760 ;
        RECT 1201.220 400.480 1201.360 400.620 ;
        RECT 1201.590 400.560 1201.910 400.620 ;
        RECT 1201.130 400.220 1201.450 400.480 ;
        RECT 1043.350 24.040 1043.670 24.100 ;
        RECT 1200.670 24.040 1200.990 24.100 ;
        RECT 1043.350 23.900 1200.990 24.040 ;
        RECT 1043.350 23.840 1043.670 23.900 ;
        RECT 1200.670 23.840 1200.990 23.900 ;
      LAYER via ;
        RECT 1201.160 496.780 1201.420 497.040 ;
        RECT 1200.700 496.440 1200.960 496.700 ;
        RECT 1200.700 476.040 1200.960 476.300 ;
        RECT 1201.620 476.040 1201.880 476.300 ;
        RECT 1201.620 400.560 1201.880 400.820 ;
        RECT 1201.160 400.220 1201.420 400.480 ;
        RECT 1043.380 23.840 1043.640 24.100 ;
        RECT 1200.700 23.840 1200.960 24.100 ;
      LAYER met2 ;
        RECT 1206.910 600.170 1207.190 604.000 ;
        RECT 1204.440 600.030 1207.190 600.170 ;
        RECT 1204.440 593.370 1204.580 600.030 ;
        RECT 1206.910 600.000 1207.190 600.030 ;
        RECT 1203.060 593.230 1204.580 593.370 ;
        RECT 1203.060 569.570 1203.200 593.230 ;
        RECT 1201.220 569.430 1203.200 569.570 ;
        RECT 1201.220 497.070 1201.360 569.430 ;
        RECT 1201.160 496.750 1201.420 497.070 ;
        RECT 1200.700 496.410 1200.960 496.730 ;
        RECT 1200.760 476.330 1200.900 496.410 ;
        RECT 1200.700 476.010 1200.960 476.330 ;
        RECT 1201.620 476.010 1201.880 476.330 ;
        RECT 1201.680 400.850 1201.820 476.010 ;
        RECT 1201.620 400.530 1201.880 400.850 ;
        RECT 1201.160 400.190 1201.420 400.510 ;
        RECT 1201.220 351.970 1201.360 400.190 ;
        RECT 1200.760 351.830 1201.360 351.970 ;
        RECT 1200.760 351.290 1200.900 351.830 ;
        RECT 1200.760 351.150 1201.360 351.290 ;
        RECT 1201.220 255.410 1201.360 351.150 ;
        RECT 1200.760 255.270 1201.360 255.410 ;
        RECT 1200.760 254.730 1200.900 255.270 ;
        RECT 1200.760 254.590 1201.360 254.730 ;
        RECT 1201.220 158.850 1201.360 254.590 ;
        RECT 1200.760 158.710 1201.360 158.850 ;
        RECT 1200.760 158.170 1200.900 158.710 ;
        RECT 1200.760 158.030 1201.360 158.170 ;
        RECT 1201.220 62.290 1201.360 158.030 ;
        RECT 1200.760 62.150 1201.360 62.290 ;
        RECT 1200.760 24.130 1200.900 62.150 ;
        RECT 1043.380 23.810 1043.640 24.130 ;
        RECT 1200.700 23.810 1200.960 24.130 ;
        RECT 1043.440 2.400 1043.580 23.810 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1061.290 24.380 1061.610 24.440 ;
        RECT 1214.930 24.380 1215.250 24.440 ;
        RECT 1061.290 24.240 1215.250 24.380 ;
        RECT 1061.290 24.180 1061.610 24.240 ;
        RECT 1214.930 24.180 1215.250 24.240 ;
      LAYER via ;
        RECT 1061.320 24.180 1061.580 24.440 ;
        RECT 1214.960 24.180 1215.220 24.440 ;
      LAYER met2 ;
        RECT 1216.110 600.170 1216.390 604.000 ;
        RECT 1215.020 600.030 1216.390 600.170 ;
        RECT 1215.020 24.470 1215.160 600.030 ;
        RECT 1216.110 600.000 1216.390 600.030 ;
        RECT 1061.320 24.150 1061.580 24.470 ;
        RECT 1214.960 24.150 1215.220 24.470 ;
        RECT 1061.380 2.400 1061.520 24.150 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1222.290 545.400 1222.610 545.660 ;
        RECT 1222.380 544.980 1222.520 545.400 ;
        RECT 1222.290 544.720 1222.610 544.980 ;
        RECT 1222.290 531.320 1222.610 531.380 ;
        RECT 1222.750 531.320 1223.070 531.380 ;
        RECT 1222.290 531.180 1223.070 531.320 ;
        RECT 1222.290 531.120 1222.610 531.180 ;
        RECT 1222.750 531.120 1223.070 531.180 ;
        RECT 1221.830 303.520 1222.150 303.580 ;
        RECT 1222.750 303.520 1223.070 303.580 ;
        RECT 1221.830 303.380 1223.070 303.520 ;
        RECT 1221.830 303.320 1222.150 303.380 ;
        RECT 1222.750 303.320 1223.070 303.380 ;
        RECT 1221.370 193.360 1221.690 193.420 ;
        RECT 1222.750 193.360 1223.070 193.420 ;
        RECT 1221.370 193.220 1223.070 193.360 ;
        RECT 1221.370 193.160 1221.690 193.220 ;
        RECT 1222.750 193.160 1223.070 193.220 ;
        RECT 1221.830 110.400 1222.150 110.460 ;
        RECT 1222.750 110.400 1223.070 110.460 ;
        RECT 1221.830 110.260 1223.070 110.400 ;
        RECT 1221.830 110.200 1222.150 110.260 ;
        RECT 1222.750 110.200 1223.070 110.260 ;
        RECT 1079.230 24.720 1079.550 24.780 ;
        RECT 1222.750 24.720 1223.070 24.780 ;
        RECT 1079.230 24.580 1223.070 24.720 ;
        RECT 1079.230 24.520 1079.550 24.580 ;
        RECT 1222.750 24.520 1223.070 24.580 ;
      LAYER via ;
        RECT 1222.320 545.400 1222.580 545.660 ;
        RECT 1222.320 544.720 1222.580 544.980 ;
        RECT 1222.320 531.120 1222.580 531.380 ;
        RECT 1222.780 531.120 1223.040 531.380 ;
        RECT 1221.860 303.320 1222.120 303.580 ;
        RECT 1222.780 303.320 1223.040 303.580 ;
        RECT 1221.400 193.160 1221.660 193.420 ;
        RECT 1222.780 193.160 1223.040 193.420 ;
        RECT 1221.860 110.200 1222.120 110.460 ;
        RECT 1222.780 110.200 1223.040 110.460 ;
        RECT 1079.260 24.520 1079.520 24.780 ;
        RECT 1222.780 24.520 1223.040 24.780 ;
      LAYER met2 ;
        RECT 1225.310 600.170 1225.590 604.000 ;
        RECT 1222.840 600.030 1225.590 600.170 ;
        RECT 1222.840 596.770 1222.980 600.030 ;
        RECT 1225.310 600.000 1225.590 600.030 ;
        RECT 1222.380 596.630 1222.980 596.770 ;
        RECT 1222.380 545.690 1222.520 596.630 ;
        RECT 1222.320 545.370 1222.580 545.690 ;
        RECT 1222.320 544.690 1222.580 545.010 ;
        RECT 1222.380 531.410 1222.520 544.690 ;
        RECT 1222.320 531.090 1222.580 531.410 ;
        RECT 1222.780 531.090 1223.040 531.410 ;
        RECT 1222.840 496.810 1222.980 531.090 ;
        RECT 1222.380 496.670 1222.980 496.810 ;
        RECT 1222.380 410.450 1222.520 496.670 ;
        RECT 1221.460 410.310 1222.520 410.450 ;
        RECT 1221.460 351.290 1221.600 410.310 ;
        RECT 1221.460 351.150 1222.060 351.290 ;
        RECT 1221.920 303.610 1222.060 351.150 ;
        RECT 1221.860 303.290 1222.120 303.610 ;
        RECT 1222.780 303.290 1223.040 303.610 ;
        RECT 1222.840 253.370 1222.980 303.290 ;
        RECT 1222.840 253.230 1223.440 253.370 ;
        RECT 1223.300 252.010 1223.440 253.230 ;
        RECT 1222.840 251.870 1223.440 252.010 ;
        RECT 1222.840 193.450 1222.980 251.870 ;
        RECT 1221.400 193.130 1221.660 193.450 ;
        RECT 1222.780 193.130 1223.040 193.450 ;
        RECT 1221.460 192.850 1221.600 193.130 ;
        RECT 1221.460 192.710 1222.060 192.850 ;
        RECT 1221.920 110.490 1222.060 192.710 ;
        RECT 1221.860 110.170 1222.120 110.490 ;
        RECT 1222.780 110.170 1223.040 110.490 ;
        RECT 1222.840 24.810 1222.980 110.170 ;
        RECT 1079.260 24.490 1079.520 24.810 ;
        RECT 1222.780 24.490 1223.040 24.810 ;
        RECT 1079.320 2.400 1079.460 24.490 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1228.730 386.480 1229.050 386.540 ;
        RECT 1229.650 386.480 1229.970 386.540 ;
        RECT 1228.730 386.340 1229.970 386.480 ;
        RECT 1228.730 386.280 1229.050 386.340 ;
        RECT 1229.650 386.280 1229.970 386.340 ;
        RECT 1229.190 303.520 1229.510 303.580 ;
        RECT 1230.110 303.520 1230.430 303.580 ;
        RECT 1229.190 303.380 1230.430 303.520 ;
        RECT 1229.190 303.320 1229.510 303.380 ;
        RECT 1230.110 303.320 1230.430 303.380 ;
        RECT 1228.730 193.360 1229.050 193.420 ;
        RECT 1230.110 193.360 1230.430 193.420 ;
        RECT 1228.730 193.220 1230.430 193.360 ;
        RECT 1228.730 193.160 1229.050 193.220 ;
        RECT 1230.110 193.160 1230.430 193.220 ;
        RECT 1229.190 110.400 1229.510 110.460 ;
        RECT 1230.110 110.400 1230.430 110.460 ;
        RECT 1229.190 110.260 1230.430 110.400 ;
        RECT 1229.190 110.200 1229.510 110.260 ;
        RECT 1230.110 110.200 1230.430 110.260 ;
        RECT 1096.710 25.060 1097.030 25.120 ;
        RECT 1230.110 25.060 1230.430 25.120 ;
        RECT 1096.710 24.920 1230.430 25.060 ;
        RECT 1096.710 24.860 1097.030 24.920 ;
        RECT 1230.110 24.860 1230.430 24.920 ;
      LAYER via ;
        RECT 1228.760 386.280 1229.020 386.540 ;
        RECT 1229.680 386.280 1229.940 386.540 ;
        RECT 1229.220 303.320 1229.480 303.580 ;
        RECT 1230.140 303.320 1230.400 303.580 ;
        RECT 1228.760 193.160 1229.020 193.420 ;
        RECT 1230.140 193.160 1230.400 193.420 ;
        RECT 1229.220 110.200 1229.480 110.460 ;
        RECT 1230.140 110.200 1230.400 110.460 ;
        RECT 1096.740 24.860 1097.000 25.120 ;
        RECT 1230.140 24.860 1230.400 25.120 ;
      LAYER met2 ;
        RECT 1234.510 600.170 1234.790 604.000 ;
        RECT 1232.500 600.030 1234.790 600.170 ;
        RECT 1232.500 596.770 1232.640 600.030 ;
        RECT 1234.510 600.000 1234.790 600.030 ;
        RECT 1230.200 596.630 1232.640 596.770 ;
        RECT 1230.200 569.570 1230.340 596.630 ;
        RECT 1229.740 569.430 1230.340 569.570 ;
        RECT 1229.740 386.570 1229.880 569.430 ;
        RECT 1228.760 386.250 1229.020 386.570 ;
        RECT 1229.680 386.250 1229.940 386.570 ;
        RECT 1228.820 351.290 1228.960 386.250 ;
        RECT 1228.820 351.150 1229.420 351.290 ;
        RECT 1229.280 303.610 1229.420 351.150 ;
        RECT 1229.220 303.290 1229.480 303.610 ;
        RECT 1230.140 303.290 1230.400 303.610 ;
        RECT 1230.200 253.370 1230.340 303.290 ;
        RECT 1230.200 253.230 1230.800 253.370 ;
        RECT 1230.660 252.010 1230.800 253.230 ;
        RECT 1230.200 251.870 1230.800 252.010 ;
        RECT 1230.200 193.450 1230.340 251.870 ;
        RECT 1228.760 193.130 1229.020 193.450 ;
        RECT 1230.140 193.130 1230.400 193.450 ;
        RECT 1228.820 192.850 1228.960 193.130 ;
        RECT 1228.820 192.710 1229.420 192.850 ;
        RECT 1229.280 110.490 1229.420 192.710 ;
        RECT 1229.220 110.170 1229.480 110.490 ;
        RECT 1230.140 110.170 1230.400 110.490 ;
        RECT 1230.200 60.250 1230.340 110.170 ;
        RECT 1230.200 60.110 1230.800 60.250 ;
        RECT 1230.660 58.890 1230.800 60.110 ;
        RECT 1230.200 58.750 1230.800 58.890 ;
        RECT 1230.200 25.150 1230.340 58.750 ;
        RECT 1096.740 24.830 1097.000 25.150 ;
        RECT 1230.140 24.830 1230.400 25.150 ;
        RECT 1096.800 2.400 1096.940 24.830 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1117.410 589.800 1117.730 589.860 ;
        RECT 1242.530 589.800 1242.850 589.860 ;
        RECT 1117.410 589.660 1242.850 589.800 ;
        RECT 1117.410 589.600 1117.730 589.660 ;
        RECT 1242.530 589.600 1242.850 589.660 ;
        RECT 1114.650 20.980 1114.970 21.040 ;
        RECT 1117.410 20.980 1117.730 21.040 ;
        RECT 1114.650 20.840 1117.730 20.980 ;
        RECT 1114.650 20.780 1114.970 20.840 ;
        RECT 1117.410 20.780 1117.730 20.840 ;
      LAYER via ;
        RECT 1117.440 589.600 1117.700 589.860 ;
        RECT 1242.560 589.600 1242.820 589.860 ;
        RECT 1114.680 20.780 1114.940 21.040 ;
        RECT 1117.440 20.780 1117.700 21.040 ;
      LAYER met2 ;
        RECT 1243.710 600.170 1243.990 604.000 ;
        RECT 1242.620 600.030 1243.990 600.170 ;
        RECT 1242.620 589.890 1242.760 600.030 ;
        RECT 1243.710 600.000 1243.990 600.030 ;
        RECT 1117.440 589.570 1117.700 589.890 ;
        RECT 1242.560 589.570 1242.820 589.890 ;
        RECT 1117.500 21.070 1117.640 589.570 ;
        RECT 1114.680 20.750 1114.940 21.070 ;
        RECT 1117.440 20.750 1117.700 21.070 ;
        RECT 1114.740 2.400 1114.880 20.750 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.110 591.500 1138.430 591.560 ;
        RECT 1251.270 591.500 1251.590 591.560 ;
        RECT 1138.110 591.360 1251.590 591.500 ;
        RECT 1138.110 591.300 1138.430 591.360 ;
        RECT 1251.270 591.300 1251.590 591.360 ;
        RECT 1132.590 20.640 1132.910 20.700 ;
        RECT 1138.110 20.640 1138.430 20.700 ;
        RECT 1132.590 20.500 1138.430 20.640 ;
        RECT 1132.590 20.440 1132.910 20.500 ;
        RECT 1138.110 20.440 1138.430 20.500 ;
      LAYER via ;
        RECT 1138.140 591.300 1138.400 591.560 ;
        RECT 1251.300 591.300 1251.560 591.560 ;
        RECT 1132.620 20.440 1132.880 20.700 ;
        RECT 1138.140 20.440 1138.400 20.700 ;
      LAYER met2 ;
        RECT 1252.910 600.170 1253.190 604.000 ;
        RECT 1251.360 600.030 1253.190 600.170 ;
        RECT 1251.360 591.590 1251.500 600.030 ;
        RECT 1252.910 600.000 1253.190 600.030 ;
        RECT 1138.140 591.270 1138.400 591.590 ;
        RECT 1251.300 591.270 1251.560 591.590 ;
        RECT 1138.200 20.730 1138.340 591.270 ;
        RECT 1132.620 20.410 1132.880 20.730 ;
        RECT 1138.140 20.410 1138.400 20.730 ;
        RECT 1132.680 2.400 1132.820 20.410 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.990 591.160 1197.310 591.220 ;
        RECT 1260.470 591.160 1260.790 591.220 ;
        RECT 1196.990 591.020 1260.790 591.160 ;
        RECT 1196.990 590.960 1197.310 591.020 ;
        RECT 1260.470 590.960 1260.790 591.020 ;
        RECT 1196.990 587.760 1197.310 587.820 ;
        RECT 1189.720 587.620 1197.310 587.760 ;
        RECT 1151.910 587.420 1152.230 587.480 ;
        RECT 1189.720 587.420 1189.860 587.620 ;
        RECT 1196.990 587.560 1197.310 587.620 ;
        RECT 1151.910 587.280 1189.860 587.420 ;
        RECT 1151.910 587.220 1152.230 587.280 ;
        RECT 1150.990 289.580 1151.310 289.640 ;
        RECT 1151.910 289.580 1152.230 289.640 ;
        RECT 1150.990 289.440 1152.230 289.580 ;
        RECT 1150.990 289.380 1151.310 289.440 ;
        RECT 1151.910 289.380 1152.230 289.440 ;
        RECT 1150.990 241.980 1151.310 242.040 ;
        RECT 1151.910 241.980 1152.230 242.040 ;
        RECT 1150.990 241.840 1152.230 241.980 ;
        RECT 1150.990 241.780 1151.310 241.840 ;
        RECT 1151.910 241.780 1152.230 241.840 ;
        RECT 1151.910 193.500 1152.230 193.760 ;
        RECT 1152.000 193.080 1152.140 193.500 ;
        RECT 1151.910 192.820 1152.230 193.080 ;
        RECT 1151.910 179.760 1152.230 179.820 ;
        RECT 1152.370 179.760 1152.690 179.820 ;
        RECT 1151.910 179.620 1152.690 179.760 ;
        RECT 1151.910 179.560 1152.230 179.620 ;
        RECT 1152.370 179.560 1152.690 179.620 ;
        RECT 1151.910 145.080 1152.230 145.140 ;
        RECT 1152.370 145.080 1152.690 145.140 ;
        RECT 1151.910 144.940 1152.690 145.080 ;
        RECT 1151.910 144.880 1152.230 144.940 ;
        RECT 1152.370 144.880 1152.690 144.940 ;
        RECT 1151.910 62.460 1152.230 62.520 ;
        RECT 1150.620 62.320 1152.230 62.460 ;
        RECT 1150.620 62.180 1150.760 62.320 ;
        RECT 1151.910 62.260 1152.230 62.320 ;
        RECT 1150.530 61.920 1150.850 62.180 ;
      LAYER via ;
        RECT 1197.020 590.960 1197.280 591.220 ;
        RECT 1260.500 590.960 1260.760 591.220 ;
        RECT 1151.940 587.220 1152.200 587.480 ;
        RECT 1197.020 587.560 1197.280 587.820 ;
        RECT 1151.020 289.380 1151.280 289.640 ;
        RECT 1151.940 289.380 1152.200 289.640 ;
        RECT 1151.020 241.780 1151.280 242.040 ;
        RECT 1151.940 241.780 1152.200 242.040 ;
        RECT 1151.940 193.500 1152.200 193.760 ;
        RECT 1151.940 192.820 1152.200 193.080 ;
        RECT 1151.940 179.560 1152.200 179.820 ;
        RECT 1152.400 179.560 1152.660 179.820 ;
        RECT 1151.940 144.880 1152.200 145.140 ;
        RECT 1152.400 144.880 1152.660 145.140 ;
        RECT 1151.940 62.260 1152.200 62.520 ;
        RECT 1150.560 61.920 1150.820 62.180 ;
      LAYER met2 ;
        RECT 1262.110 600.170 1262.390 604.000 ;
        RECT 1260.560 600.030 1262.390 600.170 ;
        RECT 1260.560 591.250 1260.700 600.030 ;
        RECT 1262.110 600.000 1262.390 600.030 ;
        RECT 1197.020 590.930 1197.280 591.250 ;
        RECT 1260.500 590.930 1260.760 591.250 ;
        RECT 1197.080 587.850 1197.220 590.930 ;
        RECT 1197.020 587.530 1197.280 587.850 ;
        RECT 1151.940 587.190 1152.200 587.510 ;
        RECT 1152.000 435.725 1152.140 587.190 ;
        RECT 1151.930 435.355 1152.210 435.725 ;
        RECT 1151.930 434.675 1152.210 435.045 ;
        RECT 1152.000 339.050 1152.140 434.675 ;
        RECT 1152.000 338.910 1152.600 339.050 ;
        RECT 1152.460 338.370 1152.600 338.910 ;
        RECT 1152.000 338.230 1152.600 338.370 ;
        RECT 1152.000 289.670 1152.140 338.230 ;
        RECT 1151.020 289.350 1151.280 289.670 ;
        RECT 1151.940 289.350 1152.200 289.670 ;
        RECT 1151.080 242.070 1151.220 289.350 ;
        RECT 1151.020 241.750 1151.280 242.070 ;
        RECT 1151.940 241.750 1152.200 242.070 ;
        RECT 1152.000 193.790 1152.140 241.750 ;
        RECT 1151.940 193.470 1152.200 193.790 ;
        RECT 1151.940 192.790 1152.200 193.110 ;
        RECT 1152.000 179.850 1152.140 192.790 ;
        RECT 1151.940 179.530 1152.200 179.850 ;
        RECT 1152.400 179.530 1152.660 179.850 ;
        RECT 1152.460 145.170 1152.600 179.530 ;
        RECT 1151.940 144.850 1152.200 145.170 ;
        RECT 1152.400 144.850 1152.660 145.170 ;
        RECT 1152.000 62.550 1152.140 144.850 ;
        RECT 1151.940 62.230 1152.200 62.550 ;
        RECT 1150.560 61.890 1150.820 62.210 ;
        RECT 1150.620 2.400 1150.760 61.890 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
      LAYER via2 ;
        RECT 1151.930 435.400 1152.210 435.680 ;
        RECT 1151.930 434.720 1152.210 435.000 ;
      LAYER met3 ;
        RECT 1151.905 435.690 1152.235 435.705 ;
        RECT 1151.905 435.375 1152.450 435.690 ;
        RECT 1152.150 435.025 1152.450 435.375 ;
        RECT 1151.905 434.710 1152.450 435.025 ;
        RECT 1151.905 434.695 1152.235 434.710 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 41.380 669.230 41.440 ;
        RECT 1015.290 41.380 1015.610 41.440 ;
        RECT 668.910 41.240 1015.610 41.380 ;
        RECT 668.910 41.180 669.230 41.240 ;
        RECT 1015.290 41.180 1015.610 41.240 ;
      LAYER via ;
        RECT 668.940 41.180 669.200 41.440 ;
        RECT 1015.320 41.180 1015.580 41.440 ;
      LAYER met2 ;
        RECT 1014.170 600.170 1014.450 604.000 ;
        RECT 1014.170 600.030 1015.520 600.170 ;
        RECT 1014.170 600.000 1014.450 600.030 ;
        RECT 1015.380 41.470 1015.520 600.030 ;
        RECT 668.940 41.150 669.200 41.470 ;
        RECT 1015.320 41.150 1015.580 41.470 ;
        RECT 669.000 2.400 669.140 41.150 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1172.610 592.180 1172.930 592.240 ;
        RECT 1269.670 592.180 1269.990 592.240 ;
        RECT 1172.610 592.040 1269.990 592.180 ;
        RECT 1172.610 591.980 1172.930 592.040 ;
        RECT 1269.670 591.980 1269.990 592.040 ;
        RECT 1168.470 20.640 1168.790 20.700 ;
        RECT 1172.610 20.640 1172.930 20.700 ;
        RECT 1168.470 20.500 1172.930 20.640 ;
        RECT 1168.470 20.440 1168.790 20.500 ;
        RECT 1172.610 20.440 1172.930 20.500 ;
      LAYER via ;
        RECT 1172.640 591.980 1172.900 592.240 ;
        RECT 1269.700 591.980 1269.960 592.240 ;
        RECT 1168.500 20.440 1168.760 20.700 ;
        RECT 1172.640 20.440 1172.900 20.700 ;
      LAYER met2 ;
        RECT 1271.310 600.170 1271.590 604.000 ;
        RECT 1269.760 600.030 1271.590 600.170 ;
        RECT 1269.760 592.270 1269.900 600.030 ;
        RECT 1271.310 600.000 1271.590 600.030 ;
        RECT 1172.640 591.950 1172.900 592.270 ;
        RECT 1269.700 591.950 1269.960 592.270 ;
        RECT 1172.700 20.730 1172.840 591.950 ;
        RECT 1168.500 20.410 1168.760 20.730 ;
        RECT 1172.640 20.410 1172.900 20.730 ;
        RECT 1168.560 2.400 1168.700 20.410 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 589.460 1186.730 589.520 ;
        RECT 1278.870 589.460 1279.190 589.520 ;
        RECT 1186.410 589.320 1279.190 589.460 ;
        RECT 1186.410 589.260 1186.730 589.320 ;
        RECT 1278.870 589.260 1279.190 589.320 ;
        RECT 1184.570 96.460 1184.890 96.520 ;
        RECT 1186.410 96.460 1186.730 96.520 ;
        RECT 1184.570 96.320 1186.730 96.460 ;
        RECT 1184.570 96.260 1184.890 96.320 ;
        RECT 1186.410 96.260 1186.730 96.320 ;
        RECT 1184.570 48.520 1184.890 48.580 ;
        RECT 1185.490 48.520 1185.810 48.580 ;
        RECT 1184.570 48.380 1185.810 48.520 ;
        RECT 1184.570 48.320 1184.890 48.380 ;
        RECT 1185.490 48.320 1185.810 48.380 ;
      LAYER via ;
        RECT 1186.440 589.260 1186.700 589.520 ;
        RECT 1278.900 589.260 1279.160 589.520 ;
        RECT 1184.600 96.260 1184.860 96.520 ;
        RECT 1186.440 96.260 1186.700 96.520 ;
        RECT 1184.600 48.320 1184.860 48.580 ;
        RECT 1185.520 48.320 1185.780 48.580 ;
      LAYER met2 ;
        RECT 1280.510 600.170 1280.790 604.000 ;
        RECT 1278.960 600.030 1280.790 600.170 ;
        RECT 1278.960 589.550 1279.100 600.030 ;
        RECT 1280.510 600.000 1280.790 600.030 ;
        RECT 1186.440 589.230 1186.700 589.550 ;
        RECT 1278.900 589.230 1279.160 589.550 ;
        RECT 1186.500 96.550 1186.640 589.230 ;
        RECT 1184.600 96.230 1184.860 96.550 ;
        RECT 1186.440 96.230 1186.700 96.550 ;
        RECT 1184.660 48.610 1184.800 96.230 ;
        RECT 1184.600 48.290 1184.860 48.610 ;
        RECT 1185.520 48.290 1185.780 48.610 ;
        RECT 1185.580 48.125 1185.720 48.290 ;
        RECT 1185.510 47.755 1185.790 48.125 ;
        RECT 1186.430 47.755 1186.710 48.125 ;
        RECT 1186.500 21.490 1186.640 47.755 ;
        RECT 1186.040 21.350 1186.640 21.490 ;
        RECT 1186.040 2.400 1186.180 21.350 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
      LAYER via2 ;
        RECT 1185.510 47.800 1185.790 48.080 ;
        RECT 1186.430 47.800 1186.710 48.080 ;
      LAYER met3 ;
        RECT 1185.485 48.090 1185.815 48.105 ;
        RECT 1186.405 48.090 1186.735 48.105 ;
        RECT 1185.485 47.790 1186.735 48.090 ;
        RECT 1185.485 47.775 1185.815 47.790 ;
        RECT 1186.405 47.775 1186.735 47.790 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.110 587.760 1207.430 587.820 ;
        RECT 1288.070 587.760 1288.390 587.820 ;
        RECT 1207.110 587.620 1288.390 587.760 ;
        RECT 1207.110 587.560 1207.430 587.620 ;
        RECT 1288.070 587.560 1288.390 587.620 ;
        RECT 1203.890 20.640 1204.210 20.700 ;
        RECT 1207.110 20.640 1207.430 20.700 ;
        RECT 1203.890 20.500 1207.430 20.640 ;
        RECT 1203.890 20.440 1204.210 20.500 ;
        RECT 1207.110 20.440 1207.430 20.500 ;
      LAYER via ;
        RECT 1207.140 587.560 1207.400 587.820 ;
        RECT 1288.100 587.560 1288.360 587.820 ;
        RECT 1203.920 20.440 1204.180 20.700 ;
        RECT 1207.140 20.440 1207.400 20.700 ;
      LAYER met2 ;
        RECT 1289.710 600.170 1289.990 604.000 ;
        RECT 1288.160 600.030 1289.990 600.170 ;
        RECT 1288.160 587.850 1288.300 600.030 ;
        RECT 1289.710 600.000 1289.990 600.030 ;
        RECT 1207.140 587.530 1207.400 587.850 ;
        RECT 1288.100 587.530 1288.360 587.850 ;
        RECT 1207.200 20.730 1207.340 587.530 ;
        RECT 1203.920 20.410 1204.180 20.730 ;
        RECT 1207.140 20.410 1207.400 20.730 ;
        RECT 1203.980 2.400 1204.120 20.410 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1227.350 588.780 1227.670 588.840 ;
        RECT 1297.270 588.780 1297.590 588.840 ;
        RECT 1227.350 588.640 1297.590 588.780 ;
        RECT 1227.350 588.580 1227.670 588.640 ;
        RECT 1297.270 588.580 1297.590 588.640 ;
        RECT 1221.830 16.560 1222.150 16.620 ;
        RECT 1227.350 16.560 1227.670 16.620 ;
        RECT 1221.830 16.420 1227.670 16.560 ;
        RECT 1221.830 16.360 1222.150 16.420 ;
        RECT 1227.350 16.360 1227.670 16.420 ;
      LAYER via ;
        RECT 1227.380 588.580 1227.640 588.840 ;
        RECT 1297.300 588.580 1297.560 588.840 ;
        RECT 1221.860 16.360 1222.120 16.620 ;
        RECT 1227.380 16.360 1227.640 16.620 ;
      LAYER met2 ;
        RECT 1298.910 600.170 1299.190 604.000 ;
        RECT 1297.360 600.030 1299.190 600.170 ;
        RECT 1297.360 588.870 1297.500 600.030 ;
        RECT 1298.910 600.000 1299.190 600.030 ;
        RECT 1227.380 588.550 1227.640 588.870 ;
        RECT 1297.300 588.550 1297.560 588.870 ;
        RECT 1227.440 16.650 1227.580 588.550 ;
        RECT 1221.860 16.330 1222.120 16.650 ;
        RECT 1227.380 16.330 1227.640 16.650 ;
        RECT 1221.920 2.400 1222.060 16.330 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.610 590.480 1241.930 590.540 ;
        RECT 1306.470 590.480 1306.790 590.540 ;
        RECT 1241.610 590.340 1306.790 590.480 ;
        RECT 1241.610 590.280 1241.930 590.340 ;
        RECT 1306.470 590.280 1306.790 590.340 ;
        RECT 1241.150 579.600 1241.470 579.660 ;
        RECT 1241.610 579.600 1241.930 579.660 ;
        RECT 1241.150 579.460 1241.930 579.600 ;
        RECT 1241.150 579.400 1241.470 579.460 ;
        RECT 1241.610 579.400 1241.930 579.460 ;
        RECT 1240.230 572.460 1240.550 572.520 ;
        RECT 1241.150 572.460 1241.470 572.520 ;
        RECT 1240.230 572.320 1241.470 572.460 ;
        RECT 1240.230 572.260 1240.550 572.320 ;
        RECT 1241.150 572.260 1241.470 572.320 ;
        RECT 1240.230 524.520 1240.550 524.580 ;
        RECT 1241.610 524.520 1241.930 524.580 ;
        RECT 1240.230 524.380 1241.930 524.520 ;
        RECT 1240.230 524.320 1240.550 524.380 ;
        RECT 1241.610 524.320 1241.930 524.380 ;
        RECT 1241.610 476.240 1241.930 476.300 ;
        RECT 1243.450 476.240 1243.770 476.300 ;
        RECT 1241.610 476.100 1243.770 476.240 ;
        RECT 1241.610 476.040 1241.930 476.100 ;
        RECT 1243.450 476.040 1243.770 476.100 ;
        RECT 1240.690 331.060 1241.010 331.120 ;
        RECT 1241.610 331.060 1241.930 331.120 ;
        RECT 1240.690 330.920 1241.930 331.060 ;
        RECT 1240.690 330.860 1241.010 330.920 ;
        RECT 1241.610 330.860 1241.930 330.920 ;
        RECT 1240.690 303.180 1241.010 303.240 ;
        RECT 1242.530 303.180 1242.850 303.240 ;
        RECT 1240.690 303.040 1242.850 303.180 ;
        RECT 1240.690 302.980 1241.010 303.040 ;
        RECT 1242.530 302.980 1242.850 303.040 ;
        RECT 1241.610 241.980 1241.930 242.040 ;
        RECT 1242.530 241.980 1242.850 242.040 ;
        RECT 1241.610 241.840 1242.850 241.980 ;
        RECT 1241.610 241.780 1241.930 241.840 ;
        RECT 1242.530 241.780 1242.850 241.840 ;
        RECT 1240.690 234.500 1241.010 234.560 ;
        RECT 1241.610 234.500 1241.930 234.560 ;
        RECT 1240.690 234.360 1241.930 234.500 ;
        RECT 1240.690 234.300 1241.010 234.360 ;
        RECT 1241.610 234.300 1241.930 234.360 ;
        RECT 1240.690 186.560 1241.010 186.620 ;
        RECT 1241.150 186.560 1241.470 186.620 ;
        RECT 1240.690 186.420 1241.470 186.560 ;
        RECT 1240.690 186.360 1241.010 186.420 ;
        RECT 1241.150 186.360 1241.470 186.420 ;
        RECT 1241.150 145.420 1241.470 145.480 ;
        RECT 1241.610 145.420 1241.930 145.480 ;
        RECT 1241.150 145.280 1241.930 145.420 ;
        RECT 1241.150 145.220 1241.470 145.280 ;
        RECT 1241.610 145.220 1241.930 145.280 ;
        RECT 1240.690 137.940 1241.010 138.000 ;
        RECT 1241.610 137.940 1241.930 138.000 ;
        RECT 1240.690 137.800 1241.930 137.940 ;
        RECT 1240.690 137.740 1241.010 137.800 ;
        RECT 1241.610 137.740 1241.930 137.800 ;
        RECT 1240.690 90.000 1241.010 90.060 ;
        RECT 1241.610 90.000 1241.930 90.060 ;
        RECT 1240.690 89.860 1241.930 90.000 ;
        RECT 1240.690 89.800 1241.010 89.860 ;
        RECT 1241.610 89.800 1241.930 89.860 ;
        RECT 1241.610 62.460 1241.930 62.520 ;
        RECT 1239.860 62.320 1241.930 62.460 ;
        RECT 1239.860 62.180 1240.000 62.320 ;
        RECT 1241.610 62.260 1241.930 62.320 ;
        RECT 1239.770 61.920 1240.090 62.180 ;
      LAYER via ;
        RECT 1241.640 590.280 1241.900 590.540 ;
        RECT 1306.500 590.280 1306.760 590.540 ;
        RECT 1241.180 579.400 1241.440 579.660 ;
        RECT 1241.640 579.400 1241.900 579.660 ;
        RECT 1240.260 572.260 1240.520 572.520 ;
        RECT 1241.180 572.260 1241.440 572.520 ;
        RECT 1240.260 524.320 1240.520 524.580 ;
        RECT 1241.640 524.320 1241.900 524.580 ;
        RECT 1241.640 476.040 1241.900 476.300 ;
        RECT 1243.480 476.040 1243.740 476.300 ;
        RECT 1240.720 330.860 1240.980 331.120 ;
        RECT 1241.640 330.860 1241.900 331.120 ;
        RECT 1240.720 302.980 1240.980 303.240 ;
        RECT 1242.560 302.980 1242.820 303.240 ;
        RECT 1241.640 241.780 1241.900 242.040 ;
        RECT 1242.560 241.780 1242.820 242.040 ;
        RECT 1240.720 234.300 1240.980 234.560 ;
        RECT 1241.640 234.300 1241.900 234.560 ;
        RECT 1240.720 186.360 1240.980 186.620 ;
        RECT 1241.180 186.360 1241.440 186.620 ;
        RECT 1241.180 145.220 1241.440 145.480 ;
        RECT 1241.640 145.220 1241.900 145.480 ;
        RECT 1240.720 137.740 1240.980 138.000 ;
        RECT 1241.640 137.740 1241.900 138.000 ;
        RECT 1240.720 89.800 1240.980 90.060 ;
        RECT 1241.640 89.800 1241.900 90.060 ;
        RECT 1241.640 62.260 1241.900 62.520 ;
        RECT 1239.800 61.920 1240.060 62.180 ;
      LAYER met2 ;
        RECT 1308.110 600.170 1308.390 604.000 ;
        RECT 1306.560 600.030 1308.390 600.170 ;
        RECT 1306.560 590.570 1306.700 600.030 ;
        RECT 1308.110 600.000 1308.390 600.030 ;
        RECT 1241.640 590.250 1241.900 590.570 ;
        RECT 1306.500 590.250 1306.760 590.570 ;
        RECT 1241.700 579.690 1241.840 590.250 ;
        RECT 1241.180 579.370 1241.440 579.690 ;
        RECT 1241.640 579.370 1241.900 579.690 ;
        RECT 1241.240 572.550 1241.380 579.370 ;
        RECT 1240.260 572.230 1240.520 572.550 ;
        RECT 1241.180 572.230 1241.440 572.550 ;
        RECT 1240.320 524.610 1240.460 572.230 ;
        RECT 1240.260 524.290 1240.520 524.610 ;
        RECT 1241.640 524.290 1241.900 524.610 ;
        RECT 1241.700 524.125 1241.840 524.290 ;
        RECT 1241.630 523.755 1241.910 524.125 ;
        RECT 1243.470 523.755 1243.750 524.125 ;
        RECT 1243.540 476.330 1243.680 523.755 ;
        RECT 1241.640 476.010 1241.900 476.330 ;
        RECT 1243.480 476.010 1243.740 476.330 ;
        RECT 1241.700 385.970 1241.840 476.010 ;
        RECT 1241.240 385.830 1241.840 385.970 ;
        RECT 1241.240 338.370 1241.380 385.830 ;
        RECT 1241.240 338.230 1241.840 338.370 ;
        RECT 1241.700 331.150 1241.840 338.230 ;
        RECT 1240.720 330.830 1240.980 331.150 ;
        RECT 1241.640 330.830 1241.900 331.150 ;
        RECT 1240.780 303.270 1240.920 330.830 ;
        RECT 1240.720 302.950 1240.980 303.270 ;
        RECT 1242.560 302.950 1242.820 303.270 ;
        RECT 1242.620 242.070 1242.760 302.950 ;
        RECT 1241.640 241.750 1241.900 242.070 ;
        RECT 1242.560 241.750 1242.820 242.070 ;
        RECT 1241.700 234.590 1241.840 241.750 ;
        RECT 1240.720 234.270 1240.980 234.590 ;
        RECT 1241.640 234.270 1241.900 234.590 ;
        RECT 1240.780 186.650 1240.920 234.270 ;
        RECT 1240.720 186.330 1240.980 186.650 ;
        RECT 1241.180 186.330 1241.440 186.650 ;
        RECT 1241.240 145.510 1241.380 186.330 ;
        RECT 1241.180 145.190 1241.440 145.510 ;
        RECT 1241.640 145.190 1241.900 145.510 ;
        RECT 1241.700 138.030 1241.840 145.190 ;
        RECT 1240.720 137.710 1240.980 138.030 ;
        RECT 1241.640 137.710 1241.900 138.030 ;
        RECT 1240.780 90.090 1240.920 137.710 ;
        RECT 1240.720 89.770 1240.980 90.090 ;
        RECT 1241.640 89.770 1241.900 90.090 ;
        RECT 1241.700 62.550 1241.840 89.770 ;
        RECT 1241.640 62.230 1241.900 62.550 ;
        RECT 1239.800 61.890 1240.060 62.210 ;
        RECT 1239.860 2.400 1240.000 61.890 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
      LAYER via2 ;
        RECT 1241.630 523.800 1241.910 524.080 ;
        RECT 1243.470 523.800 1243.750 524.080 ;
      LAYER met3 ;
        RECT 1241.605 524.090 1241.935 524.105 ;
        RECT 1243.445 524.090 1243.775 524.105 ;
        RECT 1241.605 523.790 1243.775 524.090 ;
        RECT 1241.605 523.775 1241.935 523.790 ;
        RECT 1243.445 523.775 1243.775 523.790 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 587.080 1262.630 587.140 ;
        RECT 1315.670 587.080 1315.990 587.140 ;
        RECT 1262.310 586.940 1315.990 587.080 ;
        RECT 1262.310 586.880 1262.630 586.940 ;
        RECT 1315.670 586.880 1315.990 586.940 ;
        RECT 1257.250 20.640 1257.570 20.700 ;
        RECT 1262.310 20.640 1262.630 20.700 ;
        RECT 1257.250 20.500 1262.630 20.640 ;
        RECT 1257.250 20.440 1257.570 20.500 ;
        RECT 1262.310 20.440 1262.630 20.500 ;
      LAYER via ;
        RECT 1262.340 586.880 1262.600 587.140 ;
        RECT 1315.700 586.880 1315.960 587.140 ;
        RECT 1257.280 20.440 1257.540 20.700 ;
        RECT 1262.340 20.440 1262.600 20.700 ;
      LAYER met2 ;
        RECT 1317.310 600.170 1317.590 604.000 ;
        RECT 1315.760 600.030 1317.590 600.170 ;
        RECT 1315.760 587.170 1315.900 600.030 ;
        RECT 1317.310 600.000 1317.590 600.030 ;
        RECT 1262.340 586.850 1262.600 587.170 ;
        RECT 1315.700 586.850 1315.960 587.170 ;
        RECT 1262.400 20.730 1262.540 586.850 ;
        RECT 1257.280 20.410 1257.540 20.730 ;
        RECT 1262.340 20.410 1262.600 20.730 ;
        RECT 1257.340 2.400 1257.480 20.410 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.870 590.480 1325.190 590.540 ;
        RECT 1308.400 590.340 1325.190 590.480 ;
        RECT 1276.110 590.140 1276.430 590.200 ;
        RECT 1308.400 590.140 1308.540 590.340 ;
        RECT 1324.870 590.280 1325.190 590.340 ;
        RECT 1276.110 590.000 1308.540 590.140 ;
        RECT 1276.110 589.940 1276.430 590.000 ;
      LAYER via ;
        RECT 1276.140 589.940 1276.400 590.200 ;
        RECT 1324.900 590.280 1325.160 590.540 ;
      LAYER met2 ;
        RECT 1326.510 600.170 1326.790 604.000 ;
        RECT 1324.960 600.030 1326.790 600.170 ;
        RECT 1324.960 590.570 1325.100 600.030 ;
        RECT 1326.510 600.000 1326.790 600.030 ;
        RECT 1324.900 590.250 1325.160 590.570 ;
        RECT 1276.140 589.910 1276.400 590.230 ;
        RECT 1276.200 16.730 1276.340 589.910 ;
        RECT 1275.280 16.590 1276.340 16.730 ;
        RECT 1275.280 2.400 1275.420 16.590 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 586.740 1297.130 586.800 ;
        RECT 1334.070 586.740 1334.390 586.800 ;
        RECT 1296.810 586.600 1334.390 586.740 ;
        RECT 1296.810 586.540 1297.130 586.600 ;
        RECT 1334.070 586.540 1334.390 586.600 ;
        RECT 1293.130 15.540 1293.450 15.600 ;
        RECT 1296.810 15.540 1297.130 15.600 ;
        RECT 1293.130 15.400 1297.130 15.540 ;
        RECT 1293.130 15.340 1293.450 15.400 ;
        RECT 1296.810 15.340 1297.130 15.400 ;
      LAYER via ;
        RECT 1296.840 586.540 1297.100 586.800 ;
        RECT 1334.100 586.540 1334.360 586.800 ;
        RECT 1293.160 15.340 1293.420 15.600 ;
        RECT 1296.840 15.340 1297.100 15.600 ;
      LAYER met2 ;
        RECT 1335.710 600.170 1335.990 604.000 ;
        RECT 1334.160 600.030 1335.990 600.170 ;
        RECT 1334.160 586.830 1334.300 600.030 ;
        RECT 1335.710 600.000 1335.990 600.030 ;
        RECT 1296.840 586.510 1297.100 586.830 ;
        RECT 1334.100 586.510 1334.360 586.830 ;
        RECT 1296.900 15.630 1297.040 586.510 ;
        RECT 1293.160 15.310 1293.420 15.630 ;
        RECT 1296.840 15.310 1297.100 15.630 ;
        RECT 1293.220 2.400 1293.360 15.310 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1317.510 589.800 1317.830 589.860 ;
        RECT 1343.270 589.800 1343.590 589.860 ;
        RECT 1317.510 589.660 1343.590 589.800 ;
        RECT 1317.510 589.600 1317.830 589.660 ;
        RECT 1343.270 589.600 1343.590 589.660 ;
        RECT 1311.070 17.580 1311.390 17.640 ;
        RECT 1317.510 17.580 1317.830 17.640 ;
        RECT 1311.070 17.440 1317.830 17.580 ;
        RECT 1311.070 17.380 1311.390 17.440 ;
        RECT 1317.510 17.380 1317.830 17.440 ;
      LAYER via ;
        RECT 1317.540 589.600 1317.800 589.860 ;
        RECT 1343.300 589.600 1343.560 589.860 ;
        RECT 1311.100 17.380 1311.360 17.640 ;
        RECT 1317.540 17.380 1317.800 17.640 ;
      LAYER met2 ;
        RECT 1344.910 600.170 1345.190 604.000 ;
        RECT 1343.360 600.030 1345.190 600.170 ;
        RECT 1343.360 589.890 1343.500 600.030 ;
        RECT 1344.910 600.000 1345.190 600.030 ;
        RECT 1317.540 589.570 1317.800 589.890 ;
        RECT 1343.300 589.570 1343.560 589.890 ;
        RECT 1317.600 17.670 1317.740 589.570 ;
        RECT 1311.100 17.350 1311.360 17.670 ;
        RECT 1317.540 17.350 1317.800 17.670 ;
        RECT 1311.160 2.400 1311.300 17.350 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.310 587.760 1331.630 587.820 ;
        RECT 1352.470 587.760 1352.790 587.820 ;
        RECT 1331.310 587.620 1352.790 587.760 ;
        RECT 1331.310 587.560 1331.630 587.620 ;
        RECT 1352.470 587.560 1352.790 587.620 ;
        RECT 1329.010 20.640 1329.330 20.700 ;
        RECT 1331.310 20.640 1331.630 20.700 ;
        RECT 1329.010 20.500 1331.630 20.640 ;
        RECT 1329.010 20.440 1329.330 20.500 ;
        RECT 1331.310 20.440 1331.630 20.500 ;
      LAYER via ;
        RECT 1331.340 587.560 1331.600 587.820 ;
        RECT 1352.500 587.560 1352.760 587.820 ;
        RECT 1329.040 20.440 1329.300 20.700 ;
        RECT 1331.340 20.440 1331.600 20.700 ;
      LAYER met2 ;
        RECT 1354.110 600.170 1354.390 604.000 ;
        RECT 1352.560 600.030 1354.390 600.170 ;
        RECT 1352.560 587.850 1352.700 600.030 ;
        RECT 1354.110 600.000 1354.390 600.030 ;
        RECT 1331.340 587.530 1331.600 587.850 ;
        RECT 1352.500 587.530 1352.760 587.850 ;
        RECT 1331.400 20.730 1331.540 587.530 ;
        RECT 1329.040 20.410 1329.300 20.730 ;
        RECT 1331.340 20.410 1331.600 20.730 ;
        RECT 1329.100 2.400 1329.240 20.410 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 38.320 686.710 38.380 ;
        RECT 1021.730 38.320 1022.050 38.380 ;
        RECT 686.390 38.180 1022.050 38.320 ;
        RECT 686.390 38.120 686.710 38.180 ;
        RECT 1021.730 38.120 1022.050 38.180 ;
      LAYER via ;
        RECT 686.420 38.120 686.680 38.380 ;
        RECT 1021.760 38.120 1022.020 38.380 ;
      LAYER met2 ;
        RECT 1023.370 600.170 1023.650 604.000 ;
        RECT 1021.820 600.030 1023.650 600.170 ;
        RECT 1021.820 38.410 1021.960 600.030 ;
        RECT 1023.370 600.000 1023.650 600.030 ;
        RECT 686.420 38.090 686.680 38.410 ;
        RECT 1021.760 38.090 1022.020 38.410 ;
        RECT 686.480 2.400 686.620 38.090 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1361.210 579.940 1361.530 580.000 ;
        RECT 1362.130 579.940 1362.450 580.000 ;
        RECT 1361.210 579.800 1362.450 579.940 ;
        RECT 1361.210 579.740 1361.530 579.800 ;
        RECT 1362.130 579.740 1362.450 579.800 ;
        RECT 1358.910 524.180 1359.230 524.240 ;
        RECT 1360.290 524.180 1360.610 524.240 ;
        RECT 1358.910 524.040 1360.610 524.180 ;
        RECT 1358.910 523.980 1359.230 524.040 ;
        RECT 1360.290 523.980 1360.610 524.040 ;
        RECT 1358.910 476.240 1359.230 476.300 ;
        RECT 1359.830 476.240 1360.150 476.300 ;
        RECT 1358.910 476.100 1360.150 476.240 ;
        RECT 1358.910 476.040 1359.230 476.100 ;
        RECT 1359.830 476.040 1360.150 476.100 ;
        RECT 1358.450 427.620 1358.770 427.680 ;
        RECT 1360.290 427.620 1360.610 427.680 ;
        RECT 1358.450 427.480 1360.610 427.620 ;
        RECT 1358.450 427.420 1358.770 427.480 ;
        RECT 1360.290 427.420 1360.610 427.480 ;
        RECT 1358.450 379.680 1358.770 379.740 ;
        RECT 1359.370 379.680 1359.690 379.740 ;
        RECT 1358.450 379.540 1359.690 379.680 ;
        RECT 1358.450 379.480 1358.770 379.540 ;
        RECT 1359.370 379.480 1359.690 379.540 ;
        RECT 1359.830 331.400 1360.150 331.460 ;
        RECT 1361.210 331.400 1361.530 331.460 ;
        RECT 1359.830 331.260 1361.530 331.400 ;
        RECT 1359.830 331.200 1360.150 331.260 ;
        RECT 1361.210 331.200 1361.530 331.260 ;
        RECT 1359.830 303.520 1360.150 303.580 ;
        RECT 1360.750 303.520 1361.070 303.580 ;
        RECT 1359.830 303.380 1361.070 303.520 ;
        RECT 1359.830 303.320 1360.150 303.380 ;
        RECT 1360.750 303.320 1361.070 303.380 ;
        RECT 1359.370 265.780 1359.690 265.840 ;
        RECT 1360.750 265.780 1361.070 265.840 ;
        RECT 1359.370 265.640 1361.070 265.780 ;
        RECT 1359.370 265.580 1359.690 265.640 ;
        RECT 1360.750 265.580 1361.070 265.640 ;
        RECT 1359.370 241.640 1359.690 241.700 ;
        RECT 1359.830 241.640 1360.150 241.700 ;
        RECT 1359.370 241.500 1360.150 241.640 ;
        RECT 1359.370 241.440 1359.690 241.500 ;
        RECT 1359.830 241.440 1360.150 241.500 ;
        RECT 1358.450 193.020 1358.770 193.080 ;
        RECT 1359.370 193.020 1359.690 193.080 ;
        RECT 1358.450 192.880 1359.690 193.020 ;
        RECT 1358.450 192.820 1358.770 192.880 ;
        RECT 1359.370 192.820 1359.690 192.880 ;
        RECT 1358.450 145.080 1358.770 145.140 ;
        RECT 1359.830 145.080 1360.150 145.140 ;
        RECT 1358.450 144.940 1360.150 145.080 ;
        RECT 1358.450 144.880 1358.770 144.940 ;
        RECT 1359.830 144.880 1360.150 144.940 ;
        RECT 1346.490 19.960 1346.810 20.020 ;
        RECT 1360.750 19.960 1361.070 20.020 ;
        RECT 1346.490 19.820 1361.070 19.960 ;
        RECT 1346.490 19.760 1346.810 19.820 ;
        RECT 1360.750 19.760 1361.070 19.820 ;
      LAYER via ;
        RECT 1361.240 579.740 1361.500 580.000 ;
        RECT 1362.160 579.740 1362.420 580.000 ;
        RECT 1358.940 523.980 1359.200 524.240 ;
        RECT 1360.320 523.980 1360.580 524.240 ;
        RECT 1358.940 476.040 1359.200 476.300 ;
        RECT 1359.860 476.040 1360.120 476.300 ;
        RECT 1358.480 427.420 1358.740 427.680 ;
        RECT 1360.320 427.420 1360.580 427.680 ;
        RECT 1358.480 379.480 1358.740 379.740 ;
        RECT 1359.400 379.480 1359.660 379.740 ;
        RECT 1359.860 331.200 1360.120 331.460 ;
        RECT 1361.240 331.200 1361.500 331.460 ;
        RECT 1359.860 303.320 1360.120 303.580 ;
        RECT 1360.780 303.320 1361.040 303.580 ;
        RECT 1359.400 265.580 1359.660 265.840 ;
        RECT 1360.780 265.580 1361.040 265.840 ;
        RECT 1359.400 241.440 1359.660 241.700 ;
        RECT 1359.860 241.440 1360.120 241.700 ;
        RECT 1358.480 192.820 1358.740 193.080 ;
        RECT 1359.400 192.820 1359.660 193.080 ;
        RECT 1358.480 144.880 1358.740 145.140 ;
        RECT 1359.860 144.880 1360.120 145.140 ;
        RECT 1346.520 19.760 1346.780 20.020 ;
        RECT 1360.780 19.760 1361.040 20.020 ;
      LAYER met2 ;
        RECT 1363.310 600.170 1363.590 604.000 ;
        RECT 1362.220 600.030 1363.590 600.170 ;
        RECT 1362.220 580.030 1362.360 600.030 ;
        RECT 1363.310 600.000 1363.590 600.030 ;
        RECT 1361.240 579.710 1361.500 580.030 ;
        RECT 1362.160 579.710 1362.420 580.030 ;
        RECT 1361.300 545.090 1361.440 579.710 ;
        RECT 1360.380 544.950 1361.440 545.090 ;
        RECT 1360.380 524.270 1360.520 544.950 ;
        RECT 1358.940 523.950 1359.200 524.270 ;
        RECT 1360.320 523.950 1360.580 524.270 ;
        RECT 1359.000 476.330 1359.140 523.950 ;
        RECT 1358.940 476.010 1359.200 476.330 ;
        RECT 1359.860 476.010 1360.120 476.330 ;
        RECT 1359.920 458.730 1360.060 476.010 ;
        RECT 1359.920 458.590 1360.520 458.730 ;
        RECT 1360.380 427.710 1360.520 458.590 ;
        RECT 1358.480 427.390 1358.740 427.710 ;
        RECT 1360.320 427.390 1360.580 427.710 ;
        RECT 1358.540 379.770 1358.680 427.390 ;
        RECT 1358.480 379.450 1358.740 379.770 ;
        RECT 1359.400 379.450 1359.660 379.770 ;
        RECT 1359.460 379.285 1359.600 379.450 ;
        RECT 1359.390 378.915 1359.670 379.285 ;
        RECT 1361.230 378.915 1361.510 379.285 ;
        RECT 1361.300 331.490 1361.440 378.915 ;
        RECT 1359.860 331.170 1360.120 331.490 ;
        RECT 1361.240 331.170 1361.500 331.490 ;
        RECT 1359.920 303.610 1360.060 331.170 ;
        RECT 1359.860 303.290 1360.120 303.610 ;
        RECT 1360.780 303.290 1361.040 303.610 ;
        RECT 1360.840 265.870 1360.980 303.290 ;
        RECT 1359.400 265.550 1359.660 265.870 ;
        RECT 1360.780 265.550 1361.040 265.870 ;
        RECT 1359.460 241.730 1359.600 265.550 ;
        RECT 1359.400 241.410 1359.660 241.730 ;
        RECT 1359.860 241.410 1360.120 241.730 ;
        RECT 1359.920 217.330 1360.060 241.410 ;
        RECT 1359.460 217.190 1360.060 217.330 ;
        RECT 1359.460 193.110 1359.600 217.190 ;
        RECT 1358.480 192.790 1358.740 193.110 ;
        RECT 1359.400 192.790 1359.660 193.110 ;
        RECT 1358.540 145.170 1358.680 192.790 ;
        RECT 1358.480 144.850 1358.740 145.170 ;
        RECT 1359.860 144.850 1360.120 145.170 ;
        RECT 1359.920 144.570 1360.060 144.850 ;
        RECT 1359.920 144.430 1360.980 144.570 ;
        RECT 1360.840 20.050 1360.980 144.430 ;
        RECT 1346.520 19.730 1346.780 20.050 ;
        RECT 1360.780 19.730 1361.040 20.050 ;
        RECT 1346.580 2.400 1346.720 19.730 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
      LAYER via2 ;
        RECT 1359.390 378.960 1359.670 379.240 ;
        RECT 1361.230 378.960 1361.510 379.240 ;
      LAYER met3 ;
        RECT 1359.365 379.250 1359.695 379.265 ;
        RECT 1361.205 379.250 1361.535 379.265 ;
        RECT 1359.365 378.950 1361.535 379.250 ;
        RECT 1359.365 378.935 1359.695 378.950 ;
        RECT 1361.205 378.935 1361.535 378.950 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 586.740 1366.130 586.800 ;
        RECT 1370.870 586.740 1371.190 586.800 ;
        RECT 1365.810 586.600 1371.190 586.740 ;
        RECT 1365.810 586.540 1366.130 586.600 ;
        RECT 1370.870 586.540 1371.190 586.600 ;
        RECT 1364.430 2.960 1364.750 3.020 ;
        RECT 1365.810 2.960 1366.130 3.020 ;
        RECT 1364.430 2.820 1366.130 2.960 ;
        RECT 1364.430 2.760 1364.750 2.820 ;
        RECT 1365.810 2.760 1366.130 2.820 ;
      LAYER via ;
        RECT 1365.840 586.540 1366.100 586.800 ;
        RECT 1370.900 586.540 1371.160 586.800 ;
        RECT 1364.460 2.760 1364.720 3.020 ;
        RECT 1365.840 2.760 1366.100 3.020 ;
      LAYER met2 ;
        RECT 1372.510 600.170 1372.790 604.000 ;
        RECT 1370.960 600.030 1372.790 600.170 ;
        RECT 1370.960 586.830 1371.100 600.030 ;
        RECT 1372.510 600.000 1372.790 600.030 ;
        RECT 1365.840 586.510 1366.100 586.830 ;
        RECT 1370.900 586.510 1371.160 586.830 ;
        RECT 1365.900 3.050 1366.040 586.510 ;
        RECT 1364.460 2.730 1364.720 3.050 ;
        RECT 1365.840 2.730 1366.100 3.050 ;
        RECT 1364.520 2.400 1364.660 2.730 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.070 483.040 1380.390 483.100 ;
        RECT 1380.530 483.040 1380.850 483.100 ;
        RECT 1380.070 482.900 1380.850 483.040 ;
        RECT 1380.070 482.840 1380.390 482.900 ;
        RECT 1380.530 482.840 1380.850 482.900 ;
        RECT 1380.070 435.100 1380.390 435.160 ;
        RECT 1380.530 435.100 1380.850 435.160 ;
        RECT 1380.070 434.960 1380.850 435.100 ;
        RECT 1380.070 434.900 1380.390 434.960 ;
        RECT 1380.530 434.900 1380.850 434.960 ;
        RECT 1379.610 427.620 1379.930 427.680 ;
        RECT 1380.530 427.620 1380.850 427.680 ;
        RECT 1379.610 427.480 1380.850 427.620 ;
        RECT 1379.610 427.420 1379.930 427.480 ;
        RECT 1380.530 427.420 1380.850 427.480 ;
        RECT 1379.610 379.680 1379.930 379.740 ;
        RECT 1380.530 379.680 1380.850 379.740 ;
        RECT 1379.610 379.540 1380.850 379.680 ;
        RECT 1379.610 379.480 1379.930 379.540 ;
        RECT 1380.530 379.480 1380.850 379.540 ;
        RECT 1379.610 331.060 1379.930 331.120 ;
        RECT 1380.530 331.060 1380.850 331.120 ;
        RECT 1379.610 330.920 1380.850 331.060 ;
        RECT 1379.610 330.860 1379.930 330.920 ;
        RECT 1380.530 330.860 1380.850 330.920 ;
        RECT 1379.610 283.120 1379.930 283.180 ;
        RECT 1380.070 283.120 1380.390 283.180 ;
        RECT 1379.610 282.980 1380.390 283.120 ;
        RECT 1379.610 282.920 1379.930 282.980 ;
        RECT 1380.070 282.920 1380.390 282.980 ;
        RECT 1379.610 234.500 1379.930 234.560 ;
        RECT 1380.530 234.500 1380.850 234.560 ;
        RECT 1379.610 234.360 1380.850 234.500 ;
        RECT 1379.610 234.300 1379.930 234.360 ;
        RECT 1380.530 234.300 1380.850 234.360 ;
        RECT 1379.610 186.560 1379.930 186.620 ;
        RECT 1380.070 186.560 1380.390 186.620 ;
        RECT 1379.610 186.420 1380.390 186.560 ;
        RECT 1379.610 186.360 1379.930 186.420 ;
        RECT 1380.070 186.360 1380.390 186.420 ;
        RECT 1380.530 137.940 1380.850 138.000 ;
        RECT 1380.990 137.940 1381.310 138.000 ;
        RECT 1380.530 137.800 1381.310 137.940 ;
        RECT 1380.530 137.740 1380.850 137.800 ;
        RECT 1380.990 137.740 1381.310 137.800 ;
        RECT 1380.990 48.520 1381.310 48.580 ;
        RECT 1382.370 48.520 1382.690 48.580 ;
        RECT 1380.990 48.380 1382.690 48.520 ;
        RECT 1380.990 48.320 1381.310 48.380 ;
        RECT 1382.370 48.320 1382.690 48.380 ;
      LAYER via ;
        RECT 1380.100 482.840 1380.360 483.100 ;
        RECT 1380.560 482.840 1380.820 483.100 ;
        RECT 1380.100 434.900 1380.360 435.160 ;
        RECT 1380.560 434.900 1380.820 435.160 ;
        RECT 1379.640 427.420 1379.900 427.680 ;
        RECT 1380.560 427.420 1380.820 427.680 ;
        RECT 1379.640 379.480 1379.900 379.740 ;
        RECT 1380.560 379.480 1380.820 379.740 ;
        RECT 1379.640 330.860 1379.900 331.120 ;
        RECT 1380.560 330.860 1380.820 331.120 ;
        RECT 1379.640 282.920 1379.900 283.180 ;
        RECT 1380.100 282.920 1380.360 283.180 ;
        RECT 1379.640 234.300 1379.900 234.560 ;
        RECT 1380.560 234.300 1380.820 234.560 ;
        RECT 1379.640 186.360 1379.900 186.620 ;
        RECT 1380.100 186.360 1380.360 186.620 ;
        RECT 1380.560 137.740 1380.820 138.000 ;
        RECT 1381.020 137.740 1381.280 138.000 ;
        RECT 1381.020 48.320 1381.280 48.580 ;
        RECT 1382.400 48.320 1382.660 48.580 ;
      LAYER met2 ;
        RECT 1381.250 600.170 1381.530 604.000 ;
        RECT 1380.620 600.030 1381.530 600.170 ;
        RECT 1380.620 483.130 1380.760 600.030 ;
        RECT 1381.250 600.000 1381.530 600.030 ;
        RECT 1380.100 482.810 1380.360 483.130 ;
        RECT 1380.560 482.810 1380.820 483.130 ;
        RECT 1380.160 435.190 1380.300 482.810 ;
        RECT 1380.100 434.870 1380.360 435.190 ;
        RECT 1380.560 434.870 1380.820 435.190 ;
        RECT 1380.620 427.710 1380.760 434.870 ;
        RECT 1379.640 427.390 1379.900 427.710 ;
        RECT 1380.560 427.390 1380.820 427.710 ;
        RECT 1379.700 379.770 1379.840 427.390 ;
        RECT 1379.640 379.450 1379.900 379.770 ;
        RECT 1380.560 379.450 1380.820 379.770 ;
        RECT 1380.620 331.150 1380.760 379.450 ;
        RECT 1379.640 330.830 1379.900 331.150 ;
        RECT 1380.560 330.830 1380.820 331.150 ;
        RECT 1379.700 283.210 1379.840 330.830 ;
        RECT 1379.640 282.890 1379.900 283.210 ;
        RECT 1380.100 282.890 1380.360 283.210 ;
        RECT 1380.160 241.810 1380.300 282.890 ;
        RECT 1380.160 241.670 1380.760 241.810 ;
        RECT 1380.620 234.590 1380.760 241.670 ;
        RECT 1379.640 234.270 1379.900 234.590 ;
        RECT 1380.560 234.270 1380.820 234.590 ;
        RECT 1379.700 186.650 1379.840 234.270 ;
        RECT 1379.640 186.330 1379.900 186.650 ;
        RECT 1380.100 186.330 1380.360 186.650 ;
        RECT 1380.160 145.250 1380.300 186.330 ;
        RECT 1380.160 145.110 1380.760 145.250 ;
        RECT 1380.620 138.030 1380.760 145.110 ;
        RECT 1380.560 137.710 1380.820 138.030 ;
        RECT 1381.020 137.710 1381.280 138.030 ;
        RECT 1381.080 48.610 1381.220 137.710 ;
        RECT 1381.020 48.290 1381.280 48.610 ;
        RECT 1382.400 48.290 1382.660 48.610 ;
        RECT 1382.460 2.400 1382.600 48.290 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1392.030 587.080 1392.350 587.140 ;
        RECT 1395.710 587.080 1396.030 587.140 ;
        RECT 1392.030 586.940 1396.030 587.080 ;
        RECT 1392.030 586.880 1392.350 586.940 ;
        RECT 1395.710 586.880 1396.030 586.940 ;
      LAYER via ;
        RECT 1392.060 586.880 1392.320 587.140 ;
        RECT 1395.740 586.880 1396.000 587.140 ;
      LAYER met2 ;
        RECT 1390.450 600.170 1390.730 604.000 ;
        RECT 1390.450 600.030 1392.260 600.170 ;
        RECT 1390.450 600.000 1390.730 600.030 ;
        RECT 1392.120 587.170 1392.260 600.030 ;
        RECT 1392.060 586.850 1392.320 587.170 ;
        RECT 1395.740 586.850 1396.000 587.170 ;
        RECT 1395.800 20.130 1395.940 586.850 ;
        RECT 1395.800 19.990 1400.540 20.130 ;
        RECT 1400.400 2.400 1400.540 19.990 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 587.760 1400.630 587.820 ;
        RECT 1415.030 587.760 1415.350 587.820 ;
        RECT 1400.310 587.620 1415.350 587.760 ;
        RECT 1400.310 587.560 1400.630 587.620 ;
        RECT 1415.030 587.560 1415.350 587.620 ;
        RECT 1414.570 48.520 1414.890 48.580 ;
        RECT 1416.870 48.520 1417.190 48.580 ;
        RECT 1414.570 48.380 1417.190 48.520 ;
        RECT 1414.570 48.320 1414.890 48.380 ;
        RECT 1416.870 48.320 1417.190 48.380 ;
      LAYER via ;
        RECT 1400.340 587.560 1400.600 587.820 ;
        RECT 1415.060 587.560 1415.320 587.820 ;
        RECT 1414.600 48.320 1414.860 48.580 ;
        RECT 1416.900 48.320 1417.160 48.580 ;
      LAYER met2 ;
        RECT 1399.650 600.170 1399.930 604.000 ;
        RECT 1399.650 600.030 1400.540 600.170 ;
        RECT 1399.650 600.000 1399.930 600.030 ;
        RECT 1400.400 587.850 1400.540 600.030 ;
        RECT 1400.340 587.530 1400.600 587.850 ;
        RECT 1415.060 587.530 1415.320 587.850 ;
        RECT 1415.120 72.490 1415.260 587.530 ;
        RECT 1414.660 72.350 1415.260 72.490 ;
        RECT 1414.660 48.610 1414.800 72.350 ;
        RECT 1414.600 48.290 1414.860 48.610 ;
        RECT 1416.900 48.290 1417.160 48.610 ;
        RECT 1416.960 19.450 1417.100 48.290 ;
        RECT 1416.960 19.310 1418.480 19.450 ;
        RECT 1418.340 2.400 1418.480 19.310 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1410.430 587.080 1410.750 587.140 ;
        RECT 1417.790 587.080 1418.110 587.140 ;
        RECT 1410.430 586.940 1418.110 587.080 ;
        RECT 1410.430 586.880 1410.750 586.940 ;
        RECT 1417.790 586.880 1418.110 586.940 ;
        RECT 1417.790 20.300 1418.110 20.360 ;
        RECT 1435.730 20.300 1436.050 20.360 ;
        RECT 1417.790 20.160 1436.050 20.300 ;
        RECT 1417.790 20.100 1418.110 20.160 ;
        RECT 1435.730 20.100 1436.050 20.160 ;
      LAYER via ;
        RECT 1410.460 586.880 1410.720 587.140 ;
        RECT 1417.820 586.880 1418.080 587.140 ;
        RECT 1417.820 20.100 1418.080 20.360 ;
        RECT 1435.760 20.100 1436.020 20.360 ;
      LAYER met2 ;
        RECT 1408.850 600.170 1409.130 604.000 ;
        RECT 1408.850 600.030 1410.660 600.170 ;
        RECT 1408.850 600.000 1409.130 600.030 ;
        RECT 1410.520 587.170 1410.660 600.030 ;
        RECT 1410.460 586.850 1410.720 587.170 ;
        RECT 1417.820 586.850 1418.080 587.170 ;
        RECT 1417.880 20.390 1418.020 586.850 ;
        RECT 1417.820 20.070 1418.080 20.390 ;
        RECT 1435.760 20.070 1436.020 20.390 ;
        RECT 1435.820 2.400 1435.960 20.070 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1419.630 590.820 1419.950 590.880 ;
        RECT 1450.450 590.820 1450.770 590.880 ;
        RECT 1419.630 590.680 1450.770 590.820 ;
        RECT 1419.630 590.620 1419.950 590.680 ;
        RECT 1450.450 590.620 1450.770 590.680 ;
        RECT 1450.450 2.960 1450.770 3.020 ;
        RECT 1453.670 2.960 1453.990 3.020 ;
        RECT 1450.450 2.820 1453.990 2.960 ;
        RECT 1450.450 2.760 1450.770 2.820 ;
        RECT 1453.670 2.760 1453.990 2.820 ;
      LAYER via ;
        RECT 1419.660 590.620 1419.920 590.880 ;
        RECT 1450.480 590.620 1450.740 590.880 ;
        RECT 1450.480 2.760 1450.740 3.020 ;
        RECT 1453.700 2.760 1453.960 3.020 ;
      LAYER met2 ;
        RECT 1418.050 600.170 1418.330 604.000 ;
        RECT 1418.050 600.030 1419.860 600.170 ;
        RECT 1418.050 600.000 1418.330 600.030 ;
        RECT 1419.720 590.910 1419.860 600.030 ;
        RECT 1419.660 590.590 1419.920 590.910 ;
        RECT 1450.480 590.590 1450.740 590.910 ;
        RECT 1450.540 3.050 1450.680 590.590 ;
        RECT 1450.480 2.730 1450.740 3.050 ;
        RECT 1453.700 2.730 1453.960 3.050 ;
        RECT 1453.760 2.400 1453.900 2.730 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1427.450 17.240 1427.770 17.300 ;
        RECT 1471.610 17.240 1471.930 17.300 ;
        RECT 1427.450 17.100 1471.930 17.240 ;
        RECT 1427.450 17.040 1427.770 17.100 ;
        RECT 1471.610 17.040 1471.930 17.100 ;
      LAYER via ;
        RECT 1427.480 17.040 1427.740 17.300 ;
        RECT 1471.640 17.040 1471.900 17.300 ;
      LAYER met2 ;
        RECT 1427.250 600.000 1427.530 604.000 ;
        RECT 1427.310 598.810 1427.450 600.000 ;
        RECT 1427.310 598.670 1427.680 598.810 ;
        RECT 1427.540 17.330 1427.680 598.670 ;
        RECT 1427.480 17.010 1427.740 17.330 ;
        RECT 1471.640 17.010 1471.900 17.330 ;
        RECT 1471.700 2.400 1471.840 17.010 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1438.030 586.740 1438.350 586.800 ;
        RECT 1441.710 586.740 1442.030 586.800 ;
        RECT 1438.030 586.600 1442.030 586.740 ;
        RECT 1438.030 586.540 1438.350 586.600 ;
        RECT 1441.710 586.540 1442.030 586.600 ;
        RECT 1441.250 19.620 1441.570 19.680 ;
        RECT 1489.550 19.620 1489.870 19.680 ;
        RECT 1441.250 19.480 1489.870 19.620 ;
        RECT 1441.250 19.420 1441.570 19.480 ;
        RECT 1489.550 19.420 1489.870 19.480 ;
      LAYER via ;
        RECT 1438.060 586.540 1438.320 586.800 ;
        RECT 1441.740 586.540 1442.000 586.800 ;
        RECT 1441.280 19.420 1441.540 19.680 ;
        RECT 1489.580 19.420 1489.840 19.680 ;
      LAYER met2 ;
        RECT 1436.450 600.170 1436.730 604.000 ;
        RECT 1436.450 600.030 1438.260 600.170 ;
        RECT 1436.450 600.000 1436.730 600.030 ;
        RECT 1438.120 586.830 1438.260 600.030 ;
        RECT 1438.060 586.510 1438.320 586.830 ;
        RECT 1441.740 586.510 1442.000 586.830 ;
        RECT 1441.800 41.210 1441.940 586.510 ;
        RECT 1441.340 41.070 1441.940 41.210 ;
        RECT 1441.340 19.710 1441.480 41.070 ;
        RECT 1441.280 19.390 1441.540 19.710 ;
        RECT 1489.580 19.390 1489.840 19.710 ;
        RECT 1489.640 2.400 1489.780 19.390 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1447.230 587.080 1447.550 587.140 ;
        RECT 1472.990 587.080 1473.310 587.140 ;
        RECT 1447.230 586.940 1473.310 587.080 ;
        RECT 1447.230 586.880 1447.550 586.940 ;
        RECT 1472.990 586.880 1473.310 586.940 ;
        RECT 1472.990 16.220 1473.310 16.280 ;
        RECT 1507.030 16.220 1507.350 16.280 ;
        RECT 1472.990 16.080 1507.350 16.220 ;
        RECT 1472.990 16.020 1473.310 16.080 ;
        RECT 1507.030 16.020 1507.350 16.080 ;
      LAYER via ;
        RECT 1447.260 586.880 1447.520 587.140 ;
        RECT 1473.020 586.880 1473.280 587.140 ;
        RECT 1473.020 16.020 1473.280 16.280 ;
        RECT 1507.060 16.020 1507.320 16.280 ;
      LAYER met2 ;
        RECT 1445.650 600.170 1445.930 604.000 ;
        RECT 1445.650 600.030 1447.460 600.170 ;
        RECT 1445.650 600.000 1445.930 600.030 ;
        RECT 1447.320 587.170 1447.460 600.030 ;
        RECT 1447.260 586.850 1447.520 587.170 ;
        RECT 1473.020 586.850 1473.280 587.170 ;
        RECT 1473.080 16.310 1473.220 586.850 ;
        RECT 1473.020 15.990 1473.280 16.310 ;
        RECT 1507.060 15.990 1507.320 16.310 ;
        RECT 1507.120 2.400 1507.260 15.990 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1028.170 569.400 1028.490 569.460 ;
        RECT 1030.930 569.400 1031.250 569.460 ;
        RECT 1028.170 569.260 1031.250 569.400 ;
        RECT 1028.170 569.200 1028.490 569.260 ;
        RECT 1030.930 569.200 1031.250 569.260 ;
        RECT 704.330 39.340 704.650 39.400 ;
        RECT 1028.170 39.340 1028.490 39.400 ;
        RECT 704.330 39.200 1028.490 39.340 ;
        RECT 704.330 39.140 704.650 39.200 ;
        RECT 1028.170 39.140 1028.490 39.200 ;
      LAYER via ;
        RECT 1028.200 569.200 1028.460 569.460 ;
        RECT 1030.960 569.200 1031.220 569.460 ;
        RECT 704.360 39.140 704.620 39.400 ;
        RECT 1028.200 39.140 1028.460 39.400 ;
      LAYER met2 ;
        RECT 1032.570 600.170 1032.850 604.000 ;
        RECT 1031.020 600.030 1032.850 600.170 ;
        RECT 1031.020 569.490 1031.160 600.030 ;
        RECT 1032.570 600.000 1032.850 600.030 ;
        RECT 1028.200 569.170 1028.460 569.490 ;
        RECT 1030.960 569.170 1031.220 569.490 ;
        RECT 1028.260 39.430 1028.400 569.170 ;
        RECT 704.360 39.110 704.620 39.430 ;
        RECT 1028.200 39.110 1028.460 39.430 ;
        RECT 704.420 2.400 704.560 39.110 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.050 17.580 1455.370 17.640 ;
        RECT 1524.970 17.580 1525.290 17.640 ;
        RECT 1455.050 17.440 1525.290 17.580 ;
        RECT 1455.050 17.380 1455.370 17.440 ;
        RECT 1524.970 17.380 1525.290 17.440 ;
      LAYER via ;
        RECT 1455.080 17.380 1455.340 17.640 ;
        RECT 1525.000 17.380 1525.260 17.640 ;
      LAYER met2 ;
        RECT 1454.850 600.000 1455.130 604.000 ;
        RECT 1454.910 598.810 1455.050 600.000 ;
        RECT 1454.910 598.670 1455.280 598.810 ;
        RECT 1455.140 17.670 1455.280 598.670 ;
        RECT 1455.080 17.350 1455.340 17.670 ;
        RECT 1525.000 17.350 1525.260 17.670 ;
        RECT 1525.060 2.400 1525.200 17.350 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1465.630 589.460 1465.950 589.520 ;
        RECT 1469.310 589.460 1469.630 589.520 ;
        RECT 1465.630 589.320 1469.630 589.460 ;
        RECT 1465.630 589.260 1465.950 589.320 ;
        RECT 1469.310 589.260 1469.630 589.320 ;
        RECT 1469.310 16.900 1469.630 16.960 ;
        RECT 1542.910 16.900 1543.230 16.960 ;
        RECT 1469.310 16.760 1543.230 16.900 ;
        RECT 1469.310 16.700 1469.630 16.760 ;
        RECT 1542.910 16.700 1543.230 16.760 ;
      LAYER via ;
        RECT 1465.660 589.260 1465.920 589.520 ;
        RECT 1469.340 589.260 1469.600 589.520 ;
        RECT 1469.340 16.700 1469.600 16.960 ;
        RECT 1542.940 16.700 1543.200 16.960 ;
      LAYER met2 ;
        RECT 1464.050 600.170 1464.330 604.000 ;
        RECT 1464.050 600.030 1465.860 600.170 ;
        RECT 1464.050 600.000 1464.330 600.030 ;
        RECT 1465.720 589.550 1465.860 600.030 ;
        RECT 1465.660 589.230 1465.920 589.550 ;
        RECT 1469.340 589.230 1469.600 589.550 ;
        RECT 1469.400 16.990 1469.540 589.230 ;
        RECT 1469.340 16.670 1469.600 16.990 ;
        RECT 1542.940 16.670 1543.200 16.990 ;
        RECT 1543.000 2.400 1543.140 16.670 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1474.830 588.100 1475.150 588.160 ;
        RECT 1559.470 588.100 1559.790 588.160 ;
        RECT 1474.830 587.960 1559.790 588.100 ;
        RECT 1474.830 587.900 1475.150 587.960 ;
        RECT 1559.470 587.900 1559.790 587.960 ;
      LAYER via ;
        RECT 1474.860 587.900 1475.120 588.160 ;
        RECT 1559.500 587.900 1559.760 588.160 ;
      LAYER met2 ;
        RECT 1473.250 600.170 1473.530 604.000 ;
        RECT 1473.250 600.030 1475.060 600.170 ;
        RECT 1473.250 600.000 1473.530 600.030 ;
        RECT 1474.920 588.190 1475.060 600.030 ;
        RECT 1474.860 587.870 1475.120 588.190 ;
        RECT 1559.500 587.870 1559.760 588.190 ;
        RECT 1559.560 3.130 1559.700 587.870 ;
        RECT 1559.560 2.990 1561.080 3.130 ;
        RECT 1560.940 2.400 1561.080 2.990 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1483.110 590.480 1483.430 590.540 ;
        RECT 1574.190 590.480 1574.510 590.540 ;
        RECT 1483.110 590.340 1574.510 590.480 ;
        RECT 1483.110 590.280 1483.430 590.340 ;
        RECT 1574.190 590.280 1574.510 590.340 ;
      LAYER via ;
        RECT 1483.140 590.280 1483.400 590.540 ;
        RECT 1574.220 590.280 1574.480 590.540 ;
      LAYER met2 ;
        RECT 1482.450 600.170 1482.730 604.000 ;
        RECT 1482.450 600.030 1483.340 600.170 ;
        RECT 1482.450 600.000 1482.730 600.030 ;
        RECT 1483.200 590.570 1483.340 600.030 ;
        RECT 1483.140 590.250 1483.400 590.570 ;
        RECT 1574.220 590.250 1574.480 590.570 ;
        RECT 1574.280 16.730 1574.420 590.250 ;
        RECT 1574.280 16.590 1579.020 16.730 ;
        RECT 1578.880 2.400 1579.020 16.590 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1493.230 590.140 1493.550 590.200 ;
        RECT 1594.890 590.140 1595.210 590.200 ;
        RECT 1493.230 590.000 1595.210 590.140 ;
        RECT 1493.230 589.940 1493.550 590.000 ;
        RECT 1594.890 589.940 1595.210 590.000 ;
        RECT 1594.890 2.960 1595.210 3.020 ;
        RECT 1596.270 2.960 1596.590 3.020 ;
        RECT 1594.890 2.820 1596.590 2.960 ;
        RECT 1594.890 2.760 1595.210 2.820 ;
        RECT 1596.270 2.760 1596.590 2.820 ;
      LAYER via ;
        RECT 1493.260 589.940 1493.520 590.200 ;
        RECT 1594.920 589.940 1595.180 590.200 ;
        RECT 1594.920 2.760 1595.180 3.020 ;
        RECT 1596.300 2.760 1596.560 3.020 ;
      LAYER met2 ;
        RECT 1491.650 600.170 1491.930 604.000 ;
        RECT 1491.650 600.030 1493.460 600.170 ;
        RECT 1491.650 600.000 1491.930 600.030 ;
        RECT 1493.320 590.230 1493.460 600.030 ;
        RECT 1493.260 589.910 1493.520 590.230 ;
        RECT 1594.920 589.910 1595.180 590.230 ;
        RECT 1594.980 3.050 1595.120 589.910 ;
        RECT 1594.920 2.730 1595.180 3.050 ;
        RECT 1596.300 2.730 1596.560 3.050 ;
        RECT 1596.360 2.400 1596.500 2.730 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1502.430 589.800 1502.750 589.860 ;
        RECT 1608.690 589.800 1609.010 589.860 ;
        RECT 1502.430 589.660 1609.010 589.800 ;
        RECT 1502.430 589.600 1502.750 589.660 ;
        RECT 1608.690 589.600 1609.010 589.660 ;
        RECT 1608.690 61.920 1609.010 62.180 ;
        RECT 1608.780 61.780 1608.920 61.920 ;
        RECT 1613.750 61.780 1614.070 61.840 ;
        RECT 1608.780 61.640 1614.070 61.780 ;
        RECT 1613.750 61.580 1614.070 61.640 ;
      LAYER via ;
        RECT 1502.460 589.600 1502.720 589.860 ;
        RECT 1608.720 589.600 1608.980 589.860 ;
        RECT 1608.720 61.920 1608.980 62.180 ;
        RECT 1613.780 61.580 1614.040 61.840 ;
      LAYER met2 ;
        RECT 1500.850 600.170 1501.130 604.000 ;
        RECT 1500.850 600.030 1502.660 600.170 ;
        RECT 1500.850 600.000 1501.130 600.030 ;
        RECT 1502.520 589.890 1502.660 600.030 ;
        RECT 1502.460 589.570 1502.720 589.890 ;
        RECT 1608.720 589.570 1608.980 589.890 ;
        RECT 1608.780 62.210 1608.920 589.570 ;
        RECT 1608.720 61.890 1608.980 62.210 ;
        RECT 1613.780 61.550 1614.040 61.870 ;
        RECT 1613.840 19.450 1613.980 61.550 ;
        RECT 1613.840 19.310 1614.440 19.450 ;
        RECT 1614.300 2.400 1614.440 19.310 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1510.710 588.780 1511.030 588.840 ;
        RECT 1607.770 588.780 1608.090 588.840 ;
        RECT 1510.710 588.640 1608.090 588.780 ;
        RECT 1510.710 588.580 1511.030 588.640 ;
        RECT 1607.770 588.580 1608.090 588.640 ;
        RECT 1607.770 572.800 1608.090 572.860 ;
        RECT 1628.470 572.800 1628.790 572.860 ;
        RECT 1607.770 572.660 1628.790 572.800 ;
        RECT 1607.770 572.600 1608.090 572.660 ;
        RECT 1628.470 572.600 1628.790 572.660 ;
        RECT 1628.470 524.180 1628.790 524.240 ;
        RECT 1629.390 524.180 1629.710 524.240 ;
        RECT 1628.470 524.040 1629.710 524.180 ;
        RECT 1628.470 523.980 1628.790 524.040 ;
        RECT 1629.390 523.980 1629.710 524.040 ;
        RECT 1628.470 476.240 1628.790 476.300 ;
        RECT 1629.390 476.240 1629.710 476.300 ;
        RECT 1628.470 476.100 1629.710 476.240 ;
        RECT 1628.470 476.040 1628.790 476.100 ;
        RECT 1629.390 476.040 1629.710 476.100 ;
        RECT 1628.470 427.620 1628.790 427.680 ;
        RECT 1629.390 427.620 1629.710 427.680 ;
        RECT 1628.470 427.480 1629.710 427.620 ;
        RECT 1628.470 427.420 1628.790 427.480 ;
        RECT 1629.390 427.420 1629.710 427.480 ;
        RECT 1628.470 379.680 1628.790 379.740 ;
        RECT 1629.390 379.680 1629.710 379.740 ;
        RECT 1628.470 379.540 1629.710 379.680 ;
        RECT 1628.470 379.480 1628.790 379.540 ;
        RECT 1629.390 379.480 1629.710 379.540 ;
        RECT 1627.550 331.060 1627.870 331.120 ;
        RECT 1628.470 331.060 1628.790 331.120 ;
        RECT 1627.550 330.920 1628.790 331.060 ;
        RECT 1627.550 330.860 1627.870 330.920 ;
        RECT 1628.470 330.860 1628.790 330.920 ;
        RECT 1627.550 283.120 1627.870 283.180 ;
        RECT 1628.930 283.120 1629.250 283.180 ;
        RECT 1627.550 282.980 1629.250 283.120 ;
        RECT 1627.550 282.920 1627.870 282.980 ;
        RECT 1628.930 282.920 1629.250 282.980 ;
        RECT 1627.550 234.500 1627.870 234.560 ;
        RECT 1628.470 234.500 1628.790 234.560 ;
        RECT 1627.550 234.360 1628.790 234.500 ;
        RECT 1627.550 234.300 1627.870 234.360 ;
        RECT 1628.470 234.300 1628.790 234.360 ;
        RECT 1627.550 186.560 1627.870 186.620 ;
        RECT 1628.930 186.560 1629.250 186.620 ;
        RECT 1627.550 186.420 1629.250 186.560 ;
        RECT 1627.550 186.360 1627.870 186.420 ;
        RECT 1628.930 186.360 1629.250 186.420 ;
        RECT 1627.090 137.940 1627.410 138.000 ;
        RECT 1628.470 137.940 1628.790 138.000 ;
        RECT 1627.090 137.800 1628.790 137.940 ;
        RECT 1627.090 137.740 1627.410 137.800 ;
        RECT 1628.470 137.740 1628.790 137.800 ;
        RECT 1627.090 90.000 1627.410 90.060 ;
        RECT 1628.010 90.000 1628.330 90.060 ;
        RECT 1627.090 89.860 1628.330 90.000 ;
        RECT 1627.090 89.800 1627.410 89.860 ;
        RECT 1628.010 89.800 1628.330 89.860 ;
        RECT 1628.010 48.520 1628.330 48.580 ;
        RECT 1631.230 48.520 1631.550 48.580 ;
        RECT 1628.010 48.380 1631.550 48.520 ;
        RECT 1628.010 48.320 1628.330 48.380 ;
        RECT 1631.230 48.320 1631.550 48.380 ;
        RECT 1630.770 18.940 1631.090 19.000 ;
        RECT 1631.690 18.940 1632.010 19.000 ;
        RECT 1630.770 18.800 1632.010 18.940 ;
        RECT 1630.770 18.740 1631.090 18.800 ;
        RECT 1631.690 18.740 1632.010 18.800 ;
        RECT 1631.690 2.960 1632.010 3.020 ;
        RECT 1632.150 2.960 1632.470 3.020 ;
        RECT 1631.690 2.820 1632.470 2.960 ;
        RECT 1631.690 2.760 1632.010 2.820 ;
        RECT 1632.150 2.760 1632.470 2.820 ;
      LAYER via ;
        RECT 1510.740 588.580 1511.000 588.840 ;
        RECT 1607.800 588.580 1608.060 588.840 ;
        RECT 1607.800 572.600 1608.060 572.860 ;
        RECT 1628.500 572.600 1628.760 572.860 ;
        RECT 1628.500 523.980 1628.760 524.240 ;
        RECT 1629.420 523.980 1629.680 524.240 ;
        RECT 1628.500 476.040 1628.760 476.300 ;
        RECT 1629.420 476.040 1629.680 476.300 ;
        RECT 1628.500 427.420 1628.760 427.680 ;
        RECT 1629.420 427.420 1629.680 427.680 ;
        RECT 1628.500 379.480 1628.760 379.740 ;
        RECT 1629.420 379.480 1629.680 379.740 ;
        RECT 1627.580 330.860 1627.840 331.120 ;
        RECT 1628.500 330.860 1628.760 331.120 ;
        RECT 1627.580 282.920 1627.840 283.180 ;
        RECT 1628.960 282.920 1629.220 283.180 ;
        RECT 1627.580 234.300 1627.840 234.560 ;
        RECT 1628.500 234.300 1628.760 234.560 ;
        RECT 1627.580 186.360 1627.840 186.620 ;
        RECT 1628.960 186.360 1629.220 186.620 ;
        RECT 1627.120 137.740 1627.380 138.000 ;
        RECT 1628.500 137.740 1628.760 138.000 ;
        RECT 1627.120 89.800 1627.380 90.060 ;
        RECT 1628.040 89.800 1628.300 90.060 ;
        RECT 1628.040 48.320 1628.300 48.580 ;
        RECT 1631.260 48.320 1631.520 48.580 ;
        RECT 1630.800 18.740 1631.060 19.000 ;
        RECT 1631.720 18.740 1631.980 19.000 ;
        RECT 1631.720 2.760 1631.980 3.020 ;
        RECT 1632.180 2.760 1632.440 3.020 ;
      LAYER met2 ;
        RECT 1510.050 600.170 1510.330 604.000 ;
        RECT 1510.050 600.030 1510.940 600.170 ;
        RECT 1510.050 600.000 1510.330 600.030 ;
        RECT 1510.800 588.870 1510.940 600.030 ;
        RECT 1510.740 588.550 1511.000 588.870 ;
        RECT 1607.800 588.550 1608.060 588.870 ;
        RECT 1607.860 572.890 1608.000 588.550 ;
        RECT 1607.800 572.570 1608.060 572.890 ;
        RECT 1628.500 572.570 1628.760 572.890 ;
        RECT 1628.560 524.270 1628.700 572.570 ;
        RECT 1628.500 523.950 1628.760 524.270 ;
        RECT 1629.420 523.950 1629.680 524.270 ;
        RECT 1629.480 476.330 1629.620 523.950 ;
        RECT 1628.500 476.010 1628.760 476.330 ;
        RECT 1629.420 476.010 1629.680 476.330 ;
        RECT 1628.560 427.710 1628.700 476.010 ;
        RECT 1628.500 427.390 1628.760 427.710 ;
        RECT 1629.420 427.390 1629.680 427.710 ;
        RECT 1629.480 379.770 1629.620 427.390 ;
        RECT 1628.500 379.450 1628.760 379.770 ;
        RECT 1629.420 379.450 1629.680 379.770 ;
        RECT 1628.560 331.150 1628.700 379.450 ;
        RECT 1627.580 330.830 1627.840 331.150 ;
        RECT 1628.500 330.830 1628.760 331.150 ;
        RECT 1627.640 283.210 1627.780 330.830 ;
        RECT 1627.580 282.890 1627.840 283.210 ;
        RECT 1628.960 282.890 1629.220 283.210 ;
        RECT 1629.020 241.810 1629.160 282.890 ;
        RECT 1628.560 241.670 1629.160 241.810 ;
        RECT 1628.560 234.590 1628.700 241.670 ;
        RECT 1627.580 234.270 1627.840 234.590 ;
        RECT 1628.500 234.270 1628.760 234.590 ;
        RECT 1627.640 186.650 1627.780 234.270 ;
        RECT 1627.580 186.330 1627.840 186.650 ;
        RECT 1628.960 186.330 1629.220 186.650 ;
        RECT 1629.020 145.250 1629.160 186.330 ;
        RECT 1628.560 145.110 1629.160 145.250 ;
        RECT 1628.560 138.030 1628.700 145.110 ;
        RECT 1627.120 137.710 1627.380 138.030 ;
        RECT 1628.500 137.710 1628.760 138.030 ;
        RECT 1627.180 90.090 1627.320 137.710 ;
        RECT 1627.120 89.770 1627.380 90.090 ;
        RECT 1628.040 89.770 1628.300 90.090 ;
        RECT 1628.100 48.610 1628.240 89.770 ;
        RECT 1628.040 48.290 1628.300 48.610 ;
        RECT 1631.260 48.290 1631.520 48.610 ;
        RECT 1631.320 48.010 1631.460 48.290 ;
        RECT 1630.860 47.870 1631.460 48.010 ;
        RECT 1630.860 19.030 1631.000 47.870 ;
        RECT 1630.800 18.710 1631.060 19.030 ;
        RECT 1631.720 18.710 1631.980 19.030 ;
        RECT 1631.780 3.050 1631.920 18.710 ;
        RECT 1631.720 2.730 1631.980 3.050 ;
        RECT 1632.180 2.730 1632.440 3.050 ;
        RECT 1632.240 2.400 1632.380 2.730 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1520.830 588.440 1521.150 588.500 ;
        RECT 1520.830 588.300 1617.660 588.440 ;
        RECT 1520.830 588.240 1521.150 588.300 ;
        RECT 1617.520 587.080 1617.660 588.300 ;
        RECT 1649.170 587.080 1649.490 587.140 ;
        RECT 1617.520 586.940 1649.490 587.080 ;
        RECT 1649.170 586.880 1649.490 586.940 ;
      LAYER via ;
        RECT 1520.860 588.240 1521.120 588.500 ;
        RECT 1649.200 586.880 1649.460 587.140 ;
      LAYER met2 ;
        RECT 1519.250 600.170 1519.530 604.000 ;
        RECT 1519.250 600.030 1521.060 600.170 ;
        RECT 1519.250 600.000 1519.530 600.030 ;
        RECT 1520.920 588.530 1521.060 600.030 ;
        RECT 1520.860 588.210 1521.120 588.530 ;
        RECT 1649.200 586.850 1649.460 587.170 ;
        RECT 1649.260 3.130 1649.400 586.850 ;
        RECT 1649.260 2.990 1650.320 3.130 ;
        RECT 1650.180 2.400 1650.320 2.990 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1530.030 593.200 1530.350 593.260 ;
        RECT 1664.350 593.200 1664.670 593.260 ;
        RECT 1530.030 593.060 1664.670 593.200 ;
        RECT 1530.030 593.000 1530.350 593.060 ;
        RECT 1664.350 593.000 1664.670 593.060 ;
        RECT 1664.350 2.960 1664.670 3.020 ;
        RECT 1668.030 2.960 1668.350 3.020 ;
        RECT 1664.350 2.820 1668.350 2.960 ;
        RECT 1664.350 2.760 1664.670 2.820 ;
        RECT 1668.030 2.760 1668.350 2.820 ;
      LAYER via ;
        RECT 1530.060 593.000 1530.320 593.260 ;
        RECT 1664.380 593.000 1664.640 593.260 ;
        RECT 1664.380 2.760 1664.640 3.020 ;
        RECT 1668.060 2.760 1668.320 3.020 ;
      LAYER met2 ;
        RECT 1528.450 600.170 1528.730 604.000 ;
        RECT 1528.450 600.030 1530.260 600.170 ;
        RECT 1528.450 600.000 1528.730 600.030 ;
        RECT 1530.120 593.290 1530.260 600.030 ;
        RECT 1530.060 592.970 1530.320 593.290 ;
        RECT 1664.380 592.970 1664.640 593.290 ;
        RECT 1664.440 3.050 1664.580 592.970 ;
        RECT 1664.380 2.730 1664.640 3.050 ;
        RECT 1668.060 2.730 1668.320 3.050 ;
        RECT 1668.120 2.400 1668.260 2.730 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1538.310 591.160 1538.630 591.220 ;
        RECT 1684.590 591.160 1684.910 591.220 ;
        RECT 1538.310 591.020 1684.910 591.160 ;
        RECT 1538.310 590.960 1538.630 591.020 ;
        RECT 1684.590 590.960 1684.910 591.020 ;
        RECT 1684.590 2.960 1684.910 3.020 ;
        RECT 1685.510 2.960 1685.830 3.020 ;
        RECT 1684.590 2.820 1685.830 2.960 ;
        RECT 1684.590 2.760 1684.910 2.820 ;
        RECT 1685.510 2.760 1685.830 2.820 ;
      LAYER via ;
        RECT 1538.340 590.960 1538.600 591.220 ;
        RECT 1684.620 590.960 1684.880 591.220 ;
        RECT 1684.620 2.760 1684.880 3.020 ;
        RECT 1685.540 2.760 1685.800 3.020 ;
      LAYER met2 ;
        RECT 1537.650 600.170 1537.930 604.000 ;
        RECT 1537.650 600.030 1538.540 600.170 ;
        RECT 1537.650 600.000 1537.930 600.030 ;
        RECT 1538.400 591.250 1538.540 600.030 ;
        RECT 1538.340 590.930 1538.600 591.250 ;
        RECT 1684.620 590.930 1684.880 591.250 ;
        RECT 1684.680 3.050 1684.820 590.930 ;
        RECT 1684.620 2.730 1684.880 3.050 ;
        RECT 1685.540 2.730 1685.800 3.050 ;
        RECT 1685.600 2.400 1685.740 2.730 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1043.350 110.540 1043.670 110.800 ;
        RECT 1043.440 110.120 1043.580 110.540 ;
        RECT 1043.350 109.860 1043.670 110.120 ;
        RECT 1007.470 17.920 1007.790 17.980 ;
        RECT 1042.890 17.920 1043.210 17.980 ;
        RECT 1007.470 17.780 1043.210 17.920 ;
        RECT 1007.470 17.720 1007.790 17.780 ;
        RECT 1042.890 17.720 1043.210 17.780 ;
        RECT 722.270 17.240 722.590 17.300 ;
        RECT 1007.470 17.240 1007.790 17.300 ;
        RECT 722.270 17.100 1007.790 17.240 ;
        RECT 722.270 17.040 722.590 17.100 ;
        RECT 1007.470 17.040 1007.790 17.100 ;
      LAYER via ;
        RECT 1043.380 110.540 1043.640 110.800 ;
        RECT 1043.380 109.860 1043.640 110.120 ;
        RECT 1007.500 17.720 1007.760 17.980 ;
        RECT 1042.920 17.720 1043.180 17.980 ;
        RECT 722.300 17.040 722.560 17.300 ;
        RECT 1007.500 17.040 1007.760 17.300 ;
      LAYER met2 ;
        RECT 1041.770 600.170 1042.050 604.000 ;
        RECT 1041.770 600.030 1043.580 600.170 ;
        RECT 1041.770 600.000 1042.050 600.030 ;
        RECT 1043.440 110.830 1043.580 600.030 ;
        RECT 1043.380 110.510 1043.640 110.830 ;
        RECT 1043.380 109.830 1043.640 110.150 ;
        RECT 1043.440 24.890 1043.580 109.830 ;
        RECT 1042.980 24.750 1043.580 24.890 ;
        RECT 1042.980 18.010 1043.120 24.750 ;
        RECT 1007.500 17.690 1007.760 18.010 ;
        RECT 1042.920 17.690 1043.180 18.010 ;
        RECT 1007.560 17.330 1007.700 17.690 ;
        RECT 722.300 17.010 722.560 17.330 ;
        RECT 1007.500 17.010 1007.760 17.330 ;
        RECT 722.360 2.400 722.500 17.010 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1548.430 592.180 1548.750 592.240 ;
        RECT 1697.930 592.180 1698.250 592.240 ;
        RECT 1548.430 592.040 1698.250 592.180 ;
        RECT 1548.430 591.980 1548.750 592.040 ;
        RECT 1697.930 591.980 1698.250 592.040 ;
        RECT 1697.930 62.120 1698.250 62.180 ;
        RECT 1702.990 62.120 1703.310 62.180 ;
        RECT 1697.930 61.980 1703.310 62.120 ;
        RECT 1697.930 61.920 1698.250 61.980 ;
        RECT 1702.990 61.920 1703.310 61.980 ;
      LAYER via ;
        RECT 1548.460 591.980 1548.720 592.240 ;
        RECT 1697.960 591.980 1698.220 592.240 ;
        RECT 1697.960 61.920 1698.220 62.180 ;
        RECT 1703.020 61.920 1703.280 62.180 ;
      LAYER met2 ;
        RECT 1546.850 600.170 1547.130 604.000 ;
        RECT 1546.850 600.030 1548.660 600.170 ;
        RECT 1546.850 600.000 1547.130 600.030 ;
        RECT 1548.520 592.270 1548.660 600.030 ;
        RECT 1548.460 591.950 1548.720 592.270 ;
        RECT 1697.960 591.950 1698.220 592.270 ;
        RECT 1698.020 62.210 1698.160 591.950 ;
        RECT 1697.960 61.890 1698.220 62.210 ;
        RECT 1703.020 61.890 1703.280 62.210 ;
        RECT 1703.080 26.250 1703.220 61.890 ;
        RECT 1703.080 26.110 1703.680 26.250 ;
        RECT 1703.540 2.400 1703.680 26.110 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1557.630 591.840 1557.950 591.900 ;
        RECT 1719.550 591.840 1719.870 591.900 ;
        RECT 1557.630 591.700 1719.870 591.840 ;
        RECT 1557.630 591.640 1557.950 591.700 ;
        RECT 1719.550 591.640 1719.870 591.700 ;
        RECT 1719.550 2.960 1719.870 3.020 ;
        RECT 1721.390 2.960 1721.710 3.020 ;
        RECT 1719.550 2.820 1721.710 2.960 ;
        RECT 1719.550 2.760 1719.870 2.820 ;
        RECT 1721.390 2.760 1721.710 2.820 ;
      LAYER via ;
        RECT 1557.660 591.640 1557.920 591.900 ;
        RECT 1719.580 591.640 1719.840 591.900 ;
        RECT 1719.580 2.760 1719.840 3.020 ;
        RECT 1721.420 2.760 1721.680 3.020 ;
      LAYER met2 ;
        RECT 1556.050 600.170 1556.330 604.000 ;
        RECT 1556.050 600.030 1557.860 600.170 ;
        RECT 1556.050 600.000 1556.330 600.030 ;
        RECT 1557.720 591.930 1557.860 600.030 ;
        RECT 1557.660 591.610 1557.920 591.930 ;
        RECT 1719.580 591.610 1719.840 591.930 ;
        RECT 1719.640 3.050 1719.780 591.610 ;
        RECT 1719.580 2.730 1719.840 3.050 ;
        RECT 1721.420 2.730 1721.680 3.050 ;
        RECT 1721.480 2.400 1721.620 2.730 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1565.450 24.040 1565.770 24.100 ;
        RECT 1739.330 24.040 1739.650 24.100 ;
        RECT 1565.450 23.900 1739.650 24.040 ;
        RECT 1565.450 23.840 1565.770 23.900 ;
        RECT 1739.330 23.840 1739.650 23.900 ;
      LAYER via ;
        RECT 1565.480 23.840 1565.740 24.100 ;
        RECT 1739.360 23.840 1739.620 24.100 ;
      LAYER met2 ;
        RECT 1565.250 600.000 1565.530 604.000 ;
        RECT 1565.310 598.810 1565.450 600.000 ;
        RECT 1565.310 598.670 1565.680 598.810 ;
        RECT 1565.540 24.130 1565.680 598.670 ;
        RECT 1565.480 23.810 1565.740 24.130 ;
        RECT 1739.360 23.810 1739.620 24.130 ;
        RECT 1739.420 2.400 1739.560 23.810 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1576.030 586.740 1576.350 586.800 ;
        RECT 1579.250 586.740 1579.570 586.800 ;
        RECT 1576.030 586.600 1579.570 586.740 ;
        RECT 1576.030 586.540 1576.350 586.600 ;
        RECT 1579.250 586.540 1579.570 586.600 ;
        RECT 1579.250 29.480 1579.570 29.540 ;
        RECT 1756.810 29.480 1757.130 29.540 ;
        RECT 1579.250 29.340 1757.130 29.480 ;
        RECT 1579.250 29.280 1579.570 29.340 ;
        RECT 1756.810 29.280 1757.130 29.340 ;
      LAYER via ;
        RECT 1576.060 586.540 1576.320 586.800 ;
        RECT 1579.280 586.540 1579.540 586.800 ;
        RECT 1579.280 29.280 1579.540 29.540 ;
        RECT 1756.840 29.280 1757.100 29.540 ;
      LAYER met2 ;
        RECT 1574.450 600.170 1574.730 604.000 ;
        RECT 1574.450 600.030 1576.260 600.170 ;
        RECT 1574.450 600.000 1574.730 600.030 ;
        RECT 1576.120 586.830 1576.260 600.030 ;
        RECT 1576.060 586.510 1576.320 586.830 ;
        RECT 1579.280 586.510 1579.540 586.830 ;
        RECT 1579.340 29.570 1579.480 586.510 ;
        RECT 1579.280 29.250 1579.540 29.570 ;
        RECT 1756.840 29.250 1757.100 29.570 ;
        RECT 1756.900 2.400 1757.040 29.250 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1585.690 30.160 1586.010 30.220 ;
        RECT 1774.750 30.160 1775.070 30.220 ;
        RECT 1585.690 30.020 1775.070 30.160 ;
        RECT 1585.690 29.960 1586.010 30.020 ;
        RECT 1774.750 29.960 1775.070 30.020 ;
      LAYER via ;
        RECT 1585.720 29.960 1585.980 30.220 ;
        RECT 1774.780 29.960 1775.040 30.220 ;
      LAYER met2 ;
        RECT 1583.650 600.170 1583.930 604.000 ;
        RECT 1583.650 600.030 1585.920 600.170 ;
        RECT 1583.650 600.000 1583.930 600.030 ;
        RECT 1585.780 30.250 1585.920 600.030 ;
        RECT 1585.720 29.930 1585.980 30.250 ;
        RECT 1774.780 29.930 1775.040 30.250 ;
        RECT 1774.840 2.400 1774.980 29.930 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.510 30.500 1593.830 30.560 ;
        RECT 1792.690 30.500 1793.010 30.560 ;
        RECT 1593.510 30.360 1793.010 30.500 ;
        RECT 1593.510 30.300 1593.830 30.360 ;
        RECT 1792.690 30.300 1793.010 30.360 ;
      LAYER via ;
        RECT 1593.540 30.300 1593.800 30.560 ;
        RECT 1792.720 30.300 1792.980 30.560 ;
      LAYER met2 ;
        RECT 1592.850 600.170 1593.130 604.000 ;
        RECT 1592.850 600.030 1593.740 600.170 ;
        RECT 1592.850 600.000 1593.130 600.030 ;
        RECT 1593.600 30.590 1593.740 600.030 ;
        RECT 1593.540 30.270 1593.800 30.590 ;
        RECT 1792.720 30.270 1792.980 30.590 ;
        RECT 1792.780 2.400 1792.920 30.270 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1603.630 586.740 1603.950 586.800 ;
        RECT 1606.850 586.740 1607.170 586.800 ;
        RECT 1603.630 586.600 1607.170 586.740 ;
        RECT 1603.630 586.540 1603.950 586.600 ;
        RECT 1606.850 586.540 1607.170 586.600 ;
        RECT 1606.850 20.980 1607.170 21.040 ;
        RECT 1810.630 20.980 1810.950 21.040 ;
        RECT 1606.850 20.840 1810.950 20.980 ;
        RECT 1606.850 20.780 1607.170 20.840 ;
        RECT 1810.630 20.780 1810.950 20.840 ;
      LAYER via ;
        RECT 1603.660 586.540 1603.920 586.800 ;
        RECT 1606.880 586.540 1607.140 586.800 ;
        RECT 1606.880 20.780 1607.140 21.040 ;
        RECT 1810.660 20.780 1810.920 21.040 ;
      LAYER met2 ;
        RECT 1602.050 600.170 1602.330 604.000 ;
        RECT 1602.050 600.030 1603.860 600.170 ;
        RECT 1602.050 600.000 1602.330 600.030 ;
        RECT 1603.720 586.830 1603.860 600.030 ;
        RECT 1603.660 586.510 1603.920 586.830 ;
        RECT 1606.880 586.510 1607.140 586.830 ;
        RECT 1606.940 21.070 1607.080 586.510 ;
        RECT 1606.880 20.750 1607.140 21.070 ;
        RECT 1810.660 20.750 1810.920 21.070 ;
        RECT 1810.720 2.400 1810.860 20.750 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1611.910 579.940 1612.230 580.000 ;
        RECT 1612.830 579.940 1613.150 580.000 ;
        RECT 1611.910 579.800 1613.150 579.940 ;
        RECT 1611.910 579.740 1612.230 579.800 ;
        RECT 1612.830 579.740 1613.150 579.800 ;
        RECT 1613.290 531.320 1613.610 531.380 ;
        RECT 1613.750 531.320 1614.070 531.380 ;
        RECT 1613.290 531.180 1614.070 531.320 ;
        RECT 1613.290 531.120 1613.610 531.180 ;
        RECT 1613.750 531.120 1614.070 531.180 ;
        RECT 1613.750 496.980 1614.070 497.040 ;
        RECT 1613.380 496.840 1614.070 496.980 ;
        RECT 1613.380 496.700 1613.520 496.840 ;
        RECT 1613.750 496.780 1614.070 496.840 ;
        RECT 1613.290 496.440 1613.610 496.700 ;
        RECT 1612.830 448.700 1613.150 448.760 ;
        RECT 1613.750 448.700 1614.070 448.760 ;
        RECT 1612.830 448.560 1614.070 448.700 ;
        RECT 1612.830 448.500 1613.150 448.560 ;
        RECT 1613.750 448.500 1614.070 448.560 ;
        RECT 1612.370 434.760 1612.690 434.820 ;
        RECT 1613.290 434.760 1613.610 434.820 ;
        RECT 1612.370 434.620 1613.610 434.760 ;
        RECT 1612.370 434.560 1612.690 434.620 ;
        RECT 1613.290 434.560 1613.610 434.620 ;
        RECT 1612.370 386.480 1612.690 386.540 ;
        RECT 1613.750 386.480 1614.070 386.540 ;
        RECT 1612.370 386.340 1614.070 386.480 ;
        RECT 1612.370 386.280 1612.690 386.340 ;
        RECT 1613.750 386.280 1614.070 386.340 ;
        RECT 1613.290 331.400 1613.610 331.460 ;
        RECT 1613.750 331.400 1614.070 331.460 ;
        RECT 1613.290 331.260 1614.070 331.400 ;
        RECT 1613.290 331.200 1613.610 331.260 ;
        RECT 1613.750 331.200 1614.070 331.260 ;
        RECT 1612.370 289.580 1612.690 289.640 ;
        RECT 1613.750 289.580 1614.070 289.640 ;
        RECT 1612.370 289.440 1614.070 289.580 ;
        RECT 1612.370 289.380 1612.690 289.440 ;
        RECT 1613.750 289.380 1614.070 289.440 ;
        RECT 1612.370 193.020 1612.690 193.080 ;
        RECT 1613.750 193.020 1614.070 193.080 ;
        RECT 1612.370 192.880 1614.070 193.020 ;
        RECT 1612.370 192.820 1612.690 192.880 ;
        RECT 1613.750 192.820 1614.070 192.880 ;
        RECT 1612.830 21.320 1613.150 21.380 ;
        RECT 1828.570 21.320 1828.890 21.380 ;
        RECT 1612.830 21.180 1828.890 21.320 ;
        RECT 1612.830 21.120 1613.150 21.180 ;
        RECT 1828.570 21.120 1828.890 21.180 ;
      LAYER via ;
        RECT 1611.940 579.740 1612.200 580.000 ;
        RECT 1612.860 579.740 1613.120 580.000 ;
        RECT 1613.320 531.120 1613.580 531.380 ;
        RECT 1613.780 531.120 1614.040 531.380 ;
        RECT 1613.780 496.780 1614.040 497.040 ;
        RECT 1613.320 496.440 1613.580 496.700 ;
        RECT 1612.860 448.500 1613.120 448.760 ;
        RECT 1613.780 448.500 1614.040 448.760 ;
        RECT 1612.400 434.560 1612.660 434.820 ;
        RECT 1613.320 434.560 1613.580 434.820 ;
        RECT 1612.400 386.280 1612.660 386.540 ;
        RECT 1613.780 386.280 1614.040 386.540 ;
        RECT 1613.320 331.200 1613.580 331.460 ;
        RECT 1613.780 331.200 1614.040 331.460 ;
        RECT 1612.400 289.380 1612.660 289.640 ;
        RECT 1613.780 289.380 1614.040 289.640 ;
        RECT 1612.400 192.820 1612.660 193.080 ;
        RECT 1613.780 192.820 1614.040 193.080 ;
        RECT 1612.860 21.120 1613.120 21.380 ;
        RECT 1828.600 21.120 1828.860 21.380 ;
      LAYER met2 ;
        RECT 1611.250 600.170 1611.530 604.000 ;
        RECT 1611.250 600.030 1612.140 600.170 ;
        RECT 1611.250 600.000 1611.530 600.030 ;
        RECT 1612.000 580.030 1612.140 600.030 ;
        RECT 1611.940 579.710 1612.200 580.030 ;
        RECT 1612.860 579.710 1613.120 580.030 ;
        RECT 1612.920 545.090 1613.060 579.710 ;
        RECT 1612.920 544.950 1613.520 545.090 ;
        RECT 1613.380 531.410 1613.520 544.950 ;
        RECT 1613.320 531.090 1613.580 531.410 ;
        RECT 1613.780 531.090 1614.040 531.410 ;
        RECT 1613.840 497.070 1613.980 531.090 ;
        RECT 1613.780 496.750 1614.040 497.070 ;
        RECT 1613.320 496.410 1613.580 496.730 ;
        RECT 1613.380 483.210 1613.520 496.410 ;
        RECT 1613.380 483.070 1613.980 483.210 ;
        RECT 1613.840 448.790 1613.980 483.070 ;
        RECT 1612.860 448.530 1613.120 448.790 ;
        RECT 1612.860 448.470 1613.520 448.530 ;
        RECT 1613.780 448.470 1614.040 448.790 ;
        RECT 1612.920 448.390 1613.520 448.470 ;
        RECT 1613.380 434.850 1613.520 448.390 ;
        RECT 1612.400 434.530 1612.660 434.850 ;
        RECT 1613.320 434.530 1613.580 434.850 ;
        RECT 1612.460 386.570 1612.600 434.530 ;
        RECT 1612.400 386.250 1612.660 386.570 ;
        RECT 1613.780 386.250 1614.040 386.570 ;
        RECT 1613.840 331.490 1613.980 386.250 ;
        RECT 1613.320 331.170 1613.580 331.490 ;
        RECT 1613.780 331.170 1614.040 331.490 ;
        RECT 1613.380 303.690 1613.520 331.170 ;
        RECT 1613.380 303.550 1613.980 303.690 ;
        RECT 1613.840 289.670 1613.980 303.550 ;
        RECT 1612.400 289.350 1612.660 289.670 ;
        RECT 1613.780 289.350 1614.040 289.670 ;
        RECT 1612.460 254.730 1612.600 289.350 ;
        RECT 1612.460 254.590 1613.520 254.730 ;
        RECT 1613.380 207.130 1613.520 254.590 ;
        RECT 1613.380 206.990 1613.980 207.130 ;
        RECT 1613.840 193.110 1613.980 206.990 ;
        RECT 1612.400 192.790 1612.660 193.110 ;
        RECT 1613.780 192.790 1614.040 193.110 ;
        RECT 1612.460 158.170 1612.600 192.790 ;
        RECT 1612.460 158.030 1613.520 158.170 ;
        RECT 1613.380 110.570 1613.520 158.030 ;
        RECT 1613.380 110.430 1613.980 110.570 ;
        RECT 1613.840 62.290 1613.980 110.430 ;
        RECT 1612.920 62.150 1613.980 62.290 ;
        RECT 1612.920 21.410 1613.060 62.150 ;
        RECT 1612.860 21.090 1613.120 21.410 ;
        RECT 1828.600 21.090 1828.860 21.410 ;
        RECT 1828.660 2.400 1828.800 21.090 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1620.650 21.660 1620.970 21.720 ;
        RECT 1846.050 21.660 1846.370 21.720 ;
        RECT 1620.650 21.520 1846.370 21.660 ;
        RECT 1620.650 21.460 1620.970 21.520 ;
        RECT 1846.050 21.460 1846.370 21.520 ;
      LAYER via ;
        RECT 1620.680 21.460 1620.940 21.720 ;
        RECT 1846.080 21.460 1846.340 21.720 ;
      LAYER met2 ;
        RECT 1620.450 600.000 1620.730 604.000 ;
        RECT 1620.510 598.810 1620.650 600.000 ;
        RECT 1620.510 598.670 1620.880 598.810 ;
        RECT 1620.740 21.750 1620.880 598.670 ;
        RECT 1620.680 21.430 1620.940 21.750 ;
        RECT 1846.080 21.430 1846.340 21.750 ;
        RECT 1846.140 2.400 1846.280 21.430 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1631.230 586.740 1631.550 586.800 ;
        RECT 1634.910 586.740 1635.230 586.800 ;
        RECT 1631.230 586.600 1635.230 586.740 ;
        RECT 1631.230 586.540 1631.550 586.600 ;
        RECT 1634.910 586.540 1635.230 586.600 ;
        RECT 1634.910 22.000 1635.230 22.060 ;
        RECT 1863.990 22.000 1864.310 22.060 ;
        RECT 1634.910 21.860 1864.310 22.000 ;
        RECT 1634.910 21.800 1635.230 21.860 ;
        RECT 1863.990 21.800 1864.310 21.860 ;
      LAYER via ;
        RECT 1631.260 586.540 1631.520 586.800 ;
        RECT 1634.940 586.540 1635.200 586.800 ;
        RECT 1634.940 21.800 1635.200 22.060 ;
        RECT 1864.020 21.800 1864.280 22.060 ;
      LAYER met2 ;
        RECT 1629.650 600.170 1629.930 604.000 ;
        RECT 1629.650 600.030 1631.460 600.170 ;
        RECT 1629.650 600.000 1629.930 600.030 ;
        RECT 1631.320 586.830 1631.460 600.030 ;
        RECT 1631.260 586.510 1631.520 586.830 ;
        RECT 1634.940 586.510 1635.200 586.830 ;
        RECT 1635.000 22.090 1635.140 586.510 ;
        RECT 1634.940 21.770 1635.200 22.090 ;
        RECT 1864.020 21.770 1864.280 22.090 ;
        RECT 1864.080 2.400 1864.220 21.770 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 740.210 14.180 740.530 14.240 ;
        RECT 1049.790 14.180 1050.110 14.240 ;
        RECT 740.210 14.040 1050.110 14.180 ;
        RECT 740.210 13.980 740.530 14.040 ;
        RECT 1049.790 13.980 1050.110 14.040 ;
      LAYER via ;
        RECT 740.240 13.980 740.500 14.240 ;
        RECT 1049.820 13.980 1050.080 14.240 ;
      LAYER met2 ;
        RECT 1050.970 600.170 1051.250 604.000 ;
        RECT 1049.880 600.030 1051.250 600.170 ;
        RECT 1049.880 14.270 1050.020 600.030 ;
        RECT 1050.970 600.000 1051.250 600.030 ;
        RECT 740.240 13.950 740.500 14.270 ;
        RECT 1049.820 13.950 1050.080 14.270 ;
        RECT 740.300 2.400 740.440 13.950 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1640.430 587.420 1640.750 587.480 ;
        RECT 1641.350 587.420 1641.670 587.480 ;
        RECT 1640.430 587.280 1641.670 587.420 ;
        RECT 1640.430 587.220 1640.750 587.280 ;
        RECT 1641.350 587.220 1641.670 587.280 ;
        RECT 1641.350 22.340 1641.670 22.400 ;
        RECT 1881.930 22.340 1882.250 22.400 ;
        RECT 1641.350 22.200 1882.250 22.340 ;
        RECT 1641.350 22.140 1641.670 22.200 ;
        RECT 1881.930 22.140 1882.250 22.200 ;
      LAYER via ;
        RECT 1640.460 587.220 1640.720 587.480 ;
        RECT 1641.380 587.220 1641.640 587.480 ;
        RECT 1641.380 22.140 1641.640 22.400 ;
        RECT 1881.960 22.140 1882.220 22.400 ;
      LAYER met2 ;
        RECT 1638.850 600.170 1639.130 604.000 ;
        RECT 1638.850 600.030 1640.660 600.170 ;
        RECT 1638.850 600.000 1639.130 600.030 ;
        RECT 1640.520 587.510 1640.660 600.030 ;
        RECT 1640.460 587.190 1640.720 587.510 ;
        RECT 1641.380 587.190 1641.640 587.510 ;
        RECT 1641.440 22.430 1641.580 587.190 ;
        RECT 1641.380 22.110 1641.640 22.430 ;
        RECT 1881.960 22.110 1882.220 22.430 ;
        RECT 1882.020 2.400 1882.160 22.110 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1648.710 22.680 1649.030 22.740 ;
        RECT 1899.870 22.680 1900.190 22.740 ;
        RECT 1648.710 22.540 1900.190 22.680 ;
        RECT 1648.710 22.480 1649.030 22.540 ;
        RECT 1899.870 22.480 1900.190 22.540 ;
      LAYER via ;
        RECT 1648.740 22.480 1649.000 22.740 ;
        RECT 1899.900 22.480 1900.160 22.740 ;
      LAYER met2 ;
        RECT 1647.590 600.170 1647.870 604.000 ;
        RECT 1647.590 600.030 1648.940 600.170 ;
        RECT 1647.590 600.000 1647.870 600.030 ;
        RECT 1648.800 22.770 1648.940 600.030 ;
        RECT 1648.740 22.450 1649.000 22.770 ;
        RECT 1899.900 22.450 1900.160 22.770 ;
        RECT 1899.960 2.400 1900.100 22.450 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1658.370 586.740 1658.690 586.800 ;
        RECT 1662.510 586.740 1662.830 586.800 ;
        RECT 1658.370 586.600 1662.830 586.740 ;
        RECT 1658.370 586.540 1658.690 586.600 ;
        RECT 1662.510 586.540 1662.830 586.600 ;
        RECT 1662.510 23.020 1662.830 23.080 ;
        RECT 1917.810 23.020 1918.130 23.080 ;
        RECT 1662.510 22.880 1918.130 23.020 ;
        RECT 1662.510 22.820 1662.830 22.880 ;
        RECT 1917.810 22.820 1918.130 22.880 ;
      LAYER via ;
        RECT 1658.400 586.540 1658.660 586.800 ;
        RECT 1662.540 586.540 1662.800 586.800 ;
        RECT 1662.540 22.820 1662.800 23.080 ;
        RECT 1917.840 22.820 1918.100 23.080 ;
      LAYER met2 ;
        RECT 1656.790 600.170 1657.070 604.000 ;
        RECT 1656.790 600.030 1658.600 600.170 ;
        RECT 1656.790 600.000 1657.070 600.030 ;
        RECT 1658.460 586.830 1658.600 600.030 ;
        RECT 1658.400 586.510 1658.660 586.830 ;
        RECT 1662.540 586.510 1662.800 586.830 ;
        RECT 1662.600 23.110 1662.740 586.510 ;
        RECT 1662.540 22.790 1662.800 23.110 ;
        RECT 1917.840 22.790 1918.100 23.110 ;
        RECT 1917.900 2.400 1918.040 22.790 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1667.570 586.740 1667.890 586.800 ;
        RECT 1668.950 586.740 1669.270 586.800 ;
        RECT 1667.570 586.600 1669.270 586.740 ;
        RECT 1667.570 586.540 1667.890 586.600 ;
        RECT 1668.950 586.540 1669.270 586.600 ;
        RECT 1668.950 23.360 1669.270 23.420 ;
        RECT 1935.290 23.360 1935.610 23.420 ;
        RECT 1668.950 23.220 1935.610 23.360 ;
        RECT 1668.950 23.160 1669.270 23.220 ;
        RECT 1935.290 23.160 1935.610 23.220 ;
      LAYER via ;
        RECT 1667.600 586.540 1667.860 586.800 ;
        RECT 1668.980 586.540 1669.240 586.800 ;
        RECT 1668.980 23.160 1669.240 23.420 ;
        RECT 1935.320 23.160 1935.580 23.420 ;
      LAYER met2 ;
        RECT 1665.990 600.170 1666.270 604.000 ;
        RECT 1665.990 600.030 1667.800 600.170 ;
        RECT 1665.990 600.000 1666.270 600.030 ;
        RECT 1667.660 586.830 1667.800 600.030 ;
        RECT 1667.600 586.510 1667.860 586.830 ;
        RECT 1668.980 586.510 1669.240 586.830 ;
        RECT 1669.040 23.450 1669.180 586.510 ;
        RECT 1668.980 23.130 1669.240 23.450 ;
        RECT 1935.320 23.130 1935.580 23.450 ;
        RECT 1935.380 2.400 1935.520 23.130 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1675.850 27.440 1676.170 27.500 ;
        RECT 1953.230 27.440 1953.550 27.500 ;
        RECT 1675.850 27.300 1953.550 27.440 ;
        RECT 1675.850 27.240 1676.170 27.300 ;
        RECT 1953.230 27.240 1953.550 27.300 ;
      LAYER via ;
        RECT 1675.880 27.240 1676.140 27.500 ;
        RECT 1953.260 27.240 1953.520 27.500 ;
      LAYER met2 ;
        RECT 1675.190 600.170 1675.470 604.000 ;
        RECT 1675.190 600.030 1676.080 600.170 ;
        RECT 1675.190 600.000 1675.470 600.030 ;
        RECT 1675.940 27.530 1676.080 600.030 ;
        RECT 1675.880 27.210 1676.140 27.530 ;
        RECT 1953.260 27.210 1953.520 27.530 ;
        RECT 1953.320 2.400 1953.460 27.210 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.970 586.740 1686.290 586.800 ;
        RECT 1690.110 586.740 1690.430 586.800 ;
        RECT 1685.970 586.600 1690.430 586.740 ;
        RECT 1685.970 586.540 1686.290 586.600 ;
        RECT 1690.110 586.540 1690.430 586.600 ;
        RECT 1690.110 23.700 1690.430 23.760 ;
        RECT 1971.170 23.700 1971.490 23.760 ;
        RECT 1690.110 23.560 1971.490 23.700 ;
        RECT 1690.110 23.500 1690.430 23.560 ;
        RECT 1971.170 23.500 1971.490 23.560 ;
      LAYER via ;
        RECT 1686.000 586.540 1686.260 586.800 ;
        RECT 1690.140 586.540 1690.400 586.800 ;
        RECT 1690.140 23.500 1690.400 23.760 ;
        RECT 1971.200 23.500 1971.460 23.760 ;
      LAYER met2 ;
        RECT 1684.390 600.170 1684.670 604.000 ;
        RECT 1684.390 600.030 1686.200 600.170 ;
        RECT 1684.390 600.000 1684.670 600.030 ;
        RECT 1686.060 586.830 1686.200 600.030 ;
        RECT 1686.000 586.510 1686.260 586.830 ;
        RECT 1690.140 586.510 1690.400 586.830 ;
        RECT 1690.200 23.790 1690.340 586.510 ;
        RECT 1690.140 23.470 1690.400 23.790 ;
        RECT 1971.200 23.470 1971.460 23.790 ;
        RECT 1971.260 2.400 1971.400 23.470 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1695.170 586.740 1695.490 586.800 ;
        RECT 1697.010 586.740 1697.330 586.800 ;
        RECT 1695.170 586.600 1697.330 586.740 ;
        RECT 1695.170 586.540 1695.490 586.600 ;
        RECT 1697.010 586.540 1697.330 586.600 ;
        RECT 1697.010 27.100 1697.330 27.160 ;
        RECT 1989.110 27.100 1989.430 27.160 ;
        RECT 1697.010 26.960 1989.430 27.100 ;
        RECT 1697.010 26.900 1697.330 26.960 ;
        RECT 1989.110 26.900 1989.430 26.960 ;
      LAYER via ;
        RECT 1695.200 586.540 1695.460 586.800 ;
        RECT 1697.040 586.540 1697.300 586.800 ;
        RECT 1697.040 26.900 1697.300 27.160 ;
        RECT 1989.140 26.900 1989.400 27.160 ;
      LAYER met2 ;
        RECT 1693.590 600.170 1693.870 604.000 ;
        RECT 1693.590 600.030 1695.400 600.170 ;
        RECT 1693.590 600.000 1693.870 600.030 ;
        RECT 1695.260 586.830 1695.400 600.030 ;
        RECT 1695.200 586.510 1695.460 586.830 ;
        RECT 1697.040 586.510 1697.300 586.830 ;
        RECT 1697.100 27.190 1697.240 586.510 ;
        RECT 1697.040 26.870 1697.300 27.190 ;
        RECT 1989.140 26.870 1989.400 27.190 ;
        RECT 1989.200 2.400 1989.340 26.870 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.450 26.760 1703.770 26.820 ;
        RECT 2006.590 26.760 2006.910 26.820 ;
        RECT 1703.450 26.620 2006.910 26.760 ;
        RECT 1703.450 26.560 1703.770 26.620 ;
        RECT 2006.590 26.560 2006.910 26.620 ;
      LAYER via ;
        RECT 1703.480 26.560 1703.740 26.820 ;
        RECT 2006.620 26.560 2006.880 26.820 ;
      LAYER met2 ;
        RECT 1702.790 600.170 1703.070 604.000 ;
        RECT 1702.790 600.030 1703.680 600.170 ;
        RECT 1702.790 600.000 1703.070 600.030 ;
        RECT 1703.540 26.850 1703.680 600.030 ;
        RECT 1703.480 26.530 1703.740 26.850 ;
        RECT 2006.620 26.530 2006.880 26.850 ;
        RECT 2006.680 2.400 2006.820 26.530 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1713.570 586.740 1713.890 586.800 ;
        RECT 1717.710 586.740 1718.030 586.800 ;
        RECT 1713.570 586.600 1718.030 586.740 ;
        RECT 1713.570 586.540 1713.890 586.600 ;
        RECT 1717.710 586.540 1718.030 586.600 ;
        RECT 1717.710 26.420 1718.030 26.480 ;
        RECT 2024.530 26.420 2024.850 26.480 ;
        RECT 1717.710 26.280 2024.850 26.420 ;
        RECT 1717.710 26.220 1718.030 26.280 ;
        RECT 2024.530 26.220 2024.850 26.280 ;
      LAYER via ;
        RECT 1713.600 586.540 1713.860 586.800 ;
        RECT 1717.740 586.540 1718.000 586.800 ;
        RECT 1717.740 26.220 1718.000 26.480 ;
        RECT 2024.560 26.220 2024.820 26.480 ;
      LAYER met2 ;
        RECT 1711.990 600.170 1712.270 604.000 ;
        RECT 1711.990 600.030 1713.800 600.170 ;
        RECT 1711.990 600.000 1712.270 600.030 ;
        RECT 1713.660 586.830 1713.800 600.030 ;
        RECT 1713.600 586.510 1713.860 586.830 ;
        RECT 1717.740 586.510 1718.000 586.830 ;
        RECT 1717.800 26.510 1717.940 586.510 ;
        RECT 1717.740 26.190 1718.000 26.510 ;
        RECT 2024.560 26.190 2024.820 26.510 ;
        RECT 2024.620 2.400 2024.760 26.190 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1722.770 586.740 1723.090 586.800 ;
        RECT 1724.150 586.740 1724.470 586.800 ;
        RECT 1722.770 586.600 1724.470 586.740 ;
        RECT 1722.770 586.540 1723.090 586.600 ;
        RECT 1724.150 586.540 1724.470 586.600 ;
        RECT 1724.150 26.080 1724.470 26.140 ;
        RECT 2043.390 26.080 2043.710 26.140 ;
        RECT 1724.150 25.940 2043.710 26.080 ;
        RECT 1724.150 25.880 1724.470 25.940 ;
        RECT 2043.390 25.880 2043.710 25.940 ;
      LAYER via ;
        RECT 1722.800 586.540 1723.060 586.800 ;
        RECT 1724.180 586.540 1724.440 586.800 ;
        RECT 1724.180 25.880 1724.440 26.140 ;
        RECT 2043.420 25.880 2043.680 26.140 ;
      LAYER met2 ;
        RECT 1721.190 600.170 1721.470 604.000 ;
        RECT 1721.190 600.030 1723.000 600.170 ;
        RECT 1721.190 600.000 1721.470 600.030 ;
        RECT 1722.860 586.830 1723.000 600.030 ;
        RECT 1722.800 586.510 1723.060 586.830 ;
        RECT 1724.180 586.510 1724.440 586.830 ;
        RECT 1724.240 26.170 1724.380 586.510 ;
        RECT 1724.180 25.850 1724.440 26.170 ;
        RECT 2043.420 25.850 2043.680 26.170 ;
        RECT 2043.480 17.410 2043.620 25.850 ;
        RECT 2042.560 17.270 2043.620 17.410 ;
        RECT 2042.560 2.400 2042.700 17.270 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1055.770 569.400 1056.090 569.460 ;
        RECT 1058.530 569.400 1058.850 569.460 ;
        RECT 1055.770 569.260 1058.850 569.400 ;
        RECT 1055.770 569.200 1056.090 569.260 ;
        RECT 1058.530 569.200 1058.850 569.260 ;
        RECT 858.430 27.440 858.750 27.500 ;
        RECT 1055.770 27.440 1056.090 27.500 ;
        RECT 858.430 27.300 1056.090 27.440 ;
        RECT 858.430 27.240 858.750 27.300 ;
        RECT 1055.770 27.240 1056.090 27.300 ;
        RECT 757.690 18.940 758.010 19.000 ;
        RECT 858.430 18.940 858.750 19.000 ;
        RECT 757.690 18.800 858.750 18.940 ;
        RECT 757.690 18.740 758.010 18.800 ;
        RECT 858.430 18.740 858.750 18.800 ;
      LAYER via ;
        RECT 1055.800 569.200 1056.060 569.460 ;
        RECT 1058.560 569.200 1058.820 569.460 ;
        RECT 858.460 27.240 858.720 27.500 ;
        RECT 1055.800 27.240 1056.060 27.500 ;
        RECT 757.720 18.740 757.980 19.000 ;
        RECT 858.460 18.740 858.720 19.000 ;
      LAYER met2 ;
        RECT 1060.170 600.170 1060.450 604.000 ;
        RECT 1058.620 600.030 1060.450 600.170 ;
        RECT 1058.620 569.490 1058.760 600.030 ;
        RECT 1060.170 600.000 1060.450 600.030 ;
        RECT 1055.800 569.170 1056.060 569.490 ;
        RECT 1058.560 569.170 1058.820 569.490 ;
        RECT 1055.860 27.530 1056.000 569.170 ;
        RECT 858.460 27.210 858.720 27.530 ;
        RECT 1055.800 27.210 1056.060 27.530 ;
        RECT 858.520 19.030 858.660 27.210 ;
        RECT 757.720 18.710 757.980 19.030 ;
        RECT 858.460 18.710 858.720 19.030 ;
        RECT 757.780 2.400 757.920 18.710 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1731.510 25.740 1731.830 25.800 ;
        RECT 2060.410 25.740 2060.730 25.800 ;
        RECT 1731.510 25.600 2060.730 25.740 ;
        RECT 1731.510 25.540 1731.830 25.600 ;
        RECT 2060.410 25.540 2060.730 25.600 ;
      LAYER via ;
        RECT 1731.540 25.540 1731.800 25.800 ;
        RECT 2060.440 25.540 2060.700 25.800 ;
      LAYER met2 ;
        RECT 1730.390 600.170 1730.670 604.000 ;
        RECT 1730.390 600.030 1731.740 600.170 ;
        RECT 1730.390 600.000 1730.670 600.030 ;
        RECT 1731.600 25.830 1731.740 600.030 ;
        RECT 1731.540 25.510 1731.800 25.830 ;
        RECT 2060.440 25.510 2060.700 25.830 ;
        RECT 2060.500 2.400 2060.640 25.510 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1741.170 586.740 1741.490 586.800 ;
        RECT 1745.310 586.740 1745.630 586.800 ;
        RECT 1741.170 586.600 1745.630 586.740 ;
        RECT 1741.170 586.540 1741.490 586.600 ;
        RECT 1745.310 586.540 1745.630 586.600 ;
        RECT 1745.310 25.400 1745.630 25.460 ;
        RECT 2078.350 25.400 2078.670 25.460 ;
        RECT 1745.310 25.260 2078.670 25.400 ;
        RECT 1745.310 25.200 1745.630 25.260 ;
        RECT 2078.350 25.200 2078.670 25.260 ;
      LAYER via ;
        RECT 1741.200 586.540 1741.460 586.800 ;
        RECT 1745.340 586.540 1745.600 586.800 ;
        RECT 1745.340 25.200 1745.600 25.460 ;
        RECT 2078.380 25.200 2078.640 25.460 ;
      LAYER met2 ;
        RECT 1739.590 600.170 1739.870 604.000 ;
        RECT 1739.590 600.030 1741.400 600.170 ;
        RECT 1739.590 600.000 1739.870 600.030 ;
        RECT 1741.260 586.830 1741.400 600.030 ;
        RECT 1741.200 586.510 1741.460 586.830 ;
        RECT 1745.340 586.510 1745.600 586.830 ;
        RECT 1745.400 25.490 1745.540 586.510 ;
        RECT 1745.340 25.170 1745.600 25.490 ;
        RECT 2078.380 25.170 2078.640 25.490 ;
        RECT 2078.440 2.400 2078.580 25.170 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1750.370 586.740 1750.690 586.800 ;
        RECT 1752.210 586.740 1752.530 586.800 ;
        RECT 1750.370 586.600 1752.530 586.740 ;
        RECT 1750.370 586.540 1750.690 586.600 ;
        RECT 1752.210 586.540 1752.530 586.600 ;
        RECT 2095.830 25.400 2096.150 25.460 ;
        RECT 2079.360 25.260 2096.150 25.400 ;
        RECT 1752.210 25.060 1752.530 25.120 ;
        RECT 2079.360 25.060 2079.500 25.260 ;
        RECT 2095.830 25.200 2096.150 25.260 ;
        RECT 1752.210 24.920 2079.500 25.060 ;
        RECT 1752.210 24.860 1752.530 24.920 ;
      LAYER via ;
        RECT 1750.400 586.540 1750.660 586.800 ;
        RECT 1752.240 586.540 1752.500 586.800 ;
        RECT 1752.240 24.860 1752.500 25.120 ;
        RECT 2095.860 25.200 2096.120 25.460 ;
      LAYER met2 ;
        RECT 1748.790 600.170 1749.070 604.000 ;
        RECT 1748.790 600.030 1750.600 600.170 ;
        RECT 1748.790 600.000 1749.070 600.030 ;
        RECT 1750.460 586.830 1750.600 600.030 ;
        RECT 1750.400 586.510 1750.660 586.830 ;
        RECT 1752.240 586.510 1752.500 586.830 ;
        RECT 1752.300 25.150 1752.440 586.510 ;
        RECT 2095.860 25.170 2096.120 25.490 ;
        RECT 1752.240 24.830 1752.500 25.150 ;
        RECT 2095.920 2.400 2096.060 25.170 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2066.850 25.740 2067.170 25.800 ;
        RECT 2113.770 25.740 2114.090 25.800 ;
        RECT 2066.850 25.600 2114.090 25.740 ;
        RECT 2066.850 25.540 2067.170 25.600 ;
        RECT 2113.770 25.540 2114.090 25.600 ;
        RECT 1758.650 24.720 1758.970 24.780 ;
        RECT 2066.850 24.720 2067.170 24.780 ;
        RECT 1758.650 24.580 2067.170 24.720 ;
        RECT 1758.650 24.520 1758.970 24.580 ;
        RECT 2066.850 24.520 2067.170 24.580 ;
      LAYER via ;
        RECT 2066.880 25.540 2067.140 25.800 ;
        RECT 2113.800 25.540 2114.060 25.800 ;
        RECT 1758.680 24.520 1758.940 24.780 ;
        RECT 2066.880 24.520 2067.140 24.780 ;
      LAYER met2 ;
        RECT 1757.990 600.170 1758.270 604.000 ;
        RECT 1757.990 600.030 1758.880 600.170 ;
        RECT 1757.990 600.000 1758.270 600.030 ;
        RECT 1758.740 24.810 1758.880 600.030 ;
        RECT 2066.880 25.510 2067.140 25.830 ;
        RECT 2113.800 25.510 2114.060 25.830 ;
        RECT 2066.940 24.810 2067.080 25.510 ;
        RECT 1758.680 24.490 1758.940 24.810 ;
        RECT 2066.880 24.490 2067.140 24.810 ;
        RECT 2113.860 2.400 2114.000 25.510 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.770 588.780 1769.090 588.840 ;
        RECT 1772.910 588.780 1773.230 588.840 ;
        RECT 1768.770 588.640 1773.230 588.780 ;
        RECT 1768.770 588.580 1769.090 588.640 ;
        RECT 1772.910 588.580 1773.230 588.640 ;
        RECT 1772.910 24.380 1773.230 24.440 ;
        RECT 2131.710 24.380 2132.030 24.440 ;
        RECT 1772.910 24.240 2132.030 24.380 ;
        RECT 1772.910 24.180 1773.230 24.240 ;
        RECT 2131.710 24.180 2132.030 24.240 ;
      LAYER via ;
        RECT 1768.800 588.580 1769.060 588.840 ;
        RECT 1772.940 588.580 1773.200 588.840 ;
        RECT 1772.940 24.180 1773.200 24.440 ;
        RECT 2131.740 24.180 2132.000 24.440 ;
      LAYER met2 ;
        RECT 1767.190 600.170 1767.470 604.000 ;
        RECT 1767.190 600.030 1769.000 600.170 ;
        RECT 1767.190 600.000 1767.470 600.030 ;
        RECT 1768.860 588.870 1769.000 600.030 ;
        RECT 1768.800 588.550 1769.060 588.870 ;
        RECT 1772.940 588.550 1773.200 588.870 ;
        RECT 1773.000 24.470 1773.140 588.550 ;
        RECT 1772.940 24.150 1773.200 24.470 ;
        RECT 2131.740 24.150 2132.000 24.470 ;
        RECT 2131.800 2.400 2131.940 24.150 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1777.970 586.740 1778.290 586.800 ;
        RECT 1779.810 586.740 1780.130 586.800 ;
        RECT 1777.970 586.600 1780.130 586.740 ;
        RECT 1777.970 586.540 1778.290 586.600 ;
        RECT 1779.810 586.540 1780.130 586.600 ;
        RECT 1779.810 24.040 1780.130 24.100 ;
        RECT 2149.650 24.040 2149.970 24.100 ;
        RECT 1779.810 23.900 2149.970 24.040 ;
        RECT 1779.810 23.840 1780.130 23.900 ;
        RECT 2149.650 23.840 2149.970 23.900 ;
      LAYER via ;
        RECT 1778.000 586.540 1778.260 586.800 ;
        RECT 1779.840 586.540 1780.100 586.800 ;
        RECT 1779.840 23.840 1780.100 24.100 ;
        RECT 2149.680 23.840 2149.940 24.100 ;
      LAYER met2 ;
        RECT 1776.390 600.170 1776.670 604.000 ;
        RECT 1776.390 600.030 1778.200 600.170 ;
        RECT 1776.390 600.000 1776.670 600.030 ;
        RECT 1778.060 586.830 1778.200 600.030 ;
        RECT 1778.000 586.510 1778.260 586.830 ;
        RECT 1779.840 586.510 1780.100 586.830 ;
        RECT 1779.900 24.130 1780.040 586.510 ;
        RECT 1779.840 23.810 1780.100 24.130 ;
        RECT 2149.680 23.810 2149.940 24.130 ;
        RECT 2149.740 2.400 2149.880 23.810 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1785.330 585.040 1785.650 585.100 ;
        RECT 1786.710 585.040 1787.030 585.100 ;
        RECT 1785.330 584.900 1787.030 585.040 ;
        RECT 1785.330 584.840 1785.650 584.900 ;
        RECT 1786.710 584.840 1787.030 584.900 ;
      LAYER via ;
        RECT 1785.360 584.840 1785.620 585.100 ;
        RECT 1786.740 584.840 1787.000 585.100 ;
      LAYER met2 ;
        RECT 1785.590 600.000 1785.870 604.000 ;
        RECT 1785.650 598.810 1785.790 600.000 ;
        RECT 1785.420 598.670 1785.790 598.810 ;
        RECT 1785.420 585.130 1785.560 598.670 ;
        RECT 1785.360 584.810 1785.620 585.130 ;
        RECT 1786.740 584.810 1787.000 585.130 ;
        RECT 1786.800 24.325 1786.940 584.810 ;
        RECT 1786.730 23.955 1787.010 24.325 ;
        RECT 2167.610 23.955 2167.890 24.325 ;
        RECT 2167.680 2.400 2167.820 23.955 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
      LAYER via2 ;
        RECT 1786.730 24.000 1787.010 24.280 ;
        RECT 2167.610 24.000 2167.890 24.280 ;
      LAYER met3 ;
        RECT 1786.705 24.290 1787.035 24.305 ;
        RECT 2167.585 24.290 2167.915 24.305 ;
        RECT 1786.705 23.990 2167.915 24.290 ;
        RECT 1786.705 23.975 1787.035 23.990 ;
        RECT 2167.585 23.975 2167.915 23.990 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1796.370 586.740 1796.690 586.800 ;
        RECT 1800.510 586.740 1800.830 586.800 ;
        RECT 1796.370 586.600 1800.830 586.740 ;
        RECT 1796.370 586.540 1796.690 586.600 ;
        RECT 1800.510 586.540 1800.830 586.600 ;
        RECT 1800.510 35.940 1800.830 36.000 ;
        RECT 2185.070 35.940 2185.390 36.000 ;
        RECT 1800.510 35.800 2185.390 35.940 ;
        RECT 1800.510 35.740 1800.830 35.800 ;
        RECT 2185.070 35.740 2185.390 35.800 ;
      LAYER via ;
        RECT 1796.400 586.540 1796.660 586.800 ;
        RECT 1800.540 586.540 1800.800 586.800 ;
        RECT 1800.540 35.740 1800.800 36.000 ;
        RECT 2185.100 35.740 2185.360 36.000 ;
      LAYER met2 ;
        RECT 1794.790 600.170 1795.070 604.000 ;
        RECT 1794.790 600.030 1796.600 600.170 ;
        RECT 1794.790 600.000 1795.070 600.030 ;
        RECT 1796.460 586.830 1796.600 600.030 ;
        RECT 1796.400 586.510 1796.660 586.830 ;
        RECT 1800.540 586.510 1800.800 586.830 ;
        RECT 1800.600 36.030 1800.740 586.510 ;
        RECT 1800.540 35.710 1800.800 36.030 ;
        RECT 2185.100 35.710 2185.360 36.030 ;
        RECT 2185.160 2.400 2185.300 35.710 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1805.570 586.740 1805.890 586.800 ;
        RECT 1807.410 586.740 1807.730 586.800 ;
        RECT 1805.570 586.600 1807.730 586.740 ;
        RECT 1805.570 586.540 1805.890 586.600 ;
        RECT 1807.410 586.540 1807.730 586.600 ;
        RECT 1807.410 36.280 1807.730 36.340 ;
        RECT 2203.010 36.280 2203.330 36.340 ;
        RECT 1807.410 36.140 2203.330 36.280 ;
        RECT 1807.410 36.080 1807.730 36.140 ;
        RECT 2203.010 36.080 2203.330 36.140 ;
      LAYER via ;
        RECT 1805.600 586.540 1805.860 586.800 ;
        RECT 1807.440 586.540 1807.700 586.800 ;
        RECT 1807.440 36.080 1807.700 36.340 ;
        RECT 2203.040 36.080 2203.300 36.340 ;
      LAYER met2 ;
        RECT 1803.990 600.170 1804.270 604.000 ;
        RECT 1803.990 600.030 1805.800 600.170 ;
        RECT 1803.990 600.000 1804.270 600.030 ;
        RECT 1805.660 586.830 1805.800 600.030 ;
        RECT 1805.600 586.510 1805.860 586.830 ;
        RECT 1807.440 586.510 1807.700 586.830 ;
        RECT 1807.500 36.370 1807.640 586.510 ;
        RECT 1807.440 36.050 1807.700 36.370 ;
        RECT 2203.040 36.050 2203.300 36.370 ;
        RECT 2203.100 2.400 2203.240 36.050 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.310 36.620 1814.630 36.680 ;
        RECT 2220.950 36.620 2221.270 36.680 ;
        RECT 1814.310 36.480 2221.270 36.620 ;
        RECT 1814.310 36.420 1814.630 36.480 ;
        RECT 2220.950 36.420 2221.270 36.480 ;
      LAYER via ;
        RECT 1814.340 36.420 1814.600 36.680 ;
        RECT 2220.980 36.420 2221.240 36.680 ;
      LAYER met2 ;
        RECT 1813.190 600.170 1813.470 604.000 ;
        RECT 1813.190 600.030 1814.540 600.170 ;
        RECT 1813.190 600.000 1813.470 600.030 ;
        RECT 1814.400 36.710 1814.540 600.030 ;
        RECT 1814.340 36.390 1814.600 36.710 ;
        RECT 2220.980 36.390 2221.240 36.710 ;
        RECT 2221.040 2.400 2221.180 36.390 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 775.630 25.400 775.950 25.460 ;
        RECT 1069.570 25.400 1069.890 25.460 ;
        RECT 775.630 25.260 1069.890 25.400 ;
        RECT 775.630 25.200 775.950 25.260 ;
        RECT 1069.570 25.200 1069.890 25.260 ;
      LAYER via ;
        RECT 775.660 25.200 775.920 25.460 ;
        RECT 1069.600 25.200 1069.860 25.460 ;
      LAYER met2 ;
        RECT 1069.370 600.000 1069.650 604.000 ;
        RECT 1069.430 598.810 1069.570 600.000 ;
        RECT 1069.430 598.670 1069.800 598.810 ;
        RECT 1069.660 25.490 1069.800 598.670 ;
        RECT 775.660 25.170 775.920 25.490 ;
        RECT 1069.600 25.170 1069.860 25.490 ;
        RECT 775.720 2.400 775.860 25.170 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1823.970 586.740 1824.290 586.800 ;
        RECT 1828.110 586.740 1828.430 586.800 ;
        RECT 1823.970 586.600 1828.430 586.740 ;
        RECT 1823.970 586.540 1824.290 586.600 ;
        RECT 1828.110 586.540 1828.430 586.600 ;
        RECT 1828.110 36.960 1828.430 37.020 ;
        RECT 2238.890 36.960 2239.210 37.020 ;
        RECT 1828.110 36.820 2239.210 36.960 ;
        RECT 1828.110 36.760 1828.430 36.820 ;
        RECT 2238.890 36.760 2239.210 36.820 ;
      LAYER via ;
        RECT 1824.000 586.540 1824.260 586.800 ;
        RECT 1828.140 586.540 1828.400 586.800 ;
        RECT 1828.140 36.760 1828.400 37.020 ;
        RECT 2238.920 36.760 2239.180 37.020 ;
      LAYER met2 ;
        RECT 1822.390 600.170 1822.670 604.000 ;
        RECT 1822.390 600.030 1824.200 600.170 ;
        RECT 1822.390 600.000 1822.670 600.030 ;
        RECT 1824.060 586.830 1824.200 600.030 ;
        RECT 1824.000 586.510 1824.260 586.830 ;
        RECT 1828.140 586.510 1828.400 586.830 ;
        RECT 1828.200 37.050 1828.340 586.510 ;
        RECT 1828.140 36.730 1828.400 37.050 ;
        RECT 2238.920 36.730 2239.180 37.050 ;
        RECT 2238.980 2.400 2239.120 36.730 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1833.170 586.740 1833.490 586.800 ;
        RECT 1835.010 586.740 1835.330 586.800 ;
        RECT 1833.170 586.600 1835.330 586.740 ;
        RECT 1833.170 586.540 1833.490 586.600 ;
        RECT 1835.010 586.540 1835.330 586.600 ;
        RECT 1835.010 37.300 1835.330 37.360 ;
        RECT 2256.370 37.300 2256.690 37.360 ;
        RECT 1835.010 37.160 2256.690 37.300 ;
        RECT 1835.010 37.100 1835.330 37.160 ;
        RECT 2256.370 37.100 2256.690 37.160 ;
      LAYER via ;
        RECT 1833.200 586.540 1833.460 586.800 ;
        RECT 1835.040 586.540 1835.300 586.800 ;
        RECT 1835.040 37.100 1835.300 37.360 ;
        RECT 2256.400 37.100 2256.660 37.360 ;
      LAYER met2 ;
        RECT 1831.590 600.170 1831.870 604.000 ;
        RECT 1831.590 600.030 1833.400 600.170 ;
        RECT 1831.590 600.000 1831.870 600.030 ;
        RECT 1833.260 586.830 1833.400 600.030 ;
        RECT 1833.200 586.510 1833.460 586.830 ;
        RECT 1835.040 586.510 1835.300 586.830 ;
        RECT 1835.100 37.390 1835.240 586.510 ;
        RECT 1835.040 37.070 1835.300 37.390 ;
        RECT 2256.400 37.070 2256.660 37.390 ;
        RECT 2256.460 2.400 2256.600 37.070 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1841.910 48.180 1842.230 48.240 ;
        RECT 2274.310 48.180 2274.630 48.240 ;
        RECT 1841.910 48.040 2274.630 48.180 ;
        RECT 1841.910 47.980 1842.230 48.040 ;
        RECT 2274.310 47.980 2274.630 48.040 ;
      LAYER via ;
        RECT 1841.940 47.980 1842.200 48.240 ;
        RECT 2274.340 47.980 2274.600 48.240 ;
      LAYER met2 ;
        RECT 1840.790 600.170 1841.070 604.000 ;
        RECT 1840.790 600.030 1842.140 600.170 ;
        RECT 1840.790 600.000 1841.070 600.030 ;
        RECT 1842.000 48.270 1842.140 600.030 ;
        RECT 1841.940 47.950 1842.200 48.270 ;
        RECT 2274.340 47.950 2274.600 48.270 ;
        RECT 2274.400 2.400 2274.540 47.950 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1851.570 586.740 1851.890 586.800 ;
        RECT 1855.710 586.740 1856.030 586.800 ;
        RECT 1851.570 586.600 1856.030 586.740 ;
        RECT 1851.570 586.540 1851.890 586.600 ;
        RECT 1855.710 586.540 1856.030 586.600 ;
        RECT 1855.710 47.840 1856.030 47.900 ;
        RECT 2292.250 47.840 2292.570 47.900 ;
        RECT 1855.710 47.700 2292.570 47.840 ;
        RECT 1855.710 47.640 1856.030 47.700 ;
        RECT 2292.250 47.640 2292.570 47.700 ;
      LAYER via ;
        RECT 1851.600 586.540 1851.860 586.800 ;
        RECT 1855.740 586.540 1856.000 586.800 ;
        RECT 1855.740 47.640 1856.000 47.900 ;
        RECT 2292.280 47.640 2292.540 47.900 ;
      LAYER met2 ;
        RECT 1849.990 600.170 1850.270 604.000 ;
        RECT 1849.990 600.030 1851.800 600.170 ;
        RECT 1849.990 600.000 1850.270 600.030 ;
        RECT 1851.660 586.830 1851.800 600.030 ;
        RECT 1851.600 586.510 1851.860 586.830 ;
        RECT 1855.740 586.510 1856.000 586.830 ;
        RECT 1855.800 47.930 1855.940 586.510 ;
        RECT 1855.740 47.610 1856.000 47.930 ;
        RECT 2292.280 47.610 2292.540 47.930 ;
        RECT 2292.340 2.400 2292.480 47.610 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1860.770 586.740 1861.090 586.800 ;
        RECT 1862.150 586.740 1862.470 586.800 ;
        RECT 1860.770 586.600 1862.470 586.740 ;
        RECT 1860.770 586.540 1861.090 586.600 ;
        RECT 1862.150 586.540 1862.470 586.600 ;
        RECT 1862.150 47.500 1862.470 47.560 ;
        RECT 2310.190 47.500 2310.510 47.560 ;
        RECT 1862.150 47.360 2310.510 47.500 ;
        RECT 1862.150 47.300 1862.470 47.360 ;
        RECT 2310.190 47.300 2310.510 47.360 ;
      LAYER via ;
        RECT 1860.800 586.540 1861.060 586.800 ;
        RECT 1862.180 586.540 1862.440 586.800 ;
        RECT 1862.180 47.300 1862.440 47.560 ;
        RECT 2310.220 47.300 2310.480 47.560 ;
      LAYER met2 ;
        RECT 1859.190 600.170 1859.470 604.000 ;
        RECT 1859.190 600.030 1861.000 600.170 ;
        RECT 1859.190 600.000 1859.470 600.030 ;
        RECT 1860.860 586.830 1861.000 600.030 ;
        RECT 1860.800 586.510 1861.060 586.830 ;
        RECT 1862.180 586.510 1862.440 586.830 ;
        RECT 1862.240 47.590 1862.380 586.510 ;
        RECT 1862.180 47.270 1862.440 47.590 ;
        RECT 2310.220 47.270 2310.480 47.590 ;
        RECT 2310.280 2.400 2310.420 47.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1869.510 28.120 1869.830 28.180 ;
        RECT 2328.130 28.120 2328.450 28.180 ;
        RECT 1869.510 27.980 2328.450 28.120 ;
        RECT 1869.510 27.920 1869.830 27.980 ;
        RECT 2328.130 27.920 2328.450 27.980 ;
      LAYER via ;
        RECT 1869.540 27.920 1869.800 28.180 ;
        RECT 2328.160 27.920 2328.420 28.180 ;
      LAYER met2 ;
        RECT 1868.390 600.170 1868.670 604.000 ;
        RECT 1868.390 600.030 1869.740 600.170 ;
        RECT 1868.390 600.000 1868.670 600.030 ;
        RECT 1869.600 28.210 1869.740 600.030 ;
        RECT 1869.540 27.890 1869.800 28.210 ;
        RECT 2328.160 27.890 2328.420 28.210 ;
        RECT 2328.220 2.400 2328.360 27.890 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1879.170 586.740 1879.490 586.800 ;
        RECT 1883.310 586.740 1883.630 586.800 ;
        RECT 1879.170 586.600 1883.630 586.740 ;
        RECT 1879.170 586.540 1879.490 586.600 ;
        RECT 1883.310 586.540 1883.630 586.600 ;
        RECT 1883.310 27.780 1883.630 27.840 ;
        RECT 2345.610 27.780 2345.930 27.840 ;
        RECT 1883.310 27.640 2345.930 27.780 ;
        RECT 1883.310 27.580 1883.630 27.640 ;
        RECT 2345.610 27.580 2345.930 27.640 ;
      LAYER via ;
        RECT 1879.200 586.540 1879.460 586.800 ;
        RECT 1883.340 586.540 1883.600 586.800 ;
        RECT 1883.340 27.580 1883.600 27.840 ;
        RECT 2345.640 27.580 2345.900 27.840 ;
      LAYER met2 ;
        RECT 1877.590 600.170 1877.870 604.000 ;
        RECT 1877.590 600.030 1879.400 600.170 ;
        RECT 1877.590 600.000 1877.870 600.030 ;
        RECT 1879.260 586.830 1879.400 600.030 ;
        RECT 1879.200 586.510 1879.460 586.830 ;
        RECT 1883.340 586.510 1883.600 586.830 ;
        RECT 1883.400 27.870 1883.540 586.510 ;
        RECT 1883.340 27.550 1883.600 27.870 ;
        RECT 2345.640 27.550 2345.900 27.870 ;
        RECT 2345.700 2.400 2345.840 27.550 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1888.370 586.740 1888.690 586.800 ;
        RECT 1890.210 586.740 1890.530 586.800 ;
        RECT 1888.370 586.600 1890.530 586.740 ;
        RECT 1888.370 586.540 1888.690 586.600 ;
        RECT 1890.210 586.540 1890.530 586.600 ;
        RECT 1890.210 28.460 1890.530 28.520 ;
        RECT 2363.550 28.460 2363.870 28.520 ;
        RECT 1890.210 28.320 2363.870 28.460 ;
        RECT 1890.210 28.260 1890.530 28.320 ;
        RECT 2363.550 28.260 2363.870 28.320 ;
      LAYER via ;
        RECT 1888.400 586.540 1888.660 586.800 ;
        RECT 1890.240 586.540 1890.500 586.800 ;
        RECT 1890.240 28.260 1890.500 28.520 ;
        RECT 2363.580 28.260 2363.840 28.520 ;
      LAYER met2 ;
        RECT 1886.790 600.170 1887.070 604.000 ;
        RECT 1886.790 600.030 1888.600 600.170 ;
        RECT 1886.790 600.000 1887.070 600.030 ;
        RECT 1888.460 586.830 1888.600 600.030 ;
        RECT 1888.400 586.510 1888.660 586.830 ;
        RECT 1890.240 586.510 1890.500 586.830 ;
        RECT 1890.300 28.550 1890.440 586.510 ;
        RECT 1890.240 28.230 1890.500 28.550 ;
        RECT 2363.580 28.230 2363.840 28.550 ;
        RECT 2363.640 2.400 2363.780 28.230 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1896.650 29.140 1896.970 29.200 ;
        RECT 2381.490 29.140 2381.810 29.200 ;
        RECT 1896.650 29.000 2381.810 29.140 ;
        RECT 1896.650 28.940 1896.970 29.000 ;
        RECT 2381.490 28.940 2381.810 29.000 ;
      LAYER via ;
        RECT 1896.680 28.940 1896.940 29.200 ;
        RECT 2381.520 28.940 2381.780 29.200 ;
      LAYER met2 ;
        RECT 1895.990 600.170 1896.270 604.000 ;
        RECT 1895.990 600.030 1896.880 600.170 ;
        RECT 1895.990 600.000 1896.270 600.030 ;
        RECT 1896.740 29.230 1896.880 600.030 ;
        RECT 1896.680 28.910 1896.940 29.230 ;
        RECT 2381.520 28.910 2381.780 29.230 ;
        RECT 2381.580 2.400 2381.720 28.910 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1906.770 586.740 1907.090 586.800 ;
        RECT 1910.910 586.740 1911.230 586.800 ;
        RECT 1906.770 586.600 1911.230 586.740 ;
        RECT 1906.770 586.540 1907.090 586.600 ;
        RECT 1910.910 586.540 1911.230 586.600 ;
        RECT 1910.910 28.800 1911.230 28.860 ;
        RECT 2399.430 28.800 2399.750 28.860 ;
        RECT 1910.910 28.660 2399.750 28.800 ;
        RECT 1910.910 28.600 1911.230 28.660 ;
        RECT 2399.430 28.600 2399.750 28.660 ;
      LAYER via ;
        RECT 1906.800 586.540 1907.060 586.800 ;
        RECT 1910.940 586.540 1911.200 586.800 ;
        RECT 1910.940 28.600 1911.200 28.860 ;
        RECT 2399.460 28.600 2399.720 28.860 ;
      LAYER met2 ;
        RECT 1905.190 600.170 1905.470 604.000 ;
        RECT 1905.190 600.030 1907.000 600.170 ;
        RECT 1905.190 600.000 1905.470 600.030 ;
        RECT 1906.860 586.830 1907.000 600.030 ;
        RECT 1906.800 586.510 1907.060 586.830 ;
        RECT 1910.940 586.510 1911.200 586.830 ;
        RECT 1911.000 28.890 1911.140 586.510 ;
        RECT 1910.940 28.570 1911.200 28.890 ;
        RECT 2399.460 28.570 2399.720 28.890 ;
        RECT 2399.520 2.400 2399.660 28.570 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.570 25.740 793.890 25.800 ;
        RECT 1076.470 25.740 1076.790 25.800 ;
        RECT 793.570 25.600 1076.790 25.740 ;
        RECT 793.570 25.540 793.890 25.600 ;
        RECT 1076.470 25.540 1076.790 25.600 ;
      LAYER via ;
        RECT 793.600 25.540 793.860 25.800 ;
        RECT 1076.500 25.540 1076.760 25.800 ;
      LAYER met2 ;
        RECT 1078.570 600.170 1078.850 604.000 ;
        RECT 1076.560 600.030 1078.850 600.170 ;
        RECT 1076.560 25.830 1076.700 600.030 ;
        RECT 1078.570 600.000 1078.850 600.030 ;
        RECT 793.600 25.510 793.860 25.830 ;
        RECT 1076.500 25.510 1076.760 25.830 ;
        RECT 793.660 2.400 793.800 25.510 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 993.670 583.000 993.990 583.060 ;
        RECT 997.350 583.000 997.670 583.060 ;
        RECT 993.670 582.860 997.670 583.000 ;
        RECT 993.670 582.800 993.990 582.860 ;
        RECT 997.350 582.800 997.670 582.860 ;
        RECT 639.010 36.280 639.330 36.340 ;
        RECT 993.670 36.280 993.990 36.340 ;
        RECT 639.010 36.140 993.990 36.280 ;
        RECT 639.010 36.080 639.330 36.140 ;
        RECT 993.670 36.080 993.990 36.140 ;
      LAYER via ;
        RECT 993.700 582.800 993.960 583.060 ;
        RECT 997.380 582.800 997.640 583.060 ;
        RECT 639.040 36.080 639.300 36.340 ;
        RECT 993.700 36.080 993.960 36.340 ;
      LAYER met2 ;
        RECT 998.990 600.170 999.270 604.000 ;
        RECT 997.440 600.030 999.270 600.170 ;
        RECT 997.440 583.090 997.580 600.030 ;
        RECT 998.990 600.000 999.270 600.030 ;
        RECT 993.700 582.770 993.960 583.090 ;
        RECT 997.380 582.770 997.640 583.090 ;
        RECT 993.760 36.370 993.900 582.770 ;
        RECT 639.040 36.050 639.300 36.370 ;
        RECT 993.700 36.050 993.960 36.370 ;
        RECT 639.100 2.400 639.240 36.050 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1917.350 29.820 1917.670 29.880 ;
        RECT 2422.890 29.820 2423.210 29.880 ;
        RECT 1917.350 29.680 2423.210 29.820 ;
        RECT 1917.350 29.620 1917.670 29.680 ;
        RECT 2422.890 29.620 2423.210 29.680 ;
      LAYER via ;
        RECT 1917.380 29.620 1917.640 29.880 ;
        RECT 2422.920 29.620 2423.180 29.880 ;
      LAYER met2 ;
        RECT 1917.150 600.000 1917.430 604.000 ;
        RECT 1917.210 598.810 1917.350 600.000 ;
        RECT 1917.210 598.670 1917.580 598.810 ;
        RECT 1917.440 29.910 1917.580 598.670 ;
        RECT 1917.380 29.590 1917.640 29.910 ;
        RECT 2422.920 29.590 2423.180 29.910 ;
        RECT 2422.980 2.400 2423.120 29.590 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1927.930 586.740 1928.250 586.800 ;
        RECT 1931.610 586.740 1931.930 586.800 ;
        RECT 1927.930 586.600 1931.930 586.740 ;
        RECT 1927.930 586.540 1928.250 586.600 ;
        RECT 1931.610 586.540 1931.930 586.600 ;
        RECT 1931.610 29.480 1931.930 29.540 ;
        RECT 2440.830 29.480 2441.150 29.540 ;
        RECT 1931.610 29.340 2441.150 29.480 ;
        RECT 1931.610 29.280 1931.930 29.340 ;
        RECT 2440.830 29.280 2441.150 29.340 ;
      LAYER via ;
        RECT 1927.960 586.540 1928.220 586.800 ;
        RECT 1931.640 586.540 1931.900 586.800 ;
        RECT 1931.640 29.280 1931.900 29.540 ;
        RECT 2440.860 29.280 2441.120 29.540 ;
      LAYER met2 ;
        RECT 1926.350 600.170 1926.630 604.000 ;
        RECT 1926.350 600.030 1928.160 600.170 ;
        RECT 1926.350 600.000 1926.630 600.030 ;
        RECT 1928.020 586.830 1928.160 600.030 ;
        RECT 1927.960 586.510 1928.220 586.830 ;
        RECT 1931.640 586.510 1931.900 586.830 ;
        RECT 1931.700 29.570 1931.840 586.510 ;
        RECT 1931.640 29.250 1931.900 29.570 ;
        RECT 2440.860 29.250 2441.120 29.570 ;
        RECT 2440.920 2.400 2441.060 29.250 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1937.590 545.260 1937.910 545.320 ;
        RECT 1938.510 545.260 1938.830 545.320 ;
        RECT 1937.590 545.120 1938.830 545.260 ;
        RECT 1937.590 545.060 1937.910 545.120 ;
        RECT 1938.510 545.060 1938.830 545.120 ;
        RECT 1938.510 30.160 1938.830 30.220 ;
        RECT 2458.770 30.160 2459.090 30.220 ;
        RECT 1938.510 30.020 2459.090 30.160 ;
        RECT 1938.510 29.960 1938.830 30.020 ;
        RECT 2458.770 29.960 2459.090 30.020 ;
      LAYER via ;
        RECT 1937.620 545.060 1937.880 545.320 ;
        RECT 1938.540 545.060 1938.800 545.320 ;
        RECT 1938.540 29.960 1938.800 30.220 ;
        RECT 2458.800 29.960 2459.060 30.220 ;
      LAYER met2 ;
        RECT 1935.550 600.170 1935.830 604.000 ;
        RECT 1935.550 600.030 1938.280 600.170 ;
        RECT 1935.550 600.000 1935.830 600.030 ;
        RECT 1938.140 593.370 1938.280 600.030 ;
        RECT 1937.680 593.230 1938.280 593.370 ;
        RECT 1937.680 545.350 1937.820 593.230 ;
        RECT 1937.620 545.030 1937.880 545.350 ;
        RECT 1938.540 545.030 1938.800 545.350 ;
        RECT 1938.600 30.250 1938.740 545.030 ;
        RECT 1938.540 29.930 1938.800 30.250 ;
        RECT 2458.800 29.930 2459.060 30.250 ;
        RECT 2458.860 2.400 2459.000 29.930 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1944.950 30.500 1945.270 30.560 ;
        RECT 2476.710 30.500 2477.030 30.560 ;
        RECT 1944.950 30.360 2477.030 30.500 ;
        RECT 1944.950 30.300 1945.270 30.360 ;
        RECT 2476.710 30.300 2477.030 30.360 ;
      LAYER via ;
        RECT 1944.980 30.300 1945.240 30.560 ;
        RECT 2476.740 30.300 2477.000 30.560 ;
      LAYER met2 ;
        RECT 1944.750 600.000 1945.030 604.000 ;
        RECT 1944.810 598.810 1944.950 600.000 ;
        RECT 1944.810 598.670 1945.180 598.810 ;
        RECT 1945.040 30.590 1945.180 598.670 ;
        RECT 1944.980 30.270 1945.240 30.590 ;
        RECT 2476.740 30.270 2477.000 30.590 ;
        RECT 2476.800 2.400 2476.940 30.270 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1955.530 588.100 1955.850 588.160 ;
        RECT 1958.750 588.100 1959.070 588.160 ;
        RECT 1955.530 587.960 1959.070 588.100 ;
        RECT 1955.530 587.900 1955.850 587.960 ;
        RECT 1958.750 587.900 1959.070 587.960 ;
        RECT 1958.750 34.240 1959.070 34.300 ;
        RECT 2494.650 34.240 2494.970 34.300 ;
        RECT 1958.750 34.100 2494.970 34.240 ;
        RECT 1958.750 34.040 1959.070 34.100 ;
        RECT 2494.650 34.040 2494.970 34.100 ;
      LAYER via ;
        RECT 1955.560 587.900 1955.820 588.160 ;
        RECT 1958.780 587.900 1959.040 588.160 ;
        RECT 1958.780 34.040 1959.040 34.300 ;
        RECT 2494.680 34.040 2494.940 34.300 ;
      LAYER met2 ;
        RECT 1953.950 600.170 1954.230 604.000 ;
        RECT 1953.950 600.030 1955.760 600.170 ;
        RECT 1953.950 600.000 1954.230 600.030 ;
        RECT 1955.620 588.190 1955.760 600.030 ;
        RECT 1955.560 587.870 1955.820 588.190 ;
        RECT 1958.780 587.870 1959.040 588.190 ;
        RECT 1958.840 34.330 1958.980 587.870 ;
        RECT 1958.780 34.010 1959.040 34.330 ;
        RECT 2494.680 34.010 2494.940 34.330 ;
        RECT 2494.740 2.400 2494.880 34.010 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1965.190 545.260 1965.510 545.320 ;
        RECT 1966.110 545.260 1966.430 545.320 ;
        RECT 1965.190 545.120 1966.430 545.260 ;
        RECT 1965.190 545.060 1965.510 545.120 ;
        RECT 1966.110 545.060 1966.430 545.120 ;
        RECT 1966.110 33.900 1966.430 33.960 ;
        RECT 2512.130 33.900 2512.450 33.960 ;
        RECT 1966.110 33.760 2512.450 33.900 ;
        RECT 1966.110 33.700 1966.430 33.760 ;
        RECT 2512.130 33.700 2512.450 33.760 ;
      LAYER via ;
        RECT 1965.220 545.060 1965.480 545.320 ;
        RECT 1966.140 545.060 1966.400 545.320 ;
        RECT 1966.140 33.700 1966.400 33.960 ;
        RECT 2512.160 33.700 2512.420 33.960 ;
      LAYER met2 ;
        RECT 1963.150 600.170 1963.430 604.000 ;
        RECT 1963.150 600.030 1965.880 600.170 ;
        RECT 1963.150 600.000 1963.430 600.030 ;
        RECT 1965.740 593.370 1965.880 600.030 ;
        RECT 1965.280 593.230 1965.880 593.370 ;
        RECT 1965.280 545.350 1965.420 593.230 ;
        RECT 1965.220 545.030 1965.480 545.350 ;
        RECT 1966.140 545.030 1966.400 545.350 ;
        RECT 1966.200 33.990 1966.340 545.030 ;
        RECT 1966.140 33.670 1966.400 33.990 ;
        RECT 2512.160 33.670 2512.420 33.990 ;
        RECT 2512.220 2.400 2512.360 33.670 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 33.560 1973.330 33.620 ;
        RECT 2530.070 33.560 2530.390 33.620 ;
        RECT 1973.010 33.420 2530.390 33.560 ;
        RECT 1973.010 33.360 1973.330 33.420 ;
        RECT 2530.070 33.360 2530.390 33.420 ;
      LAYER via ;
        RECT 1973.040 33.360 1973.300 33.620 ;
        RECT 2530.100 33.360 2530.360 33.620 ;
      LAYER met2 ;
        RECT 1972.350 600.170 1972.630 604.000 ;
        RECT 1972.350 600.030 1973.240 600.170 ;
        RECT 1972.350 600.000 1972.630 600.030 ;
        RECT 1973.100 33.650 1973.240 600.030 ;
        RECT 1973.040 33.330 1973.300 33.650 ;
        RECT 2530.100 33.330 2530.360 33.650 ;
        RECT 2530.160 2.400 2530.300 33.330 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1983.130 586.740 1983.450 586.800 ;
        RECT 1986.810 586.740 1987.130 586.800 ;
        RECT 1983.130 586.600 1987.130 586.740 ;
        RECT 1983.130 586.540 1983.450 586.600 ;
        RECT 1986.810 586.540 1987.130 586.600 ;
        RECT 1986.810 33.220 1987.130 33.280 ;
        RECT 2548.010 33.220 2548.330 33.280 ;
        RECT 1986.810 33.080 2548.330 33.220 ;
        RECT 1986.810 33.020 1987.130 33.080 ;
        RECT 2548.010 33.020 2548.330 33.080 ;
      LAYER via ;
        RECT 1983.160 586.540 1983.420 586.800 ;
        RECT 1986.840 586.540 1987.100 586.800 ;
        RECT 1986.840 33.020 1987.100 33.280 ;
        RECT 2548.040 33.020 2548.300 33.280 ;
      LAYER met2 ;
        RECT 1981.550 600.170 1981.830 604.000 ;
        RECT 1981.550 600.030 1983.360 600.170 ;
        RECT 1981.550 600.000 1981.830 600.030 ;
        RECT 1983.220 586.830 1983.360 600.030 ;
        RECT 1983.160 586.510 1983.420 586.830 ;
        RECT 1986.840 586.510 1987.100 586.830 ;
        RECT 1986.900 33.310 1987.040 586.510 ;
        RECT 1986.840 32.990 1987.100 33.310 ;
        RECT 2548.040 32.990 2548.300 33.310 ;
        RECT 2548.100 2.400 2548.240 32.990 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1993.250 32.880 1993.570 32.940 ;
        RECT 2565.950 32.880 2566.270 32.940 ;
        RECT 1993.250 32.740 2566.270 32.880 ;
        RECT 1993.250 32.680 1993.570 32.740 ;
        RECT 2565.950 32.680 2566.270 32.740 ;
      LAYER via ;
        RECT 1993.280 32.680 1993.540 32.940 ;
        RECT 2565.980 32.680 2566.240 32.940 ;
      LAYER met2 ;
        RECT 1990.750 600.170 1991.030 604.000 ;
        RECT 1990.750 600.030 1993.480 600.170 ;
        RECT 1990.750 600.000 1991.030 600.030 ;
        RECT 1993.340 32.970 1993.480 600.030 ;
        RECT 1993.280 32.650 1993.540 32.970 ;
        RECT 2565.980 32.650 2566.240 32.970 ;
        RECT 2566.040 2.400 2566.180 32.650 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1999.690 32.540 2000.010 32.600 ;
        RECT 2583.890 32.540 2584.210 32.600 ;
        RECT 1999.690 32.400 2584.210 32.540 ;
        RECT 1999.690 32.340 2000.010 32.400 ;
        RECT 2583.890 32.340 2584.210 32.400 ;
      LAYER via ;
        RECT 1999.720 32.340 1999.980 32.600 ;
        RECT 2583.920 32.340 2584.180 32.600 ;
      LAYER met2 ;
        RECT 1999.950 600.000 2000.230 604.000 ;
        RECT 2000.010 598.810 2000.150 600.000 ;
        RECT 1999.780 598.670 2000.150 598.810 ;
        RECT 1999.780 32.630 1999.920 598.670 ;
        RECT 1999.720 32.310 1999.980 32.630 ;
        RECT 2583.920 32.310 2584.180 32.630 ;
        RECT 2583.980 2.400 2584.120 32.310 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.490 26.080 817.810 26.140 ;
        RECT 1090.730 26.080 1091.050 26.140 ;
        RECT 817.490 25.940 1091.050 26.080 ;
        RECT 817.490 25.880 817.810 25.940 ;
        RECT 1090.730 25.880 1091.050 25.940 ;
      LAYER via ;
        RECT 817.520 25.880 817.780 26.140 ;
        RECT 1090.760 25.880 1091.020 26.140 ;
      LAYER met2 ;
        RECT 1090.530 600.000 1090.810 604.000 ;
        RECT 1090.590 598.810 1090.730 600.000 ;
        RECT 1090.590 598.670 1090.960 598.810 ;
        RECT 1090.820 26.170 1090.960 598.670 ;
        RECT 817.520 25.850 817.780 26.170 ;
        RECT 1090.760 25.850 1091.020 26.170 ;
        RECT 817.580 2.400 817.720 25.850 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2010.730 586.740 2011.050 586.800 ;
        RECT 2013.950 586.740 2014.270 586.800 ;
        RECT 2010.730 586.600 2014.270 586.740 ;
        RECT 2010.730 586.540 2011.050 586.600 ;
        RECT 2013.950 586.540 2014.270 586.600 ;
        RECT 2013.950 32.200 2014.270 32.260 ;
        RECT 2601.370 32.200 2601.690 32.260 ;
        RECT 2013.950 32.060 2601.690 32.200 ;
        RECT 2013.950 32.000 2014.270 32.060 ;
        RECT 2601.370 32.000 2601.690 32.060 ;
      LAYER via ;
        RECT 2010.760 586.540 2011.020 586.800 ;
        RECT 2013.980 586.540 2014.240 586.800 ;
        RECT 2013.980 32.000 2014.240 32.260 ;
        RECT 2601.400 32.000 2601.660 32.260 ;
      LAYER met2 ;
        RECT 2009.150 600.170 2009.430 604.000 ;
        RECT 2009.150 600.030 2010.960 600.170 ;
        RECT 2009.150 600.000 2009.430 600.030 ;
        RECT 2010.820 586.830 2010.960 600.030 ;
        RECT 2010.760 586.510 2011.020 586.830 ;
        RECT 2013.980 586.510 2014.240 586.830 ;
        RECT 2014.040 32.290 2014.180 586.510 ;
        RECT 2013.980 31.970 2014.240 32.290 ;
        RECT 2601.400 31.970 2601.660 32.290 ;
        RECT 2601.460 2.400 2601.600 31.970 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2019.010 579.600 2019.330 579.660 ;
        RECT 2020.390 579.600 2020.710 579.660 ;
        RECT 2019.010 579.460 2020.710 579.600 ;
        RECT 2019.010 579.400 2019.330 579.460 ;
        RECT 2020.390 579.400 2020.710 579.460 ;
        RECT 2019.010 531.660 2019.330 531.720 ;
        RECT 2019.470 531.660 2019.790 531.720 ;
        RECT 2019.010 531.520 2019.790 531.660 ;
        RECT 2019.010 531.460 2019.330 531.520 ;
        RECT 2019.470 531.460 2019.790 531.520 ;
        RECT 2019.470 496.780 2019.790 497.040 ;
        RECT 2019.560 496.640 2019.700 496.780 ;
        RECT 2019.930 496.640 2020.250 496.700 ;
        RECT 2019.560 496.500 2020.250 496.640 ;
        RECT 2019.930 496.440 2020.250 496.500 ;
        RECT 2018.550 483.040 2018.870 483.100 ;
        RECT 2019.930 483.040 2020.250 483.100 ;
        RECT 2018.550 482.900 2020.250 483.040 ;
        RECT 2018.550 482.840 2018.870 482.900 ;
        RECT 2019.930 482.840 2020.250 482.900 ;
        RECT 2018.550 435.100 2018.870 435.160 ;
        RECT 2019.470 435.100 2019.790 435.160 ;
        RECT 2018.550 434.960 2019.790 435.100 ;
        RECT 2018.550 434.900 2018.870 434.960 ;
        RECT 2019.470 434.900 2019.790 434.960 ;
        RECT 2019.010 379.340 2019.330 379.400 ;
        RECT 2019.930 379.340 2020.250 379.400 ;
        RECT 2019.010 379.200 2020.250 379.340 ;
        RECT 2019.010 379.140 2019.330 379.200 ;
        RECT 2019.930 379.140 2020.250 379.200 ;
        RECT 2019.010 331.400 2019.330 331.460 ;
        RECT 2020.390 331.400 2020.710 331.460 ;
        RECT 2019.010 331.260 2020.710 331.400 ;
        RECT 2019.010 331.200 2019.330 331.260 ;
        RECT 2020.390 331.200 2020.710 331.260 ;
        RECT 2020.390 304.200 2020.710 304.260 ;
        RECT 2020.020 304.060 2020.710 304.200 ;
        RECT 2020.020 303.580 2020.160 304.060 ;
        RECT 2020.390 304.000 2020.710 304.060 ;
        RECT 2019.930 303.320 2020.250 303.580 ;
        RECT 2019.010 282.780 2019.330 282.840 ;
        RECT 2019.930 282.780 2020.250 282.840 ;
        RECT 2019.010 282.640 2020.250 282.780 ;
        RECT 2019.010 282.580 2019.330 282.640 ;
        RECT 2019.930 282.580 2020.250 282.640 ;
        RECT 2019.010 234.840 2019.330 234.900 ;
        RECT 2020.390 234.840 2020.710 234.900 ;
        RECT 2019.010 234.700 2020.710 234.840 ;
        RECT 2019.010 234.640 2019.330 234.700 ;
        RECT 2020.390 234.640 2020.710 234.700 ;
        RECT 2019.010 186.560 2019.330 186.620 ;
        RECT 2019.930 186.560 2020.250 186.620 ;
        RECT 2019.010 186.420 2020.250 186.560 ;
        RECT 2019.010 186.360 2019.330 186.420 ;
        RECT 2019.930 186.360 2020.250 186.420 ;
        RECT 2019.010 145.080 2019.330 145.140 ;
        RECT 2020.390 145.080 2020.710 145.140 ;
        RECT 2019.010 144.940 2020.710 145.080 ;
        RECT 2019.010 144.880 2019.330 144.940 ;
        RECT 2020.390 144.880 2020.710 144.940 ;
        RECT 2020.390 110.740 2020.710 110.800 ;
        RECT 2020.020 110.600 2020.710 110.740 ;
        RECT 2020.020 110.460 2020.160 110.600 ;
        RECT 2020.390 110.540 2020.710 110.600 ;
        RECT 2019.930 110.200 2020.250 110.460 ;
        RECT 2020.850 31.860 2021.170 31.920 ;
        RECT 2619.310 31.860 2619.630 31.920 ;
        RECT 2020.850 31.720 2619.630 31.860 ;
        RECT 2020.850 31.660 2021.170 31.720 ;
        RECT 2619.310 31.660 2619.630 31.720 ;
      LAYER via ;
        RECT 2019.040 579.400 2019.300 579.660 ;
        RECT 2020.420 579.400 2020.680 579.660 ;
        RECT 2019.040 531.460 2019.300 531.720 ;
        RECT 2019.500 531.460 2019.760 531.720 ;
        RECT 2019.500 496.780 2019.760 497.040 ;
        RECT 2019.960 496.440 2020.220 496.700 ;
        RECT 2018.580 482.840 2018.840 483.100 ;
        RECT 2019.960 482.840 2020.220 483.100 ;
        RECT 2018.580 434.900 2018.840 435.160 ;
        RECT 2019.500 434.900 2019.760 435.160 ;
        RECT 2019.040 379.140 2019.300 379.400 ;
        RECT 2019.960 379.140 2020.220 379.400 ;
        RECT 2019.040 331.200 2019.300 331.460 ;
        RECT 2020.420 331.200 2020.680 331.460 ;
        RECT 2020.420 304.000 2020.680 304.260 ;
        RECT 2019.960 303.320 2020.220 303.580 ;
        RECT 2019.040 282.580 2019.300 282.840 ;
        RECT 2019.960 282.580 2020.220 282.840 ;
        RECT 2019.040 234.640 2019.300 234.900 ;
        RECT 2020.420 234.640 2020.680 234.900 ;
        RECT 2019.040 186.360 2019.300 186.620 ;
        RECT 2019.960 186.360 2020.220 186.620 ;
        RECT 2019.040 144.880 2019.300 145.140 ;
        RECT 2020.420 144.880 2020.680 145.140 ;
        RECT 2020.420 110.540 2020.680 110.800 ;
        RECT 2019.960 110.200 2020.220 110.460 ;
        RECT 2020.880 31.660 2021.140 31.920 ;
        RECT 2619.340 31.660 2619.600 31.920 ;
      LAYER met2 ;
        RECT 2018.350 600.850 2018.630 604.000 ;
        RECT 2018.350 600.710 2020.620 600.850 ;
        RECT 2018.350 600.000 2018.630 600.710 ;
        RECT 2020.480 579.690 2020.620 600.710 ;
        RECT 2019.040 579.370 2019.300 579.690 ;
        RECT 2020.420 579.370 2020.680 579.690 ;
        RECT 2019.100 531.750 2019.240 579.370 ;
        RECT 2019.040 531.430 2019.300 531.750 ;
        RECT 2019.500 531.430 2019.760 531.750 ;
        RECT 2019.560 497.070 2019.700 531.430 ;
        RECT 2019.500 496.750 2019.760 497.070 ;
        RECT 2019.960 496.410 2020.220 496.730 ;
        RECT 2020.020 483.130 2020.160 496.410 ;
        RECT 2018.580 482.810 2018.840 483.130 ;
        RECT 2019.960 482.810 2020.220 483.130 ;
        RECT 2018.640 435.190 2018.780 482.810 ;
        RECT 2018.580 434.870 2018.840 435.190 ;
        RECT 2019.500 434.870 2019.760 435.190 ;
        RECT 2019.560 399.570 2019.700 434.870 ;
        RECT 2019.560 399.430 2020.160 399.570 ;
        RECT 2020.020 379.430 2020.160 399.430 ;
        RECT 2019.040 379.110 2019.300 379.430 ;
        RECT 2019.960 379.110 2020.220 379.430 ;
        RECT 2019.100 331.490 2019.240 379.110 ;
        RECT 2019.040 331.170 2019.300 331.490 ;
        RECT 2020.420 331.170 2020.680 331.490 ;
        RECT 2020.480 304.290 2020.620 331.170 ;
        RECT 2020.420 303.970 2020.680 304.290 ;
        RECT 2019.960 303.290 2020.220 303.610 ;
        RECT 2020.020 282.870 2020.160 303.290 ;
        RECT 2019.040 282.550 2019.300 282.870 ;
        RECT 2019.960 282.550 2020.220 282.870 ;
        RECT 2019.100 234.930 2019.240 282.550 ;
        RECT 2019.040 234.610 2019.300 234.930 ;
        RECT 2020.420 234.610 2020.680 234.930 ;
        RECT 2020.480 218.010 2020.620 234.610 ;
        RECT 2020.020 217.870 2020.620 218.010 ;
        RECT 2020.020 186.650 2020.160 217.870 ;
        RECT 2019.040 186.330 2019.300 186.650 ;
        RECT 2019.960 186.330 2020.220 186.650 ;
        RECT 2019.100 145.170 2019.240 186.330 ;
        RECT 2019.040 144.850 2019.300 145.170 ;
        RECT 2020.420 144.850 2020.680 145.170 ;
        RECT 2020.480 110.830 2020.620 144.850 ;
        RECT 2020.420 110.510 2020.680 110.830 ;
        RECT 2019.960 110.170 2020.220 110.490 ;
        RECT 2020.020 62.290 2020.160 110.170 ;
        RECT 2020.020 62.150 2021.080 62.290 ;
        RECT 2020.940 31.950 2021.080 62.150 ;
        RECT 2020.880 31.630 2021.140 31.950 ;
        RECT 2619.340 31.630 2619.600 31.950 ;
        RECT 2619.400 2.400 2619.540 31.630 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2027.750 31.180 2028.070 31.240 ;
        RECT 2637.250 31.180 2637.570 31.240 ;
        RECT 2027.750 31.040 2637.570 31.180 ;
        RECT 2027.750 30.980 2028.070 31.040 ;
        RECT 2637.250 30.980 2637.570 31.040 ;
      LAYER via ;
        RECT 2027.780 30.980 2028.040 31.240 ;
        RECT 2637.280 30.980 2637.540 31.240 ;
      LAYER met2 ;
        RECT 2027.550 600.000 2027.830 604.000 ;
        RECT 2027.610 598.810 2027.750 600.000 ;
        RECT 2027.610 598.670 2027.980 598.810 ;
        RECT 2027.840 31.270 2027.980 598.670 ;
        RECT 2027.780 30.950 2028.040 31.270 ;
        RECT 2637.280 30.950 2637.540 31.270 ;
        RECT 2637.340 2.400 2637.480 30.950 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2038.330 586.740 2038.650 586.800 ;
        RECT 2042.010 586.740 2042.330 586.800 ;
        RECT 2038.330 586.600 2042.330 586.740 ;
        RECT 2038.330 586.540 2038.650 586.600 ;
        RECT 2042.010 586.540 2042.330 586.600 ;
        RECT 2042.010 31.520 2042.330 31.580 ;
        RECT 2655.190 31.520 2655.510 31.580 ;
        RECT 2042.010 31.380 2655.510 31.520 ;
        RECT 2042.010 31.320 2042.330 31.380 ;
        RECT 2655.190 31.320 2655.510 31.380 ;
      LAYER via ;
        RECT 2038.360 586.540 2038.620 586.800 ;
        RECT 2042.040 586.540 2042.300 586.800 ;
        RECT 2042.040 31.320 2042.300 31.580 ;
        RECT 2655.220 31.320 2655.480 31.580 ;
      LAYER met2 ;
        RECT 2036.750 600.170 2037.030 604.000 ;
        RECT 2036.750 600.030 2038.560 600.170 ;
        RECT 2036.750 600.000 2037.030 600.030 ;
        RECT 2038.420 586.830 2038.560 600.030 ;
        RECT 2038.360 586.510 2038.620 586.830 ;
        RECT 2042.040 586.510 2042.300 586.830 ;
        RECT 2042.100 31.610 2042.240 586.510 ;
        RECT 2042.040 31.290 2042.300 31.610 ;
        RECT 2655.220 31.290 2655.480 31.610 ;
        RECT 2655.280 2.400 2655.420 31.290 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2047.990 30.840 2048.310 30.900 ;
        RECT 2672.670 30.840 2672.990 30.900 ;
        RECT 2047.990 30.700 2672.990 30.840 ;
        RECT 2047.990 30.640 2048.310 30.700 ;
        RECT 2672.670 30.640 2672.990 30.700 ;
      LAYER via ;
        RECT 2048.020 30.640 2048.280 30.900 ;
        RECT 2672.700 30.640 2672.960 30.900 ;
      LAYER met2 ;
        RECT 2045.950 600.170 2046.230 604.000 ;
        RECT 2045.950 600.030 2048.220 600.170 ;
        RECT 2045.950 600.000 2046.230 600.030 ;
        RECT 2048.080 30.930 2048.220 600.030 ;
        RECT 2048.020 30.610 2048.280 30.930 ;
        RECT 2672.700 30.610 2672.960 30.930 ;
        RECT 2672.760 2.400 2672.900 30.610 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2055.150 600.000 2055.430 604.000 ;
        RECT 2055.210 598.810 2055.350 600.000 ;
        RECT 2055.210 598.670 2055.580 598.810 ;
        RECT 2055.440 31.125 2055.580 598.670 ;
        RECT 2055.370 30.755 2055.650 31.125 ;
        RECT 2690.630 30.755 2690.910 31.125 ;
        RECT 2690.700 2.400 2690.840 30.755 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
      LAYER via2 ;
        RECT 2055.370 30.800 2055.650 31.080 ;
        RECT 2690.630 30.800 2690.910 31.080 ;
      LAYER met3 ;
        RECT 2055.345 31.090 2055.675 31.105 ;
        RECT 2690.605 31.090 2690.935 31.105 ;
        RECT 2055.345 30.790 2690.935 31.090 ;
        RECT 2055.345 30.775 2055.675 30.790 ;
        RECT 2690.605 30.775 2690.935 30.790 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2065.930 586.740 2066.250 586.800 ;
        RECT 2069.610 586.740 2069.930 586.800 ;
        RECT 2065.930 586.600 2069.930 586.740 ;
        RECT 2065.930 586.540 2066.250 586.600 ;
        RECT 2069.610 586.540 2069.930 586.600 ;
        RECT 2069.610 39.000 2069.930 39.060 ;
        RECT 2708.550 39.000 2708.870 39.060 ;
        RECT 2069.610 38.860 2708.870 39.000 ;
        RECT 2069.610 38.800 2069.930 38.860 ;
        RECT 2708.550 38.800 2708.870 38.860 ;
      LAYER via ;
        RECT 2065.960 586.540 2066.220 586.800 ;
        RECT 2069.640 586.540 2069.900 586.800 ;
        RECT 2069.640 38.800 2069.900 39.060 ;
        RECT 2708.580 38.800 2708.840 39.060 ;
      LAYER met2 ;
        RECT 2064.350 600.170 2064.630 604.000 ;
        RECT 2064.350 600.030 2066.160 600.170 ;
        RECT 2064.350 600.000 2064.630 600.030 ;
        RECT 2066.020 586.830 2066.160 600.030 ;
        RECT 2065.960 586.510 2066.220 586.830 ;
        RECT 2069.640 586.510 2069.900 586.830 ;
        RECT 2069.700 39.090 2069.840 586.510 ;
        RECT 2069.640 38.770 2069.900 39.090 ;
        RECT 2708.580 38.770 2708.840 39.090 ;
        RECT 2708.640 2.400 2708.780 38.770 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2074.210 579.600 2074.530 579.660 ;
        RECT 2074.670 579.600 2074.990 579.660 ;
        RECT 2074.210 579.460 2074.990 579.600 ;
        RECT 2074.210 579.400 2074.530 579.460 ;
        RECT 2074.670 579.400 2074.990 579.460 ;
        RECT 2074.210 524.180 2074.530 524.240 ;
        RECT 2075.130 524.180 2075.450 524.240 ;
        RECT 2074.210 524.040 2075.450 524.180 ;
        RECT 2074.210 523.980 2074.530 524.040 ;
        RECT 2075.130 523.980 2075.450 524.040 ;
        RECT 2074.210 476.240 2074.530 476.300 ;
        RECT 2076.050 476.240 2076.370 476.300 ;
        RECT 2074.210 476.100 2076.370 476.240 ;
        RECT 2074.210 476.040 2074.530 476.100 ;
        RECT 2076.050 476.040 2076.370 476.100 ;
        RECT 2076.050 448.840 2076.370 449.100 ;
        RECT 2076.140 448.420 2076.280 448.840 ;
        RECT 2076.050 448.160 2076.370 448.420 ;
        RECT 2074.670 434.760 2074.990 434.820 ;
        RECT 2075.590 434.760 2075.910 434.820 ;
        RECT 2074.670 434.620 2075.910 434.760 ;
        RECT 2074.670 434.560 2074.990 434.620 ;
        RECT 2075.590 434.560 2075.910 434.620 ;
        RECT 2074.210 427.620 2074.530 427.680 ;
        RECT 2074.670 427.620 2074.990 427.680 ;
        RECT 2074.210 427.480 2074.990 427.620 ;
        RECT 2074.210 427.420 2074.530 427.480 ;
        RECT 2074.670 427.420 2074.990 427.480 ;
        RECT 2074.210 379.680 2074.530 379.740 ;
        RECT 2075.130 379.680 2075.450 379.740 ;
        RECT 2074.210 379.540 2075.450 379.680 ;
        RECT 2074.210 379.480 2074.530 379.540 ;
        RECT 2075.130 379.480 2075.450 379.540 ;
        RECT 2074.210 331.060 2074.530 331.120 ;
        RECT 2075.130 331.060 2075.450 331.120 ;
        RECT 2074.210 330.920 2075.450 331.060 ;
        RECT 2074.210 330.860 2074.530 330.920 ;
        RECT 2075.130 330.860 2075.450 330.920 ;
        RECT 2074.210 283.120 2074.530 283.180 ;
        RECT 2075.130 283.120 2075.450 283.180 ;
        RECT 2074.210 282.980 2075.450 283.120 ;
        RECT 2074.210 282.920 2074.530 282.980 ;
        RECT 2075.130 282.920 2075.450 282.980 ;
        RECT 2074.210 234.840 2074.530 234.900 ;
        RECT 2074.670 234.840 2074.990 234.900 ;
        RECT 2074.210 234.700 2074.990 234.840 ;
        RECT 2074.210 234.640 2074.530 234.700 ;
        RECT 2074.670 234.640 2074.990 234.700 ;
        RECT 2073.750 227.700 2074.070 227.760 ;
        RECT 2074.210 227.700 2074.530 227.760 ;
        RECT 2073.750 227.560 2074.530 227.700 ;
        RECT 2073.750 227.500 2074.070 227.560 ;
        RECT 2074.210 227.500 2074.530 227.560 ;
        RECT 2074.210 179.760 2074.530 179.820 ;
        RECT 2075.130 179.760 2075.450 179.820 ;
        RECT 2074.210 179.620 2075.450 179.760 ;
        RECT 2074.210 179.560 2074.530 179.620 ;
        RECT 2075.130 179.560 2075.450 179.620 ;
        RECT 2074.210 131.140 2074.530 131.200 ;
        RECT 2075.130 131.140 2075.450 131.200 ;
        RECT 2074.210 131.000 2075.450 131.140 ;
        RECT 2074.210 130.940 2074.530 131.000 ;
        RECT 2075.130 130.940 2075.450 131.000 ;
        RECT 2074.210 83.200 2074.530 83.260 ;
        RECT 2075.130 83.200 2075.450 83.260 ;
        RECT 2074.210 83.060 2075.450 83.200 ;
        RECT 2074.210 83.000 2074.530 83.060 ;
        RECT 2075.130 83.000 2075.450 83.060 ;
        RECT 2075.130 62.460 2075.450 62.520 ;
        RECT 2074.760 62.320 2075.450 62.460 ;
        RECT 2074.760 62.180 2074.900 62.320 ;
        RECT 2075.130 62.260 2075.450 62.320 ;
        RECT 2074.670 61.920 2074.990 62.180 ;
        RECT 2074.670 38.660 2074.990 38.720 ;
        RECT 2726.490 38.660 2726.810 38.720 ;
        RECT 2074.670 38.520 2726.810 38.660 ;
        RECT 2074.670 38.460 2074.990 38.520 ;
        RECT 2726.490 38.460 2726.810 38.520 ;
      LAYER via ;
        RECT 2074.240 579.400 2074.500 579.660 ;
        RECT 2074.700 579.400 2074.960 579.660 ;
        RECT 2074.240 523.980 2074.500 524.240 ;
        RECT 2075.160 523.980 2075.420 524.240 ;
        RECT 2074.240 476.040 2074.500 476.300 ;
        RECT 2076.080 476.040 2076.340 476.300 ;
        RECT 2076.080 448.840 2076.340 449.100 ;
        RECT 2076.080 448.160 2076.340 448.420 ;
        RECT 2074.700 434.560 2074.960 434.820 ;
        RECT 2075.620 434.560 2075.880 434.820 ;
        RECT 2074.240 427.420 2074.500 427.680 ;
        RECT 2074.700 427.420 2074.960 427.680 ;
        RECT 2074.240 379.480 2074.500 379.740 ;
        RECT 2075.160 379.480 2075.420 379.740 ;
        RECT 2074.240 330.860 2074.500 331.120 ;
        RECT 2075.160 330.860 2075.420 331.120 ;
        RECT 2074.240 282.920 2074.500 283.180 ;
        RECT 2075.160 282.920 2075.420 283.180 ;
        RECT 2074.240 234.640 2074.500 234.900 ;
        RECT 2074.700 234.640 2074.960 234.900 ;
        RECT 2073.780 227.500 2074.040 227.760 ;
        RECT 2074.240 227.500 2074.500 227.760 ;
        RECT 2074.240 179.560 2074.500 179.820 ;
        RECT 2075.160 179.560 2075.420 179.820 ;
        RECT 2074.240 130.940 2074.500 131.200 ;
        RECT 2075.160 130.940 2075.420 131.200 ;
        RECT 2074.240 83.000 2074.500 83.260 ;
        RECT 2075.160 83.000 2075.420 83.260 ;
        RECT 2075.160 62.260 2075.420 62.520 ;
        RECT 2074.700 61.920 2074.960 62.180 ;
        RECT 2074.700 38.460 2074.960 38.720 ;
        RECT 2726.520 38.460 2726.780 38.720 ;
      LAYER met2 ;
        RECT 2073.550 600.850 2073.830 604.000 ;
        RECT 2073.550 600.710 2074.440 600.850 ;
        RECT 2073.550 600.000 2073.830 600.710 ;
        RECT 2074.300 579.690 2074.440 600.710 ;
        RECT 2074.240 579.370 2074.500 579.690 ;
        RECT 2074.700 579.370 2074.960 579.690 ;
        RECT 2074.760 544.410 2074.900 579.370 ;
        RECT 2074.760 544.270 2075.360 544.410 ;
        RECT 2075.220 524.270 2075.360 544.270 ;
        RECT 2074.240 523.950 2074.500 524.270 ;
        RECT 2075.160 523.950 2075.420 524.270 ;
        RECT 2074.300 476.330 2074.440 523.950 ;
        RECT 2074.240 476.010 2074.500 476.330 ;
        RECT 2076.080 476.010 2076.340 476.330 ;
        RECT 2076.140 449.130 2076.280 476.010 ;
        RECT 2076.080 448.810 2076.340 449.130 ;
        RECT 2076.080 448.130 2076.340 448.450 ;
        RECT 2076.140 434.930 2076.280 448.130 ;
        RECT 2075.680 434.850 2076.280 434.930 ;
        RECT 2074.700 434.530 2074.960 434.850 ;
        RECT 2075.620 434.790 2076.280 434.850 ;
        RECT 2075.620 434.530 2075.880 434.790 ;
        RECT 2074.760 427.710 2074.900 434.530 ;
        RECT 2074.240 427.390 2074.500 427.710 ;
        RECT 2074.700 427.390 2074.960 427.710 ;
        RECT 2074.300 379.770 2074.440 427.390 ;
        RECT 2074.240 379.450 2074.500 379.770 ;
        RECT 2075.160 379.450 2075.420 379.770 ;
        RECT 2075.220 331.150 2075.360 379.450 ;
        RECT 2074.240 330.830 2074.500 331.150 ;
        RECT 2075.160 330.830 2075.420 331.150 ;
        RECT 2074.300 283.210 2074.440 330.830 ;
        RECT 2074.240 282.890 2074.500 283.210 ;
        RECT 2075.160 282.890 2075.420 283.210 ;
        RECT 2075.220 258.810 2075.360 282.890 ;
        RECT 2074.300 258.670 2075.360 258.810 ;
        RECT 2074.300 234.930 2074.440 258.670 ;
        RECT 2074.240 234.610 2074.500 234.930 ;
        RECT 2074.700 234.610 2074.960 234.930 ;
        RECT 2074.760 234.445 2074.900 234.610 ;
        RECT 2073.770 234.075 2074.050 234.445 ;
        RECT 2074.690 234.075 2074.970 234.445 ;
        RECT 2073.840 227.790 2073.980 234.075 ;
        RECT 2073.780 227.470 2074.040 227.790 ;
        RECT 2074.240 227.470 2074.500 227.790 ;
        RECT 2074.300 179.850 2074.440 227.470 ;
        RECT 2074.240 179.530 2074.500 179.850 ;
        RECT 2075.160 179.530 2075.420 179.850 ;
        RECT 2075.220 131.230 2075.360 179.530 ;
        RECT 2074.240 130.910 2074.500 131.230 ;
        RECT 2075.160 130.910 2075.420 131.230 ;
        RECT 2074.300 83.290 2074.440 130.910 ;
        RECT 2074.240 82.970 2074.500 83.290 ;
        RECT 2075.160 82.970 2075.420 83.290 ;
        RECT 2075.220 62.550 2075.360 82.970 ;
        RECT 2075.160 62.230 2075.420 62.550 ;
        RECT 2074.700 61.890 2074.960 62.210 ;
        RECT 2074.760 38.750 2074.900 61.890 ;
        RECT 2074.700 38.430 2074.960 38.750 ;
        RECT 2726.520 38.430 2726.780 38.750 ;
        RECT 2726.580 2.400 2726.720 38.430 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
      LAYER via2 ;
        RECT 2073.770 234.120 2074.050 234.400 ;
        RECT 2074.690 234.120 2074.970 234.400 ;
      LAYER met3 ;
        RECT 2073.745 234.410 2074.075 234.425 ;
        RECT 2074.665 234.410 2074.995 234.425 ;
        RECT 2073.745 234.110 2074.995 234.410 ;
        RECT 2073.745 234.095 2074.075 234.110 ;
        RECT 2074.665 234.095 2074.995 234.110 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2082.950 38.320 2083.270 38.380 ;
        RECT 2744.430 38.320 2744.750 38.380 ;
        RECT 2082.950 38.180 2744.750 38.320 ;
        RECT 2082.950 38.120 2083.270 38.180 ;
        RECT 2744.430 38.120 2744.750 38.180 ;
      LAYER via ;
        RECT 2082.980 38.120 2083.240 38.380 ;
        RECT 2744.460 38.120 2744.720 38.380 ;
      LAYER met2 ;
        RECT 2082.750 600.000 2083.030 604.000 ;
        RECT 2082.810 598.810 2082.950 600.000 ;
        RECT 2082.810 598.670 2083.180 598.810 ;
        RECT 2083.040 38.410 2083.180 598.670 ;
        RECT 2082.980 38.090 2083.240 38.410 ;
        RECT 2744.460 38.090 2744.720 38.410 ;
        RECT 2744.520 2.400 2744.660 38.090 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2093.070 587.420 2093.390 587.480 ;
        RECT 2097.210 587.420 2097.530 587.480 ;
        RECT 2093.070 587.280 2097.530 587.420 ;
        RECT 2093.070 587.220 2093.390 587.280 ;
        RECT 2097.210 587.220 2097.530 587.280 ;
        RECT 2097.210 47.160 2097.530 47.220 ;
        RECT 2761.910 47.160 2762.230 47.220 ;
        RECT 2097.210 47.020 2762.230 47.160 ;
        RECT 2097.210 46.960 2097.530 47.020 ;
        RECT 2761.910 46.960 2762.230 47.020 ;
      LAYER via ;
        RECT 2093.100 587.220 2093.360 587.480 ;
        RECT 2097.240 587.220 2097.500 587.480 ;
        RECT 2097.240 46.960 2097.500 47.220 ;
        RECT 2761.940 46.960 2762.200 47.220 ;
      LAYER met2 ;
        RECT 2091.490 600.170 2091.770 604.000 ;
        RECT 2091.490 600.030 2093.300 600.170 ;
        RECT 2091.490 600.000 2091.770 600.030 ;
        RECT 2093.160 587.510 2093.300 600.030 ;
        RECT 2093.100 587.190 2093.360 587.510 ;
        RECT 2097.240 587.190 2097.500 587.510 ;
        RECT 2097.300 47.250 2097.440 587.190 ;
        RECT 2097.240 46.930 2097.500 47.250 ;
        RECT 2761.940 46.930 2762.200 47.250 ;
        RECT 2762.000 2.400 2762.140 46.930 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1097.630 569.400 1097.950 569.460 ;
        RECT 1098.550 569.400 1098.870 569.460 ;
        RECT 1097.630 569.260 1098.870 569.400 ;
        RECT 1097.630 569.200 1097.950 569.260 ;
        RECT 1098.550 569.200 1098.870 569.260 ;
        RECT 835.430 26.420 835.750 26.480 ;
        RECT 1097.630 26.420 1097.950 26.480 ;
        RECT 835.430 26.280 1097.950 26.420 ;
        RECT 835.430 26.220 835.750 26.280 ;
        RECT 1097.630 26.220 1097.950 26.280 ;
      LAYER via ;
        RECT 1097.660 569.200 1097.920 569.460 ;
        RECT 1098.580 569.200 1098.840 569.460 ;
        RECT 835.460 26.220 835.720 26.480 ;
        RECT 1097.660 26.220 1097.920 26.480 ;
      LAYER met2 ;
        RECT 1099.730 600.170 1100.010 604.000 ;
        RECT 1098.640 600.030 1100.010 600.170 ;
        RECT 1098.640 569.490 1098.780 600.030 ;
        RECT 1099.730 600.000 1100.010 600.030 ;
        RECT 1097.660 569.170 1097.920 569.490 ;
        RECT 1098.580 569.170 1098.840 569.490 ;
        RECT 1097.720 26.510 1097.860 569.170 ;
        RECT 835.460 26.190 835.720 26.510 ;
        RECT 1097.660 26.190 1097.920 26.510 ;
        RECT 835.520 2.400 835.660 26.190 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2102.730 579.600 2103.050 579.660 ;
        RECT 2103.190 579.600 2103.510 579.660 ;
        RECT 2102.730 579.460 2103.510 579.600 ;
        RECT 2102.730 579.400 2103.050 579.460 ;
        RECT 2103.190 579.400 2103.510 579.460 ;
        RECT 2103.190 545.260 2103.510 545.320 ;
        RECT 2102.820 545.120 2103.510 545.260 ;
        RECT 2102.820 544.980 2102.960 545.120 ;
        RECT 2103.190 545.060 2103.510 545.120 ;
        RECT 2102.730 544.720 2103.050 544.980 ;
        RECT 2102.730 531.320 2103.050 531.380 ;
        RECT 2103.190 531.320 2103.510 531.380 ;
        RECT 2102.730 531.180 2103.510 531.320 ;
        RECT 2102.730 531.120 2103.050 531.180 ;
        RECT 2103.190 531.120 2103.510 531.180 ;
        RECT 2102.730 483.040 2103.050 483.100 ;
        RECT 2103.650 483.040 2103.970 483.100 ;
        RECT 2102.730 482.900 2103.970 483.040 ;
        RECT 2102.730 482.840 2103.050 482.900 ;
        RECT 2103.650 482.840 2103.970 482.900 ;
        RECT 2102.730 435.100 2103.050 435.160 ;
        RECT 2103.190 435.100 2103.510 435.160 ;
        RECT 2102.730 434.960 2103.510 435.100 ;
        RECT 2102.730 434.900 2103.050 434.960 ;
        RECT 2103.190 434.900 2103.510 434.960 ;
        RECT 2102.730 387.160 2103.050 387.220 ;
        RECT 2102.730 387.020 2103.420 387.160 ;
        RECT 2102.730 386.960 2103.050 387.020 ;
        RECT 2103.280 386.540 2103.420 387.020 ;
        RECT 2103.190 386.280 2103.510 386.540 ;
        RECT 2102.730 338.540 2103.050 338.600 ;
        RECT 2103.190 338.540 2103.510 338.600 ;
        RECT 2102.730 338.400 2103.510 338.540 ;
        RECT 2102.730 338.340 2103.050 338.400 ;
        RECT 2103.190 338.340 2103.510 338.400 ;
        RECT 2101.350 282.780 2101.670 282.840 ;
        RECT 2102.730 282.780 2103.050 282.840 ;
        RECT 2101.350 282.640 2103.050 282.780 ;
        RECT 2101.350 282.580 2101.670 282.640 ;
        RECT 2102.730 282.580 2103.050 282.640 ;
        RECT 2101.350 234.840 2101.670 234.900 ;
        RECT 2102.270 234.840 2102.590 234.900 ;
        RECT 2101.350 234.700 2102.590 234.840 ;
        RECT 2101.350 234.640 2101.670 234.700 ;
        RECT 2102.270 234.640 2102.590 234.700 ;
        RECT 2101.350 137.940 2101.670 138.000 ;
        RECT 2102.270 137.940 2102.590 138.000 ;
        RECT 2101.350 137.800 2102.590 137.940 ;
        RECT 2101.350 137.740 2101.670 137.800 ;
        RECT 2102.270 137.740 2102.590 137.800 ;
        RECT 2101.350 90.000 2101.670 90.060 ;
        RECT 2102.730 90.000 2103.050 90.060 ;
        RECT 2101.350 89.860 2103.050 90.000 ;
        RECT 2101.350 89.800 2101.670 89.860 ;
        RECT 2102.730 89.800 2103.050 89.860 ;
        RECT 2102.730 62.460 2103.050 62.520 ;
        RECT 2102.360 62.320 2103.050 62.460 ;
        RECT 2102.360 62.180 2102.500 62.320 ;
        RECT 2102.730 62.260 2103.050 62.320 ;
        RECT 2102.270 61.920 2102.590 62.180 ;
        RECT 2102.270 46.820 2102.590 46.880 ;
        RECT 2779.850 46.820 2780.170 46.880 ;
        RECT 2102.270 46.680 2780.170 46.820 ;
        RECT 2102.270 46.620 2102.590 46.680 ;
        RECT 2779.850 46.620 2780.170 46.680 ;
      LAYER via ;
        RECT 2102.760 579.400 2103.020 579.660 ;
        RECT 2103.220 579.400 2103.480 579.660 ;
        RECT 2103.220 545.060 2103.480 545.320 ;
        RECT 2102.760 544.720 2103.020 544.980 ;
        RECT 2102.760 531.120 2103.020 531.380 ;
        RECT 2103.220 531.120 2103.480 531.380 ;
        RECT 2102.760 482.840 2103.020 483.100 ;
        RECT 2103.680 482.840 2103.940 483.100 ;
        RECT 2102.760 434.900 2103.020 435.160 ;
        RECT 2103.220 434.900 2103.480 435.160 ;
        RECT 2102.760 386.960 2103.020 387.220 ;
        RECT 2103.220 386.280 2103.480 386.540 ;
        RECT 2102.760 338.340 2103.020 338.600 ;
        RECT 2103.220 338.340 2103.480 338.600 ;
        RECT 2101.380 282.580 2101.640 282.840 ;
        RECT 2102.760 282.580 2103.020 282.840 ;
        RECT 2101.380 234.640 2101.640 234.900 ;
        RECT 2102.300 234.640 2102.560 234.900 ;
        RECT 2101.380 137.740 2101.640 138.000 ;
        RECT 2102.300 137.740 2102.560 138.000 ;
        RECT 2101.380 89.800 2101.640 90.060 ;
        RECT 2102.760 89.800 2103.020 90.060 ;
        RECT 2102.760 62.260 2103.020 62.520 ;
        RECT 2102.300 61.920 2102.560 62.180 ;
        RECT 2102.300 46.620 2102.560 46.880 ;
        RECT 2779.880 46.620 2780.140 46.880 ;
      LAYER met2 ;
        RECT 2100.690 600.850 2100.970 604.000 ;
        RECT 2100.690 600.710 2102.040 600.850 ;
        RECT 2100.690 600.000 2100.970 600.710 ;
        RECT 2101.900 589.970 2102.040 600.710 ;
        RECT 2101.900 589.830 2102.960 589.970 ;
        RECT 2102.820 579.690 2102.960 589.830 ;
        RECT 2102.760 579.370 2103.020 579.690 ;
        RECT 2103.220 579.370 2103.480 579.690 ;
        RECT 2103.280 545.350 2103.420 579.370 ;
        RECT 2103.220 545.030 2103.480 545.350 ;
        RECT 2102.760 544.690 2103.020 545.010 ;
        RECT 2102.820 531.490 2102.960 544.690 ;
        RECT 2102.820 531.410 2103.420 531.490 ;
        RECT 2102.760 531.350 2103.480 531.410 ;
        RECT 2102.760 531.090 2103.020 531.350 ;
        RECT 2103.220 531.090 2103.480 531.350 ;
        RECT 2102.820 496.810 2102.960 531.090 ;
        RECT 2102.820 496.670 2103.420 496.810 ;
        RECT 2103.280 483.210 2103.420 496.670 ;
        RECT 2103.280 483.130 2103.880 483.210 ;
        RECT 2102.760 482.810 2103.020 483.130 ;
        RECT 2103.280 483.070 2103.940 483.130 ;
        RECT 2103.680 482.810 2103.940 483.070 ;
        RECT 2102.820 435.190 2102.960 482.810 ;
        RECT 2103.740 482.655 2103.880 482.810 ;
        RECT 2102.760 434.870 2103.020 435.190 ;
        RECT 2103.220 434.870 2103.480 435.190 ;
        RECT 2103.280 410.450 2103.420 434.870 ;
        RECT 2102.820 410.310 2103.420 410.450 ;
        RECT 2102.820 387.250 2102.960 410.310 ;
        RECT 2102.760 386.930 2103.020 387.250 ;
        RECT 2103.220 386.480 2103.480 386.570 ;
        RECT 2102.820 386.340 2103.480 386.480 ;
        RECT 2102.820 352.650 2102.960 386.340 ;
        RECT 2103.220 386.250 2103.480 386.340 ;
        RECT 2102.820 352.510 2103.420 352.650 ;
        RECT 2103.280 338.630 2103.420 352.510 ;
        RECT 2102.760 338.370 2103.020 338.630 ;
        RECT 2102.360 338.310 2103.020 338.370 ;
        RECT 2103.220 338.310 2103.480 338.630 ;
        RECT 2102.360 338.230 2102.960 338.310 ;
        RECT 2102.360 307.090 2102.500 338.230 ;
        RECT 2102.360 306.950 2103.420 307.090 ;
        RECT 2103.280 284.085 2103.420 306.950 ;
        RECT 2103.210 283.715 2103.490 284.085 ;
        RECT 2102.750 283.035 2103.030 283.405 ;
        RECT 2102.820 282.870 2102.960 283.035 ;
        RECT 2101.380 282.550 2101.640 282.870 ;
        RECT 2102.760 282.550 2103.020 282.870 ;
        RECT 2101.440 234.930 2101.580 282.550 ;
        RECT 2101.380 234.610 2101.640 234.930 ;
        RECT 2102.300 234.610 2102.560 234.930 ;
        RECT 2102.360 210.530 2102.500 234.610 ;
        RECT 2102.360 210.390 2102.960 210.530 ;
        RECT 2102.820 159.645 2102.960 210.390 ;
        RECT 2102.750 159.275 2103.030 159.645 ;
        RECT 2102.290 144.995 2102.570 145.365 ;
        RECT 2102.360 138.030 2102.500 144.995 ;
        RECT 2101.380 137.710 2101.640 138.030 ;
        RECT 2102.300 137.710 2102.560 138.030 ;
        RECT 2101.440 90.090 2101.580 137.710 ;
        RECT 2101.380 89.770 2101.640 90.090 ;
        RECT 2102.760 89.770 2103.020 90.090 ;
        RECT 2102.820 62.550 2102.960 89.770 ;
        RECT 2102.760 62.230 2103.020 62.550 ;
        RECT 2102.300 61.890 2102.560 62.210 ;
        RECT 2102.360 46.910 2102.500 61.890 ;
        RECT 2102.300 46.590 2102.560 46.910 ;
        RECT 2779.880 46.590 2780.140 46.910 ;
        RECT 2779.940 2.400 2780.080 46.590 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
      LAYER via2 ;
        RECT 2103.210 283.760 2103.490 284.040 ;
        RECT 2102.750 283.080 2103.030 283.360 ;
        RECT 2102.750 159.320 2103.030 159.600 ;
        RECT 2102.290 145.040 2102.570 145.320 ;
      LAYER met3 ;
        RECT 2103.185 284.050 2103.515 284.065 ;
        RECT 2103.185 283.735 2103.730 284.050 ;
        RECT 2102.725 283.370 2103.055 283.385 ;
        RECT 2103.430 283.370 2103.730 283.735 ;
        RECT 2102.725 283.070 2103.730 283.370 ;
        RECT 2102.725 283.055 2103.055 283.070 ;
        RECT 2102.725 159.620 2103.055 159.625 ;
        RECT 2102.470 159.610 2103.055 159.620 ;
        RECT 2102.270 159.310 2103.055 159.610 ;
        RECT 2102.470 159.300 2103.055 159.310 ;
        RECT 2102.725 159.295 2103.055 159.300 ;
        RECT 2102.265 145.340 2102.595 145.345 ;
        RECT 2102.265 145.330 2102.850 145.340 ;
        RECT 2102.265 145.030 2103.050 145.330 ;
        RECT 2102.265 145.020 2102.850 145.030 ;
        RECT 2102.265 145.015 2102.595 145.020 ;
      LAYER via3 ;
        RECT 2102.500 159.300 2102.820 159.620 ;
        RECT 2102.500 145.020 2102.820 145.340 ;
      LAYER met4 ;
        RECT 2102.495 159.295 2102.825 159.625 ;
        RECT 2102.510 145.345 2102.810 159.295 ;
        RECT 2102.495 145.015 2102.825 145.345 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2110.550 46.480 2110.870 46.540 ;
        RECT 2797.790 46.480 2798.110 46.540 ;
        RECT 2110.550 46.340 2798.110 46.480 ;
        RECT 2110.550 46.280 2110.870 46.340 ;
        RECT 2797.790 46.280 2798.110 46.340 ;
      LAYER via ;
        RECT 2110.580 46.280 2110.840 46.540 ;
        RECT 2797.820 46.280 2798.080 46.540 ;
      LAYER met2 ;
        RECT 2109.890 600.170 2110.170 604.000 ;
        RECT 2109.890 600.030 2110.780 600.170 ;
        RECT 2109.890 600.000 2110.170 600.030 ;
        RECT 2110.640 46.570 2110.780 600.030 ;
        RECT 2110.580 46.250 2110.840 46.570 ;
        RECT 2797.820 46.250 2798.080 46.570 ;
        RECT 2797.880 2.400 2798.020 46.250 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2120.670 587.420 2120.990 587.480 ;
        RECT 2124.810 587.420 2125.130 587.480 ;
        RECT 2120.670 587.280 2125.130 587.420 ;
        RECT 2120.670 587.220 2120.990 587.280 ;
        RECT 2124.810 587.220 2125.130 587.280 ;
        RECT 2124.810 46.140 2125.130 46.200 ;
        RECT 2815.730 46.140 2816.050 46.200 ;
        RECT 2124.810 46.000 2816.050 46.140 ;
        RECT 2124.810 45.940 2125.130 46.000 ;
        RECT 2815.730 45.940 2816.050 46.000 ;
      LAYER via ;
        RECT 2120.700 587.220 2120.960 587.480 ;
        RECT 2124.840 587.220 2125.100 587.480 ;
        RECT 2124.840 45.940 2125.100 46.200 ;
        RECT 2815.760 45.940 2816.020 46.200 ;
      LAYER met2 ;
        RECT 2119.090 600.170 2119.370 604.000 ;
        RECT 2119.090 600.030 2120.900 600.170 ;
        RECT 2119.090 600.000 2119.370 600.030 ;
        RECT 2120.760 587.510 2120.900 600.030 ;
        RECT 2120.700 587.190 2120.960 587.510 ;
        RECT 2124.840 587.190 2125.100 587.510 ;
        RECT 2124.900 46.230 2125.040 587.190 ;
        RECT 2124.840 45.910 2125.100 46.230 ;
        RECT 2815.760 45.910 2816.020 46.230 ;
        RECT 2815.820 2.400 2815.960 45.910 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2129.410 579.600 2129.730 579.660 ;
        RECT 2130.330 579.600 2130.650 579.660 ;
        RECT 2129.410 579.460 2130.650 579.600 ;
        RECT 2129.410 579.400 2129.730 579.460 ;
        RECT 2130.330 579.400 2130.650 579.460 ;
        RECT 2130.330 531.320 2130.650 531.380 ;
        RECT 2130.330 531.180 2131.480 531.320 ;
        RECT 2130.330 531.120 2130.650 531.180 ;
        RECT 2131.340 531.040 2131.480 531.180 ;
        RECT 2131.250 530.780 2131.570 531.040 ;
        RECT 2129.410 458.900 2129.730 458.960 ;
        RECT 2130.790 458.900 2131.110 458.960 ;
        RECT 2129.410 458.760 2131.110 458.900 ;
        RECT 2129.410 458.700 2129.730 458.760 ;
        RECT 2130.790 458.700 2131.110 458.760 ;
        RECT 2129.410 435.440 2129.730 435.500 ;
        RECT 2130.790 435.440 2131.110 435.500 ;
        RECT 2129.410 435.300 2131.110 435.440 ;
        RECT 2129.410 435.240 2129.730 435.300 ;
        RECT 2130.790 435.240 2131.110 435.300 ;
        RECT 2130.330 379.340 2130.650 379.400 ;
        RECT 2131.250 379.340 2131.570 379.400 ;
        RECT 2130.330 379.200 2131.570 379.340 ;
        RECT 2130.330 379.140 2130.650 379.200 ;
        RECT 2131.250 379.140 2131.570 379.200 ;
        RECT 2130.330 324.260 2130.650 324.320 ;
        RECT 2130.790 324.260 2131.110 324.320 ;
        RECT 2130.330 324.120 2131.110 324.260 ;
        RECT 2130.330 324.060 2130.650 324.120 ;
        RECT 2130.790 324.060 2131.110 324.120 ;
        RECT 2130.330 276.320 2130.650 276.380 ;
        RECT 2130.790 276.320 2131.110 276.380 ;
        RECT 2130.330 276.180 2131.110 276.320 ;
        RECT 2130.330 276.120 2130.650 276.180 ;
        RECT 2130.790 276.120 2131.110 276.180 ;
        RECT 2129.870 255.580 2130.190 255.640 ;
        RECT 2129.870 255.440 2130.560 255.580 ;
        RECT 2129.870 255.380 2130.190 255.440 ;
        RECT 2130.420 255.300 2130.560 255.440 ;
        RECT 2130.330 255.040 2130.650 255.300 ;
        RECT 2129.870 228.040 2130.190 228.100 ;
        RECT 2130.330 228.040 2130.650 228.100 ;
        RECT 2129.870 227.900 2130.650 228.040 ;
        RECT 2129.870 227.840 2130.190 227.900 ;
        RECT 2130.330 227.840 2130.650 227.900 ;
        RECT 2130.330 138.280 2130.650 138.340 ;
        RECT 2130.790 138.280 2131.110 138.340 ;
        RECT 2130.330 138.140 2131.110 138.280 ;
        RECT 2130.330 138.080 2130.650 138.140 ;
        RECT 2130.790 138.080 2131.110 138.140 ;
        RECT 2130.330 131.140 2130.650 131.200 ;
        RECT 2140.910 131.140 2141.230 131.200 ;
        RECT 2130.330 131.000 2141.230 131.140 ;
        RECT 2130.330 130.940 2130.650 131.000 ;
        RECT 2140.910 130.940 2141.230 131.000 ;
        RECT 2140.910 45.800 2141.230 45.860 ;
        RECT 2833.670 45.800 2833.990 45.860 ;
        RECT 2140.910 45.660 2833.990 45.800 ;
        RECT 2140.910 45.600 2141.230 45.660 ;
        RECT 2833.670 45.600 2833.990 45.660 ;
      LAYER via ;
        RECT 2129.440 579.400 2129.700 579.660 ;
        RECT 2130.360 579.400 2130.620 579.660 ;
        RECT 2130.360 531.120 2130.620 531.380 ;
        RECT 2131.280 530.780 2131.540 531.040 ;
        RECT 2129.440 458.700 2129.700 458.960 ;
        RECT 2130.820 458.700 2131.080 458.960 ;
        RECT 2129.440 435.240 2129.700 435.500 ;
        RECT 2130.820 435.240 2131.080 435.500 ;
        RECT 2130.360 379.140 2130.620 379.400 ;
        RECT 2131.280 379.140 2131.540 379.400 ;
        RECT 2130.360 324.060 2130.620 324.320 ;
        RECT 2130.820 324.060 2131.080 324.320 ;
        RECT 2130.360 276.120 2130.620 276.380 ;
        RECT 2130.820 276.120 2131.080 276.380 ;
        RECT 2129.900 255.380 2130.160 255.640 ;
        RECT 2130.360 255.040 2130.620 255.300 ;
        RECT 2129.900 227.840 2130.160 228.100 ;
        RECT 2130.360 227.840 2130.620 228.100 ;
        RECT 2130.360 138.080 2130.620 138.340 ;
        RECT 2130.820 138.080 2131.080 138.340 ;
        RECT 2130.360 130.940 2130.620 131.200 ;
        RECT 2140.940 130.940 2141.200 131.200 ;
        RECT 2140.940 45.600 2141.200 45.860 ;
        RECT 2833.700 45.600 2833.960 45.860 ;
      LAYER met2 ;
        RECT 2128.290 600.000 2128.570 604.000 ;
        RECT 2128.350 598.810 2128.490 600.000 ;
        RECT 2128.350 598.670 2128.720 598.810 ;
        RECT 2128.580 580.565 2128.720 598.670 ;
        RECT 2128.510 580.195 2128.790 580.565 ;
        RECT 2129.440 579.370 2129.700 579.690 ;
        RECT 2130.350 579.515 2130.630 579.885 ;
        RECT 2130.360 579.370 2130.620 579.515 ;
        RECT 2129.500 544.410 2129.640 579.370 ;
        RECT 2129.500 544.270 2130.560 544.410 ;
        RECT 2130.420 531.410 2130.560 544.270 ;
        RECT 2130.360 531.090 2130.620 531.410 ;
        RECT 2131.280 530.750 2131.540 531.070 ;
        RECT 2131.340 496.810 2131.480 530.750 ;
        RECT 2130.880 496.670 2131.480 496.810 ;
        RECT 2130.880 458.990 2131.020 496.670 ;
        RECT 2129.440 458.670 2129.700 458.990 ;
        RECT 2130.820 458.670 2131.080 458.990 ;
        RECT 2129.500 435.530 2129.640 458.670 ;
        RECT 2129.440 435.210 2129.700 435.530 ;
        RECT 2130.820 435.210 2131.080 435.530 ;
        RECT 2130.880 403.650 2131.020 435.210 ;
        RECT 2130.420 403.510 2131.020 403.650 ;
        RECT 2130.420 379.430 2130.560 403.510 ;
        RECT 2130.360 379.110 2130.620 379.430 ;
        RECT 2131.280 379.110 2131.540 379.430 ;
        RECT 2131.340 331.685 2131.480 379.110 ;
        RECT 2130.350 331.315 2130.630 331.685 ;
        RECT 2131.270 331.315 2131.550 331.685 ;
        RECT 2130.420 324.350 2130.560 331.315 ;
        RECT 2130.360 324.030 2130.620 324.350 ;
        RECT 2130.820 324.030 2131.080 324.350 ;
        RECT 2130.880 276.410 2131.020 324.030 ;
        RECT 2130.360 276.090 2130.620 276.410 ;
        RECT 2130.820 276.090 2131.080 276.410 ;
        RECT 2130.420 275.810 2130.560 276.090 ;
        RECT 2129.960 275.670 2130.560 275.810 ;
        RECT 2129.960 255.670 2130.100 275.670 ;
        RECT 2129.900 255.350 2130.160 255.670 ;
        RECT 2130.360 255.010 2130.620 255.330 ;
        RECT 2130.420 228.130 2130.560 255.010 ;
        RECT 2129.900 227.810 2130.160 228.130 ;
        RECT 2130.360 227.810 2130.620 228.130 ;
        RECT 2129.960 227.530 2130.100 227.810 ;
        RECT 2129.960 227.390 2131.020 227.530 ;
        RECT 2130.880 206.450 2131.020 227.390 ;
        RECT 2130.420 206.310 2131.020 206.450 ;
        RECT 2130.420 159.530 2130.560 206.310 ;
        RECT 2130.420 159.390 2131.020 159.530 ;
        RECT 2130.880 138.370 2131.020 159.390 ;
        RECT 2130.360 138.050 2130.620 138.370 ;
        RECT 2130.820 138.050 2131.080 138.370 ;
        RECT 2130.420 131.230 2130.560 138.050 ;
        RECT 2130.360 130.910 2130.620 131.230 ;
        RECT 2140.940 130.910 2141.200 131.230 ;
        RECT 2141.000 45.890 2141.140 130.910 ;
        RECT 2140.940 45.570 2141.200 45.890 ;
        RECT 2833.700 45.570 2833.960 45.890 ;
        RECT 2833.760 2.400 2833.900 45.570 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
      LAYER via2 ;
        RECT 2128.510 580.240 2128.790 580.520 ;
        RECT 2130.350 579.560 2130.630 579.840 ;
        RECT 2130.350 331.360 2130.630 331.640 ;
        RECT 2131.270 331.360 2131.550 331.640 ;
      LAYER met3 ;
        RECT 2128.485 580.530 2128.815 580.545 ;
        RECT 2128.485 580.230 2131.330 580.530 ;
        RECT 2128.485 580.215 2128.815 580.230 ;
        RECT 2130.325 579.850 2130.655 579.865 ;
        RECT 2131.030 579.850 2131.330 580.230 ;
        RECT 2130.325 579.550 2131.330 579.850 ;
        RECT 2130.325 579.535 2130.655 579.550 ;
        RECT 2130.325 331.650 2130.655 331.665 ;
        RECT 2131.245 331.650 2131.575 331.665 ;
        RECT 2130.325 331.350 2131.575 331.650 ;
        RECT 2130.325 331.335 2130.655 331.350 ;
        RECT 2131.245 331.335 2131.575 331.350 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2138.150 45.460 2138.470 45.520 ;
        RECT 2851.150 45.460 2851.470 45.520 ;
        RECT 2138.150 45.320 2851.470 45.460 ;
        RECT 2138.150 45.260 2138.470 45.320 ;
        RECT 2851.150 45.260 2851.470 45.320 ;
      LAYER via ;
        RECT 2138.180 45.260 2138.440 45.520 ;
        RECT 2851.180 45.260 2851.440 45.520 ;
      LAYER met2 ;
        RECT 2137.490 600.170 2137.770 604.000 ;
        RECT 2137.490 600.030 2138.380 600.170 ;
        RECT 2137.490 600.000 2137.770 600.030 ;
        RECT 2138.240 45.550 2138.380 600.030 ;
        RECT 2138.180 45.230 2138.440 45.550 ;
        RECT 2851.180 45.230 2851.440 45.550 ;
        RECT 2851.240 2.400 2851.380 45.230 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2148.270 588.440 2148.590 588.500 ;
        RECT 2152.410 588.440 2152.730 588.500 ;
        RECT 2148.270 588.300 2152.730 588.440 ;
        RECT 2148.270 588.240 2148.590 588.300 ;
        RECT 2152.410 588.240 2152.730 588.300 ;
        RECT 2152.410 37.980 2152.730 38.040 ;
        RECT 2869.090 37.980 2869.410 38.040 ;
        RECT 2152.410 37.840 2869.410 37.980 ;
        RECT 2152.410 37.780 2152.730 37.840 ;
        RECT 2869.090 37.780 2869.410 37.840 ;
      LAYER via ;
        RECT 2148.300 588.240 2148.560 588.500 ;
        RECT 2152.440 588.240 2152.700 588.500 ;
        RECT 2152.440 37.780 2152.700 38.040 ;
        RECT 2869.120 37.780 2869.380 38.040 ;
      LAYER met2 ;
        RECT 2146.690 600.170 2146.970 604.000 ;
        RECT 2146.690 600.030 2148.500 600.170 ;
        RECT 2146.690 600.000 2146.970 600.030 ;
        RECT 2148.360 588.530 2148.500 600.030 ;
        RECT 2148.300 588.210 2148.560 588.530 ;
        RECT 2152.440 588.210 2152.700 588.530 ;
        RECT 2152.500 38.070 2152.640 588.210 ;
        RECT 2152.440 37.750 2152.700 38.070 ;
        RECT 2869.120 37.750 2869.380 38.070 ;
        RECT 2869.180 2.400 2869.320 37.750 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2158.390 531.320 2158.710 531.380 ;
        RECT 2158.850 531.320 2159.170 531.380 ;
        RECT 2158.390 531.180 2159.170 531.320 ;
        RECT 2158.390 531.120 2158.710 531.180 ;
        RECT 2158.850 531.120 2159.170 531.180 ;
        RECT 2158.850 496.980 2159.170 497.040 ;
        RECT 2158.480 496.840 2159.170 496.980 ;
        RECT 2158.480 496.700 2158.620 496.840 ;
        RECT 2158.850 496.780 2159.170 496.840 ;
        RECT 2158.390 496.440 2158.710 496.700 ;
        RECT 2157.930 427.960 2158.250 428.020 ;
        RECT 2158.850 427.960 2159.170 428.020 ;
        RECT 2157.930 427.820 2159.170 427.960 ;
        RECT 2157.930 427.760 2158.250 427.820 ;
        RECT 2158.850 427.760 2159.170 427.820 ;
        RECT 2157.010 400.760 2157.330 400.820 ;
        RECT 2157.930 400.760 2158.250 400.820 ;
        RECT 2157.010 400.620 2158.250 400.760 ;
        RECT 2157.010 400.560 2157.330 400.620 ;
        RECT 2157.930 400.560 2158.250 400.620 ;
        RECT 2157.010 372.880 2157.330 372.940 ;
        RECT 2157.930 372.880 2158.250 372.940 ;
        RECT 2157.010 372.740 2158.250 372.880 ;
        RECT 2157.010 372.680 2157.330 372.740 ;
        RECT 2157.930 372.680 2158.250 372.740 ;
        RECT 2157.010 324.260 2157.330 324.320 ;
        RECT 2157.930 324.260 2158.250 324.320 ;
        RECT 2157.010 324.120 2158.250 324.260 ;
        RECT 2157.010 324.060 2157.330 324.120 ;
        RECT 2157.930 324.060 2158.250 324.120 ;
        RECT 2157.010 276.320 2157.330 276.380 ;
        RECT 2157.930 276.320 2158.250 276.380 ;
        RECT 2157.010 276.180 2158.250 276.320 ;
        RECT 2157.010 276.120 2157.330 276.180 ;
        RECT 2157.930 276.120 2158.250 276.180 ;
        RECT 2157.470 227.700 2157.790 227.760 ;
        RECT 2157.930 227.700 2158.250 227.760 ;
        RECT 2157.470 227.560 2158.250 227.700 ;
        RECT 2157.470 227.500 2157.790 227.560 ;
        RECT 2157.930 227.500 2158.250 227.560 ;
        RECT 2157.010 179.760 2157.330 179.820 ;
        RECT 2157.470 179.760 2157.790 179.820 ;
        RECT 2157.010 179.620 2157.790 179.760 ;
        RECT 2157.010 179.560 2157.330 179.620 ;
        RECT 2157.470 179.560 2157.790 179.620 ;
        RECT 2157.010 138.280 2157.330 138.340 ;
        RECT 2158.390 138.280 2158.710 138.340 ;
        RECT 2157.010 138.140 2158.710 138.280 ;
        RECT 2157.010 138.080 2157.330 138.140 ;
        RECT 2158.390 138.080 2158.710 138.140 ;
        RECT 2158.390 110.740 2158.710 110.800 ;
        RECT 2158.020 110.600 2158.710 110.740 ;
        RECT 2158.020 110.460 2158.160 110.600 ;
        RECT 2158.390 110.540 2158.710 110.600 ;
        RECT 2157.930 110.200 2158.250 110.460 ;
        RECT 2157.930 89.660 2158.250 89.720 ;
        RECT 2162.530 89.660 2162.850 89.720 ;
        RECT 2157.930 89.520 2162.850 89.660 ;
        RECT 2157.930 89.460 2158.250 89.520 ;
        RECT 2162.530 89.460 2162.850 89.520 ;
        RECT 2162.530 45.120 2162.850 45.180 ;
        RECT 2887.030 45.120 2887.350 45.180 ;
        RECT 2162.530 44.980 2887.350 45.120 ;
        RECT 2162.530 44.920 2162.850 44.980 ;
        RECT 2887.030 44.920 2887.350 44.980 ;
      LAYER via ;
        RECT 2158.420 531.120 2158.680 531.380 ;
        RECT 2158.880 531.120 2159.140 531.380 ;
        RECT 2158.880 496.780 2159.140 497.040 ;
        RECT 2158.420 496.440 2158.680 496.700 ;
        RECT 2157.960 427.760 2158.220 428.020 ;
        RECT 2158.880 427.760 2159.140 428.020 ;
        RECT 2157.040 400.560 2157.300 400.820 ;
        RECT 2157.960 400.560 2158.220 400.820 ;
        RECT 2157.040 372.680 2157.300 372.940 ;
        RECT 2157.960 372.680 2158.220 372.940 ;
        RECT 2157.040 324.060 2157.300 324.320 ;
        RECT 2157.960 324.060 2158.220 324.320 ;
        RECT 2157.040 276.120 2157.300 276.380 ;
        RECT 2157.960 276.120 2158.220 276.380 ;
        RECT 2157.500 227.500 2157.760 227.760 ;
        RECT 2157.960 227.500 2158.220 227.760 ;
        RECT 2157.040 179.560 2157.300 179.820 ;
        RECT 2157.500 179.560 2157.760 179.820 ;
        RECT 2157.040 138.080 2157.300 138.340 ;
        RECT 2158.420 138.080 2158.680 138.340 ;
        RECT 2158.420 110.540 2158.680 110.800 ;
        RECT 2157.960 110.200 2158.220 110.460 ;
        RECT 2157.960 89.460 2158.220 89.720 ;
        RECT 2162.560 89.460 2162.820 89.720 ;
        RECT 2162.560 44.920 2162.820 45.180 ;
        RECT 2887.060 44.920 2887.320 45.180 ;
      LAYER met2 ;
        RECT 2155.890 600.170 2156.170 604.000 ;
        RECT 2155.890 600.030 2158.620 600.170 ;
        RECT 2155.890 600.000 2156.170 600.030 ;
        RECT 2158.480 570.250 2158.620 600.030 ;
        RECT 2157.560 570.110 2158.620 570.250 ;
        RECT 2157.560 545.090 2157.700 570.110 ;
        RECT 2157.560 544.950 2158.620 545.090 ;
        RECT 2158.480 531.410 2158.620 544.950 ;
        RECT 2158.420 531.090 2158.680 531.410 ;
        RECT 2158.880 531.090 2159.140 531.410 ;
        RECT 2158.940 497.070 2159.080 531.090 ;
        RECT 2158.880 496.750 2159.140 497.070 ;
        RECT 2158.420 496.410 2158.680 496.730 ;
        RECT 2158.480 483.210 2158.620 496.410 ;
        RECT 2158.480 483.070 2159.080 483.210 ;
        RECT 2158.940 428.050 2159.080 483.070 ;
        RECT 2157.960 427.730 2158.220 428.050 ;
        RECT 2158.880 427.730 2159.140 428.050 ;
        RECT 2158.020 400.850 2158.160 427.730 ;
        RECT 2157.040 400.530 2157.300 400.850 ;
        RECT 2157.960 400.530 2158.220 400.850 ;
        RECT 2157.100 372.970 2157.240 400.530 ;
        RECT 2157.040 372.650 2157.300 372.970 ;
        RECT 2157.960 372.650 2158.220 372.970 ;
        RECT 2158.020 324.350 2158.160 372.650 ;
        RECT 2157.040 324.030 2157.300 324.350 ;
        RECT 2157.960 324.030 2158.220 324.350 ;
        RECT 2157.100 276.410 2157.240 324.030 ;
        RECT 2157.040 276.090 2157.300 276.410 ;
        RECT 2157.960 276.090 2158.220 276.410 ;
        RECT 2158.020 227.790 2158.160 276.090 ;
        RECT 2157.500 227.470 2157.760 227.790 ;
        RECT 2157.960 227.470 2158.220 227.790 ;
        RECT 2157.560 179.850 2157.700 227.470 ;
        RECT 2157.040 179.530 2157.300 179.850 ;
        RECT 2157.500 179.530 2157.760 179.850 ;
        RECT 2157.100 138.370 2157.240 179.530 ;
        RECT 2157.040 138.050 2157.300 138.370 ;
        RECT 2158.420 138.050 2158.680 138.370 ;
        RECT 2158.480 110.830 2158.620 138.050 ;
        RECT 2158.420 110.510 2158.680 110.830 ;
        RECT 2157.960 110.170 2158.220 110.490 ;
        RECT 2158.020 89.750 2158.160 110.170 ;
        RECT 2157.960 89.430 2158.220 89.750 ;
        RECT 2162.560 89.430 2162.820 89.750 ;
        RECT 2162.620 45.210 2162.760 89.430 ;
        RECT 2162.560 44.890 2162.820 45.210 ;
        RECT 2887.060 44.890 2887.320 45.210 ;
        RECT 2887.120 2.400 2887.260 44.890 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2165.750 44.780 2166.070 44.840 ;
        RECT 2904.970 44.780 2905.290 44.840 ;
        RECT 2165.750 44.640 2905.290 44.780 ;
        RECT 2165.750 44.580 2166.070 44.640 ;
        RECT 2904.970 44.580 2905.290 44.640 ;
      LAYER via ;
        RECT 2165.780 44.580 2166.040 44.840 ;
        RECT 2905.000 44.580 2905.260 44.840 ;
      LAYER met2 ;
        RECT 2165.090 600.170 2165.370 604.000 ;
        RECT 2165.090 600.030 2165.980 600.170 ;
        RECT 2165.090 600.000 2165.370 600.030 ;
        RECT 2165.840 44.870 2165.980 600.030 ;
        RECT 2165.780 44.550 2166.040 44.870 ;
        RECT 2905.000 44.550 2905.260 44.870 ;
        RECT 2905.060 2.400 2905.200 44.550 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1104.990 531.320 1105.310 531.380 ;
        RECT 1105.910 531.320 1106.230 531.380 ;
        RECT 1104.990 531.180 1106.230 531.320 ;
        RECT 1104.990 531.120 1105.310 531.180 ;
        RECT 1105.910 531.120 1106.230 531.180 ;
        RECT 1104.990 483.380 1105.310 483.440 ;
        RECT 1105.910 483.380 1106.230 483.440 ;
        RECT 1104.990 483.240 1106.230 483.380 ;
        RECT 1104.990 483.180 1105.310 483.240 ;
        RECT 1105.910 483.180 1106.230 483.240 ;
        RECT 1104.990 337.860 1105.310 337.920 ;
        RECT 1105.450 337.860 1105.770 337.920 ;
        RECT 1104.990 337.720 1105.770 337.860 ;
        RECT 1104.990 337.660 1105.310 337.720 ;
        RECT 1105.450 337.660 1105.770 337.720 ;
        RECT 1104.990 290.260 1105.310 290.320 ;
        RECT 1105.450 290.260 1105.770 290.320 ;
        RECT 1104.990 290.120 1105.770 290.260 ;
        RECT 1104.990 290.060 1105.310 290.120 ;
        RECT 1105.450 290.060 1105.770 290.120 ;
        RECT 1104.990 289.580 1105.310 289.640 ;
        RECT 1105.910 289.580 1106.230 289.640 ;
        RECT 1104.990 289.440 1106.230 289.580 ;
        RECT 1104.990 289.380 1105.310 289.440 ;
        RECT 1105.910 289.380 1106.230 289.440 ;
        RECT 1104.990 241.640 1105.310 241.700 ;
        RECT 1105.910 241.640 1106.230 241.700 ;
        RECT 1104.990 241.500 1106.230 241.640 ;
        RECT 1104.990 241.440 1105.310 241.500 ;
        RECT 1105.910 241.440 1106.230 241.500 ;
        RECT 1104.990 193.020 1105.310 193.080 ;
        RECT 1105.910 193.020 1106.230 193.080 ;
        RECT 1104.990 192.880 1106.230 193.020 ;
        RECT 1104.990 192.820 1105.310 192.880 ;
        RECT 1105.910 192.820 1106.230 192.880 ;
        RECT 1104.990 145.080 1105.310 145.140 ;
        RECT 1105.910 145.080 1106.230 145.140 ;
        RECT 1104.990 144.940 1106.230 145.080 ;
        RECT 1104.990 144.880 1105.310 144.940 ;
        RECT 1105.910 144.880 1106.230 144.940 ;
        RECT 1104.990 110.540 1105.310 110.800 ;
        RECT 1105.080 110.120 1105.220 110.540 ;
        RECT 1104.990 109.860 1105.310 110.120 ;
        RECT 852.910 26.760 853.230 26.820 ;
        RECT 1104.990 26.760 1105.310 26.820 ;
        RECT 852.910 26.620 1105.310 26.760 ;
        RECT 852.910 26.560 853.230 26.620 ;
        RECT 1104.990 26.560 1105.310 26.620 ;
      LAYER via ;
        RECT 1105.020 531.120 1105.280 531.380 ;
        RECT 1105.940 531.120 1106.200 531.380 ;
        RECT 1105.020 483.180 1105.280 483.440 ;
        RECT 1105.940 483.180 1106.200 483.440 ;
        RECT 1105.020 337.660 1105.280 337.920 ;
        RECT 1105.480 337.660 1105.740 337.920 ;
        RECT 1105.020 290.060 1105.280 290.320 ;
        RECT 1105.480 290.060 1105.740 290.320 ;
        RECT 1105.020 289.380 1105.280 289.640 ;
        RECT 1105.940 289.380 1106.200 289.640 ;
        RECT 1105.020 241.440 1105.280 241.700 ;
        RECT 1105.940 241.440 1106.200 241.700 ;
        RECT 1105.020 192.820 1105.280 193.080 ;
        RECT 1105.940 192.820 1106.200 193.080 ;
        RECT 1105.020 144.880 1105.280 145.140 ;
        RECT 1105.940 144.880 1106.200 145.140 ;
        RECT 1105.020 110.540 1105.280 110.800 ;
        RECT 1105.020 109.860 1105.280 110.120 ;
        RECT 852.940 26.560 853.200 26.820 ;
        RECT 1105.020 26.560 1105.280 26.820 ;
      LAYER met2 ;
        RECT 1108.930 600.170 1109.210 604.000 ;
        RECT 1107.380 600.030 1109.210 600.170 ;
        RECT 1107.380 579.885 1107.520 600.030 ;
        RECT 1108.930 600.000 1109.210 600.030 ;
        RECT 1105.010 579.515 1105.290 579.885 ;
        RECT 1107.310 579.515 1107.590 579.885 ;
        RECT 1105.080 531.410 1105.220 579.515 ;
        RECT 1105.020 531.090 1105.280 531.410 ;
        RECT 1105.940 531.090 1106.200 531.410 ;
        RECT 1106.000 483.470 1106.140 531.090 ;
        RECT 1105.020 483.150 1105.280 483.470 ;
        RECT 1105.940 483.150 1106.200 483.470 ;
        RECT 1105.080 337.950 1105.220 483.150 ;
        RECT 1105.020 337.630 1105.280 337.950 ;
        RECT 1105.480 337.630 1105.740 337.950 ;
        RECT 1105.540 290.350 1105.680 337.630 ;
        RECT 1105.020 290.030 1105.280 290.350 ;
        RECT 1105.480 290.030 1105.740 290.350 ;
        RECT 1105.080 289.670 1105.220 290.030 ;
        RECT 1105.020 289.350 1105.280 289.670 ;
        RECT 1105.940 289.350 1106.200 289.670 ;
        RECT 1106.000 241.730 1106.140 289.350 ;
        RECT 1105.020 241.410 1105.280 241.730 ;
        RECT 1105.940 241.410 1106.200 241.730 ;
        RECT 1105.080 193.110 1105.220 241.410 ;
        RECT 1105.020 192.790 1105.280 193.110 ;
        RECT 1105.940 192.790 1106.200 193.110 ;
        RECT 1106.000 145.170 1106.140 192.790 ;
        RECT 1105.020 144.850 1105.280 145.170 ;
        RECT 1105.940 144.850 1106.200 145.170 ;
        RECT 1105.080 110.830 1105.220 144.850 ;
        RECT 1105.020 110.510 1105.280 110.830 ;
        RECT 1105.020 109.830 1105.280 110.150 ;
        RECT 1105.080 26.850 1105.220 109.830 ;
        RECT 852.940 26.530 853.200 26.850 ;
        RECT 1105.020 26.530 1105.280 26.850 ;
        RECT 853.000 2.400 853.140 26.530 ;
        RECT 852.790 -4.800 853.350 2.400 ;
      LAYER via2 ;
        RECT 1105.010 579.560 1105.290 579.840 ;
        RECT 1107.310 579.560 1107.590 579.840 ;
      LAYER met3 ;
        RECT 1104.985 579.850 1105.315 579.865 ;
        RECT 1107.285 579.850 1107.615 579.865 ;
        RECT 1104.985 579.550 1107.615 579.850 ;
        RECT 1104.985 579.535 1105.315 579.550 ;
        RECT 1107.285 579.535 1107.615 579.550 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1097.170 592.520 1097.490 592.580 ;
        RECT 1118.330 592.520 1118.650 592.580 ;
        RECT 1097.170 592.380 1118.650 592.520 ;
        RECT 1097.170 592.320 1097.490 592.380 ;
        RECT 1118.330 592.320 1118.650 592.380 ;
        RECT 927.890 588.780 928.210 588.840 ;
        RECT 1097.170 588.780 1097.490 588.840 ;
        RECT 927.890 588.640 1097.490 588.780 ;
        RECT 927.890 588.580 928.210 588.640 ;
        RECT 1097.170 588.580 1097.490 588.640 ;
        RECT 870.850 20.300 871.170 20.360 ;
        RECT 927.890 20.300 928.210 20.360 ;
        RECT 870.850 20.160 928.210 20.300 ;
        RECT 870.850 20.100 871.170 20.160 ;
        RECT 927.890 20.100 928.210 20.160 ;
      LAYER via ;
        RECT 1097.200 592.320 1097.460 592.580 ;
        RECT 1118.360 592.320 1118.620 592.580 ;
        RECT 927.920 588.580 928.180 588.840 ;
        RECT 1097.200 588.580 1097.460 588.840 ;
        RECT 870.880 20.100 871.140 20.360 ;
        RECT 927.920 20.100 928.180 20.360 ;
      LAYER met2 ;
        RECT 1118.130 600.000 1118.410 604.000 ;
        RECT 1118.190 598.810 1118.330 600.000 ;
        RECT 1118.190 598.670 1118.560 598.810 ;
        RECT 1118.420 592.610 1118.560 598.670 ;
        RECT 1097.200 592.290 1097.460 592.610 ;
        RECT 1118.360 592.290 1118.620 592.610 ;
        RECT 1097.260 588.870 1097.400 592.290 ;
        RECT 927.920 588.550 928.180 588.870 ;
        RECT 1097.200 588.550 1097.460 588.870 ;
        RECT 927.980 20.390 928.120 588.550 ;
        RECT 870.880 20.070 871.140 20.390 ;
        RECT 927.920 20.070 928.180 20.390 ;
        RECT 870.940 2.400 871.080 20.070 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 928.350 589.460 928.670 589.520 ;
        RECT 1125.690 589.460 1126.010 589.520 ;
        RECT 928.350 589.320 1126.010 589.460 ;
        RECT 928.350 589.260 928.670 589.320 ;
        RECT 1125.690 589.260 1126.010 589.320 ;
        RECT 888.790 20.640 889.110 20.700 ;
        RECT 928.350 20.640 928.670 20.700 ;
        RECT 888.790 20.500 928.670 20.640 ;
        RECT 888.790 20.440 889.110 20.500 ;
        RECT 928.350 20.440 928.670 20.500 ;
      LAYER via ;
        RECT 928.380 589.260 928.640 589.520 ;
        RECT 1125.720 589.260 1125.980 589.520 ;
        RECT 888.820 20.440 889.080 20.700 ;
        RECT 928.380 20.440 928.640 20.700 ;
      LAYER met2 ;
        RECT 1127.330 600.170 1127.610 604.000 ;
        RECT 1125.780 600.030 1127.610 600.170 ;
        RECT 1125.780 589.550 1125.920 600.030 ;
        RECT 1127.330 600.000 1127.610 600.030 ;
        RECT 928.380 589.230 928.640 589.550 ;
        RECT 1125.720 589.230 1125.980 589.550 ;
        RECT 928.440 20.730 928.580 589.230 ;
        RECT 888.820 20.410 889.080 20.730 ;
        RECT 928.380 20.410 928.640 20.730 ;
        RECT 888.880 2.400 889.020 20.410 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1072.790 586.740 1073.110 586.800 ;
        RECT 1134.890 586.740 1135.210 586.800 ;
        RECT 1072.790 586.600 1135.210 586.740 ;
        RECT 1072.790 586.540 1073.110 586.600 ;
        RECT 1134.890 586.540 1135.210 586.600 ;
        RECT 1036.450 17.240 1036.770 17.300 ;
        RECT 1072.790 17.240 1073.110 17.300 ;
        RECT 1036.450 17.100 1073.110 17.240 ;
        RECT 1036.450 17.040 1036.770 17.100 ;
        RECT 1072.790 17.040 1073.110 17.100 ;
        RECT 906.730 16.220 907.050 16.280 ;
        RECT 989.530 16.220 989.850 16.280 ;
        RECT 906.730 16.080 989.850 16.220 ;
        RECT 906.730 16.020 907.050 16.080 ;
        RECT 989.530 16.020 989.850 16.080 ;
        RECT 1027.710 16.220 1028.030 16.280 ;
        RECT 1036.450 16.220 1036.770 16.280 ;
        RECT 1027.710 16.080 1036.770 16.220 ;
        RECT 1027.710 16.020 1028.030 16.080 ;
        RECT 1036.450 16.020 1036.770 16.080 ;
        RECT 1013.910 14.520 1014.230 14.580 ;
        RECT 1027.710 14.520 1028.030 14.580 ;
        RECT 1013.910 14.380 1028.030 14.520 ;
        RECT 1013.910 14.320 1014.230 14.380 ;
        RECT 1027.710 14.320 1028.030 14.380 ;
        RECT 989.530 13.500 989.850 13.560 ;
        RECT 1013.910 13.500 1014.230 13.560 ;
        RECT 989.530 13.360 1014.230 13.500 ;
        RECT 989.530 13.300 989.850 13.360 ;
        RECT 1013.910 13.300 1014.230 13.360 ;
      LAYER via ;
        RECT 1072.820 586.540 1073.080 586.800 ;
        RECT 1134.920 586.540 1135.180 586.800 ;
        RECT 1036.480 17.040 1036.740 17.300 ;
        RECT 1072.820 17.040 1073.080 17.300 ;
        RECT 906.760 16.020 907.020 16.280 ;
        RECT 989.560 16.020 989.820 16.280 ;
        RECT 1027.740 16.020 1028.000 16.280 ;
        RECT 1036.480 16.020 1036.740 16.280 ;
        RECT 1013.940 14.320 1014.200 14.580 ;
        RECT 1027.740 14.320 1028.000 14.580 ;
        RECT 989.560 13.300 989.820 13.560 ;
        RECT 1013.940 13.300 1014.200 13.560 ;
      LAYER met2 ;
        RECT 1136.530 600.170 1136.810 604.000 ;
        RECT 1134.980 600.030 1136.810 600.170 ;
        RECT 1134.980 586.830 1135.120 600.030 ;
        RECT 1136.530 600.000 1136.810 600.030 ;
        RECT 1072.820 586.510 1073.080 586.830 ;
        RECT 1134.920 586.510 1135.180 586.830 ;
        RECT 1072.880 17.330 1073.020 586.510 ;
        RECT 1036.480 17.010 1036.740 17.330 ;
        RECT 1072.820 17.010 1073.080 17.330 ;
        RECT 1036.540 16.310 1036.680 17.010 ;
        RECT 906.760 15.990 907.020 16.310 ;
        RECT 989.560 15.990 989.820 16.310 ;
        RECT 1027.740 15.990 1028.000 16.310 ;
        RECT 1036.480 15.990 1036.740 16.310 ;
        RECT 906.820 2.400 906.960 15.990 ;
        RECT 989.620 13.590 989.760 15.990 ;
        RECT 1027.800 14.610 1027.940 15.990 ;
        RECT 1013.940 14.290 1014.200 14.610 ;
        RECT 1027.740 14.290 1028.000 14.610 ;
        RECT 1014.000 13.590 1014.140 14.290 ;
        RECT 989.560 13.270 989.820 13.590 ;
        RECT 1013.940 13.270 1014.200 13.590 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.930 588.780 1146.250 588.840 ;
        RECT 1100.020 588.640 1146.250 588.780 ;
        RECT 1100.020 588.100 1100.160 588.640 ;
        RECT 1145.930 588.580 1146.250 588.640 ;
        RECT 1002.500 587.960 1100.160 588.100 ;
        RECT 969.290 587.760 969.610 587.820 ;
        RECT 1002.500 587.760 1002.640 587.960 ;
        RECT 969.290 587.620 1002.640 587.760 ;
        RECT 969.290 587.560 969.610 587.620 ;
        RECT 924.210 15.880 924.530 15.940 ;
        RECT 924.210 15.740 950.660 15.880 ;
        RECT 924.210 15.680 924.530 15.740 ;
        RECT 950.520 15.540 950.660 15.740 ;
        RECT 969.290 15.540 969.610 15.600 ;
        RECT 950.520 15.400 969.610 15.540 ;
        RECT 969.290 15.340 969.610 15.400 ;
      LAYER via ;
        RECT 1145.960 588.580 1146.220 588.840 ;
        RECT 969.320 587.560 969.580 587.820 ;
        RECT 924.240 15.680 924.500 15.940 ;
        RECT 969.320 15.340 969.580 15.600 ;
      LAYER met2 ;
        RECT 1145.730 600.000 1146.010 604.000 ;
        RECT 1145.790 598.810 1145.930 600.000 ;
        RECT 1145.790 598.670 1146.160 598.810 ;
        RECT 1146.020 588.870 1146.160 598.670 ;
        RECT 1145.960 588.550 1146.220 588.870 ;
        RECT 969.320 587.530 969.580 587.850 ;
        RECT 924.240 15.650 924.500 15.970 ;
        RECT 924.300 2.400 924.440 15.650 ;
        RECT 969.380 15.630 969.520 587.530 ;
        RECT 969.320 15.310 969.580 15.630 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 942.150 20.300 942.470 20.360 ;
        RECT 1152.830 20.300 1153.150 20.360 ;
        RECT 942.150 20.160 1153.150 20.300 ;
        RECT 942.150 20.100 942.470 20.160 ;
        RECT 1152.830 20.100 1153.150 20.160 ;
      LAYER via ;
        RECT 942.180 20.100 942.440 20.360 ;
        RECT 1152.860 20.100 1153.120 20.360 ;
      LAYER met2 ;
        RECT 1154.930 600.170 1155.210 604.000 ;
        RECT 1152.920 600.030 1155.210 600.170 ;
        RECT 1152.920 20.390 1153.060 600.030 ;
        RECT 1154.930 600.000 1155.210 600.030 ;
        RECT 942.180 20.070 942.440 20.390 ;
        RECT 1152.860 20.070 1153.120 20.390 ;
        RECT 942.240 2.400 942.380 20.070 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1161.110 572.800 1161.430 572.860 ;
        RECT 1162.950 572.800 1163.270 572.860 ;
        RECT 1161.110 572.660 1163.270 572.800 ;
        RECT 1161.110 572.600 1161.430 572.660 ;
        RECT 1162.950 572.600 1163.270 572.660 ;
        RECT 1161.110 497.320 1161.430 497.380 ;
        RECT 1160.740 497.180 1161.430 497.320 ;
        RECT 1160.740 497.040 1160.880 497.180 ;
        RECT 1161.110 497.120 1161.430 497.180 ;
        RECT 1160.650 496.780 1160.970 497.040 ;
        RECT 1160.650 420.820 1160.970 420.880 ;
        RECT 1161.570 420.820 1161.890 420.880 ;
        RECT 1160.650 420.680 1161.890 420.820 ;
        RECT 1160.650 420.620 1160.970 420.680 ;
        RECT 1161.570 420.620 1161.890 420.680 ;
        RECT 1160.650 396.680 1160.970 396.740 ;
        RECT 1161.570 396.680 1161.890 396.740 ;
        RECT 1160.650 396.540 1161.890 396.680 ;
        RECT 1160.650 396.480 1160.970 396.540 ;
        RECT 1161.570 396.480 1161.890 396.540 ;
        RECT 990.450 16.560 990.770 16.620 ;
        RECT 1160.650 16.560 1160.970 16.620 ;
        RECT 990.450 16.420 1160.970 16.560 ;
        RECT 990.450 16.360 990.770 16.420 ;
        RECT 1160.650 16.360 1160.970 16.420 ;
        RECT 960.090 15.200 960.410 15.260 ;
        RECT 990.450 15.200 990.770 15.260 ;
        RECT 960.090 15.060 990.770 15.200 ;
        RECT 960.090 15.000 960.410 15.060 ;
        RECT 990.450 15.000 990.770 15.060 ;
      LAYER via ;
        RECT 1161.140 572.600 1161.400 572.860 ;
        RECT 1162.980 572.600 1163.240 572.860 ;
        RECT 1161.140 497.120 1161.400 497.380 ;
        RECT 1160.680 496.780 1160.940 497.040 ;
        RECT 1160.680 420.620 1160.940 420.880 ;
        RECT 1161.600 420.620 1161.860 420.880 ;
        RECT 1160.680 396.480 1160.940 396.740 ;
        RECT 1161.600 396.480 1161.860 396.740 ;
        RECT 990.480 16.360 990.740 16.620 ;
        RECT 1160.680 16.360 1160.940 16.620 ;
        RECT 960.120 15.000 960.380 15.260 ;
        RECT 990.480 15.000 990.740 15.260 ;
      LAYER met2 ;
        RECT 1164.130 600.170 1164.410 604.000 ;
        RECT 1163.040 600.030 1164.410 600.170 ;
        RECT 1163.040 572.890 1163.180 600.030 ;
        RECT 1164.130 600.000 1164.410 600.030 ;
        RECT 1161.140 572.570 1161.400 572.890 ;
        RECT 1162.980 572.570 1163.240 572.890 ;
        RECT 1161.200 497.410 1161.340 572.570 ;
        RECT 1161.140 497.090 1161.400 497.410 ;
        RECT 1160.680 496.750 1160.940 497.070 ;
        RECT 1160.740 420.910 1160.880 496.750 ;
        RECT 1160.680 420.590 1160.940 420.910 ;
        RECT 1161.600 420.590 1161.860 420.910 ;
        RECT 1161.660 396.770 1161.800 420.590 ;
        RECT 1160.680 396.450 1160.940 396.770 ;
        RECT 1161.600 396.450 1161.860 396.770 ;
        RECT 1160.740 303.690 1160.880 396.450 ;
        RECT 1160.280 303.550 1160.880 303.690 ;
        RECT 1160.280 303.010 1160.420 303.550 ;
        RECT 1160.280 302.870 1160.880 303.010 ;
        RECT 1160.740 207.130 1160.880 302.870 ;
        RECT 1160.280 206.990 1160.880 207.130 ;
        RECT 1160.280 206.450 1160.420 206.990 ;
        RECT 1160.280 206.310 1160.880 206.450 ;
        RECT 1160.740 110.570 1160.880 206.310 ;
        RECT 1160.280 110.430 1160.880 110.570 ;
        RECT 1160.280 109.890 1160.420 110.430 ;
        RECT 1160.280 109.750 1160.880 109.890 ;
        RECT 1160.740 16.650 1160.880 109.750 ;
        RECT 990.480 16.330 990.740 16.650 ;
        RECT 1160.680 16.330 1160.940 16.650 ;
        RECT 990.540 15.290 990.680 16.330 ;
        RECT 960.120 14.970 960.380 15.290 ;
        RECT 990.480 14.970 990.740 15.290 ;
        RECT 960.180 2.400 960.320 14.970 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1001.950 589.120 1002.270 589.180 ;
        RECT 1173.530 589.120 1173.850 589.180 ;
        RECT 1001.950 588.980 1173.850 589.120 ;
        RECT 1001.950 588.920 1002.270 588.980 ;
        RECT 1173.530 588.920 1173.850 588.980 ;
        RECT 979.410 588.100 979.730 588.160 ;
        RECT 1001.950 588.100 1002.270 588.160 ;
        RECT 979.410 587.960 1002.270 588.100 ;
        RECT 979.410 587.900 979.730 587.960 ;
        RECT 1001.950 587.900 1002.270 587.960 ;
      LAYER via ;
        RECT 1001.980 588.920 1002.240 589.180 ;
        RECT 1173.560 588.920 1173.820 589.180 ;
        RECT 979.440 587.900 979.700 588.160 ;
        RECT 1001.980 587.900 1002.240 588.160 ;
      LAYER met2 ;
        RECT 1173.330 600.000 1173.610 604.000 ;
        RECT 1173.390 598.810 1173.530 600.000 ;
        RECT 1173.390 598.670 1173.760 598.810 ;
        RECT 1173.620 589.210 1173.760 598.670 ;
        RECT 1001.980 588.890 1002.240 589.210 ;
        RECT 1173.560 588.890 1173.820 589.210 ;
        RECT 1002.040 588.190 1002.180 588.890 ;
        RECT 979.440 587.870 979.700 588.190 ;
        RECT 1001.980 587.870 1002.240 588.190 ;
        RECT 979.500 3.130 979.640 587.870 ;
        RECT 978.120 2.990 979.640 3.130 ;
        RECT 978.120 2.400 978.260 2.990 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 35.940 657.270 36.000 ;
        RECT 1007.930 35.940 1008.250 36.000 ;
        RECT 656.950 35.800 1008.250 35.940 ;
        RECT 656.950 35.740 657.270 35.800 ;
        RECT 1007.930 35.740 1008.250 35.800 ;
      LAYER via ;
        RECT 656.980 35.740 657.240 36.000 ;
        RECT 1007.960 35.740 1008.220 36.000 ;
      LAYER met2 ;
        RECT 1008.190 600.000 1008.470 604.000 ;
        RECT 1008.250 598.810 1008.390 600.000 ;
        RECT 1008.020 598.670 1008.390 598.810 ;
        RECT 1008.020 36.030 1008.160 598.670 ;
        RECT 656.980 35.710 657.240 36.030 ;
        RECT 1007.960 35.710 1008.220 36.030 ;
        RECT 657.040 2.400 657.180 35.710 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1127.990 589.460 1128.310 589.520 ;
        RECT 1180.890 589.460 1181.210 589.520 ;
        RECT 1127.990 589.320 1181.210 589.460 ;
        RECT 1127.990 589.260 1128.310 589.320 ;
        RECT 1180.890 589.260 1181.210 589.320 ;
        RECT 995.970 15.200 996.290 15.260 ;
        RECT 1127.990 15.200 1128.310 15.260 ;
        RECT 995.970 15.060 1128.310 15.200 ;
        RECT 995.970 15.000 996.290 15.060 ;
        RECT 1127.990 15.000 1128.310 15.060 ;
      LAYER via ;
        RECT 1128.020 589.260 1128.280 589.520 ;
        RECT 1180.920 589.260 1181.180 589.520 ;
        RECT 996.000 15.000 996.260 15.260 ;
        RECT 1128.020 15.000 1128.280 15.260 ;
      LAYER met2 ;
        RECT 1182.530 600.170 1182.810 604.000 ;
        RECT 1180.980 600.030 1182.810 600.170 ;
        RECT 1180.980 589.550 1181.120 600.030 ;
        RECT 1182.530 600.000 1182.810 600.030 ;
        RECT 1128.020 589.230 1128.280 589.550 ;
        RECT 1180.920 589.230 1181.180 589.550 ;
        RECT 1128.080 15.290 1128.220 589.230 ;
        RECT 996.000 14.970 996.260 15.290 ;
        RECT 1128.020 14.970 1128.280 15.290 ;
        RECT 996.060 2.400 996.200 14.970 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1155.590 591.160 1155.910 591.220 ;
        RECT 1190.090 591.160 1190.410 591.220 ;
        RECT 1155.590 591.020 1190.410 591.160 ;
        RECT 1155.590 590.960 1155.910 591.020 ;
        RECT 1190.090 590.960 1190.410 591.020 ;
        RECT 1013.450 15.540 1013.770 15.600 ;
        RECT 1155.590 15.540 1155.910 15.600 ;
        RECT 1013.450 15.400 1155.910 15.540 ;
        RECT 1013.450 15.340 1013.770 15.400 ;
        RECT 1155.590 15.340 1155.910 15.400 ;
      LAYER via ;
        RECT 1155.620 590.960 1155.880 591.220 ;
        RECT 1190.120 590.960 1190.380 591.220 ;
        RECT 1013.480 15.340 1013.740 15.600 ;
        RECT 1155.620 15.340 1155.880 15.600 ;
      LAYER met2 ;
        RECT 1191.730 600.170 1192.010 604.000 ;
        RECT 1190.180 600.030 1192.010 600.170 ;
        RECT 1190.180 591.250 1190.320 600.030 ;
        RECT 1191.730 600.000 1192.010 600.030 ;
        RECT 1155.620 590.930 1155.880 591.250 ;
        RECT 1190.120 590.930 1190.380 591.250 ;
        RECT 1155.680 15.630 1155.820 590.930 ;
        RECT 1013.480 15.310 1013.740 15.630 ;
        RECT 1155.620 15.310 1155.880 15.630 ;
        RECT 1013.540 2.400 1013.680 15.310 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1162.490 592.520 1162.810 592.580 ;
        RECT 1201.130 592.520 1201.450 592.580 ;
        RECT 1162.490 592.380 1201.450 592.520 ;
        RECT 1162.490 592.320 1162.810 592.380 ;
        RECT 1201.130 592.320 1201.450 592.380 ;
        RECT 1031.390 14.860 1031.710 14.920 ;
        RECT 1162.030 14.860 1162.350 14.920 ;
        RECT 1031.390 14.720 1162.350 14.860 ;
        RECT 1031.390 14.660 1031.710 14.720 ;
        RECT 1162.030 14.660 1162.350 14.720 ;
      LAYER via ;
        RECT 1162.520 592.320 1162.780 592.580 ;
        RECT 1201.160 592.320 1201.420 592.580 ;
        RECT 1031.420 14.660 1031.680 14.920 ;
        RECT 1162.060 14.660 1162.320 14.920 ;
      LAYER met2 ;
        RECT 1200.930 600.000 1201.210 604.000 ;
        RECT 1200.990 598.810 1201.130 600.000 ;
        RECT 1200.990 598.670 1201.360 598.810 ;
        RECT 1201.220 592.610 1201.360 598.670 ;
        RECT 1162.520 592.290 1162.780 592.610 ;
        RECT 1201.160 592.290 1201.420 592.610 ;
        RECT 1162.580 21.490 1162.720 592.290 ;
        RECT 1162.120 21.350 1162.720 21.490 ;
        RECT 1162.120 14.950 1162.260 21.350 ;
        RECT 1031.420 14.630 1031.680 14.950 ;
        RECT 1162.060 14.630 1162.320 14.950 ;
        RECT 1031.480 2.400 1031.620 14.630 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1182.730 592.860 1183.050 592.920 ;
        RECT 1208.490 592.860 1208.810 592.920 ;
        RECT 1182.730 592.720 1208.810 592.860 ;
        RECT 1182.730 592.660 1183.050 592.720 ;
        RECT 1208.490 592.660 1208.810 592.720 ;
        RECT 1118.790 592.520 1119.110 592.580 ;
        RECT 1149.150 592.520 1149.470 592.580 ;
        RECT 1118.790 592.380 1149.470 592.520 ;
        RECT 1118.790 592.320 1119.110 592.380 ;
        RECT 1149.150 592.320 1149.470 592.380 ;
        RECT 1055.310 587.080 1055.630 587.140 ;
        RECT 1118.790 587.080 1119.110 587.140 ;
        RECT 1055.310 586.940 1119.110 587.080 ;
        RECT 1055.310 586.880 1055.630 586.940 ;
        RECT 1118.790 586.880 1119.110 586.940 ;
        RECT 1149.150 587.080 1149.470 587.140 ;
        RECT 1182.730 587.080 1183.050 587.140 ;
        RECT 1149.150 586.940 1183.050 587.080 ;
        RECT 1149.150 586.880 1149.470 586.940 ;
        RECT 1182.730 586.880 1183.050 586.940 ;
        RECT 1049.330 18.600 1049.650 18.660 ;
        RECT 1055.310 18.600 1055.630 18.660 ;
        RECT 1049.330 18.460 1055.630 18.600 ;
        RECT 1049.330 18.400 1049.650 18.460 ;
        RECT 1055.310 18.400 1055.630 18.460 ;
      LAYER via ;
        RECT 1182.760 592.660 1183.020 592.920 ;
        RECT 1208.520 592.660 1208.780 592.920 ;
        RECT 1118.820 592.320 1119.080 592.580 ;
        RECT 1149.180 592.320 1149.440 592.580 ;
        RECT 1055.340 586.880 1055.600 587.140 ;
        RECT 1118.820 586.880 1119.080 587.140 ;
        RECT 1149.180 586.880 1149.440 587.140 ;
        RECT 1182.760 586.880 1183.020 587.140 ;
        RECT 1049.360 18.400 1049.620 18.660 ;
        RECT 1055.340 18.400 1055.600 18.660 ;
      LAYER met2 ;
        RECT 1210.130 600.170 1210.410 604.000 ;
        RECT 1208.580 600.030 1210.410 600.170 ;
        RECT 1208.580 592.950 1208.720 600.030 ;
        RECT 1210.130 600.000 1210.410 600.030 ;
        RECT 1182.760 592.630 1183.020 592.950 ;
        RECT 1208.520 592.630 1208.780 592.950 ;
        RECT 1118.820 592.290 1119.080 592.610 ;
        RECT 1149.180 592.290 1149.440 592.610 ;
        RECT 1118.880 587.170 1119.020 592.290 ;
        RECT 1149.240 587.170 1149.380 592.290 ;
        RECT 1182.820 587.170 1182.960 592.630 ;
        RECT 1055.340 586.850 1055.600 587.170 ;
        RECT 1118.820 586.850 1119.080 587.170 ;
        RECT 1149.180 586.850 1149.440 587.170 ;
        RECT 1182.760 586.850 1183.020 587.170 ;
        RECT 1055.400 18.690 1055.540 586.850 ;
        RECT 1049.360 18.370 1049.620 18.690 ;
        RECT 1055.340 18.370 1055.600 18.690 ;
        RECT 1049.420 2.400 1049.560 18.370 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 593.200 1069.430 593.260 ;
        RECT 1217.690 593.200 1218.010 593.260 ;
        RECT 1069.110 593.060 1218.010 593.200 ;
        RECT 1069.110 593.000 1069.430 593.060 ;
        RECT 1217.690 593.000 1218.010 593.060 ;
      LAYER via ;
        RECT 1069.140 593.000 1069.400 593.260 ;
        RECT 1217.720 593.000 1217.980 593.260 ;
      LAYER met2 ;
        RECT 1219.330 600.170 1219.610 604.000 ;
        RECT 1217.780 600.030 1219.610 600.170 ;
        RECT 1217.780 593.290 1217.920 600.030 ;
        RECT 1219.330 600.000 1219.610 600.030 ;
        RECT 1069.140 592.970 1069.400 593.290 ;
        RECT 1217.720 592.970 1217.980 593.290 ;
        RECT 1069.200 3.130 1069.340 592.970 ;
        RECT 1067.360 2.990 1069.340 3.130 ;
        RECT 1067.360 2.400 1067.500 2.990 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1085.210 17.240 1085.530 17.300 ;
        RECT 1172.610 17.240 1172.930 17.300 ;
        RECT 1085.210 17.100 1172.930 17.240 ;
        RECT 1085.210 17.040 1085.530 17.100 ;
        RECT 1172.610 17.040 1172.930 17.100 ;
        RECT 1173.530 17.240 1173.850 17.300 ;
        RECT 1218.150 17.240 1218.470 17.300 ;
        RECT 1173.530 17.100 1218.470 17.240 ;
        RECT 1173.530 17.040 1173.850 17.100 ;
        RECT 1218.150 17.040 1218.470 17.100 ;
      LAYER via ;
        RECT 1085.240 17.040 1085.500 17.300 ;
        RECT 1172.640 17.040 1172.900 17.300 ;
        RECT 1173.560 17.040 1173.820 17.300 ;
        RECT 1218.180 17.040 1218.440 17.300 ;
      LAYER met2 ;
        RECT 1228.530 600.000 1228.810 604.000 ;
        RECT 1228.590 598.810 1228.730 600.000 ;
        RECT 1228.590 598.670 1228.960 598.810 ;
        RECT 1228.820 586.685 1228.960 598.670 ;
        RECT 1218.170 586.315 1218.450 586.685 ;
        RECT 1228.750 586.315 1229.030 586.685 ;
        RECT 1172.700 17.330 1173.760 17.410 ;
        RECT 1218.240 17.330 1218.380 586.315 ;
        RECT 1085.240 17.010 1085.500 17.330 ;
        RECT 1172.640 17.270 1173.820 17.330 ;
        RECT 1172.640 17.010 1172.900 17.270 ;
        RECT 1173.560 17.010 1173.820 17.270 ;
        RECT 1218.180 17.010 1218.440 17.330 ;
        RECT 1085.300 2.400 1085.440 17.010 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
      LAYER via2 ;
        RECT 1218.170 586.360 1218.450 586.640 ;
        RECT 1228.750 586.360 1229.030 586.640 ;
      LAYER met3 ;
        RECT 1218.145 586.650 1218.475 586.665 ;
        RECT 1228.725 586.650 1229.055 586.665 ;
        RECT 1218.145 586.350 1229.055 586.650 ;
        RECT 1218.145 586.335 1218.475 586.350 ;
        RECT 1228.725 586.335 1229.055 586.350 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1190.090 587.420 1190.410 587.480 ;
        RECT 1190.090 587.280 1227.580 587.420 ;
        RECT 1190.090 587.220 1190.410 587.280 ;
        RECT 1227.440 587.080 1227.580 587.280 ;
        RECT 1236.090 587.080 1236.410 587.140 ;
        RECT 1227.440 586.940 1236.410 587.080 ;
        RECT 1236.090 586.880 1236.410 586.940 ;
        RECT 1102.690 16.220 1103.010 16.280 ;
        RECT 1190.090 16.220 1190.410 16.280 ;
        RECT 1102.690 16.080 1190.410 16.220 ;
        RECT 1102.690 16.020 1103.010 16.080 ;
        RECT 1190.090 16.020 1190.410 16.080 ;
      LAYER via ;
        RECT 1190.120 587.220 1190.380 587.480 ;
        RECT 1236.120 586.880 1236.380 587.140 ;
        RECT 1102.720 16.020 1102.980 16.280 ;
        RECT 1190.120 16.020 1190.380 16.280 ;
      LAYER met2 ;
        RECT 1237.730 600.170 1238.010 604.000 ;
        RECT 1236.180 600.030 1238.010 600.170 ;
        RECT 1190.120 587.190 1190.380 587.510 ;
        RECT 1190.180 16.310 1190.320 587.190 ;
        RECT 1236.180 587.170 1236.320 600.030 ;
        RECT 1237.730 600.000 1238.010 600.030 ;
        RECT 1236.120 586.850 1236.380 587.170 ;
        RECT 1102.720 15.990 1102.980 16.310 ;
        RECT 1190.120 15.990 1190.380 16.310 ;
        RECT 1102.780 2.400 1102.920 15.990 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1242.530 496.780 1242.850 497.040 ;
        RECT 1242.070 496.640 1242.390 496.700 ;
        RECT 1242.620 496.640 1242.760 496.780 ;
        RECT 1242.070 496.500 1242.760 496.640 ;
        RECT 1242.070 496.440 1242.390 496.500 ;
        RECT 1242.990 434.900 1243.310 435.160 ;
        RECT 1243.080 434.420 1243.220 434.900 ;
        RECT 1243.450 434.420 1243.770 434.480 ;
        RECT 1243.080 434.280 1243.770 434.420 ;
        RECT 1243.450 434.220 1243.770 434.280 ;
        RECT 1242.530 420.820 1242.850 420.880 ;
        RECT 1243.450 420.820 1243.770 420.880 ;
        RECT 1242.530 420.680 1243.770 420.820 ;
        RECT 1242.530 420.620 1242.850 420.680 ;
        RECT 1243.450 420.620 1243.770 420.680 ;
        RECT 1242.530 372.880 1242.850 372.940 ;
        RECT 1243.910 372.880 1244.230 372.940 ;
        RECT 1242.530 372.740 1244.230 372.880 ;
        RECT 1242.530 372.680 1242.850 372.740 ;
        RECT 1243.910 372.680 1244.230 372.740 ;
        RECT 1242.530 331.400 1242.850 331.460 ;
        RECT 1243.910 331.400 1244.230 331.460 ;
        RECT 1242.530 331.260 1244.230 331.400 ;
        RECT 1242.530 331.200 1242.850 331.260 ;
        RECT 1243.910 331.200 1244.230 331.260 ;
        RECT 1242.070 303.520 1242.390 303.580 ;
        RECT 1242.990 303.520 1243.310 303.580 ;
        RECT 1242.070 303.380 1243.310 303.520 ;
        RECT 1242.070 303.320 1242.390 303.380 ;
        RECT 1242.990 303.320 1243.310 303.380 ;
        RECT 1242.990 217.500 1243.310 217.560 ;
        RECT 1243.910 217.500 1244.230 217.560 ;
        RECT 1242.990 217.360 1244.230 217.500 ;
        RECT 1242.990 217.300 1243.310 217.360 ;
        RECT 1243.910 217.300 1244.230 217.360 ;
        RECT 1243.450 193.360 1243.770 193.420 ;
        RECT 1243.910 193.360 1244.230 193.420 ;
        RECT 1243.450 193.220 1244.230 193.360 ;
        RECT 1243.450 193.160 1243.770 193.220 ;
        RECT 1243.910 193.160 1244.230 193.220 ;
        RECT 1242.530 145.080 1242.850 145.140 ;
        RECT 1243.450 145.080 1243.770 145.140 ;
        RECT 1242.530 144.940 1243.770 145.080 ;
        RECT 1242.530 144.880 1242.850 144.940 ;
        RECT 1243.450 144.880 1243.770 144.940 ;
        RECT 1242.070 110.400 1242.390 110.460 ;
        RECT 1242.990 110.400 1243.310 110.460 ;
        RECT 1242.070 110.260 1243.310 110.400 ;
        RECT 1242.070 110.200 1242.390 110.260 ;
        RECT 1242.990 110.200 1243.310 110.260 ;
        RECT 1120.630 18.260 1120.950 18.320 ;
        RECT 1144.090 18.260 1144.410 18.320 ;
        RECT 1120.630 18.120 1144.410 18.260 ;
        RECT 1120.630 18.060 1120.950 18.120 ;
        RECT 1144.090 18.060 1144.410 18.120 ;
        RECT 1242.990 17.920 1243.310 17.980 ;
        RECT 1173.160 17.780 1243.310 17.920 ;
        RECT 1144.090 16.900 1144.410 16.960 ;
        RECT 1144.090 16.760 1172.840 16.900 ;
        RECT 1144.090 16.700 1144.410 16.760 ;
        RECT 1172.700 16.560 1172.840 16.760 ;
        RECT 1173.160 16.560 1173.300 17.780 ;
        RECT 1242.990 17.720 1243.310 17.780 ;
        RECT 1172.700 16.420 1173.300 16.560 ;
      LAYER via ;
        RECT 1242.560 496.780 1242.820 497.040 ;
        RECT 1242.100 496.440 1242.360 496.700 ;
        RECT 1243.020 434.900 1243.280 435.160 ;
        RECT 1243.480 434.220 1243.740 434.480 ;
        RECT 1242.560 420.620 1242.820 420.880 ;
        RECT 1243.480 420.620 1243.740 420.880 ;
        RECT 1242.560 372.680 1242.820 372.940 ;
        RECT 1243.940 372.680 1244.200 372.940 ;
        RECT 1242.560 331.200 1242.820 331.460 ;
        RECT 1243.940 331.200 1244.200 331.460 ;
        RECT 1242.100 303.320 1242.360 303.580 ;
        RECT 1243.020 303.320 1243.280 303.580 ;
        RECT 1243.020 217.300 1243.280 217.560 ;
        RECT 1243.940 217.300 1244.200 217.560 ;
        RECT 1243.480 193.160 1243.740 193.420 ;
        RECT 1243.940 193.160 1244.200 193.420 ;
        RECT 1242.560 144.880 1242.820 145.140 ;
        RECT 1243.480 144.880 1243.740 145.140 ;
        RECT 1242.100 110.200 1242.360 110.460 ;
        RECT 1243.020 110.200 1243.280 110.460 ;
        RECT 1120.660 18.060 1120.920 18.320 ;
        RECT 1144.120 18.060 1144.380 18.320 ;
        RECT 1144.120 16.700 1144.380 16.960 ;
        RECT 1243.020 17.720 1243.280 17.980 ;
      LAYER met2 ;
        RECT 1246.930 600.850 1247.210 604.000 ;
        RECT 1244.460 600.710 1247.210 600.850 ;
        RECT 1244.460 596.770 1244.600 600.710 ;
        RECT 1246.930 600.000 1247.210 600.710 ;
        RECT 1243.080 596.630 1244.600 596.770 ;
        RECT 1243.080 545.090 1243.220 596.630 ;
        RECT 1242.620 544.950 1243.220 545.090 ;
        RECT 1242.620 497.070 1242.760 544.950 ;
        RECT 1242.560 496.750 1242.820 497.070 ;
        RECT 1242.100 496.410 1242.360 496.730 ;
        RECT 1242.160 483.325 1242.300 496.410 ;
        RECT 1242.090 482.955 1242.370 483.325 ;
        RECT 1243.010 482.955 1243.290 483.325 ;
        RECT 1243.080 435.190 1243.220 482.955 ;
        RECT 1243.020 434.870 1243.280 435.190 ;
        RECT 1243.480 434.190 1243.740 434.510 ;
        RECT 1243.540 420.910 1243.680 434.190 ;
        RECT 1242.560 420.590 1242.820 420.910 ;
        RECT 1243.480 420.590 1243.740 420.910 ;
        RECT 1242.620 372.970 1242.760 420.590 ;
        RECT 1242.560 372.650 1242.820 372.970 ;
        RECT 1243.940 372.650 1244.200 372.970 ;
        RECT 1244.000 331.490 1244.140 372.650 ;
        RECT 1242.560 331.170 1242.820 331.490 ;
        RECT 1243.940 331.170 1244.200 331.490 ;
        RECT 1242.620 303.690 1242.760 331.170 ;
        RECT 1242.160 303.610 1242.760 303.690 ;
        RECT 1242.100 303.550 1242.760 303.610 ;
        RECT 1242.100 303.290 1242.360 303.550 ;
        RECT 1243.020 303.290 1243.280 303.610 ;
        RECT 1243.080 265.610 1243.220 303.290 ;
        RECT 1243.080 265.470 1244.140 265.610 ;
        RECT 1244.000 254.730 1244.140 265.470 ;
        RECT 1243.540 254.590 1244.140 254.730 ;
        RECT 1243.540 241.130 1243.680 254.590 ;
        RECT 1243.080 240.990 1243.680 241.130 ;
        RECT 1243.080 217.590 1243.220 240.990 ;
        RECT 1243.020 217.270 1243.280 217.590 ;
        RECT 1243.940 217.270 1244.200 217.590 ;
        RECT 1244.000 193.450 1244.140 217.270 ;
        RECT 1243.480 193.130 1243.740 193.450 ;
        RECT 1243.940 193.130 1244.200 193.450 ;
        RECT 1243.540 145.170 1243.680 193.130 ;
        RECT 1242.560 144.850 1242.820 145.170 ;
        RECT 1243.480 144.850 1243.740 145.170 ;
        RECT 1242.620 110.570 1242.760 144.850 ;
        RECT 1242.160 110.490 1242.760 110.570 ;
        RECT 1242.100 110.430 1242.760 110.490 ;
        RECT 1242.100 110.170 1242.360 110.430 ;
        RECT 1243.020 110.170 1243.280 110.490 ;
        RECT 1243.080 60.250 1243.220 110.170 ;
        RECT 1243.080 60.110 1243.680 60.250 ;
        RECT 1243.540 58.890 1243.680 60.110 ;
        RECT 1243.080 58.750 1243.680 58.890 ;
        RECT 1120.660 18.030 1120.920 18.350 ;
        RECT 1144.120 18.030 1144.380 18.350 ;
        RECT 1120.720 2.400 1120.860 18.030 ;
        RECT 1144.180 16.990 1144.320 18.030 ;
        RECT 1243.080 18.010 1243.220 58.750 ;
        RECT 1243.020 17.690 1243.280 18.010 ;
        RECT 1144.120 16.670 1144.380 16.990 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
      LAYER via2 ;
        RECT 1242.090 483.000 1242.370 483.280 ;
        RECT 1243.010 483.000 1243.290 483.280 ;
      LAYER met3 ;
        RECT 1242.065 483.290 1242.395 483.305 ;
        RECT 1242.985 483.290 1243.315 483.305 ;
        RECT 1242.065 482.990 1243.315 483.290 ;
        RECT 1242.065 482.975 1242.395 482.990 ;
        RECT 1242.985 482.975 1243.315 482.990 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 590.140 1145.330 590.200 ;
        RECT 1256.330 590.140 1256.650 590.200 ;
        RECT 1145.010 590.000 1256.650 590.140 ;
        RECT 1145.010 589.940 1145.330 590.000 ;
        RECT 1256.330 589.940 1256.650 590.000 ;
        RECT 1138.570 20.640 1138.890 20.700 ;
        RECT 1145.010 20.640 1145.330 20.700 ;
        RECT 1138.570 20.500 1145.330 20.640 ;
        RECT 1138.570 20.440 1138.890 20.500 ;
        RECT 1145.010 20.440 1145.330 20.500 ;
      LAYER via ;
        RECT 1145.040 589.940 1145.300 590.200 ;
        RECT 1256.360 589.940 1256.620 590.200 ;
        RECT 1138.600 20.440 1138.860 20.700 ;
        RECT 1145.040 20.440 1145.300 20.700 ;
      LAYER met2 ;
        RECT 1256.130 600.000 1256.410 604.000 ;
        RECT 1256.190 598.810 1256.330 600.000 ;
        RECT 1256.190 598.670 1256.560 598.810 ;
        RECT 1256.420 590.230 1256.560 598.670 ;
        RECT 1145.040 589.910 1145.300 590.230 ;
        RECT 1256.360 589.910 1256.620 590.230 ;
        RECT 1145.100 20.730 1145.240 589.910 ;
        RECT 1138.600 20.410 1138.860 20.730 ;
        RECT 1145.040 20.410 1145.300 20.730 ;
        RECT 1138.660 2.400 1138.800 20.410 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.810 591.840 1159.130 591.900 ;
        RECT 1263.690 591.840 1264.010 591.900 ;
        RECT 1158.810 591.700 1264.010 591.840 ;
        RECT 1158.810 591.640 1159.130 591.700 ;
        RECT 1263.690 591.640 1264.010 591.700 ;
        RECT 1156.510 20.640 1156.830 20.700 ;
        RECT 1158.810 20.640 1159.130 20.700 ;
        RECT 1156.510 20.500 1159.130 20.640 ;
        RECT 1156.510 20.440 1156.830 20.500 ;
        RECT 1158.810 20.440 1159.130 20.500 ;
      LAYER via ;
        RECT 1158.840 591.640 1159.100 591.900 ;
        RECT 1263.720 591.640 1263.980 591.900 ;
        RECT 1156.540 20.440 1156.800 20.700 ;
        RECT 1158.840 20.440 1159.100 20.700 ;
      LAYER met2 ;
        RECT 1265.330 600.170 1265.610 604.000 ;
        RECT 1263.780 600.030 1265.610 600.170 ;
        RECT 1263.780 591.930 1263.920 600.030 ;
        RECT 1265.330 600.000 1265.610 600.030 ;
        RECT 1158.840 591.610 1159.100 591.930 ;
        RECT 1263.720 591.610 1263.980 591.930 ;
        RECT 1158.900 20.730 1159.040 591.610 ;
        RECT 1156.540 20.410 1156.800 20.730 ;
        RECT 1158.840 20.410 1159.100 20.730 ;
        RECT 1156.600 2.400 1156.740 20.410 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1014.370 572.800 1014.690 572.860 ;
        RECT 1015.750 572.800 1016.070 572.860 ;
        RECT 1014.370 572.660 1016.070 572.800 ;
        RECT 1014.370 572.600 1014.690 572.660 ;
        RECT 1015.750 572.600 1016.070 572.660 ;
        RECT 674.430 37.980 674.750 38.040 ;
        RECT 1014.370 37.980 1014.690 38.040 ;
        RECT 674.430 37.840 1014.690 37.980 ;
        RECT 674.430 37.780 674.750 37.840 ;
        RECT 1014.370 37.780 1014.690 37.840 ;
      LAYER via ;
        RECT 1014.400 572.600 1014.660 572.860 ;
        RECT 1015.780 572.600 1016.040 572.860 ;
        RECT 674.460 37.780 674.720 38.040 ;
        RECT 1014.400 37.780 1014.660 38.040 ;
      LAYER met2 ;
        RECT 1017.390 600.170 1017.670 604.000 ;
        RECT 1015.840 600.030 1017.670 600.170 ;
        RECT 1015.840 572.890 1015.980 600.030 ;
        RECT 1017.390 600.000 1017.670 600.030 ;
        RECT 1014.400 572.570 1014.660 572.890 ;
        RECT 1015.780 572.570 1016.040 572.890 ;
        RECT 1014.460 38.070 1014.600 572.570 ;
        RECT 674.460 37.750 674.720 38.070 ;
        RECT 1014.400 37.750 1014.660 38.070 ;
        RECT 674.520 2.400 674.660 37.750 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1252.190 586.740 1252.510 586.800 ;
        RECT 1272.890 586.740 1273.210 586.800 ;
        RECT 1252.190 586.600 1273.210 586.740 ;
        RECT 1252.190 586.540 1252.510 586.600 ;
        RECT 1272.890 586.540 1273.210 586.600 ;
        RECT 1173.990 18.940 1174.310 19.000 ;
        RECT 1252.190 18.940 1252.510 19.000 ;
        RECT 1173.990 18.800 1252.510 18.940 ;
        RECT 1173.990 18.740 1174.310 18.800 ;
        RECT 1252.190 18.740 1252.510 18.800 ;
      LAYER via ;
        RECT 1252.220 586.540 1252.480 586.800 ;
        RECT 1272.920 586.540 1273.180 586.800 ;
        RECT 1174.020 18.740 1174.280 19.000 ;
        RECT 1252.220 18.740 1252.480 19.000 ;
      LAYER met2 ;
        RECT 1274.530 600.170 1274.810 604.000 ;
        RECT 1272.980 600.030 1274.810 600.170 ;
        RECT 1272.980 586.830 1273.120 600.030 ;
        RECT 1274.530 600.000 1274.810 600.030 ;
        RECT 1252.220 586.510 1252.480 586.830 ;
        RECT 1272.920 586.510 1273.180 586.830 ;
        RECT 1252.280 19.030 1252.420 586.510 ;
        RECT 1174.020 18.710 1174.280 19.030 ;
        RECT 1252.220 18.710 1252.480 19.030 ;
        RECT 1174.080 2.400 1174.220 18.710 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1193.310 589.120 1193.630 589.180 ;
        RECT 1283.470 589.120 1283.790 589.180 ;
        RECT 1193.310 588.980 1283.790 589.120 ;
        RECT 1193.310 588.920 1193.630 588.980 ;
        RECT 1283.470 588.920 1283.790 588.980 ;
        RECT 1191.010 96.460 1191.330 96.520 ;
        RECT 1193.310 96.460 1193.630 96.520 ;
        RECT 1191.010 96.320 1193.630 96.460 ;
        RECT 1191.010 96.260 1191.330 96.320 ;
        RECT 1193.310 96.260 1193.630 96.320 ;
        RECT 1191.010 48.520 1191.330 48.580 ;
        RECT 1191.930 48.520 1192.250 48.580 ;
        RECT 1191.010 48.380 1192.250 48.520 ;
        RECT 1191.010 48.320 1191.330 48.380 ;
        RECT 1191.930 48.320 1192.250 48.380 ;
      LAYER via ;
        RECT 1193.340 588.920 1193.600 589.180 ;
        RECT 1283.500 588.920 1283.760 589.180 ;
        RECT 1191.040 96.260 1191.300 96.520 ;
        RECT 1193.340 96.260 1193.600 96.520 ;
        RECT 1191.040 48.320 1191.300 48.580 ;
        RECT 1191.960 48.320 1192.220 48.580 ;
      LAYER met2 ;
        RECT 1283.730 600.000 1284.010 604.000 ;
        RECT 1283.790 598.810 1283.930 600.000 ;
        RECT 1283.560 598.670 1283.930 598.810 ;
        RECT 1283.560 589.210 1283.700 598.670 ;
        RECT 1193.340 588.890 1193.600 589.210 ;
        RECT 1283.500 588.890 1283.760 589.210 ;
        RECT 1193.400 96.550 1193.540 588.890 ;
        RECT 1191.040 96.230 1191.300 96.550 ;
        RECT 1193.340 96.230 1193.600 96.550 ;
        RECT 1191.100 48.610 1191.240 96.230 ;
        RECT 1191.040 48.290 1191.300 48.610 ;
        RECT 1191.960 48.290 1192.220 48.610 ;
        RECT 1192.020 2.400 1192.160 48.290 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1266.910 593.200 1267.230 593.260 ;
        RECT 1291.290 593.200 1291.610 593.260 ;
        RECT 1266.910 593.060 1291.610 593.200 ;
        RECT 1266.910 593.000 1267.230 593.060 ;
        RECT 1291.290 593.000 1291.610 593.060 ;
        RECT 1256.790 590.140 1257.110 590.200 ;
        RECT 1266.910 590.140 1267.230 590.200 ;
        RECT 1256.790 590.000 1267.230 590.140 ;
        RECT 1256.790 589.940 1257.110 590.000 ;
        RECT 1266.910 589.940 1267.230 590.000 ;
        RECT 1217.690 587.080 1218.010 587.140 ;
        RECT 1217.690 586.940 1227.120 587.080 ;
        RECT 1217.690 586.880 1218.010 586.940 ;
        RECT 1226.980 586.740 1227.120 586.940 ;
        RECT 1226.980 586.600 1251.960 586.740 ;
        RECT 1251.820 586.400 1251.960 586.600 ;
        RECT 1256.790 586.400 1257.110 586.460 ;
        RECT 1251.820 586.260 1257.110 586.400 ;
        RECT 1256.790 586.200 1257.110 586.260 ;
        RECT 1209.870 20.300 1210.190 20.360 ;
        RECT 1217.690 20.300 1218.010 20.360 ;
        RECT 1209.870 20.160 1218.010 20.300 ;
        RECT 1209.870 20.100 1210.190 20.160 ;
        RECT 1217.690 20.100 1218.010 20.160 ;
      LAYER via ;
        RECT 1266.940 593.000 1267.200 593.260 ;
        RECT 1291.320 593.000 1291.580 593.260 ;
        RECT 1256.820 589.940 1257.080 590.200 ;
        RECT 1266.940 589.940 1267.200 590.200 ;
        RECT 1217.720 586.880 1217.980 587.140 ;
        RECT 1256.820 586.200 1257.080 586.460 ;
        RECT 1209.900 20.100 1210.160 20.360 ;
        RECT 1217.720 20.100 1217.980 20.360 ;
      LAYER met2 ;
        RECT 1292.470 600.170 1292.750 604.000 ;
        RECT 1291.380 600.030 1292.750 600.170 ;
        RECT 1291.380 593.290 1291.520 600.030 ;
        RECT 1292.470 600.000 1292.750 600.030 ;
        RECT 1266.940 592.970 1267.200 593.290 ;
        RECT 1291.320 592.970 1291.580 593.290 ;
        RECT 1267.000 590.230 1267.140 592.970 ;
        RECT 1256.820 589.910 1257.080 590.230 ;
        RECT 1266.940 589.910 1267.200 590.230 ;
        RECT 1217.720 586.850 1217.980 587.170 ;
        RECT 1217.780 20.390 1217.920 586.850 ;
        RECT 1256.880 586.490 1257.020 589.910 ;
        RECT 1256.820 586.170 1257.080 586.490 ;
        RECT 1209.900 20.070 1210.160 20.390 ;
        RECT 1217.720 20.070 1217.980 20.390 ;
        RECT 1209.960 2.400 1210.100 20.070 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 587.420 1228.130 587.480 ;
        RECT 1300.030 587.420 1300.350 587.480 ;
        RECT 1227.810 587.280 1300.350 587.420 ;
        RECT 1227.810 587.220 1228.130 587.280 ;
        RECT 1300.030 587.220 1300.350 587.280 ;
      LAYER via ;
        RECT 1227.840 587.220 1228.100 587.480 ;
        RECT 1300.060 587.220 1300.320 587.480 ;
      LAYER met2 ;
        RECT 1301.670 600.170 1301.950 604.000 ;
        RECT 1300.120 600.030 1301.950 600.170 ;
        RECT 1300.120 587.510 1300.260 600.030 ;
        RECT 1301.670 600.000 1301.950 600.030 ;
        RECT 1227.840 587.190 1228.100 587.510 ;
        RECT 1300.060 587.190 1300.320 587.510 ;
        RECT 1227.900 2.400 1228.040 587.190 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 589.800 1248.830 589.860 ;
        RECT 1311.070 589.800 1311.390 589.860 ;
        RECT 1248.510 589.660 1311.390 589.800 ;
        RECT 1248.510 589.600 1248.830 589.660 ;
        RECT 1311.070 589.600 1311.390 589.660 ;
        RECT 1245.750 16.560 1246.070 16.620 ;
        RECT 1248.510 16.560 1248.830 16.620 ;
        RECT 1245.750 16.420 1248.830 16.560 ;
        RECT 1245.750 16.360 1246.070 16.420 ;
        RECT 1248.510 16.360 1248.830 16.420 ;
      LAYER via ;
        RECT 1248.540 589.600 1248.800 589.860 ;
        RECT 1311.100 589.600 1311.360 589.860 ;
        RECT 1245.780 16.360 1246.040 16.620 ;
        RECT 1248.540 16.360 1248.800 16.620 ;
      LAYER met2 ;
        RECT 1310.870 600.000 1311.150 604.000 ;
        RECT 1310.930 598.810 1311.070 600.000 ;
        RECT 1310.930 598.670 1311.300 598.810 ;
        RECT 1311.160 589.890 1311.300 598.670 ;
        RECT 1248.540 589.570 1248.800 589.890 ;
        RECT 1311.100 589.570 1311.360 589.890 ;
        RECT 1248.600 16.650 1248.740 589.570 ;
        RECT 1245.780 16.330 1246.040 16.650 ;
        RECT 1248.540 16.330 1248.800 16.650 ;
        RECT 1245.840 2.400 1245.980 16.330 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1273.350 591.160 1273.670 591.220 ;
        RECT 1318.430 591.160 1318.750 591.220 ;
        RECT 1273.350 591.020 1318.750 591.160 ;
        RECT 1273.350 590.960 1273.670 591.020 ;
        RECT 1318.430 590.960 1318.750 591.020 ;
        RECT 1263.230 15.200 1263.550 15.260 ;
        RECT 1272.890 15.200 1273.210 15.260 ;
        RECT 1263.230 15.060 1273.210 15.200 ;
        RECT 1263.230 15.000 1263.550 15.060 ;
        RECT 1272.890 15.000 1273.210 15.060 ;
      LAYER via ;
        RECT 1273.380 590.960 1273.640 591.220 ;
        RECT 1318.460 590.960 1318.720 591.220 ;
        RECT 1263.260 15.000 1263.520 15.260 ;
        RECT 1272.920 15.000 1273.180 15.260 ;
      LAYER met2 ;
        RECT 1320.070 600.170 1320.350 604.000 ;
        RECT 1318.520 600.030 1320.350 600.170 ;
        RECT 1318.520 591.250 1318.660 600.030 ;
        RECT 1320.070 600.000 1320.350 600.030 ;
        RECT 1273.380 590.930 1273.640 591.250 ;
        RECT 1318.460 590.930 1318.720 591.250 ;
        RECT 1273.440 578.410 1273.580 590.930 ;
        RECT 1272.980 578.270 1273.580 578.410 ;
        RECT 1272.980 15.290 1273.120 578.270 ;
        RECT 1263.260 14.970 1263.520 15.290 ;
        RECT 1272.920 14.970 1273.180 15.290 ;
        RECT 1263.320 2.400 1263.460 14.970 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 592.180 1283.330 592.240 ;
        RECT 1327.630 592.180 1327.950 592.240 ;
        RECT 1283.010 592.040 1327.950 592.180 ;
        RECT 1283.010 591.980 1283.330 592.040 ;
        RECT 1327.630 591.980 1327.950 592.040 ;
      LAYER via ;
        RECT 1283.040 591.980 1283.300 592.240 ;
        RECT 1327.660 591.980 1327.920 592.240 ;
      LAYER met2 ;
        RECT 1329.270 600.170 1329.550 604.000 ;
        RECT 1327.720 600.030 1329.550 600.170 ;
        RECT 1327.720 592.270 1327.860 600.030 ;
        RECT 1329.270 600.000 1329.550 600.030 ;
        RECT 1283.040 591.950 1283.300 592.270 ;
        RECT 1327.660 591.950 1327.920 592.270 ;
        RECT 1283.100 16.730 1283.240 591.950 ;
        RECT 1281.260 16.590 1283.240 16.730 ;
        RECT 1281.260 2.400 1281.400 16.590 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1307.390 588.440 1307.710 588.500 ;
        RECT 1338.670 588.440 1338.990 588.500 ;
        RECT 1307.390 588.300 1338.990 588.440 ;
        RECT 1307.390 588.240 1307.710 588.300 ;
        RECT 1338.670 588.240 1338.990 588.300 ;
        RECT 1299.110 17.580 1299.430 17.640 ;
        RECT 1307.390 17.580 1307.710 17.640 ;
        RECT 1299.110 17.440 1307.710 17.580 ;
        RECT 1299.110 17.380 1299.430 17.440 ;
        RECT 1307.390 17.380 1307.710 17.440 ;
      LAYER via ;
        RECT 1307.420 588.240 1307.680 588.500 ;
        RECT 1338.700 588.240 1338.960 588.500 ;
        RECT 1299.140 17.380 1299.400 17.640 ;
        RECT 1307.420 17.380 1307.680 17.640 ;
      LAYER met2 ;
        RECT 1338.470 600.000 1338.750 604.000 ;
        RECT 1338.530 598.810 1338.670 600.000 ;
        RECT 1338.530 598.670 1338.900 598.810 ;
        RECT 1338.760 588.530 1338.900 598.670 ;
        RECT 1307.420 588.210 1307.680 588.530 ;
        RECT 1338.700 588.210 1338.960 588.530 ;
        RECT 1307.480 17.670 1307.620 588.210 ;
        RECT 1299.140 17.350 1299.400 17.670 ;
        RECT 1307.420 17.350 1307.680 17.670 ;
        RECT 1299.200 2.400 1299.340 17.350 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.050 589.460 1317.370 589.520 ;
        RECT 1346.030 589.460 1346.350 589.520 ;
        RECT 1317.050 589.320 1346.350 589.460 ;
        RECT 1317.050 589.260 1317.370 589.320 ;
        RECT 1346.030 589.260 1346.350 589.320 ;
      LAYER via ;
        RECT 1317.080 589.260 1317.340 589.520 ;
        RECT 1346.060 589.260 1346.320 589.520 ;
      LAYER met2 ;
        RECT 1347.670 600.170 1347.950 604.000 ;
        RECT 1346.120 600.030 1347.950 600.170 ;
        RECT 1346.120 589.550 1346.260 600.030 ;
        RECT 1347.670 600.000 1347.950 600.030 ;
        RECT 1317.080 589.230 1317.340 589.550 ;
        RECT 1346.060 589.230 1346.320 589.550 ;
        RECT 1317.140 2.400 1317.280 589.230 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 587.420 1338.530 587.480 ;
        RECT 1355.230 587.420 1355.550 587.480 ;
        RECT 1338.210 587.280 1355.550 587.420 ;
        RECT 1338.210 587.220 1338.530 587.280 ;
        RECT 1355.230 587.220 1355.550 587.280 ;
        RECT 1334.990 16.560 1335.310 16.620 ;
        RECT 1338.210 16.560 1338.530 16.620 ;
        RECT 1334.990 16.420 1338.530 16.560 ;
        RECT 1334.990 16.360 1335.310 16.420 ;
        RECT 1338.210 16.360 1338.530 16.420 ;
      LAYER via ;
        RECT 1338.240 587.220 1338.500 587.480 ;
        RECT 1355.260 587.220 1355.520 587.480 ;
        RECT 1335.020 16.360 1335.280 16.620 ;
        RECT 1338.240 16.360 1338.500 16.620 ;
      LAYER met2 ;
        RECT 1356.870 600.170 1357.150 604.000 ;
        RECT 1355.320 600.030 1357.150 600.170 ;
        RECT 1355.320 587.510 1355.460 600.030 ;
        RECT 1356.870 600.000 1357.150 600.030 ;
        RECT 1338.240 587.190 1338.500 587.510 ;
        RECT 1355.260 587.190 1355.520 587.510 ;
        RECT 1338.300 16.650 1338.440 587.190 ;
        RECT 1335.020 16.330 1335.280 16.650 ;
        RECT 1338.240 16.330 1338.500 16.650 ;
        RECT 1335.080 2.400 1335.220 16.330 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1021.270 583.000 1021.590 583.060 ;
        RECT 1024.490 583.000 1024.810 583.060 ;
        RECT 1021.270 582.860 1024.810 583.000 ;
        RECT 1021.270 582.800 1021.590 582.860 ;
        RECT 1024.490 582.800 1024.810 582.860 ;
        RECT 692.370 22.340 692.690 22.400 ;
        RECT 1021.270 22.340 1021.590 22.400 ;
        RECT 692.370 22.200 1021.590 22.340 ;
        RECT 692.370 22.140 692.690 22.200 ;
        RECT 1021.270 22.140 1021.590 22.200 ;
      LAYER via ;
        RECT 1021.300 582.800 1021.560 583.060 ;
        RECT 1024.520 582.800 1024.780 583.060 ;
        RECT 692.400 22.140 692.660 22.400 ;
        RECT 1021.300 22.140 1021.560 22.400 ;
      LAYER met2 ;
        RECT 1026.130 600.170 1026.410 604.000 ;
        RECT 1024.580 600.030 1026.410 600.170 ;
        RECT 1024.580 583.090 1024.720 600.030 ;
        RECT 1026.130 600.000 1026.410 600.030 ;
        RECT 1021.300 582.770 1021.560 583.090 ;
        RECT 1024.520 582.770 1024.780 583.090 ;
        RECT 1021.360 22.430 1021.500 582.770 ;
        RECT 692.400 22.110 692.660 22.430 ;
        RECT 1021.300 22.110 1021.560 22.430 ;
        RECT 692.460 2.400 692.600 22.110 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.470 17.240 1352.790 17.300 ;
        RECT 1366.730 17.240 1367.050 17.300 ;
        RECT 1352.470 17.100 1367.050 17.240 ;
        RECT 1352.470 17.040 1352.790 17.100 ;
        RECT 1366.730 17.040 1367.050 17.100 ;
      LAYER via ;
        RECT 1352.500 17.040 1352.760 17.300 ;
        RECT 1366.760 17.040 1367.020 17.300 ;
      LAYER met2 ;
        RECT 1366.070 600.170 1366.350 604.000 ;
        RECT 1366.070 600.030 1366.960 600.170 ;
        RECT 1366.070 600.000 1366.350 600.030 ;
        RECT 1366.820 17.330 1366.960 600.030 ;
        RECT 1352.500 17.010 1352.760 17.330 ;
        RECT 1366.760 17.010 1367.020 17.330 ;
        RECT 1352.560 2.400 1352.700 17.010 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.410 20.640 1370.730 20.700 ;
        RECT 1372.710 20.640 1373.030 20.700 ;
        RECT 1370.410 20.500 1373.030 20.640 ;
        RECT 1370.410 20.440 1370.730 20.500 ;
        RECT 1372.710 20.440 1373.030 20.500 ;
      LAYER via ;
        RECT 1370.440 20.440 1370.700 20.700 ;
        RECT 1372.740 20.440 1373.000 20.700 ;
      LAYER met2 ;
        RECT 1375.270 600.170 1375.550 604.000 ;
        RECT 1373.260 600.030 1375.550 600.170 ;
        RECT 1373.260 586.570 1373.400 600.030 ;
        RECT 1375.270 600.000 1375.550 600.030 ;
        RECT 1372.800 586.430 1373.400 586.570 ;
        RECT 1372.800 20.730 1372.940 586.430 ;
        RECT 1370.440 20.410 1370.700 20.730 ;
        RECT 1372.740 20.410 1373.000 20.730 ;
        RECT 1370.500 2.400 1370.640 20.410 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1384.470 600.170 1384.750 604.000 ;
        RECT 1384.470 600.030 1386.740 600.170 ;
        RECT 1384.470 600.000 1384.750 600.030 ;
        RECT 1386.600 19.450 1386.740 600.030 ;
        RECT 1386.600 19.310 1388.580 19.450 ;
        RECT 1388.440 2.400 1388.580 19.310 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1395.250 586.740 1395.570 586.800 ;
        RECT 1401.690 586.740 1402.010 586.800 ;
        RECT 1395.250 586.600 1402.010 586.740 ;
        RECT 1395.250 586.540 1395.570 586.600 ;
        RECT 1401.690 586.540 1402.010 586.600 ;
        RECT 1402.150 48.520 1402.470 48.580 ;
        RECT 1406.290 48.520 1406.610 48.580 ;
        RECT 1402.150 48.380 1406.610 48.520 ;
        RECT 1402.150 48.320 1402.470 48.380 ;
        RECT 1406.290 48.320 1406.610 48.380 ;
      LAYER via ;
        RECT 1395.280 586.540 1395.540 586.800 ;
        RECT 1401.720 586.540 1401.980 586.800 ;
        RECT 1402.180 48.320 1402.440 48.580 ;
        RECT 1406.320 48.320 1406.580 48.580 ;
      LAYER met2 ;
        RECT 1393.670 600.170 1393.950 604.000 ;
        RECT 1393.670 600.030 1395.480 600.170 ;
        RECT 1393.670 600.000 1393.950 600.030 ;
        RECT 1395.340 586.830 1395.480 600.030 ;
        RECT 1395.280 586.510 1395.540 586.830 ;
        RECT 1401.720 586.510 1401.980 586.830 ;
        RECT 1401.780 72.490 1401.920 586.510 ;
        RECT 1401.780 72.350 1402.380 72.490 ;
        RECT 1402.240 48.610 1402.380 72.350 ;
        RECT 1402.180 48.290 1402.440 48.610 ;
        RECT 1406.320 48.290 1406.580 48.610 ;
        RECT 1406.380 2.400 1406.520 48.290 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1404.450 586.740 1404.770 586.800 ;
        RECT 1406.750 586.740 1407.070 586.800 ;
        RECT 1404.450 586.600 1407.070 586.740 ;
        RECT 1404.450 586.540 1404.770 586.600 ;
        RECT 1406.750 586.540 1407.070 586.600 ;
        RECT 1406.750 15.880 1407.070 15.940 ;
        RECT 1423.770 15.880 1424.090 15.940 ;
        RECT 1406.750 15.740 1424.090 15.880 ;
        RECT 1406.750 15.680 1407.070 15.740 ;
        RECT 1423.770 15.680 1424.090 15.740 ;
      LAYER via ;
        RECT 1404.480 586.540 1404.740 586.800 ;
        RECT 1406.780 586.540 1407.040 586.800 ;
        RECT 1406.780 15.680 1407.040 15.940 ;
        RECT 1423.800 15.680 1424.060 15.940 ;
      LAYER met2 ;
        RECT 1402.870 600.170 1403.150 604.000 ;
        RECT 1402.870 600.030 1404.680 600.170 ;
        RECT 1402.870 600.000 1403.150 600.030 ;
        RECT 1404.540 586.830 1404.680 600.030 ;
        RECT 1404.480 586.510 1404.740 586.830 ;
        RECT 1406.780 586.510 1407.040 586.830 ;
        RECT 1406.840 15.970 1406.980 586.510 ;
        RECT 1406.780 15.650 1407.040 15.970 ;
        RECT 1423.800 15.650 1424.060 15.970 ;
        RECT 1423.860 2.400 1424.000 15.650 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1413.650 587.420 1413.970 587.480 ;
        RECT 1424.690 587.420 1425.010 587.480 ;
        RECT 1413.650 587.280 1425.010 587.420 ;
        RECT 1413.650 587.220 1413.970 587.280 ;
        RECT 1424.690 587.220 1425.010 587.280 ;
        RECT 1424.690 20.640 1425.010 20.700 ;
        RECT 1441.710 20.640 1442.030 20.700 ;
        RECT 1424.690 20.500 1442.030 20.640 ;
        RECT 1424.690 20.440 1425.010 20.500 ;
        RECT 1441.710 20.440 1442.030 20.500 ;
      LAYER via ;
        RECT 1413.680 587.220 1413.940 587.480 ;
        RECT 1424.720 587.220 1424.980 587.480 ;
        RECT 1424.720 20.440 1424.980 20.700 ;
        RECT 1441.740 20.440 1442.000 20.700 ;
      LAYER met2 ;
        RECT 1412.070 600.170 1412.350 604.000 ;
        RECT 1412.070 600.030 1413.880 600.170 ;
        RECT 1412.070 600.000 1412.350 600.030 ;
        RECT 1413.740 587.510 1413.880 600.030 ;
        RECT 1413.680 587.190 1413.940 587.510 ;
        RECT 1424.720 587.190 1424.980 587.510 ;
        RECT 1424.780 20.730 1424.920 587.190 ;
        RECT 1424.720 20.410 1424.980 20.730 ;
        RECT 1441.740 20.410 1442.000 20.730 ;
        RECT 1441.800 2.400 1441.940 20.410 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1422.850 590.480 1423.170 590.540 ;
        RECT 1456.890 590.480 1457.210 590.540 ;
        RECT 1422.850 590.340 1457.210 590.480 ;
        RECT 1422.850 590.280 1423.170 590.340 ;
        RECT 1456.890 590.280 1457.210 590.340 ;
        RECT 1456.890 2.960 1457.210 3.020 ;
        RECT 1459.650 2.960 1459.970 3.020 ;
        RECT 1456.890 2.820 1459.970 2.960 ;
        RECT 1456.890 2.760 1457.210 2.820 ;
        RECT 1459.650 2.760 1459.970 2.820 ;
      LAYER via ;
        RECT 1422.880 590.280 1423.140 590.540 ;
        RECT 1456.920 590.280 1457.180 590.540 ;
        RECT 1456.920 2.760 1457.180 3.020 ;
        RECT 1459.680 2.760 1459.940 3.020 ;
      LAYER met2 ;
        RECT 1421.270 600.170 1421.550 604.000 ;
        RECT 1421.270 600.030 1423.080 600.170 ;
        RECT 1421.270 600.000 1421.550 600.030 ;
        RECT 1422.940 590.570 1423.080 600.030 ;
        RECT 1422.880 590.250 1423.140 590.570 ;
        RECT 1456.920 590.250 1457.180 590.570 ;
        RECT 1456.980 3.050 1457.120 590.250 ;
        RECT 1456.920 2.730 1457.180 3.050 ;
        RECT 1459.680 2.730 1459.940 3.050 ;
        RECT 1459.740 2.400 1459.880 2.730 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1432.050 586.740 1432.370 586.800 ;
        RECT 1434.810 586.740 1435.130 586.800 ;
        RECT 1432.050 586.600 1435.130 586.740 ;
        RECT 1432.050 586.540 1432.370 586.600 ;
        RECT 1434.810 586.540 1435.130 586.600 ;
        RECT 1434.810 19.280 1435.130 19.340 ;
        RECT 1477.590 19.280 1477.910 19.340 ;
        RECT 1434.810 19.140 1477.910 19.280 ;
        RECT 1434.810 19.080 1435.130 19.140 ;
        RECT 1477.590 19.080 1477.910 19.140 ;
      LAYER via ;
        RECT 1432.080 586.540 1432.340 586.800 ;
        RECT 1434.840 586.540 1435.100 586.800 ;
        RECT 1434.840 19.080 1435.100 19.340 ;
        RECT 1477.620 19.080 1477.880 19.340 ;
      LAYER met2 ;
        RECT 1430.470 600.170 1430.750 604.000 ;
        RECT 1430.470 600.030 1432.280 600.170 ;
        RECT 1430.470 600.000 1430.750 600.030 ;
        RECT 1432.140 586.830 1432.280 600.030 ;
        RECT 1432.080 586.510 1432.340 586.830 ;
        RECT 1434.840 586.510 1435.100 586.830 ;
        RECT 1434.900 19.370 1435.040 586.510 ;
        RECT 1434.840 19.050 1435.100 19.370 ;
        RECT 1477.620 19.050 1477.880 19.370 ;
        RECT 1477.680 2.400 1477.820 19.050 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1440.330 18.940 1440.650 19.000 ;
        RECT 1495.530 18.940 1495.850 19.000 ;
        RECT 1440.330 18.800 1495.850 18.940 ;
        RECT 1440.330 18.740 1440.650 18.800 ;
        RECT 1495.530 18.740 1495.850 18.800 ;
      LAYER via ;
        RECT 1440.360 18.740 1440.620 19.000 ;
        RECT 1495.560 18.740 1495.820 19.000 ;
      LAYER met2 ;
        RECT 1439.670 600.170 1439.950 604.000 ;
        RECT 1439.670 600.030 1441.480 600.170 ;
        RECT 1439.670 600.000 1439.950 600.030 ;
        RECT 1441.340 41.890 1441.480 600.030 ;
        RECT 1440.420 41.750 1441.480 41.890 ;
        RECT 1440.420 19.030 1440.560 41.750 ;
        RECT 1440.360 18.710 1440.620 19.030 ;
        RECT 1495.560 18.710 1495.820 19.030 ;
        RECT 1495.620 2.400 1495.760 18.710 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1449.990 586.740 1450.310 586.800 ;
        RECT 1455.510 586.740 1455.830 586.800 ;
        RECT 1449.990 586.600 1455.830 586.740 ;
        RECT 1449.990 586.540 1450.310 586.600 ;
        RECT 1455.510 586.540 1455.830 586.600 ;
        RECT 1455.510 17.920 1455.830 17.980 ;
        RECT 1513.010 17.920 1513.330 17.980 ;
        RECT 1455.510 17.780 1513.330 17.920 ;
        RECT 1455.510 17.720 1455.830 17.780 ;
        RECT 1513.010 17.720 1513.330 17.780 ;
      LAYER via ;
        RECT 1450.020 586.540 1450.280 586.800 ;
        RECT 1455.540 586.540 1455.800 586.800 ;
        RECT 1455.540 17.720 1455.800 17.980 ;
        RECT 1513.040 17.720 1513.300 17.980 ;
      LAYER met2 ;
        RECT 1448.870 600.170 1449.150 604.000 ;
        RECT 1448.870 600.030 1450.220 600.170 ;
        RECT 1448.870 600.000 1449.150 600.030 ;
        RECT 1450.080 586.830 1450.220 600.030 ;
        RECT 1450.020 586.510 1450.280 586.830 ;
        RECT 1455.540 586.510 1455.800 586.830 ;
        RECT 1455.600 18.010 1455.740 586.510 ;
        RECT 1455.540 17.690 1455.800 18.010 ;
        RECT 1513.040 17.690 1513.300 18.010 ;
        RECT 1513.100 2.400 1513.240 17.690 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1035.070 290.060 1035.390 290.320 ;
        RECT 1035.160 289.640 1035.300 290.060 ;
        RECT 1035.070 289.380 1035.390 289.640 ;
        RECT 710.310 24.380 710.630 24.440 ;
        RECT 1035.070 24.380 1035.390 24.440 ;
        RECT 710.310 24.240 1035.390 24.380 ;
        RECT 710.310 24.180 710.630 24.240 ;
        RECT 1035.070 24.180 1035.390 24.240 ;
      LAYER via ;
        RECT 1035.100 290.060 1035.360 290.320 ;
        RECT 1035.100 289.380 1035.360 289.640 ;
        RECT 710.340 24.180 710.600 24.440 ;
        RECT 1035.100 24.180 1035.360 24.440 ;
      LAYER met2 ;
        RECT 1035.330 600.000 1035.610 604.000 ;
        RECT 1035.390 598.810 1035.530 600.000 ;
        RECT 1035.160 598.670 1035.530 598.810 ;
        RECT 1035.160 290.350 1035.300 598.670 ;
        RECT 1035.100 290.030 1035.360 290.350 ;
        RECT 1035.100 289.350 1035.360 289.670 ;
        RECT 1035.160 24.470 1035.300 289.350 ;
        RECT 710.340 24.150 710.600 24.470 ;
        RECT 1035.100 24.150 1035.360 24.470 ;
        RECT 710.400 2.400 710.540 24.150 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1459.650 586.740 1459.970 586.800 ;
        RECT 1462.410 586.740 1462.730 586.800 ;
        RECT 1459.650 586.600 1462.730 586.740 ;
        RECT 1459.650 586.540 1459.970 586.600 ;
        RECT 1462.410 586.540 1462.730 586.600 ;
        RECT 1462.410 16.560 1462.730 16.620 ;
        RECT 1530.950 16.560 1531.270 16.620 ;
        RECT 1462.410 16.420 1531.270 16.560 ;
        RECT 1462.410 16.360 1462.730 16.420 ;
        RECT 1530.950 16.360 1531.270 16.420 ;
      LAYER via ;
        RECT 1459.680 586.540 1459.940 586.800 ;
        RECT 1462.440 586.540 1462.700 586.800 ;
        RECT 1462.440 16.360 1462.700 16.620 ;
        RECT 1530.980 16.360 1531.240 16.620 ;
      LAYER met2 ;
        RECT 1458.070 600.170 1458.350 604.000 ;
        RECT 1458.070 600.030 1459.880 600.170 ;
        RECT 1458.070 600.000 1458.350 600.030 ;
        RECT 1459.740 586.830 1459.880 600.030 ;
        RECT 1459.680 586.510 1459.940 586.830 ;
        RECT 1462.440 586.510 1462.700 586.830 ;
        RECT 1462.500 16.650 1462.640 586.510 ;
        RECT 1462.440 16.330 1462.700 16.650 ;
        RECT 1530.980 16.330 1531.240 16.650 ;
        RECT 1531.040 2.400 1531.180 16.330 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1468.850 591.160 1469.170 591.220 ;
        RECT 1514.390 591.160 1514.710 591.220 ;
        RECT 1468.850 591.020 1514.710 591.160 ;
        RECT 1468.850 590.960 1469.170 591.020 ;
        RECT 1514.390 590.960 1514.710 591.020 ;
        RECT 1514.390 15.880 1514.710 15.940 ;
        RECT 1548.890 15.880 1549.210 15.940 ;
        RECT 1514.390 15.740 1549.210 15.880 ;
        RECT 1514.390 15.680 1514.710 15.740 ;
        RECT 1548.890 15.680 1549.210 15.740 ;
      LAYER via ;
        RECT 1468.880 590.960 1469.140 591.220 ;
        RECT 1514.420 590.960 1514.680 591.220 ;
        RECT 1514.420 15.680 1514.680 15.940 ;
        RECT 1548.920 15.680 1549.180 15.940 ;
      LAYER met2 ;
        RECT 1467.270 600.170 1467.550 604.000 ;
        RECT 1467.270 600.030 1469.080 600.170 ;
        RECT 1467.270 600.000 1467.550 600.030 ;
        RECT 1468.940 591.250 1469.080 600.030 ;
        RECT 1468.880 590.930 1469.140 591.250 ;
        RECT 1514.420 590.930 1514.680 591.250 ;
        RECT 1514.480 15.970 1514.620 590.930 ;
        RECT 1514.420 15.650 1514.680 15.970 ;
        RECT 1548.920 15.650 1549.180 15.970 ;
        RECT 1548.980 2.400 1549.120 15.650 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1478.050 590.820 1478.370 590.880 ;
        RECT 1541.990 590.820 1542.310 590.880 ;
        RECT 1478.050 590.680 1542.310 590.820 ;
        RECT 1478.050 590.620 1478.370 590.680 ;
        RECT 1541.990 590.620 1542.310 590.680 ;
        RECT 1541.990 14.860 1542.310 14.920 ;
        RECT 1566.830 14.860 1567.150 14.920 ;
        RECT 1541.990 14.720 1567.150 14.860 ;
        RECT 1541.990 14.660 1542.310 14.720 ;
        RECT 1566.830 14.660 1567.150 14.720 ;
      LAYER via ;
        RECT 1478.080 590.620 1478.340 590.880 ;
        RECT 1542.020 590.620 1542.280 590.880 ;
        RECT 1542.020 14.660 1542.280 14.920 ;
        RECT 1566.860 14.660 1567.120 14.920 ;
      LAYER met2 ;
        RECT 1476.470 600.170 1476.750 604.000 ;
        RECT 1476.470 600.030 1478.280 600.170 ;
        RECT 1476.470 600.000 1476.750 600.030 ;
        RECT 1478.140 590.910 1478.280 600.030 ;
        RECT 1478.080 590.590 1478.340 590.910 ;
        RECT 1542.020 590.590 1542.280 590.910 ;
        RECT 1542.080 14.950 1542.220 590.590 ;
        RECT 1542.020 14.630 1542.280 14.950 ;
        RECT 1566.860 14.630 1567.120 14.950 ;
        RECT 1566.920 2.400 1567.060 14.630 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1487.250 589.800 1487.570 589.860 ;
        RECT 1490.010 589.800 1490.330 589.860 ;
        RECT 1487.250 589.660 1490.330 589.800 ;
        RECT 1487.250 589.600 1487.570 589.660 ;
        RECT 1490.010 589.600 1490.330 589.660 ;
        RECT 1490.010 20.300 1490.330 20.360 ;
        RECT 1584.770 20.300 1585.090 20.360 ;
        RECT 1490.010 20.160 1585.090 20.300 ;
        RECT 1490.010 20.100 1490.330 20.160 ;
        RECT 1584.770 20.100 1585.090 20.160 ;
      LAYER via ;
        RECT 1487.280 589.600 1487.540 589.860 ;
        RECT 1490.040 589.600 1490.300 589.860 ;
        RECT 1490.040 20.100 1490.300 20.360 ;
        RECT 1584.800 20.100 1585.060 20.360 ;
      LAYER met2 ;
        RECT 1485.670 600.170 1485.950 604.000 ;
        RECT 1485.670 600.030 1487.480 600.170 ;
        RECT 1485.670 600.000 1485.950 600.030 ;
        RECT 1487.340 589.890 1487.480 600.030 ;
        RECT 1487.280 589.570 1487.540 589.890 ;
        RECT 1490.040 589.570 1490.300 589.890 ;
        RECT 1490.100 20.390 1490.240 589.570 ;
        RECT 1490.040 20.070 1490.300 20.390 ;
        RECT 1584.800 20.070 1585.060 20.390 ;
        RECT 1584.860 2.400 1585.000 20.070 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1496.910 19.280 1497.230 19.340 ;
        RECT 1602.250 19.280 1602.570 19.340 ;
        RECT 1496.910 19.140 1602.570 19.280 ;
        RECT 1496.910 19.080 1497.230 19.140 ;
        RECT 1602.250 19.080 1602.570 19.140 ;
      LAYER via ;
        RECT 1496.940 19.080 1497.200 19.340 ;
        RECT 1602.280 19.080 1602.540 19.340 ;
      LAYER met2 ;
        RECT 1494.870 600.170 1495.150 604.000 ;
        RECT 1494.870 600.030 1497.140 600.170 ;
        RECT 1494.870 600.000 1495.150 600.030 ;
        RECT 1497.000 19.370 1497.140 600.030 ;
        RECT 1496.940 19.050 1497.200 19.370 ;
        RECT 1602.280 19.050 1602.540 19.370 ;
        RECT 1602.340 2.400 1602.480 19.050 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1505.650 586.740 1505.970 586.800 ;
        RECT 1510.710 586.740 1511.030 586.800 ;
        RECT 1505.650 586.600 1511.030 586.740 ;
        RECT 1505.650 586.540 1505.970 586.600 ;
        RECT 1510.710 586.540 1511.030 586.600 ;
        RECT 1510.710 19.620 1511.030 19.680 ;
        RECT 1620.190 19.620 1620.510 19.680 ;
        RECT 1510.710 19.480 1620.510 19.620 ;
        RECT 1510.710 19.420 1511.030 19.480 ;
        RECT 1620.190 19.420 1620.510 19.480 ;
      LAYER via ;
        RECT 1505.680 586.540 1505.940 586.800 ;
        RECT 1510.740 586.540 1511.000 586.800 ;
        RECT 1510.740 19.420 1511.000 19.680 ;
        RECT 1620.220 19.420 1620.480 19.680 ;
      LAYER met2 ;
        RECT 1504.070 600.170 1504.350 604.000 ;
        RECT 1504.070 600.030 1505.880 600.170 ;
        RECT 1504.070 600.000 1504.350 600.030 ;
        RECT 1505.740 586.830 1505.880 600.030 ;
        RECT 1505.680 586.510 1505.940 586.830 ;
        RECT 1510.740 586.510 1511.000 586.830 ;
        RECT 1510.800 19.710 1510.940 586.510 ;
        RECT 1510.740 19.390 1511.000 19.710 ;
        RECT 1620.220 19.390 1620.480 19.710 ;
        RECT 1620.280 2.400 1620.420 19.390 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1514.850 586.740 1515.170 586.800 ;
        RECT 1517.610 586.740 1517.930 586.800 ;
        RECT 1514.850 586.600 1517.930 586.740 ;
        RECT 1514.850 586.540 1515.170 586.600 ;
        RECT 1517.610 586.540 1517.930 586.600 ;
        RECT 1517.610 18.600 1517.930 18.660 ;
        RECT 1638.130 18.600 1638.450 18.660 ;
        RECT 1517.610 18.460 1638.450 18.600 ;
        RECT 1517.610 18.400 1517.930 18.460 ;
        RECT 1638.130 18.400 1638.450 18.460 ;
      LAYER via ;
        RECT 1514.880 586.540 1515.140 586.800 ;
        RECT 1517.640 586.540 1517.900 586.800 ;
        RECT 1517.640 18.400 1517.900 18.660 ;
        RECT 1638.160 18.400 1638.420 18.660 ;
      LAYER met2 ;
        RECT 1513.270 600.170 1513.550 604.000 ;
        RECT 1513.270 600.030 1515.080 600.170 ;
        RECT 1513.270 600.000 1513.550 600.030 ;
        RECT 1514.940 586.830 1515.080 600.030 ;
        RECT 1514.880 586.510 1515.140 586.830 ;
        RECT 1517.640 586.510 1517.900 586.830 ;
        RECT 1517.700 18.690 1517.840 586.510 ;
        RECT 1517.640 18.370 1517.900 18.690 ;
        RECT 1638.160 18.370 1638.420 18.690 ;
        RECT 1638.220 2.400 1638.360 18.370 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1524.050 589.460 1524.370 589.520 ;
        RECT 1656.530 589.460 1656.850 589.520 ;
        RECT 1524.050 589.320 1656.850 589.460 ;
        RECT 1524.050 589.260 1524.370 589.320 ;
        RECT 1656.530 589.260 1656.850 589.320 ;
      LAYER via ;
        RECT 1524.080 589.260 1524.340 589.520 ;
        RECT 1656.560 589.260 1656.820 589.520 ;
      LAYER met2 ;
        RECT 1522.470 600.170 1522.750 604.000 ;
        RECT 1522.470 600.030 1524.280 600.170 ;
        RECT 1522.470 600.000 1522.750 600.030 ;
        RECT 1524.140 589.550 1524.280 600.030 ;
        RECT 1524.080 589.230 1524.340 589.550 ;
        RECT 1656.560 589.230 1656.820 589.550 ;
        RECT 1656.620 3.130 1656.760 589.230 ;
        RECT 1656.160 2.990 1656.760 3.130 ;
        RECT 1656.160 2.400 1656.300 2.990 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1533.250 589.120 1533.570 589.180 ;
        RECT 1533.250 588.980 1622.720 589.120 ;
        RECT 1533.250 588.920 1533.570 588.980 ;
        RECT 1622.580 588.440 1622.720 588.980 ;
        RECT 1646.410 588.440 1646.730 588.500 ;
        RECT 1622.580 588.300 1646.730 588.440 ;
        RECT 1646.410 588.240 1646.730 588.300 ;
        RECT 1646.410 572.800 1646.730 572.860 ;
        RECT 1669.870 572.800 1670.190 572.860 ;
        RECT 1646.410 572.660 1670.190 572.800 ;
        RECT 1646.410 572.600 1646.730 572.660 ;
        RECT 1669.870 572.600 1670.190 572.660 ;
        RECT 1669.870 524.180 1670.190 524.240 ;
        RECT 1670.790 524.180 1671.110 524.240 ;
        RECT 1669.870 524.040 1671.110 524.180 ;
        RECT 1669.870 523.980 1670.190 524.040 ;
        RECT 1670.790 523.980 1671.110 524.040 ;
        RECT 1669.870 476.240 1670.190 476.300 ;
        RECT 1670.790 476.240 1671.110 476.300 ;
        RECT 1669.870 476.100 1671.110 476.240 ;
        RECT 1669.870 476.040 1670.190 476.100 ;
        RECT 1670.790 476.040 1671.110 476.100 ;
        RECT 1669.870 427.620 1670.190 427.680 ;
        RECT 1670.790 427.620 1671.110 427.680 ;
        RECT 1669.870 427.480 1671.110 427.620 ;
        RECT 1669.870 427.420 1670.190 427.480 ;
        RECT 1670.790 427.420 1671.110 427.480 ;
        RECT 1669.870 379.680 1670.190 379.740 ;
        RECT 1670.790 379.680 1671.110 379.740 ;
        RECT 1669.870 379.540 1671.110 379.680 ;
        RECT 1669.870 379.480 1670.190 379.540 ;
        RECT 1670.790 379.480 1671.110 379.540 ;
        RECT 1669.870 331.060 1670.190 331.120 ;
        RECT 1670.790 331.060 1671.110 331.120 ;
        RECT 1669.870 330.920 1671.110 331.060 ;
        RECT 1669.870 330.860 1670.190 330.920 ;
        RECT 1670.790 330.860 1671.110 330.920 ;
        RECT 1669.870 283.120 1670.190 283.180 ;
        RECT 1670.790 283.120 1671.110 283.180 ;
        RECT 1669.870 282.980 1671.110 283.120 ;
        RECT 1669.870 282.920 1670.190 282.980 ;
        RECT 1670.790 282.920 1671.110 282.980 ;
        RECT 1669.870 234.500 1670.190 234.560 ;
        RECT 1670.790 234.500 1671.110 234.560 ;
        RECT 1669.870 234.360 1671.110 234.500 ;
        RECT 1669.870 234.300 1670.190 234.360 ;
        RECT 1670.790 234.300 1671.110 234.360 ;
        RECT 1669.870 186.560 1670.190 186.620 ;
        RECT 1670.790 186.560 1671.110 186.620 ;
        RECT 1669.870 186.420 1671.110 186.560 ;
        RECT 1669.870 186.360 1670.190 186.420 ;
        RECT 1670.790 186.360 1671.110 186.420 ;
        RECT 1669.870 137.940 1670.190 138.000 ;
        RECT 1671.710 137.940 1672.030 138.000 ;
        RECT 1669.870 137.800 1672.030 137.940 ;
        RECT 1669.870 137.740 1670.190 137.800 ;
        RECT 1671.710 137.740 1672.030 137.800 ;
        RECT 1672.170 23.700 1672.490 23.760 ;
        RECT 1673.090 23.700 1673.410 23.760 ;
        RECT 1672.170 23.560 1673.410 23.700 ;
        RECT 1672.170 23.500 1672.490 23.560 ;
        RECT 1673.090 23.500 1673.410 23.560 ;
        RECT 1673.090 2.960 1673.410 3.020 ;
        RECT 1673.550 2.960 1673.870 3.020 ;
        RECT 1673.090 2.820 1673.870 2.960 ;
        RECT 1673.090 2.760 1673.410 2.820 ;
        RECT 1673.550 2.760 1673.870 2.820 ;
      LAYER via ;
        RECT 1533.280 588.920 1533.540 589.180 ;
        RECT 1646.440 588.240 1646.700 588.500 ;
        RECT 1646.440 572.600 1646.700 572.860 ;
        RECT 1669.900 572.600 1670.160 572.860 ;
        RECT 1669.900 523.980 1670.160 524.240 ;
        RECT 1670.820 523.980 1671.080 524.240 ;
        RECT 1669.900 476.040 1670.160 476.300 ;
        RECT 1670.820 476.040 1671.080 476.300 ;
        RECT 1669.900 427.420 1670.160 427.680 ;
        RECT 1670.820 427.420 1671.080 427.680 ;
        RECT 1669.900 379.480 1670.160 379.740 ;
        RECT 1670.820 379.480 1671.080 379.740 ;
        RECT 1669.900 330.860 1670.160 331.120 ;
        RECT 1670.820 330.860 1671.080 331.120 ;
        RECT 1669.900 282.920 1670.160 283.180 ;
        RECT 1670.820 282.920 1671.080 283.180 ;
        RECT 1669.900 234.300 1670.160 234.560 ;
        RECT 1670.820 234.300 1671.080 234.560 ;
        RECT 1669.900 186.360 1670.160 186.620 ;
        RECT 1670.820 186.360 1671.080 186.620 ;
        RECT 1669.900 137.740 1670.160 138.000 ;
        RECT 1671.740 137.740 1672.000 138.000 ;
        RECT 1672.200 23.500 1672.460 23.760 ;
        RECT 1673.120 23.500 1673.380 23.760 ;
        RECT 1673.120 2.760 1673.380 3.020 ;
        RECT 1673.580 2.760 1673.840 3.020 ;
      LAYER met2 ;
        RECT 1531.670 600.170 1531.950 604.000 ;
        RECT 1531.670 600.030 1533.480 600.170 ;
        RECT 1531.670 600.000 1531.950 600.030 ;
        RECT 1533.340 589.210 1533.480 600.030 ;
        RECT 1533.280 588.890 1533.540 589.210 ;
        RECT 1646.440 588.210 1646.700 588.530 ;
        RECT 1646.500 572.890 1646.640 588.210 ;
        RECT 1646.440 572.570 1646.700 572.890 ;
        RECT 1669.900 572.570 1670.160 572.890 ;
        RECT 1669.960 524.270 1670.100 572.570 ;
        RECT 1669.900 523.950 1670.160 524.270 ;
        RECT 1670.820 523.950 1671.080 524.270 ;
        RECT 1670.880 476.330 1671.020 523.950 ;
        RECT 1669.900 476.010 1670.160 476.330 ;
        RECT 1670.820 476.010 1671.080 476.330 ;
        RECT 1669.960 427.710 1670.100 476.010 ;
        RECT 1669.900 427.390 1670.160 427.710 ;
        RECT 1670.820 427.390 1671.080 427.710 ;
        RECT 1670.880 379.770 1671.020 427.390 ;
        RECT 1669.900 379.450 1670.160 379.770 ;
        RECT 1670.820 379.450 1671.080 379.770 ;
        RECT 1669.960 331.150 1670.100 379.450 ;
        RECT 1669.900 330.830 1670.160 331.150 ;
        RECT 1670.820 330.830 1671.080 331.150 ;
        RECT 1670.880 283.210 1671.020 330.830 ;
        RECT 1669.900 282.890 1670.160 283.210 ;
        RECT 1670.820 282.890 1671.080 283.210 ;
        RECT 1669.960 234.590 1670.100 282.890 ;
        RECT 1669.900 234.270 1670.160 234.590 ;
        RECT 1670.820 234.270 1671.080 234.590 ;
        RECT 1670.880 186.650 1671.020 234.270 ;
        RECT 1669.900 186.330 1670.160 186.650 ;
        RECT 1670.820 186.330 1671.080 186.650 ;
        RECT 1669.960 138.030 1670.100 186.330 ;
        RECT 1669.900 137.710 1670.160 138.030 ;
        RECT 1671.740 137.710 1672.000 138.030 ;
        RECT 1671.800 61.610 1671.940 137.710 ;
        RECT 1671.800 61.470 1672.860 61.610 ;
        RECT 1672.720 48.010 1672.860 61.470 ;
        RECT 1672.260 47.870 1672.860 48.010 ;
        RECT 1672.260 23.790 1672.400 47.870 ;
        RECT 1672.200 23.470 1672.460 23.790 ;
        RECT 1673.120 23.470 1673.380 23.790 ;
        RECT 1673.180 3.050 1673.320 23.470 ;
        RECT 1673.120 2.730 1673.380 3.050 ;
        RECT 1673.580 2.730 1673.840 3.050 ;
        RECT 1673.640 2.400 1673.780 2.730 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1542.450 592.860 1542.770 592.920 ;
        RECT 1691.950 592.860 1692.270 592.920 ;
        RECT 1542.450 592.720 1692.270 592.860 ;
        RECT 1542.450 592.660 1542.770 592.720 ;
        RECT 1691.950 592.660 1692.270 592.720 ;
      LAYER via ;
        RECT 1542.480 592.660 1542.740 592.920 ;
        RECT 1691.980 592.660 1692.240 592.920 ;
      LAYER met2 ;
        RECT 1540.870 600.170 1541.150 604.000 ;
        RECT 1540.870 600.030 1542.680 600.170 ;
        RECT 1540.870 600.000 1541.150 600.030 ;
        RECT 1542.540 592.950 1542.680 600.030 ;
        RECT 1542.480 592.630 1542.740 592.950 ;
        RECT 1691.980 592.630 1692.240 592.950 ;
        RECT 1692.040 3.130 1692.180 592.630 ;
        RECT 1691.580 2.990 1692.180 3.130 ;
        RECT 1691.580 2.400 1691.720 2.990 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1043.810 497.320 1044.130 497.380 ;
        RECT 1042.980 497.180 1044.130 497.320 ;
        RECT 1042.980 497.040 1043.120 497.180 ;
        RECT 1043.810 497.120 1044.130 497.180 ;
        RECT 1042.890 496.780 1043.210 497.040 ;
        RECT 1042.890 168.880 1043.210 168.940 ;
        RECT 1043.810 168.880 1044.130 168.940 ;
        RECT 1042.890 168.740 1044.130 168.880 ;
        RECT 1042.890 168.680 1043.210 168.740 ;
        RECT 1043.810 168.680 1044.130 168.740 ;
        RECT 1043.810 111.080 1044.130 111.140 ;
        RECT 1042.980 110.940 1044.130 111.080 ;
        RECT 1042.980 110.460 1043.120 110.940 ;
        RECT 1043.810 110.880 1044.130 110.940 ;
        RECT 1042.890 110.200 1043.210 110.460 ;
        RECT 1041.970 62.460 1042.290 62.520 ;
        RECT 1042.890 62.460 1043.210 62.520 ;
        RECT 1041.970 62.320 1043.210 62.460 ;
        RECT 1041.970 62.260 1042.290 62.320 ;
        RECT 1042.890 62.260 1043.210 62.320 ;
        RECT 728.250 24.040 728.570 24.100 ;
        RECT 1041.970 24.040 1042.290 24.100 ;
        RECT 728.250 23.900 1042.290 24.040 ;
        RECT 728.250 23.840 728.570 23.900 ;
        RECT 1041.970 23.840 1042.290 23.900 ;
      LAYER via ;
        RECT 1043.840 497.120 1044.100 497.380 ;
        RECT 1042.920 496.780 1043.180 497.040 ;
        RECT 1042.920 168.680 1043.180 168.940 ;
        RECT 1043.840 168.680 1044.100 168.940 ;
        RECT 1043.840 110.880 1044.100 111.140 ;
        RECT 1042.920 110.200 1043.180 110.460 ;
        RECT 1042.000 62.260 1042.260 62.520 ;
        RECT 1042.920 62.260 1043.180 62.520 ;
        RECT 728.280 23.840 728.540 24.100 ;
        RECT 1042.000 23.840 1042.260 24.100 ;
      LAYER met2 ;
        RECT 1044.530 600.170 1044.810 604.000 ;
        RECT 1043.900 600.030 1044.810 600.170 ;
        RECT 1043.900 497.410 1044.040 600.030 ;
        RECT 1044.530 600.000 1044.810 600.030 ;
        RECT 1043.840 497.090 1044.100 497.410 ;
        RECT 1042.920 496.750 1043.180 497.070 ;
        RECT 1042.980 168.970 1043.120 496.750 ;
        RECT 1042.920 168.650 1043.180 168.970 ;
        RECT 1043.840 168.650 1044.100 168.970 ;
        RECT 1043.900 111.170 1044.040 168.650 ;
        RECT 1043.840 110.850 1044.100 111.170 ;
        RECT 1042.920 110.170 1043.180 110.490 ;
        RECT 1042.980 62.550 1043.120 110.170 ;
        RECT 1042.000 62.230 1042.260 62.550 ;
        RECT 1042.920 62.230 1043.180 62.550 ;
        RECT 1042.060 24.130 1042.200 62.230 ;
        RECT 728.280 23.810 728.540 24.130 ;
        RECT 1042.000 23.810 1042.260 24.130 ;
        RECT 728.340 2.400 728.480 23.810 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1552.110 24.720 1552.430 24.780 ;
        RECT 1709.430 24.720 1709.750 24.780 ;
        RECT 1552.110 24.580 1709.750 24.720 ;
        RECT 1552.110 24.520 1552.430 24.580 ;
        RECT 1709.430 24.520 1709.750 24.580 ;
      LAYER via ;
        RECT 1552.140 24.520 1552.400 24.780 ;
        RECT 1709.460 24.520 1709.720 24.780 ;
      LAYER met2 ;
        RECT 1550.070 600.170 1550.350 604.000 ;
        RECT 1550.070 600.030 1552.340 600.170 ;
        RECT 1550.070 600.000 1550.350 600.030 ;
        RECT 1552.200 24.810 1552.340 600.030 ;
        RECT 1552.140 24.490 1552.400 24.810 ;
        RECT 1709.460 24.490 1709.720 24.810 ;
        RECT 1709.520 2.400 1709.660 24.490 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1558.550 590.820 1558.870 590.880 ;
        RECT 1725.990 590.820 1726.310 590.880 ;
        RECT 1558.550 590.680 1726.310 590.820 ;
        RECT 1558.550 590.620 1558.870 590.680 ;
        RECT 1725.990 590.620 1726.310 590.680 ;
      LAYER via ;
        RECT 1558.580 590.620 1558.840 590.880 ;
        RECT 1726.020 590.620 1726.280 590.880 ;
      LAYER met2 ;
        RECT 1558.810 600.000 1559.090 604.000 ;
        RECT 1558.870 598.810 1559.010 600.000 ;
        RECT 1558.640 598.670 1559.010 598.810 ;
        RECT 1558.640 590.910 1558.780 598.670 ;
        RECT 1558.580 590.590 1558.840 590.910 ;
        RECT 1726.020 590.590 1726.280 590.910 ;
        RECT 1726.080 3.130 1726.220 590.590 ;
        RECT 1726.080 2.990 1727.600 3.130 ;
        RECT 1727.460 2.400 1727.600 2.990 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1569.590 586.740 1569.910 586.800 ;
        RECT 1572.810 586.740 1573.130 586.800 ;
        RECT 1569.590 586.600 1573.130 586.740 ;
        RECT 1569.590 586.540 1569.910 586.600 ;
        RECT 1572.810 586.540 1573.130 586.600 ;
        RECT 1572.810 24.380 1573.130 24.440 ;
        RECT 1745.310 24.380 1745.630 24.440 ;
        RECT 1572.810 24.240 1745.630 24.380 ;
        RECT 1572.810 24.180 1573.130 24.240 ;
        RECT 1745.310 24.180 1745.630 24.240 ;
      LAYER via ;
        RECT 1569.620 586.540 1569.880 586.800 ;
        RECT 1572.840 586.540 1573.100 586.800 ;
        RECT 1572.840 24.180 1573.100 24.440 ;
        RECT 1745.340 24.180 1745.600 24.440 ;
      LAYER met2 ;
        RECT 1568.010 600.170 1568.290 604.000 ;
        RECT 1568.010 600.030 1569.820 600.170 ;
        RECT 1568.010 600.000 1568.290 600.030 ;
        RECT 1569.680 586.830 1569.820 600.030 ;
        RECT 1569.620 586.510 1569.880 586.830 ;
        RECT 1572.840 586.510 1573.100 586.830 ;
        RECT 1572.900 24.470 1573.040 586.510 ;
        RECT 1572.840 24.150 1573.100 24.470 ;
        RECT 1745.340 24.150 1745.600 24.470 ;
        RECT 1745.400 2.400 1745.540 24.150 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1579.710 29.820 1580.030 29.880 ;
        RECT 1762.790 29.820 1763.110 29.880 ;
        RECT 1579.710 29.680 1763.110 29.820 ;
        RECT 1579.710 29.620 1580.030 29.680 ;
        RECT 1762.790 29.620 1763.110 29.680 ;
      LAYER via ;
        RECT 1579.740 29.620 1580.000 29.880 ;
        RECT 1762.820 29.620 1763.080 29.880 ;
      LAYER met2 ;
        RECT 1577.210 600.170 1577.490 604.000 ;
        RECT 1577.210 600.030 1579.940 600.170 ;
        RECT 1577.210 600.000 1577.490 600.030 ;
        RECT 1579.800 29.910 1579.940 600.030 ;
        RECT 1579.740 29.590 1580.000 29.910 ;
        RECT 1762.820 29.590 1763.080 29.910 ;
        RECT 1762.880 2.400 1763.020 29.590 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1586.150 34.240 1586.470 34.300 ;
        RECT 1780.730 34.240 1781.050 34.300 ;
        RECT 1586.150 34.100 1781.050 34.240 ;
        RECT 1586.150 34.040 1586.470 34.100 ;
        RECT 1780.730 34.040 1781.050 34.100 ;
      LAYER via ;
        RECT 1586.180 34.040 1586.440 34.300 ;
        RECT 1780.760 34.040 1781.020 34.300 ;
      LAYER met2 ;
        RECT 1586.410 600.000 1586.690 604.000 ;
        RECT 1586.470 598.810 1586.610 600.000 ;
        RECT 1586.240 598.670 1586.610 598.810 ;
        RECT 1586.240 34.330 1586.380 598.670 ;
        RECT 1586.180 34.010 1586.440 34.330 ;
        RECT 1780.760 34.010 1781.020 34.330 ;
        RECT 1780.820 2.400 1780.960 34.010 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1597.190 586.740 1597.510 586.800 ;
        RECT 1600.410 586.740 1600.730 586.800 ;
        RECT 1597.190 586.600 1600.730 586.740 ;
        RECT 1597.190 586.540 1597.510 586.600 ;
        RECT 1600.410 586.540 1600.730 586.600 ;
        RECT 1600.410 16.900 1600.730 16.960 ;
        RECT 1798.670 16.900 1798.990 16.960 ;
        RECT 1600.410 16.760 1798.990 16.900 ;
        RECT 1600.410 16.700 1600.730 16.760 ;
        RECT 1798.670 16.700 1798.990 16.760 ;
      LAYER via ;
        RECT 1597.220 586.540 1597.480 586.800 ;
        RECT 1600.440 586.540 1600.700 586.800 ;
        RECT 1600.440 16.700 1600.700 16.960 ;
        RECT 1798.700 16.700 1798.960 16.960 ;
      LAYER met2 ;
        RECT 1595.610 600.170 1595.890 604.000 ;
        RECT 1595.610 600.030 1597.420 600.170 ;
        RECT 1595.610 600.000 1595.890 600.030 ;
        RECT 1597.280 586.830 1597.420 600.030 ;
        RECT 1597.220 586.510 1597.480 586.830 ;
        RECT 1600.440 586.510 1600.700 586.830 ;
        RECT 1600.500 16.990 1600.640 586.510 ;
        RECT 1600.440 16.670 1600.700 16.990 ;
        RECT 1798.700 16.670 1798.960 16.990 ;
        RECT 1798.760 2.400 1798.900 16.670 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 20.640 1607.630 20.700 ;
        RECT 1769.690 20.640 1770.010 20.700 ;
        RECT 1607.310 20.500 1770.010 20.640 ;
        RECT 1607.310 20.440 1607.630 20.500 ;
        RECT 1769.690 20.440 1770.010 20.500 ;
        RECT 1770.610 19.960 1770.930 20.020 ;
        RECT 1816.610 19.960 1816.930 20.020 ;
        RECT 1770.610 19.820 1816.930 19.960 ;
        RECT 1770.610 19.760 1770.930 19.820 ;
        RECT 1816.610 19.760 1816.930 19.820 ;
      LAYER via ;
        RECT 1607.340 20.440 1607.600 20.700 ;
        RECT 1769.720 20.440 1769.980 20.700 ;
        RECT 1770.640 19.760 1770.900 20.020 ;
        RECT 1816.640 19.760 1816.900 20.020 ;
      LAYER met2 ;
        RECT 1604.810 600.170 1605.090 604.000 ;
        RECT 1604.810 600.030 1607.540 600.170 ;
        RECT 1604.810 600.000 1605.090 600.030 ;
        RECT 1607.400 20.730 1607.540 600.030 ;
        RECT 1769.780 20.730 1770.840 20.810 ;
        RECT 1607.340 20.410 1607.600 20.730 ;
        RECT 1769.720 20.670 1770.840 20.730 ;
        RECT 1769.720 20.410 1769.980 20.670 ;
        RECT 1770.700 20.050 1770.840 20.670 ;
        RECT 1770.640 19.730 1770.900 20.050 ;
        RECT 1816.640 19.730 1816.900 20.050 ;
        RECT 1816.700 2.400 1816.840 19.730 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1614.210 19.960 1614.530 20.020 ;
        RECT 1770.150 19.960 1770.470 20.020 ;
        RECT 1614.210 19.820 1770.470 19.960 ;
        RECT 1614.210 19.760 1614.530 19.820 ;
        RECT 1770.150 19.760 1770.470 19.820 ;
        RECT 1770.150 17.920 1770.470 17.980 ;
        RECT 1834.550 17.920 1834.870 17.980 ;
        RECT 1770.150 17.780 1834.870 17.920 ;
        RECT 1770.150 17.720 1770.470 17.780 ;
        RECT 1834.550 17.720 1834.870 17.780 ;
      LAYER via ;
        RECT 1614.240 19.760 1614.500 20.020 ;
        RECT 1770.180 19.760 1770.440 20.020 ;
        RECT 1770.180 17.720 1770.440 17.980 ;
        RECT 1834.580 17.720 1834.840 17.980 ;
      LAYER met2 ;
        RECT 1614.010 600.000 1614.290 604.000 ;
        RECT 1614.070 598.810 1614.210 600.000 ;
        RECT 1614.070 598.670 1614.440 598.810 ;
        RECT 1614.300 20.050 1614.440 598.670 ;
        RECT 1614.240 19.730 1614.500 20.050 ;
        RECT 1770.180 19.730 1770.440 20.050 ;
        RECT 1770.240 18.010 1770.380 19.730 ;
        RECT 1770.180 17.690 1770.440 18.010 ;
        RECT 1834.580 17.690 1834.840 18.010 ;
        RECT 1834.640 2.400 1834.780 17.690 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1624.790 587.420 1625.110 587.480 ;
        RECT 1631.690 587.420 1632.010 587.480 ;
        RECT 1624.790 587.280 1632.010 587.420 ;
        RECT 1624.790 587.220 1625.110 587.280 ;
        RECT 1631.690 587.220 1632.010 587.280 ;
        RECT 1631.690 19.620 1632.010 19.680 ;
        RECT 1852.030 19.620 1852.350 19.680 ;
        RECT 1631.690 19.480 1852.350 19.620 ;
        RECT 1631.690 19.420 1632.010 19.480 ;
        RECT 1852.030 19.420 1852.350 19.480 ;
      LAYER via ;
        RECT 1624.820 587.220 1625.080 587.480 ;
        RECT 1631.720 587.220 1631.980 587.480 ;
        RECT 1631.720 19.420 1631.980 19.680 ;
        RECT 1852.060 19.420 1852.320 19.680 ;
      LAYER met2 ;
        RECT 1623.210 600.170 1623.490 604.000 ;
        RECT 1623.210 600.030 1625.020 600.170 ;
        RECT 1623.210 600.000 1623.490 600.030 ;
        RECT 1624.880 587.510 1625.020 600.030 ;
        RECT 1624.820 587.190 1625.080 587.510 ;
        RECT 1631.720 587.190 1631.980 587.510 ;
        RECT 1631.780 19.710 1631.920 587.190 ;
        RECT 1631.720 19.390 1631.980 19.710 ;
        RECT 1852.060 19.390 1852.320 19.710 ;
        RECT 1852.120 2.400 1852.260 19.390 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1634.450 33.900 1634.770 33.960 ;
        RECT 1869.970 33.900 1870.290 33.960 ;
        RECT 1634.450 33.760 1870.290 33.900 ;
        RECT 1634.450 33.700 1634.770 33.760 ;
        RECT 1869.970 33.700 1870.290 33.760 ;
      LAYER via ;
        RECT 1634.480 33.700 1634.740 33.960 ;
        RECT 1870.000 33.700 1870.260 33.960 ;
      LAYER met2 ;
        RECT 1632.410 600.170 1632.690 604.000 ;
        RECT 1632.410 600.030 1634.680 600.170 ;
        RECT 1632.410 600.000 1632.690 600.030 ;
        RECT 1634.540 33.990 1634.680 600.030 ;
        RECT 1634.480 33.670 1634.740 33.990 ;
        RECT 1870.000 33.670 1870.260 33.990 ;
        RECT 1870.060 2.400 1870.200 33.670 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1049.330 569.400 1049.650 569.460 ;
        RECT 1052.090 569.400 1052.410 569.460 ;
        RECT 1049.330 569.260 1052.410 569.400 ;
        RECT 1049.330 569.200 1049.650 569.260 ;
        RECT 1052.090 569.200 1052.410 569.260 ;
        RECT 746.190 24.720 746.510 24.780 ;
        RECT 1049.330 24.720 1049.650 24.780 ;
        RECT 746.190 24.580 1049.650 24.720 ;
        RECT 746.190 24.520 746.510 24.580 ;
        RECT 1049.330 24.520 1049.650 24.580 ;
      LAYER via ;
        RECT 1049.360 569.200 1049.620 569.460 ;
        RECT 1052.120 569.200 1052.380 569.460 ;
        RECT 746.220 24.520 746.480 24.780 ;
        RECT 1049.360 24.520 1049.620 24.780 ;
      LAYER met2 ;
        RECT 1053.730 600.170 1054.010 604.000 ;
        RECT 1052.180 600.030 1054.010 600.170 ;
        RECT 1052.180 569.490 1052.320 600.030 ;
        RECT 1053.730 600.000 1054.010 600.030 ;
        RECT 1049.360 569.170 1049.620 569.490 ;
        RECT 1052.120 569.170 1052.380 569.490 ;
        RECT 1049.420 24.810 1049.560 569.170 ;
        RECT 746.220 24.490 746.480 24.810 ;
        RECT 1049.360 24.490 1049.620 24.810 ;
        RECT 746.280 2.400 746.420 24.490 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1640.890 33.560 1641.210 33.620 ;
        RECT 1887.910 33.560 1888.230 33.620 ;
        RECT 1640.890 33.420 1888.230 33.560 ;
        RECT 1640.890 33.360 1641.210 33.420 ;
        RECT 1887.910 33.360 1888.230 33.420 ;
      LAYER via ;
        RECT 1640.920 33.360 1641.180 33.620 ;
        RECT 1887.940 33.360 1888.200 33.620 ;
      LAYER met2 ;
        RECT 1641.610 600.170 1641.890 604.000 ;
        RECT 1640.980 600.030 1641.890 600.170 ;
        RECT 1640.980 33.650 1641.120 600.030 ;
        RECT 1641.610 600.000 1641.890 600.030 ;
        RECT 1640.920 33.330 1641.180 33.650 ;
        RECT 1887.940 33.330 1888.200 33.650 ;
        RECT 1888.000 2.400 1888.140 33.330 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1652.390 586.740 1652.710 586.800 ;
        RECT 1655.150 586.740 1655.470 586.800 ;
        RECT 1652.390 586.600 1655.470 586.740 ;
        RECT 1652.390 586.540 1652.710 586.600 ;
        RECT 1655.150 586.540 1655.470 586.600 ;
        RECT 1655.150 33.220 1655.470 33.280 ;
        RECT 1905.850 33.220 1906.170 33.280 ;
        RECT 1655.150 33.080 1906.170 33.220 ;
        RECT 1655.150 33.020 1655.470 33.080 ;
        RECT 1905.850 33.020 1906.170 33.080 ;
      LAYER via ;
        RECT 1652.420 586.540 1652.680 586.800 ;
        RECT 1655.180 586.540 1655.440 586.800 ;
        RECT 1655.180 33.020 1655.440 33.280 ;
        RECT 1905.880 33.020 1906.140 33.280 ;
      LAYER met2 ;
        RECT 1650.810 600.170 1651.090 604.000 ;
        RECT 1650.810 600.030 1652.620 600.170 ;
        RECT 1650.810 600.000 1651.090 600.030 ;
        RECT 1652.480 586.830 1652.620 600.030 ;
        RECT 1652.420 586.510 1652.680 586.830 ;
        RECT 1655.180 586.510 1655.440 586.830 ;
        RECT 1655.240 33.310 1655.380 586.510 ;
        RECT 1655.180 32.990 1655.440 33.310 ;
        RECT 1905.880 32.990 1906.140 33.310 ;
        RECT 1905.940 2.400 1906.080 32.990 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.050 32.880 1662.370 32.940 ;
        RECT 1923.330 32.880 1923.650 32.940 ;
        RECT 1662.050 32.740 1923.650 32.880 ;
        RECT 1662.050 32.680 1662.370 32.740 ;
        RECT 1923.330 32.680 1923.650 32.740 ;
      LAYER via ;
        RECT 1662.080 32.680 1662.340 32.940 ;
        RECT 1923.360 32.680 1923.620 32.940 ;
      LAYER met2 ;
        RECT 1660.010 600.170 1660.290 604.000 ;
        RECT 1660.010 600.030 1662.280 600.170 ;
        RECT 1660.010 600.000 1660.290 600.030 ;
        RECT 1662.140 32.970 1662.280 600.030 ;
        RECT 1662.080 32.650 1662.340 32.970 ;
        RECT 1923.360 32.650 1923.620 32.970 ;
        RECT 1923.420 2.400 1923.560 32.650 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1668.490 32.200 1668.810 32.260 ;
        RECT 1941.270 32.200 1941.590 32.260 ;
        RECT 1668.490 32.060 1941.590 32.200 ;
        RECT 1668.490 32.000 1668.810 32.060 ;
        RECT 1941.270 32.000 1941.590 32.060 ;
      LAYER via ;
        RECT 1668.520 32.000 1668.780 32.260 ;
        RECT 1941.300 32.000 1941.560 32.260 ;
      LAYER met2 ;
        RECT 1669.210 600.170 1669.490 604.000 ;
        RECT 1668.580 600.030 1669.490 600.170 ;
        RECT 1668.580 32.290 1668.720 600.030 ;
        RECT 1669.210 600.000 1669.490 600.030 ;
        RECT 1668.520 31.970 1668.780 32.290 ;
        RECT 1941.300 31.970 1941.560 32.290 ;
        RECT 1941.360 2.400 1941.500 31.970 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1679.990 586.740 1680.310 586.800 ;
        RECT 1683.210 586.740 1683.530 586.800 ;
        RECT 1679.990 586.600 1683.530 586.740 ;
        RECT 1679.990 586.540 1680.310 586.600 ;
        RECT 1683.210 586.540 1683.530 586.600 ;
        RECT 1683.210 32.540 1683.530 32.600 ;
        RECT 1959.210 32.540 1959.530 32.600 ;
        RECT 1683.210 32.400 1959.530 32.540 ;
        RECT 1683.210 32.340 1683.530 32.400 ;
        RECT 1959.210 32.340 1959.530 32.400 ;
      LAYER via ;
        RECT 1680.020 586.540 1680.280 586.800 ;
        RECT 1683.240 586.540 1683.500 586.800 ;
        RECT 1683.240 32.340 1683.500 32.600 ;
        RECT 1959.240 32.340 1959.500 32.600 ;
      LAYER met2 ;
        RECT 1678.410 600.170 1678.690 604.000 ;
        RECT 1678.410 600.030 1680.220 600.170 ;
        RECT 1678.410 600.000 1678.690 600.030 ;
        RECT 1680.080 586.830 1680.220 600.030 ;
        RECT 1680.020 586.510 1680.280 586.830 ;
        RECT 1683.240 586.510 1683.500 586.830 ;
        RECT 1683.300 32.630 1683.440 586.510 ;
        RECT 1683.240 32.310 1683.500 32.630 ;
        RECT 1959.240 32.310 1959.500 32.630 ;
        RECT 1959.300 2.400 1959.440 32.310 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1689.650 31.860 1689.970 31.920 ;
        RECT 1977.150 31.860 1977.470 31.920 ;
        RECT 1689.650 31.720 1977.470 31.860 ;
        RECT 1689.650 31.660 1689.970 31.720 ;
        RECT 1977.150 31.660 1977.470 31.720 ;
      LAYER via ;
        RECT 1689.680 31.660 1689.940 31.920 ;
        RECT 1977.180 31.660 1977.440 31.920 ;
      LAYER met2 ;
        RECT 1687.610 600.170 1687.890 604.000 ;
        RECT 1687.610 600.030 1689.880 600.170 ;
        RECT 1687.610 600.000 1687.890 600.030 ;
        RECT 1689.740 31.950 1689.880 600.030 ;
        RECT 1689.680 31.630 1689.940 31.950 ;
        RECT 1977.180 31.630 1977.440 31.950 ;
        RECT 1977.240 2.400 1977.380 31.630 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1696.550 31.180 1696.870 31.240 ;
        RECT 1995.090 31.180 1995.410 31.240 ;
        RECT 1696.550 31.040 1995.410 31.180 ;
        RECT 1696.550 30.980 1696.870 31.040 ;
        RECT 1995.090 30.980 1995.410 31.040 ;
      LAYER via ;
        RECT 1696.580 30.980 1696.840 31.240 ;
        RECT 1995.120 30.980 1995.380 31.240 ;
      LAYER met2 ;
        RECT 1696.810 600.000 1697.090 604.000 ;
        RECT 1696.870 598.810 1697.010 600.000 ;
        RECT 1696.640 598.670 1697.010 598.810 ;
        RECT 1696.640 31.270 1696.780 598.670 ;
        RECT 1696.580 30.950 1696.840 31.270 ;
        RECT 1995.120 30.950 1995.380 31.270 ;
        RECT 1995.180 2.400 1995.320 30.950 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1707.590 586.740 1707.910 586.800 ;
        RECT 1710.810 586.740 1711.130 586.800 ;
        RECT 1707.590 586.600 1711.130 586.740 ;
        RECT 1707.590 586.540 1707.910 586.600 ;
        RECT 1710.810 586.540 1711.130 586.600 ;
        RECT 1710.810 31.520 1711.130 31.580 ;
        RECT 2012.570 31.520 2012.890 31.580 ;
        RECT 1710.810 31.380 2012.890 31.520 ;
        RECT 1710.810 31.320 1711.130 31.380 ;
        RECT 2012.570 31.320 2012.890 31.380 ;
      LAYER via ;
        RECT 1707.620 586.540 1707.880 586.800 ;
        RECT 1710.840 586.540 1711.100 586.800 ;
        RECT 1710.840 31.320 1711.100 31.580 ;
        RECT 2012.600 31.320 2012.860 31.580 ;
      LAYER met2 ;
        RECT 1706.010 600.170 1706.290 604.000 ;
        RECT 1706.010 600.030 1707.820 600.170 ;
        RECT 1706.010 600.000 1706.290 600.030 ;
        RECT 1707.680 586.830 1707.820 600.030 ;
        RECT 1707.620 586.510 1707.880 586.830 ;
        RECT 1710.840 586.510 1711.100 586.830 ;
        RECT 1710.900 31.610 1711.040 586.510 ;
        RECT 1710.840 31.290 1711.100 31.610 ;
        RECT 2012.600 31.290 2012.860 31.610 ;
        RECT 2012.660 2.400 2012.800 31.290 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1717.250 30.840 1717.570 30.900 ;
        RECT 2030.510 30.840 2030.830 30.900 ;
        RECT 1717.250 30.700 2030.830 30.840 ;
        RECT 1717.250 30.640 1717.570 30.700 ;
        RECT 2030.510 30.640 2030.830 30.700 ;
      LAYER via ;
        RECT 1717.280 30.640 1717.540 30.900 ;
        RECT 2030.540 30.640 2030.800 30.900 ;
      LAYER met2 ;
        RECT 1715.210 600.170 1715.490 604.000 ;
        RECT 1715.210 600.030 1717.480 600.170 ;
        RECT 1715.210 600.000 1715.490 600.030 ;
        RECT 1717.340 30.930 1717.480 600.030 ;
        RECT 1717.280 30.610 1717.540 30.930 ;
        RECT 2030.540 30.610 2030.800 30.930 ;
        RECT 2030.600 2.400 2030.740 30.610 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1723.690 38.660 1724.010 38.720 ;
        RECT 2048.450 38.660 2048.770 38.720 ;
        RECT 1723.690 38.520 2048.770 38.660 ;
        RECT 1723.690 38.460 1724.010 38.520 ;
        RECT 2048.450 38.460 2048.770 38.520 ;
      LAYER via ;
        RECT 1723.720 38.460 1723.980 38.720 ;
        RECT 2048.480 38.460 2048.740 38.720 ;
      LAYER met2 ;
        RECT 1724.410 600.170 1724.690 604.000 ;
        RECT 1723.780 600.030 1724.690 600.170 ;
        RECT 1723.780 38.750 1723.920 600.030 ;
        RECT 1724.410 600.000 1724.690 600.030 ;
        RECT 1723.720 38.430 1723.980 38.750 ;
        RECT 2048.480 38.430 2048.740 38.750 ;
        RECT 2048.540 2.400 2048.680 38.430 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 763.670 25.060 763.990 25.120 ;
        RECT 1063.130 25.060 1063.450 25.120 ;
        RECT 763.670 24.920 1063.450 25.060 ;
        RECT 763.670 24.860 763.990 24.920 ;
        RECT 1063.130 24.860 1063.450 24.920 ;
      LAYER via ;
        RECT 763.700 24.860 763.960 25.120 ;
        RECT 1063.160 24.860 1063.420 25.120 ;
      LAYER met2 ;
        RECT 1062.930 600.000 1063.210 604.000 ;
        RECT 1062.990 598.810 1063.130 600.000 ;
        RECT 1062.990 598.670 1063.360 598.810 ;
        RECT 1063.220 25.150 1063.360 598.670 ;
        RECT 763.700 24.830 763.960 25.150 ;
        RECT 1063.160 24.830 1063.420 25.150 ;
        RECT 763.760 2.400 763.900 24.830 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1735.190 586.740 1735.510 586.800 ;
        RECT 1738.410 586.740 1738.730 586.800 ;
        RECT 1735.190 586.600 1738.730 586.740 ;
        RECT 1735.190 586.540 1735.510 586.600 ;
        RECT 1738.410 586.540 1738.730 586.600 ;
        RECT 1738.410 38.320 1738.730 38.380 ;
        RECT 2066.390 38.320 2066.710 38.380 ;
        RECT 1738.410 38.180 2066.710 38.320 ;
        RECT 1738.410 38.120 1738.730 38.180 ;
        RECT 2066.390 38.120 2066.710 38.180 ;
      LAYER via ;
        RECT 1735.220 586.540 1735.480 586.800 ;
        RECT 1738.440 586.540 1738.700 586.800 ;
        RECT 1738.440 38.120 1738.700 38.380 ;
        RECT 2066.420 38.120 2066.680 38.380 ;
      LAYER met2 ;
        RECT 1733.610 600.170 1733.890 604.000 ;
        RECT 1733.610 600.030 1735.420 600.170 ;
        RECT 1733.610 600.000 1733.890 600.030 ;
        RECT 1735.280 586.830 1735.420 600.030 ;
        RECT 1735.220 586.510 1735.480 586.830 ;
        RECT 1738.440 586.510 1738.700 586.830 ;
        RECT 1738.500 38.410 1738.640 586.510 ;
        RECT 1738.440 38.090 1738.700 38.410 ;
        RECT 2066.420 38.090 2066.680 38.410 ;
        RECT 2066.480 2.400 2066.620 38.090 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1744.850 37.980 1745.170 38.040 ;
        RECT 2063.170 37.980 2063.490 38.040 ;
        RECT 1744.850 37.840 2063.490 37.980 ;
        RECT 1744.850 37.780 1745.170 37.840 ;
        RECT 2063.170 37.780 2063.490 37.840 ;
        RECT 2063.170 35.260 2063.490 35.320 ;
        RECT 2084.330 35.260 2084.650 35.320 ;
        RECT 2063.170 35.120 2084.650 35.260 ;
        RECT 2063.170 35.060 2063.490 35.120 ;
        RECT 2084.330 35.060 2084.650 35.120 ;
      LAYER via ;
        RECT 1744.880 37.780 1745.140 38.040 ;
        RECT 2063.200 37.780 2063.460 38.040 ;
        RECT 2063.200 35.060 2063.460 35.320 ;
        RECT 2084.360 35.060 2084.620 35.320 ;
      LAYER met2 ;
        RECT 1742.810 600.170 1743.090 604.000 ;
        RECT 1742.810 600.030 1745.080 600.170 ;
        RECT 1742.810 600.000 1743.090 600.030 ;
        RECT 1744.940 38.070 1745.080 600.030 ;
        RECT 1744.880 37.750 1745.140 38.070 ;
        RECT 2063.200 37.750 2063.460 38.070 ;
        RECT 2063.260 35.350 2063.400 37.750 ;
        RECT 2063.200 35.030 2063.460 35.350 ;
        RECT 2084.360 35.030 2084.620 35.350 ;
        RECT 2084.420 2.400 2084.560 35.030 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1751.750 45.800 1752.070 45.860 ;
        RECT 2101.810 45.800 2102.130 45.860 ;
        RECT 1751.750 45.660 2102.130 45.800 ;
        RECT 1751.750 45.600 1752.070 45.660 ;
        RECT 2101.810 45.600 2102.130 45.660 ;
      LAYER via ;
        RECT 1751.780 45.600 1752.040 45.860 ;
        RECT 2101.840 45.600 2102.100 45.860 ;
      LAYER met2 ;
        RECT 1752.010 600.000 1752.290 604.000 ;
        RECT 1752.070 598.810 1752.210 600.000 ;
        RECT 1751.840 598.670 1752.210 598.810 ;
        RECT 1751.840 45.890 1751.980 598.670 ;
        RECT 1751.780 45.570 1752.040 45.890 ;
        RECT 2101.840 45.570 2102.100 45.890 ;
        RECT 2101.900 2.400 2102.040 45.570 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1762.790 592.860 1763.110 592.920 ;
        RECT 1766.010 592.860 1766.330 592.920 ;
        RECT 1762.790 592.720 1766.330 592.860 ;
        RECT 1762.790 592.660 1763.110 592.720 ;
        RECT 1766.010 592.660 1766.330 592.720 ;
        RECT 1766.010 45.460 1766.330 45.520 ;
        RECT 2119.750 45.460 2120.070 45.520 ;
        RECT 1766.010 45.320 2120.070 45.460 ;
        RECT 1766.010 45.260 1766.330 45.320 ;
        RECT 2119.750 45.260 2120.070 45.320 ;
      LAYER via ;
        RECT 1762.820 592.660 1763.080 592.920 ;
        RECT 1766.040 592.660 1766.300 592.920 ;
        RECT 1766.040 45.260 1766.300 45.520 ;
        RECT 2119.780 45.260 2120.040 45.520 ;
      LAYER met2 ;
        RECT 1761.210 600.170 1761.490 604.000 ;
        RECT 1761.210 600.030 1763.020 600.170 ;
        RECT 1761.210 600.000 1761.490 600.030 ;
        RECT 1762.880 592.950 1763.020 600.030 ;
        RECT 1762.820 592.630 1763.080 592.950 ;
        RECT 1766.040 592.630 1766.300 592.950 ;
        RECT 1766.100 45.550 1766.240 592.630 ;
        RECT 1766.040 45.230 1766.300 45.550 ;
        RECT 2119.780 45.230 2120.040 45.550 ;
        RECT 2119.840 2.400 2119.980 45.230 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.450 45.120 1772.770 45.180 ;
        RECT 2137.690 45.120 2138.010 45.180 ;
        RECT 1772.450 44.980 2138.010 45.120 ;
        RECT 1772.450 44.920 1772.770 44.980 ;
        RECT 2137.690 44.920 2138.010 44.980 ;
      LAYER via ;
        RECT 1772.480 44.920 1772.740 45.180 ;
        RECT 2137.720 44.920 2137.980 45.180 ;
      LAYER met2 ;
        RECT 1770.410 600.170 1770.690 604.000 ;
        RECT 1770.410 600.030 1772.680 600.170 ;
        RECT 1770.410 600.000 1770.690 600.030 ;
        RECT 1772.540 45.210 1772.680 600.030 ;
        RECT 1772.480 44.890 1772.740 45.210 ;
        RECT 2137.720 44.890 2137.980 45.210 ;
        RECT 2137.780 2.400 2137.920 44.890 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.350 44.780 1779.670 44.840 ;
        RECT 2155.630 44.780 2155.950 44.840 ;
        RECT 1779.350 44.640 2155.950 44.780 ;
        RECT 1779.350 44.580 1779.670 44.640 ;
        RECT 2155.630 44.580 2155.950 44.640 ;
      LAYER via ;
        RECT 1779.380 44.580 1779.640 44.840 ;
        RECT 2155.660 44.580 2155.920 44.840 ;
      LAYER met2 ;
        RECT 1779.610 600.000 1779.890 604.000 ;
        RECT 1779.670 598.810 1779.810 600.000 ;
        RECT 1779.440 598.670 1779.810 598.810 ;
        RECT 1779.440 44.870 1779.580 598.670 ;
        RECT 1779.380 44.550 1779.640 44.870 ;
        RECT 2155.660 44.550 2155.920 44.870 ;
        RECT 2155.720 2.400 2155.860 44.550 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1790.390 587.760 1790.710 587.820 ;
        RECT 1793.150 587.760 1793.470 587.820 ;
        RECT 1790.390 587.620 1793.470 587.760 ;
        RECT 1790.390 587.560 1790.710 587.620 ;
        RECT 1793.150 587.560 1793.470 587.620 ;
        RECT 1793.150 42.400 1793.470 42.460 ;
        RECT 2173.110 42.400 2173.430 42.460 ;
        RECT 1793.150 42.260 2173.430 42.400 ;
        RECT 1793.150 42.200 1793.470 42.260 ;
        RECT 2173.110 42.200 2173.430 42.260 ;
      LAYER via ;
        RECT 1790.420 587.560 1790.680 587.820 ;
        RECT 1793.180 587.560 1793.440 587.820 ;
        RECT 1793.180 42.200 1793.440 42.460 ;
        RECT 2173.140 42.200 2173.400 42.460 ;
      LAYER met2 ;
        RECT 1788.810 600.170 1789.090 604.000 ;
        RECT 1788.810 600.030 1790.620 600.170 ;
        RECT 1788.810 600.000 1789.090 600.030 ;
        RECT 1790.480 587.850 1790.620 600.030 ;
        RECT 1790.420 587.530 1790.680 587.850 ;
        RECT 1793.180 587.530 1793.440 587.850 ;
        RECT 1793.240 42.490 1793.380 587.530 ;
        RECT 1793.180 42.170 1793.440 42.490 ;
        RECT 2173.140 42.170 2173.400 42.490 ;
        RECT 2173.200 2.400 2173.340 42.170 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.050 42.740 1800.370 42.800 ;
        RECT 2191.050 42.740 2191.370 42.800 ;
        RECT 1800.050 42.600 2191.370 42.740 ;
        RECT 1800.050 42.540 1800.370 42.600 ;
        RECT 2191.050 42.540 2191.370 42.600 ;
      LAYER via ;
        RECT 1800.080 42.540 1800.340 42.800 ;
        RECT 2191.080 42.540 2191.340 42.800 ;
      LAYER met2 ;
        RECT 1798.010 600.170 1798.290 604.000 ;
        RECT 1798.010 600.030 1800.280 600.170 ;
        RECT 1798.010 600.000 1798.290 600.030 ;
        RECT 1800.140 42.830 1800.280 600.030 ;
        RECT 1800.080 42.510 1800.340 42.830 ;
        RECT 2191.080 42.510 2191.340 42.830 ;
        RECT 2191.140 2.400 2191.280 42.510 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1806.950 43.420 1807.270 43.480 ;
        RECT 2208.990 43.420 2209.310 43.480 ;
        RECT 1806.950 43.280 2209.310 43.420 ;
        RECT 1806.950 43.220 1807.270 43.280 ;
        RECT 2208.990 43.220 2209.310 43.280 ;
      LAYER via ;
        RECT 1806.980 43.220 1807.240 43.480 ;
        RECT 2209.020 43.220 2209.280 43.480 ;
      LAYER met2 ;
        RECT 1807.210 600.000 1807.490 604.000 ;
        RECT 1807.270 598.810 1807.410 600.000 ;
        RECT 1807.040 598.670 1807.410 598.810 ;
        RECT 1807.040 43.510 1807.180 598.670 ;
        RECT 1806.980 43.190 1807.240 43.510 ;
        RECT 2209.020 43.190 2209.280 43.510 ;
        RECT 2209.080 2.400 2209.220 43.190 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1817.990 586.740 1818.310 586.800 ;
        RECT 1821.210 586.740 1821.530 586.800 ;
        RECT 1817.990 586.600 1821.530 586.740 ;
        RECT 1817.990 586.540 1818.310 586.600 ;
        RECT 1821.210 586.540 1821.530 586.600 ;
        RECT 1821.210 43.080 1821.530 43.140 ;
        RECT 2226.930 43.080 2227.250 43.140 ;
        RECT 1821.210 42.940 2227.250 43.080 ;
        RECT 1821.210 42.880 1821.530 42.940 ;
        RECT 2226.930 42.880 2227.250 42.940 ;
      LAYER via ;
        RECT 1818.020 586.540 1818.280 586.800 ;
        RECT 1821.240 586.540 1821.500 586.800 ;
        RECT 1821.240 42.880 1821.500 43.140 ;
        RECT 2226.960 42.880 2227.220 43.140 ;
      LAYER met2 ;
        RECT 1816.410 600.170 1816.690 604.000 ;
        RECT 1816.410 600.030 1818.220 600.170 ;
        RECT 1816.410 600.000 1816.690 600.030 ;
        RECT 1818.080 586.830 1818.220 600.030 ;
        RECT 1818.020 586.510 1818.280 586.830 ;
        RECT 1821.240 586.510 1821.500 586.830 ;
        RECT 1821.300 43.170 1821.440 586.510 ;
        RECT 1821.240 42.850 1821.500 43.170 ;
        RECT 2226.960 42.850 2227.220 43.170 ;
        RECT 2227.020 2.400 2227.160 42.850 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1070.030 22.000 1070.350 22.060 ;
        RECT 814.360 21.860 1070.350 22.000 ;
        RECT 781.610 20.640 781.930 20.700 ;
        RECT 814.360 20.640 814.500 21.860 ;
        RECT 1070.030 21.800 1070.350 21.860 ;
        RECT 781.610 20.500 814.500 20.640 ;
        RECT 781.610 20.440 781.930 20.500 ;
      LAYER via ;
        RECT 781.640 20.440 781.900 20.700 ;
        RECT 1070.060 21.800 1070.320 22.060 ;
      LAYER met2 ;
        RECT 1072.130 600.170 1072.410 604.000 ;
        RECT 1070.120 600.030 1072.410 600.170 ;
        RECT 1070.120 22.090 1070.260 600.030 ;
        RECT 1072.130 600.000 1072.410 600.030 ;
        RECT 1070.060 21.770 1070.320 22.090 ;
        RECT 781.640 20.410 781.900 20.730 ;
        RECT 781.700 2.400 781.840 20.410 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1827.650 43.760 1827.970 43.820 ;
        RECT 2244.870 43.760 2245.190 43.820 ;
        RECT 1827.650 43.620 2245.190 43.760 ;
        RECT 1827.650 43.560 1827.970 43.620 ;
        RECT 2244.870 43.560 2245.190 43.620 ;
      LAYER via ;
        RECT 1827.680 43.560 1827.940 43.820 ;
        RECT 2244.900 43.560 2245.160 43.820 ;
      LAYER met2 ;
        RECT 1825.150 600.170 1825.430 604.000 ;
        RECT 1825.150 600.030 1827.880 600.170 ;
        RECT 1825.150 600.000 1825.430 600.030 ;
        RECT 1827.740 43.850 1827.880 600.030 ;
        RECT 1827.680 43.530 1827.940 43.850 ;
        RECT 2244.900 43.530 2245.160 43.850 ;
        RECT 2244.960 2.400 2245.100 43.530 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1834.550 44.100 1834.870 44.160 ;
        RECT 2262.350 44.100 2262.670 44.160 ;
        RECT 1834.550 43.960 2262.670 44.100 ;
        RECT 1834.550 43.900 1834.870 43.960 ;
        RECT 2262.350 43.900 2262.670 43.960 ;
      LAYER via ;
        RECT 1834.580 43.900 1834.840 44.160 ;
        RECT 2262.380 43.900 2262.640 44.160 ;
      LAYER met2 ;
        RECT 1834.350 600.000 1834.630 604.000 ;
        RECT 1834.410 598.810 1834.550 600.000 ;
        RECT 1834.410 598.670 1834.780 598.810 ;
        RECT 1834.640 44.190 1834.780 598.670 ;
        RECT 1834.580 43.870 1834.840 44.190 ;
        RECT 2262.380 43.870 2262.640 44.190 ;
        RECT 2262.440 2.400 2262.580 43.870 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1845.130 586.740 1845.450 586.800 ;
        RECT 1848.810 586.740 1849.130 586.800 ;
        RECT 1845.130 586.600 1849.130 586.740 ;
        RECT 1845.130 586.540 1845.450 586.600 ;
        RECT 1848.810 586.540 1849.130 586.600 ;
        RECT 1848.810 44.440 1849.130 44.500 ;
        RECT 2280.290 44.440 2280.610 44.500 ;
        RECT 1848.810 44.300 2280.610 44.440 ;
        RECT 1848.810 44.240 1849.130 44.300 ;
        RECT 2280.290 44.240 2280.610 44.300 ;
      LAYER via ;
        RECT 1845.160 586.540 1845.420 586.800 ;
        RECT 1848.840 586.540 1849.100 586.800 ;
        RECT 1848.840 44.240 1849.100 44.500 ;
        RECT 2280.320 44.240 2280.580 44.500 ;
      LAYER met2 ;
        RECT 1843.550 600.170 1843.830 604.000 ;
        RECT 1843.550 600.030 1845.360 600.170 ;
        RECT 1843.550 600.000 1843.830 600.030 ;
        RECT 1845.220 586.830 1845.360 600.030 ;
        RECT 1845.160 586.510 1845.420 586.830 ;
        RECT 1848.840 586.510 1849.100 586.830 ;
        RECT 1848.900 44.530 1849.040 586.510 ;
        RECT 1848.840 44.210 1849.100 44.530 ;
        RECT 2280.320 44.210 2280.580 44.530 ;
        RECT 2280.380 2.400 2280.520 44.210 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.250 53.620 1855.570 53.680 ;
        RECT 2298.230 53.620 2298.550 53.680 ;
        RECT 1855.250 53.480 2298.550 53.620 ;
        RECT 1855.250 53.420 1855.570 53.480 ;
        RECT 2298.230 53.420 2298.550 53.480 ;
      LAYER via ;
        RECT 1855.280 53.420 1855.540 53.680 ;
        RECT 2298.260 53.420 2298.520 53.680 ;
      LAYER met2 ;
        RECT 1852.750 600.170 1853.030 604.000 ;
        RECT 1852.750 600.030 1855.480 600.170 ;
        RECT 1852.750 600.000 1853.030 600.030 ;
        RECT 1855.340 53.710 1855.480 600.030 ;
        RECT 1855.280 53.390 1855.540 53.710 ;
        RECT 2298.260 53.390 2298.520 53.710 ;
        RECT 2298.320 2.400 2298.460 53.390 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1861.690 53.280 1862.010 53.340 ;
        RECT 2316.170 53.280 2316.490 53.340 ;
        RECT 1861.690 53.140 2316.490 53.280 ;
        RECT 1861.690 53.080 1862.010 53.140 ;
        RECT 2316.170 53.080 2316.490 53.140 ;
      LAYER via ;
        RECT 1861.720 53.080 1861.980 53.340 ;
        RECT 2316.200 53.080 2316.460 53.340 ;
      LAYER met2 ;
        RECT 1861.950 600.000 1862.230 604.000 ;
        RECT 1862.010 598.810 1862.150 600.000 ;
        RECT 1861.780 598.670 1862.150 598.810 ;
        RECT 1861.780 53.370 1861.920 598.670 ;
        RECT 1861.720 53.050 1861.980 53.370 ;
        RECT 2316.200 53.050 2316.460 53.370 ;
        RECT 2316.260 2.400 2316.400 53.050 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1872.730 586.740 1873.050 586.800 ;
        RECT 1875.950 586.740 1876.270 586.800 ;
        RECT 1872.730 586.600 1876.270 586.740 ;
        RECT 1872.730 586.540 1873.050 586.600 ;
        RECT 1875.950 586.540 1876.270 586.600 ;
        RECT 1875.950 52.940 1876.270 53.000 ;
        RECT 2334.110 52.940 2334.430 53.000 ;
        RECT 1875.950 52.800 2334.430 52.940 ;
        RECT 1875.950 52.740 1876.270 52.800 ;
        RECT 2334.110 52.740 2334.430 52.800 ;
      LAYER via ;
        RECT 1872.760 586.540 1873.020 586.800 ;
        RECT 1875.980 586.540 1876.240 586.800 ;
        RECT 1875.980 52.740 1876.240 53.000 ;
        RECT 2334.140 52.740 2334.400 53.000 ;
      LAYER met2 ;
        RECT 1871.150 600.170 1871.430 604.000 ;
        RECT 1871.150 600.030 1872.960 600.170 ;
        RECT 1871.150 600.000 1871.430 600.030 ;
        RECT 1872.820 586.830 1872.960 600.030 ;
        RECT 1872.760 586.510 1873.020 586.830 ;
        RECT 1875.980 586.510 1876.240 586.830 ;
        RECT 1876.040 53.030 1876.180 586.510 ;
        RECT 1875.980 52.710 1876.240 53.030 ;
        RECT 2334.140 52.710 2334.400 53.030 ;
        RECT 2334.200 2.400 2334.340 52.710 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1882.850 52.600 1883.170 52.660 ;
        RECT 2351.590 52.600 2351.910 52.660 ;
        RECT 1882.850 52.460 2351.910 52.600 ;
        RECT 1882.850 52.400 1883.170 52.460 ;
        RECT 2351.590 52.400 2351.910 52.460 ;
      LAYER via ;
        RECT 1882.880 52.400 1883.140 52.660 ;
        RECT 2351.620 52.400 2351.880 52.660 ;
      LAYER met2 ;
        RECT 1880.350 600.170 1880.630 604.000 ;
        RECT 1880.350 600.030 1883.080 600.170 ;
        RECT 1880.350 600.000 1880.630 600.030 ;
        RECT 1882.940 52.690 1883.080 600.030 ;
        RECT 1882.880 52.370 1883.140 52.690 ;
        RECT 2351.620 52.370 2351.880 52.690 ;
        RECT 2351.680 2.400 2351.820 52.370 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1889.750 52.260 1890.070 52.320 ;
        RECT 2366.770 52.260 2367.090 52.320 ;
        RECT 1889.750 52.120 2367.090 52.260 ;
        RECT 1889.750 52.060 1890.070 52.120 ;
        RECT 2366.770 52.060 2367.090 52.120 ;
        RECT 2366.770 2.960 2367.090 3.020 ;
        RECT 2369.530 2.960 2369.850 3.020 ;
        RECT 2366.770 2.820 2369.850 2.960 ;
        RECT 2366.770 2.760 2367.090 2.820 ;
        RECT 2369.530 2.760 2369.850 2.820 ;
      LAYER via ;
        RECT 1889.780 52.060 1890.040 52.320 ;
        RECT 2366.800 52.060 2367.060 52.320 ;
        RECT 2366.800 2.760 2367.060 3.020 ;
        RECT 2369.560 2.760 2369.820 3.020 ;
      LAYER met2 ;
        RECT 1889.550 600.000 1889.830 604.000 ;
        RECT 1889.610 598.810 1889.750 600.000 ;
        RECT 1889.610 598.670 1889.980 598.810 ;
        RECT 1889.840 52.350 1889.980 598.670 ;
        RECT 1889.780 52.030 1890.040 52.350 ;
        RECT 2366.800 52.030 2367.060 52.350 ;
        RECT 2366.860 3.050 2367.000 52.030 ;
        RECT 2366.800 2.730 2367.060 3.050 ;
        RECT 2369.560 2.730 2369.820 3.050 ;
        RECT 2369.620 2.400 2369.760 2.730 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1900.330 586.740 1900.650 586.800 ;
        RECT 1904.010 586.740 1904.330 586.800 ;
        RECT 1900.330 586.600 1904.330 586.740 ;
        RECT 1900.330 586.540 1900.650 586.600 ;
        RECT 1904.010 586.540 1904.330 586.600 ;
        RECT 1904.010 51.920 1904.330 51.980 ;
        RECT 2388.390 51.920 2388.710 51.980 ;
        RECT 1904.010 51.780 2388.710 51.920 ;
        RECT 1904.010 51.720 1904.330 51.780 ;
        RECT 2388.390 51.720 2388.710 51.780 ;
      LAYER via ;
        RECT 1900.360 586.540 1900.620 586.800 ;
        RECT 1904.040 586.540 1904.300 586.800 ;
        RECT 1904.040 51.720 1904.300 51.980 ;
        RECT 2388.420 51.720 2388.680 51.980 ;
      LAYER met2 ;
        RECT 1898.750 600.170 1899.030 604.000 ;
        RECT 1898.750 600.030 1900.560 600.170 ;
        RECT 1898.750 600.000 1899.030 600.030 ;
        RECT 1900.420 586.830 1900.560 600.030 ;
        RECT 1900.360 586.510 1900.620 586.830 ;
        RECT 1904.040 586.510 1904.300 586.830 ;
        RECT 1904.100 52.010 1904.240 586.510 ;
        RECT 1904.040 51.690 1904.300 52.010 ;
        RECT 2388.420 51.690 2388.680 52.010 ;
        RECT 2388.480 37.130 2388.620 51.690 ;
        RECT 2387.560 36.990 2388.620 37.130 ;
        RECT 2387.560 2.400 2387.700 36.990 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1910.450 51.580 1910.770 51.640 ;
        RECT 2405.410 51.580 2405.730 51.640 ;
        RECT 1910.450 51.440 2405.730 51.580 ;
        RECT 1910.450 51.380 1910.770 51.440 ;
        RECT 2405.410 51.380 2405.730 51.440 ;
      LAYER via ;
        RECT 1910.480 51.380 1910.740 51.640 ;
        RECT 2405.440 51.380 2405.700 51.640 ;
      LAYER met2 ;
        RECT 1907.950 600.170 1908.230 604.000 ;
        RECT 1907.950 600.030 1910.680 600.170 ;
        RECT 1907.950 600.000 1908.230 600.030 ;
        RECT 1910.540 51.670 1910.680 600.030 ;
        RECT 1910.480 51.350 1910.740 51.670 ;
        RECT 2405.440 51.350 2405.700 51.670 ;
        RECT 2405.500 2.400 2405.640 51.350 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1076.010 579.600 1076.330 579.660 ;
        RECT 1076.930 579.600 1077.250 579.660 ;
        RECT 1076.010 579.460 1077.250 579.600 ;
        RECT 1076.010 579.400 1076.330 579.460 ;
        RECT 1076.930 579.400 1077.250 579.460 ;
        RECT 1076.010 531.660 1076.330 531.720 ;
        RECT 1076.930 531.660 1077.250 531.720 ;
        RECT 1076.010 531.520 1077.250 531.660 ;
        RECT 1076.010 531.460 1076.330 531.520 ;
        RECT 1076.930 531.460 1077.250 531.520 ;
        RECT 1076.930 524.180 1077.250 524.240 ;
        RECT 1077.850 524.180 1078.170 524.240 ;
        RECT 1076.930 524.040 1078.170 524.180 ;
        RECT 1076.930 523.980 1077.250 524.040 ;
        RECT 1077.850 523.980 1078.170 524.040 ;
        RECT 1076.930 476.240 1077.250 476.300 ;
        RECT 1077.850 476.240 1078.170 476.300 ;
        RECT 1076.930 476.100 1078.170 476.240 ;
        RECT 1076.930 476.040 1077.250 476.100 ;
        RECT 1077.850 476.040 1078.170 476.100 ;
        RECT 1076.930 427.620 1077.250 427.680 ;
        RECT 1077.850 427.620 1078.170 427.680 ;
        RECT 1076.930 427.480 1078.170 427.620 ;
        RECT 1076.930 427.420 1077.250 427.480 ;
        RECT 1077.850 427.420 1078.170 427.480 ;
        RECT 1076.930 379.680 1077.250 379.740 ;
        RECT 1077.850 379.680 1078.170 379.740 ;
        RECT 1076.930 379.540 1078.170 379.680 ;
        RECT 1076.930 379.480 1077.250 379.540 ;
        RECT 1077.850 379.480 1078.170 379.540 ;
        RECT 1076.930 331.060 1077.250 331.120 ;
        RECT 1077.850 331.060 1078.170 331.120 ;
        RECT 1076.930 330.920 1078.170 331.060 ;
        RECT 1076.930 330.860 1077.250 330.920 ;
        RECT 1077.850 330.860 1078.170 330.920 ;
        RECT 1076.930 241.980 1077.250 242.040 ;
        RECT 1077.850 241.980 1078.170 242.040 ;
        RECT 1076.930 241.840 1078.170 241.980 ;
        RECT 1076.930 241.780 1077.250 241.840 ;
        RECT 1077.850 241.780 1078.170 241.840 ;
        RECT 1076.930 234.500 1077.250 234.560 ;
        RECT 1077.850 234.500 1078.170 234.560 ;
        RECT 1076.930 234.360 1078.170 234.500 ;
        RECT 1076.930 234.300 1077.250 234.360 ;
        RECT 1077.850 234.300 1078.170 234.360 ;
        RECT 1076.930 145.420 1077.250 145.480 ;
        RECT 1077.850 145.420 1078.170 145.480 ;
        RECT 1076.930 145.280 1078.170 145.420 ;
        RECT 1076.930 145.220 1077.250 145.280 ;
        RECT 1077.850 145.220 1078.170 145.280 ;
        RECT 1075.090 137.940 1075.410 138.000 ;
        RECT 1076.930 137.940 1077.250 138.000 ;
        RECT 1075.090 137.800 1077.250 137.940 ;
        RECT 1075.090 137.740 1075.410 137.800 ;
        RECT 1076.930 137.740 1077.250 137.800 ;
        RECT 1075.090 90.000 1075.410 90.060 ;
        RECT 1076.010 90.000 1076.330 90.060 ;
        RECT 1075.090 89.860 1076.330 90.000 ;
        RECT 1075.090 89.800 1075.410 89.860 ;
        RECT 1076.010 89.800 1076.330 89.860 ;
        RECT 1076.010 48.520 1076.330 48.580 ;
        RECT 1077.390 48.520 1077.710 48.580 ;
        RECT 1076.010 48.380 1077.710 48.520 ;
        RECT 1076.010 48.320 1076.330 48.380 ;
        RECT 1077.390 48.320 1077.710 48.380 ;
        RECT 828.070 21.660 828.390 21.720 ;
        RECT 1077.390 21.660 1077.710 21.720 ;
        RECT 828.070 21.520 1077.710 21.660 ;
        RECT 828.070 21.460 828.390 21.520 ;
        RECT 1077.390 21.460 1077.710 21.520 ;
        RECT 799.550 17.580 799.870 17.640 ;
        RECT 828.070 17.580 828.390 17.640 ;
        RECT 799.550 17.440 828.390 17.580 ;
        RECT 799.550 17.380 799.870 17.440 ;
        RECT 828.070 17.380 828.390 17.440 ;
      LAYER via ;
        RECT 1076.040 579.400 1076.300 579.660 ;
        RECT 1076.960 579.400 1077.220 579.660 ;
        RECT 1076.040 531.460 1076.300 531.720 ;
        RECT 1076.960 531.460 1077.220 531.720 ;
        RECT 1076.960 523.980 1077.220 524.240 ;
        RECT 1077.880 523.980 1078.140 524.240 ;
        RECT 1076.960 476.040 1077.220 476.300 ;
        RECT 1077.880 476.040 1078.140 476.300 ;
        RECT 1076.960 427.420 1077.220 427.680 ;
        RECT 1077.880 427.420 1078.140 427.680 ;
        RECT 1076.960 379.480 1077.220 379.740 ;
        RECT 1077.880 379.480 1078.140 379.740 ;
        RECT 1076.960 330.860 1077.220 331.120 ;
        RECT 1077.880 330.860 1078.140 331.120 ;
        RECT 1076.960 241.780 1077.220 242.040 ;
        RECT 1077.880 241.780 1078.140 242.040 ;
        RECT 1076.960 234.300 1077.220 234.560 ;
        RECT 1077.880 234.300 1078.140 234.560 ;
        RECT 1076.960 145.220 1077.220 145.480 ;
        RECT 1077.880 145.220 1078.140 145.480 ;
        RECT 1075.120 137.740 1075.380 138.000 ;
        RECT 1076.960 137.740 1077.220 138.000 ;
        RECT 1075.120 89.800 1075.380 90.060 ;
        RECT 1076.040 89.800 1076.300 90.060 ;
        RECT 1076.040 48.320 1076.300 48.580 ;
        RECT 1077.420 48.320 1077.680 48.580 ;
        RECT 828.100 21.460 828.360 21.720 ;
        RECT 1077.420 21.460 1077.680 21.720 ;
        RECT 799.580 17.380 799.840 17.640 ;
        RECT 828.100 17.380 828.360 17.640 ;
      LAYER met2 ;
        RECT 1081.330 600.850 1081.610 604.000 ;
        RECT 1079.320 600.710 1081.610 600.850 ;
        RECT 1079.320 596.770 1079.460 600.710 ;
        RECT 1081.330 600.000 1081.610 600.710 ;
        RECT 1077.020 596.630 1079.460 596.770 ;
        RECT 1077.020 579.690 1077.160 596.630 ;
        RECT 1076.040 579.370 1076.300 579.690 ;
        RECT 1076.960 579.370 1077.220 579.690 ;
        RECT 1076.100 531.750 1076.240 579.370 ;
        RECT 1076.040 531.430 1076.300 531.750 ;
        RECT 1076.960 531.430 1077.220 531.750 ;
        RECT 1077.020 524.270 1077.160 531.430 ;
        RECT 1076.960 523.950 1077.220 524.270 ;
        RECT 1077.880 523.950 1078.140 524.270 ;
        RECT 1077.940 476.330 1078.080 523.950 ;
        RECT 1076.960 476.010 1077.220 476.330 ;
        RECT 1077.880 476.010 1078.140 476.330 ;
        RECT 1077.020 427.710 1077.160 476.010 ;
        RECT 1076.960 427.390 1077.220 427.710 ;
        RECT 1077.880 427.390 1078.140 427.710 ;
        RECT 1077.940 379.770 1078.080 427.390 ;
        RECT 1076.960 379.450 1077.220 379.770 ;
        RECT 1077.880 379.450 1078.140 379.770 ;
        RECT 1077.020 331.150 1077.160 379.450 ;
        RECT 1076.960 330.830 1077.220 331.150 ;
        RECT 1077.880 330.830 1078.140 331.150 ;
        RECT 1077.940 242.070 1078.080 330.830 ;
        RECT 1076.960 241.750 1077.220 242.070 ;
        RECT 1077.880 241.750 1078.140 242.070 ;
        RECT 1077.020 234.590 1077.160 241.750 ;
        RECT 1076.960 234.270 1077.220 234.590 ;
        RECT 1077.880 234.270 1078.140 234.590 ;
        RECT 1077.940 145.510 1078.080 234.270 ;
        RECT 1076.960 145.190 1077.220 145.510 ;
        RECT 1077.880 145.190 1078.140 145.510 ;
        RECT 1077.020 138.030 1077.160 145.190 ;
        RECT 1075.120 137.710 1075.380 138.030 ;
        RECT 1076.960 137.710 1077.220 138.030 ;
        RECT 1075.180 90.090 1075.320 137.710 ;
        RECT 1075.120 89.770 1075.380 90.090 ;
        RECT 1076.040 89.770 1076.300 90.090 ;
        RECT 1076.100 48.610 1076.240 89.770 ;
        RECT 1076.040 48.290 1076.300 48.610 ;
        RECT 1077.420 48.290 1077.680 48.610 ;
        RECT 1077.480 21.750 1077.620 48.290 ;
        RECT 828.100 21.430 828.360 21.750 ;
        RECT 1077.420 21.430 1077.680 21.750 ;
        RECT 828.160 17.670 828.300 21.430 ;
        RECT 799.580 17.350 799.840 17.670 ;
        RECT 828.100 17.350 828.360 17.670 ;
        RECT 799.640 2.400 799.780 17.350 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 36.620 645.310 36.680 ;
        RECT 1001.030 36.620 1001.350 36.680 ;
        RECT 644.990 36.480 1001.350 36.620 ;
        RECT 644.990 36.420 645.310 36.480 ;
        RECT 1001.030 36.420 1001.350 36.480 ;
      LAYER via ;
        RECT 645.020 36.420 645.280 36.680 ;
        RECT 1001.060 36.420 1001.320 36.680 ;
      LAYER met2 ;
        RECT 1001.750 600.170 1002.030 604.000 ;
        RECT 1001.120 600.030 1002.030 600.170 ;
        RECT 1001.120 36.710 1001.260 600.030 ;
        RECT 1001.750 600.000 1002.030 600.030 ;
        RECT 645.020 36.390 645.280 36.710 ;
        RECT 1001.060 36.390 1001.320 36.710 ;
        RECT 645.080 2.400 645.220 36.390 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1921.950 587.760 1922.270 587.820 ;
        RECT 1993.710 587.760 1994.030 587.820 ;
        RECT 1921.950 587.620 1994.030 587.760 ;
        RECT 1921.950 587.560 1922.270 587.620 ;
        RECT 1993.710 587.560 1994.030 587.620 ;
        RECT 1994.170 587.760 1994.490 587.820 ;
        RECT 2066.390 587.760 2066.710 587.820 ;
        RECT 1994.170 587.620 2066.710 587.760 ;
        RECT 1994.170 587.560 1994.490 587.620 ;
        RECT 2066.390 587.560 2066.710 587.620 ;
        RECT 2065.930 18.600 2066.250 18.660 ;
        RECT 2090.310 18.600 2090.630 18.660 ;
        RECT 2065.930 18.460 2090.630 18.600 ;
        RECT 2065.930 18.400 2066.250 18.460 ;
        RECT 2090.310 18.400 2090.630 18.460 ;
        RECT 2090.770 18.260 2091.090 18.320 ;
        RECT 2111.470 18.260 2111.790 18.320 ;
        RECT 2090.770 18.120 2111.790 18.260 ;
        RECT 2090.770 18.060 2091.090 18.120 ;
        RECT 2111.470 18.060 2111.790 18.120 ;
        RECT 2090.310 17.580 2090.630 17.640 ;
        RECT 2090.770 17.580 2091.090 17.640 ;
        RECT 2090.310 17.440 2091.090 17.580 ;
        RECT 2090.310 17.380 2090.630 17.440 ;
        RECT 2090.770 17.380 2091.090 17.440 ;
        RECT 2410.930 14.860 2411.250 14.920 ;
        RECT 2428.870 14.860 2429.190 14.920 ;
        RECT 2235.760 14.720 2284.200 14.860 ;
        RECT 2173.570 14.520 2173.890 14.580 ;
        RECT 2186.910 14.520 2187.230 14.580 ;
        RECT 2173.570 14.380 2187.230 14.520 ;
        RECT 2173.570 14.320 2173.890 14.380 ;
        RECT 2186.910 14.320 2187.230 14.380 ;
        RECT 2187.370 14.520 2187.690 14.580 ;
        RECT 2235.760 14.520 2235.900 14.720 ;
        RECT 2187.370 14.380 2235.900 14.520 ;
        RECT 2284.060 14.520 2284.200 14.720 ;
        RECT 2410.930 14.720 2429.190 14.860 ;
        RECT 2410.930 14.660 2411.250 14.720 ;
        RECT 2428.870 14.660 2429.190 14.720 ;
        RECT 2318.470 14.520 2318.790 14.580 ;
        RECT 2284.060 14.380 2318.790 14.520 ;
        RECT 2187.370 14.320 2187.690 14.380 ;
        RECT 2318.470 14.320 2318.790 14.380 ;
        RECT 2366.310 14.180 2366.630 14.240 ;
        RECT 2410.010 14.180 2410.330 14.240 ;
        RECT 2366.310 14.040 2410.330 14.180 ;
        RECT 2366.310 13.980 2366.630 14.040 ;
        RECT 2410.010 13.980 2410.330 14.040 ;
        RECT 2111.470 13.840 2111.790 13.900 ;
        RECT 2173.570 13.840 2173.890 13.900 ;
        RECT 2111.470 13.700 2173.890 13.840 ;
        RECT 2111.470 13.640 2111.790 13.700 ;
        RECT 2173.570 13.640 2173.890 13.700 ;
      LAYER via ;
        RECT 1921.980 587.560 1922.240 587.820 ;
        RECT 1993.740 587.560 1994.000 587.820 ;
        RECT 1994.200 587.560 1994.460 587.820 ;
        RECT 2066.420 587.560 2066.680 587.820 ;
        RECT 2065.960 18.400 2066.220 18.660 ;
        RECT 2090.340 18.400 2090.600 18.660 ;
        RECT 2090.800 18.060 2091.060 18.320 ;
        RECT 2111.500 18.060 2111.760 18.320 ;
        RECT 2090.340 17.380 2090.600 17.640 ;
        RECT 2090.800 17.380 2091.060 17.640 ;
        RECT 2173.600 14.320 2173.860 14.580 ;
        RECT 2186.940 14.320 2187.200 14.580 ;
        RECT 2187.400 14.320 2187.660 14.580 ;
        RECT 2410.960 14.660 2411.220 14.920 ;
        RECT 2428.900 14.660 2429.160 14.920 ;
        RECT 2318.500 14.320 2318.760 14.580 ;
        RECT 2366.340 13.980 2366.600 14.240 ;
        RECT 2410.040 13.980 2410.300 14.240 ;
        RECT 2111.500 13.640 2111.760 13.900 ;
        RECT 2173.600 13.640 2173.860 13.900 ;
      LAYER met2 ;
        RECT 1920.370 600.170 1920.650 604.000 ;
        RECT 1920.370 600.030 1922.180 600.170 ;
        RECT 1920.370 600.000 1920.650 600.030 ;
        RECT 1922.040 587.850 1922.180 600.030 ;
        RECT 1993.800 587.850 1994.400 587.930 ;
        RECT 1921.980 587.530 1922.240 587.850 ;
        RECT 1993.740 587.790 1994.460 587.850 ;
        RECT 1993.740 587.530 1994.000 587.790 ;
        RECT 1994.200 587.530 1994.460 587.790 ;
        RECT 2066.420 587.530 2066.680 587.850 ;
        RECT 2066.480 39.850 2066.620 587.530 ;
        RECT 2066.020 39.710 2066.620 39.850 ;
        RECT 2066.020 18.690 2066.160 39.710 ;
        RECT 2065.960 18.370 2066.220 18.690 ;
        RECT 2090.340 18.370 2090.600 18.690 ;
        RECT 2090.400 17.670 2090.540 18.370 ;
        RECT 2090.800 18.030 2091.060 18.350 ;
        RECT 2111.500 18.030 2111.760 18.350 ;
        RECT 2090.860 17.670 2091.000 18.030 ;
        RECT 2090.340 17.350 2090.600 17.670 ;
        RECT 2090.800 17.350 2091.060 17.670 ;
        RECT 2111.560 13.930 2111.700 18.030 ;
        RECT 2187.000 14.610 2187.600 14.690 ;
        RECT 2173.600 14.290 2173.860 14.610 ;
        RECT 2186.940 14.550 2187.660 14.610 ;
        RECT 2186.940 14.290 2187.200 14.550 ;
        RECT 2187.400 14.290 2187.660 14.550 ;
        RECT 2318.490 14.435 2318.770 14.805 ;
        RECT 2366.330 14.435 2366.610 14.805 ;
        RECT 2410.960 14.630 2411.220 14.950 ;
        RECT 2428.900 14.630 2429.160 14.950 ;
        RECT 2318.500 14.290 2318.760 14.435 ;
        RECT 2173.660 13.930 2173.800 14.290 ;
        RECT 2366.400 14.270 2366.540 14.435 ;
        RECT 2366.340 13.950 2366.600 14.270 ;
        RECT 2410.040 14.180 2410.300 14.270 ;
        RECT 2411.020 14.180 2411.160 14.630 ;
        RECT 2410.040 14.040 2411.160 14.180 ;
        RECT 2410.040 13.950 2410.300 14.040 ;
        RECT 2111.500 13.610 2111.760 13.930 ;
        RECT 2173.600 13.610 2173.860 13.930 ;
        RECT 2428.960 2.400 2429.100 14.630 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
      LAYER via2 ;
        RECT 2318.490 14.480 2318.770 14.760 ;
        RECT 2366.330 14.480 2366.610 14.760 ;
      LAYER met3 ;
        RECT 2318.465 14.770 2318.795 14.785 ;
        RECT 2366.305 14.770 2366.635 14.785 ;
        RECT 2318.465 14.470 2366.635 14.770 ;
        RECT 2318.465 14.455 2318.795 14.470 ;
        RECT 2366.305 14.455 2366.635 14.470 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1931.150 591.160 1931.470 591.220 ;
        RECT 2349.290 591.160 2349.610 591.220 ;
        RECT 1931.150 591.020 2349.610 591.160 ;
        RECT 1931.150 590.960 1931.470 591.020 ;
        RECT 2349.290 590.960 2349.610 591.020 ;
        RECT 2349.290 15.540 2349.610 15.600 ;
        RECT 2446.810 15.540 2447.130 15.600 ;
        RECT 2349.290 15.400 2447.130 15.540 ;
        RECT 2349.290 15.340 2349.610 15.400 ;
        RECT 2446.810 15.340 2447.130 15.400 ;
      LAYER via ;
        RECT 1931.180 590.960 1931.440 591.220 ;
        RECT 2349.320 590.960 2349.580 591.220 ;
        RECT 2349.320 15.340 2349.580 15.600 ;
        RECT 2446.840 15.340 2447.100 15.600 ;
      LAYER met2 ;
        RECT 1929.570 600.170 1929.850 604.000 ;
        RECT 1929.570 600.030 1931.380 600.170 ;
        RECT 1929.570 600.000 1929.850 600.030 ;
        RECT 1931.240 591.250 1931.380 600.030 ;
        RECT 1931.180 590.930 1931.440 591.250 ;
        RECT 2349.320 590.930 2349.580 591.250 ;
        RECT 2349.380 15.630 2349.520 590.930 ;
        RECT 2349.320 15.310 2349.580 15.630 ;
        RECT 2446.840 15.310 2447.100 15.630 ;
        RECT 2446.900 2.400 2447.040 15.310 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1940.350 586.740 1940.670 586.800 ;
        RECT 1945.410 586.740 1945.730 586.800 ;
        RECT 1940.350 586.600 1945.730 586.740 ;
        RECT 1940.350 586.540 1940.670 586.600 ;
        RECT 1945.410 586.540 1945.730 586.600 ;
        RECT 1945.410 16.900 1945.730 16.960 ;
        RECT 2464.750 16.900 2465.070 16.960 ;
        RECT 1945.410 16.760 2465.070 16.900 ;
        RECT 1945.410 16.700 1945.730 16.760 ;
        RECT 2464.750 16.700 2465.070 16.760 ;
      LAYER via ;
        RECT 1940.380 586.540 1940.640 586.800 ;
        RECT 1945.440 586.540 1945.700 586.800 ;
        RECT 1945.440 16.700 1945.700 16.960 ;
        RECT 2464.780 16.700 2465.040 16.960 ;
      LAYER met2 ;
        RECT 1938.770 600.170 1939.050 604.000 ;
        RECT 1938.770 600.030 1940.580 600.170 ;
        RECT 1938.770 600.000 1939.050 600.030 ;
        RECT 1940.440 586.830 1940.580 600.030 ;
        RECT 1940.380 586.510 1940.640 586.830 ;
        RECT 1945.440 586.510 1945.700 586.830 ;
        RECT 1945.500 16.990 1945.640 586.510 ;
        RECT 1945.440 16.670 1945.700 16.990 ;
        RECT 2464.780 16.670 2465.040 16.990 ;
        RECT 2464.840 2.400 2464.980 16.670 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1949.550 591.500 1949.870 591.560 ;
        RECT 2369.990 591.500 2370.310 591.560 ;
        RECT 1949.550 591.360 2370.310 591.500 ;
        RECT 1949.550 591.300 1949.870 591.360 ;
        RECT 2369.990 591.300 2370.310 591.360 ;
        RECT 2369.990 15.880 2370.310 15.940 ;
        RECT 2482.690 15.880 2483.010 15.940 ;
        RECT 2369.990 15.740 2483.010 15.880 ;
        RECT 2369.990 15.680 2370.310 15.740 ;
        RECT 2482.690 15.680 2483.010 15.740 ;
      LAYER via ;
        RECT 1949.580 591.300 1949.840 591.560 ;
        RECT 2370.020 591.300 2370.280 591.560 ;
        RECT 2370.020 15.680 2370.280 15.940 ;
        RECT 2482.720 15.680 2482.980 15.940 ;
      LAYER met2 ;
        RECT 1947.970 600.170 1948.250 604.000 ;
        RECT 1947.970 600.030 1949.780 600.170 ;
        RECT 1947.970 600.000 1948.250 600.030 ;
        RECT 1949.640 591.590 1949.780 600.030 ;
        RECT 1949.580 591.270 1949.840 591.590 ;
        RECT 2370.020 591.270 2370.280 591.590 ;
        RECT 2370.080 15.970 2370.220 591.270 ;
        RECT 2370.020 15.650 2370.280 15.970 ;
        RECT 2482.720 15.650 2482.980 15.970 ;
        RECT 2482.780 2.400 2482.920 15.650 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1958.750 20.640 1959.070 20.700 ;
        RECT 2500.630 20.640 2500.950 20.700 ;
        RECT 1958.750 20.500 2500.950 20.640 ;
        RECT 1958.750 20.440 1959.070 20.500 ;
        RECT 2500.630 20.440 2500.950 20.500 ;
      LAYER via ;
        RECT 1958.780 20.440 1959.040 20.700 ;
        RECT 2500.660 20.440 2500.920 20.700 ;
      LAYER met2 ;
        RECT 1957.170 600.170 1957.450 604.000 ;
        RECT 1957.170 600.030 1959.440 600.170 ;
        RECT 1957.170 600.000 1957.450 600.030 ;
        RECT 1959.300 33.730 1959.440 600.030 ;
        RECT 1958.840 33.590 1959.440 33.730 ;
        RECT 1958.840 20.730 1958.980 33.590 ;
        RECT 1958.780 20.410 1959.040 20.730 ;
        RECT 2500.660 20.410 2500.920 20.730 ;
        RECT 2500.720 2.400 2500.860 20.410 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1967.950 592.520 1968.270 592.580 ;
        RECT 2376.890 592.520 2377.210 592.580 ;
        RECT 1967.950 592.380 2377.210 592.520 ;
        RECT 1967.950 592.320 1968.270 592.380 ;
        RECT 2376.890 592.320 2377.210 592.380 ;
        RECT 2376.890 34.580 2377.210 34.640 ;
        RECT 2412.310 34.580 2412.630 34.640 ;
        RECT 2376.890 34.440 2412.630 34.580 ;
        RECT 2376.890 34.380 2377.210 34.440 ;
        RECT 2412.310 34.380 2412.630 34.440 ;
        RECT 2451.870 16.220 2452.190 16.280 ;
        RECT 2518.110 16.220 2518.430 16.280 ;
        RECT 2451.870 16.080 2518.430 16.220 ;
        RECT 2451.870 16.020 2452.190 16.080 ;
        RECT 2518.110 16.020 2518.430 16.080 ;
        RECT 2412.310 15.200 2412.630 15.260 ;
        RECT 2412.310 15.060 2431.860 15.200 ;
        RECT 2412.310 15.000 2412.630 15.060 ;
        RECT 2431.720 14.520 2431.860 15.060 ;
        RECT 2451.870 14.520 2452.190 14.580 ;
        RECT 2431.720 14.380 2452.190 14.520 ;
        RECT 2451.870 14.320 2452.190 14.380 ;
      LAYER via ;
        RECT 1967.980 592.320 1968.240 592.580 ;
        RECT 2376.920 592.320 2377.180 592.580 ;
        RECT 2376.920 34.380 2377.180 34.640 ;
        RECT 2412.340 34.380 2412.600 34.640 ;
        RECT 2451.900 16.020 2452.160 16.280 ;
        RECT 2518.140 16.020 2518.400 16.280 ;
        RECT 2412.340 15.000 2412.600 15.260 ;
        RECT 2451.900 14.320 2452.160 14.580 ;
      LAYER met2 ;
        RECT 1966.370 600.170 1966.650 604.000 ;
        RECT 1966.370 600.030 1968.180 600.170 ;
        RECT 1966.370 600.000 1966.650 600.030 ;
        RECT 1968.040 592.610 1968.180 600.030 ;
        RECT 1967.980 592.290 1968.240 592.610 ;
        RECT 2376.920 592.290 2377.180 592.610 ;
        RECT 2376.980 34.670 2377.120 592.290 ;
        RECT 2376.920 34.350 2377.180 34.670 ;
        RECT 2412.340 34.350 2412.600 34.670 ;
        RECT 2412.400 15.290 2412.540 34.350 ;
        RECT 2451.900 15.990 2452.160 16.310 ;
        RECT 2518.140 15.990 2518.400 16.310 ;
        RECT 2412.340 14.970 2412.600 15.290 ;
        RECT 2451.960 14.610 2452.100 15.990 ;
        RECT 2451.900 14.290 2452.160 14.610 ;
        RECT 2518.200 2.400 2518.340 15.990 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1975.540 598.980 1975.860 599.040 ;
        RECT 1979.910 598.980 1980.230 599.040 ;
        RECT 1975.540 598.840 1980.230 598.980 ;
        RECT 1975.540 598.780 1975.860 598.840 ;
        RECT 1979.910 598.780 1980.230 598.840 ;
        RECT 1979.910 20.300 1980.230 20.360 ;
        RECT 2536.050 20.300 2536.370 20.360 ;
        RECT 1979.910 20.160 2536.370 20.300 ;
        RECT 1979.910 20.100 1980.230 20.160 ;
        RECT 2536.050 20.100 2536.370 20.160 ;
      LAYER via ;
        RECT 1975.570 598.780 1975.830 599.040 ;
        RECT 1979.940 598.780 1980.200 599.040 ;
        RECT 1979.940 20.100 1980.200 20.360 ;
        RECT 2536.080 20.100 2536.340 20.360 ;
      LAYER met2 ;
        RECT 1975.570 600.000 1975.850 604.000 ;
        RECT 1975.630 599.070 1975.770 600.000 ;
        RECT 1975.570 598.750 1975.830 599.070 ;
        RECT 1979.940 598.750 1980.200 599.070 ;
        RECT 1980.000 20.390 1980.140 598.750 ;
        RECT 1979.940 20.070 1980.200 20.390 ;
        RECT 2536.080 20.070 2536.340 20.390 ;
        RECT 2536.140 2.400 2536.280 20.070 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1986.350 592.180 1986.670 592.240 ;
        RECT 2390.690 592.180 2391.010 592.240 ;
        RECT 1986.350 592.040 2391.010 592.180 ;
        RECT 1986.350 591.980 1986.670 592.040 ;
        RECT 2390.690 591.980 2391.010 592.040 ;
        RECT 2410.470 16.220 2410.790 16.280 ;
        RECT 2451.410 16.220 2451.730 16.280 ;
        RECT 2410.470 16.080 2451.730 16.220 ;
        RECT 2410.470 16.020 2410.790 16.080 ;
        RECT 2451.410 16.020 2451.730 16.080 ;
        RECT 2390.690 14.860 2391.010 14.920 ;
        RECT 2410.470 14.860 2410.790 14.920 ;
        RECT 2390.690 14.720 2410.790 14.860 ;
        RECT 2390.690 14.660 2391.010 14.720 ;
        RECT 2410.470 14.660 2410.790 14.720 ;
        RECT 2454.170 14.860 2454.490 14.920 ;
        RECT 2553.990 14.860 2554.310 14.920 ;
        RECT 2454.170 14.720 2554.310 14.860 ;
        RECT 2454.170 14.660 2454.490 14.720 ;
        RECT 2553.990 14.660 2554.310 14.720 ;
      LAYER via ;
        RECT 1986.380 591.980 1986.640 592.240 ;
        RECT 2390.720 591.980 2390.980 592.240 ;
        RECT 2410.500 16.020 2410.760 16.280 ;
        RECT 2451.440 16.020 2451.700 16.280 ;
        RECT 2390.720 14.660 2390.980 14.920 ;
        RECT 2410.500 14.660 2410.760 14.920 ;
        RECT 2454.200 14.660 2454.460 14.920 ;
        RECT 2554.020 14.660 2554.280 14.920 ;
      LAYER met2 ;
        RECT 1984.770 600.170 1985.050 604.000 ;
        RECT 1984.770 600.030 1986.580 600.170 ;
        RECT 1984.770 600.000 1985.050 600.030 ;
        RECT 1986.440 592.270 1986.580 600.030 ;
        RECT 1986.380 591.950 1986.640 592.270 ;
        RECT 2390.720 591.950 2390.980 592.270 ;
        RECT 2390.780 14.950 2390.920 591.950 ;
        RECT 2410.500 15.990 2410.760 16.310 ;
        RECT 2451.440 15.990 2451.700 16.310 ;
        RECT 2410.560 14.950 2410.700 15.990 ;
        RECT 2451.500 15.485 2451.640 15.990 ;
        RECT 2451.430 15.115 2451.710 15.485 ;
        RECT 2454.190 15.115 2454.470 15.485 ;
        RECT 2454.260 14.950 2454.400 15.115 ;
        RECT 2390.720 14.630 2390.980 14.950 ;
        RECT 2410.500 14.630 2410.760 14.950 ;
        RECT 2454.200 14.630 2454.460 14.950 ;
        RECT 2554.020 14.630 2554.280 14.950 ;
        RECT 2554.080 2.400 2554.220 14.630 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
      LAYER via2 ;
        RECT 2451.430 15.160 2451.710 15.440 ;
        RECT 2454.190 15.160 2454.470 15.440 ;
      LAYER met3 ;
        RECT 2451.405 15.450 2451.735 15.465 ;
        RECT 2454.165 15.450 2454.495 15.465 ;
        RECT 2451.405 15.150 2454.495 15.450 ;
        RECT 2451.405 15.135 2451.735 15.150 ;
        RECT 2454.165 15.135 2454.495 15.150 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1995.550 586.740 1995.870 586.800 ;
        RECT 2000.610 586.740 2000.930 586.800 ;
        RECT 1995.550 586.600 2000.930 586.740 ;
        RECT 1995.550 586.540 1995.870 586.600 ;
        RECT 2000.610 586.540 2000.930 586.600 ;
        RECT 2000.610 19.960 2000.930 20.020 ;
        RECT 2571.930 19.960 2572.250 20.020 ;
        RECT 2000.610 19.820 2572.250 19.960 ;
        RECT 2000.610 19.760 2000.930 19.820 ;
        RECT 2571.930 19.760 2572.250 19.820 ;
      LAYER via ;
        RECT 1995.580 586.540 1995.840 586.800 ;
        RECT 2000.640 586.540 2000.900 586.800 ;
        RECT 2000.640 19.760 2000.900 20.020 ;
        RECT 2571.960 19.760 2572.220 20.020 ;
      LAYER met2 ;
        RECT 1993.970 600.170 1994.250 604.000 ;
        RECT 1993.970 600.030 1995.780 600.170 ;
        RECT 1993.970 600.000 1994.250 600.030 ;
        RECT 1995.640 586.830 1995.780 600.030 ;
        RECT 1995.580 586.510 1995.840 586.830 ;
        RECT 2000.640 586.510 2000.900 586.830 ;
        RECT 2000.700 20.050 2000.840 586.510 ;
        RECT 2000.640 19.730 2000.900 20.050 ;
        RECT 2571.960 19.730 2572.220 20.050 ;
        RECT 2572.020 2.400 2572.160 19.730 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2084.790 589.460 2085.110 589.520 ;
        RECT 2103.650 589.460 2103.970 589.520 ;
        RECT 2084.790 589.320 2103.970 589.460 ;
        RECT 2084.790 589.260 2085.110 589.320 ;
        RECT 2103.650 589.260 2103.970 589.320 ;
        RECT 2318.930 589.120 2319.250 589.180 ;
        RECT 2138.700 588.980 2319.250 589.120 ;
        RECT 2004.290 588.780 2004.610 588.840 ;
        RECT 2065.470 588.780 2065.790 588.840 ;
        RECT 2004.290 588.640 2065.790 588.780 ;
        RECT 2004.290 588.580 2004.610 588.640 ;
        RECT 2065.470 588.580 2065.790 588.640 ;
        RECT 2122.050 588.440 2122.370 588.500 ;
        RECT 2138.700 588.440 2138.840 588.980 ;
        RECT 2318.930 588.920 2319.250 588.980 ;
        RECT 2320.770 589.120 2321.090 589.180 ;
        RECT 2404.490 589.120 2404.810 589.180 ;
        RECT 2320.770 588.980 2404.810 589.120 ;
        RECT 2320.770 588.920 2321.090 588.980 ;
        RECT 2404.490 588.920 2404.810 588.980 ;
        RECT 2122.050 588.300 2138.840 588.440 ;
        RECT 2122.050 588.240 2122.370 588.300 ;
        RECT 2084.790 587.760 2085.110 587.820 ;
        RECT 2066.940 587.620 2085.110 587.760 ;
        RECT 2065.470 587.420 2065.790 587.480 ;
        RECT 2066.940 587.420 2067.080 587.620 ;
        RECT 2084.790 587.560 2085.110 587.620 ;
        RECT 2103.650 587.760 2103.970 587.820 ;
        RECT 2103.650 587.620 2111.700 587.760 ;
        RECT 2103.650 587.560 2103.970 587.620 ;
        RECT 2065.470 587.280 2067.080 587.420 ;
        RECT 2111.560 587.420 2111.700 587.620 ;
        RECT 2120.210 587.420 2120.530 587.480 ;
        RECT 2111.560 587.280 2120.530 587.420 ;
        RECT 2065.470 587.220 2065.790 587.280 ;
        RECT 2120.210 587.220 2120.530 587.280 ;
        RECT 2411.850 16.560 2412.170 16.620 ;
        RECT 2453.250 16.560 2453.570 16.620 ;
        RECT 2411.850 16.420 2453.570 16.560 ;
        RECT 2411.850 16.360 2412.170 16.420 ;
        RECT 2453.250 16.360 2453.570 16.420 ;
        RECT 2404.490 15.200 2404.810 15.260 ;
        RECT 2411.850 15.200 2412.170 15.260 ;
        RECT 2404.490 15.060 2412.170 15.200 ;
        RECT 2404.490 15.000 2404.810 15.060 ;
        RECT 2411.850 15.000 2412.170 15.060 ;
        RECT 2453.250 14.180 2453.570 14.240 ;
        RECT 2589.410 14.180 2589.730 14.240 ;
        RECT 2453.250 14.040 2589.730 14.180 ;
        RECT 2453.250 13.980 2453.570 14.040 ;
        RECT 2589.410 13.980 2589.730 14.040 ;
      LAYER via ;
        RECT 2084.820 589.260 2085.080 589.520 ;
        RECT 2103.680 589.260 2103.940 589.520 ;
        RECT 2004.320 588.580 2004.580 588.840 ;
        RECT 2065.500 588.580 2065.760 588.840 ;
        RECT 2122.080 588.240 2122.340 588.500 ;
        RECT 2318.960 588.920 2319.220 589.180 ;
        RECT 2320.800 588.920 2321.060 589.180 ;
        RECT 2404.520 588.920 2404.780 589.180 ;
        RECT 2065.500 587.220 2065.760 587.480 ;
        RECT 2084.820 587.560 2085.080 587.820 ;
        RECT 2103.680 587.560 2103.940 587.820 ;
        RECT 2120.240 587.220 2120.500 587.480 ;
        RECT 2411.880 16.360 2412.140 16.620 ;
        RECT 2453.280 16.360 2453.540 16.620 ;
        RECT 2404.520 15.000 2404.780 15.260 ;
        RECT 2411.880 15.000 2412.140 15.260 ;
        RECT 2453.280 13.980 2453.540 14.240 ;
        RECT 2589.440 13.980 2589.700 14.240 ;
      LAYER met2 ;
        RECT 2002.710 600.170 2002.990 604.000 ;
        RECT 2002.710 600.030 2004.520 600.170 ;
        RECT 2002.710 600.000 2002.990 600.030 ;
        RECT 2004.380 588.870 2004.520 600.030 ;
        RECT 2084.820 589.230 2085.080 589.550 ;
        RECT 2103.680 589.230 2103.940 589.550 ;
        RECT 2004.320 588.550 2004.580 588.870 ;
        RECT 2065.500 588.550 2065.760 588.870 ;
        RECT 2065.560 587.510 2065.700 588.550 ;
        RECT 2084.880 587.850 2085.020 589.230 ;
        RECT 2103.740 587.850 2103.880 589.230 ;
        RECT 2121.220 589.150 2122.280 589.290 ;
        RECT 2084.820 587.530 2085.080 587.850 ;
        RECT 2103.680 587.530 2103.940 587.850 ;
        RECT 2065.500 587.190 2065.760 587.510 ;
        RECT 2120.240 587.190 2120.500 587.510 ;
        RECT 2120.300 586.570 2120.440 587.190 ;
        RECT 2121.220 586.570 2121.360 589.150 ;
        RECT 2122.140 588.530 2122.280 589.150 ;
        RECT 2318.950 589.035 2319.230 589.405 ;
        RECT 2320.790 589.035 2321.070 589.405 ;
        RECT 2318.960 588.890 2319.220 589.035 ;
        RECT 2320.800 588.890 2321.060 589.035 ;
        RECT 2404.520 588.890 2404.780 589.210 ;
        RECT 2122.080 588.210 2122.340 588.530 ;
        RECT 2120.300 586.430 2121.360 586.570 ;
        RECT 2404.580 15.290 2404.720 588.890 ;
        RECT 2411.880 16.330 2412.140 16.650 ;
        RECT 2453.280 16.330 2453.540 16.650 ;
        RECT 2411.940 15.290 2412.080 16.330 ;
        RECT 2404.520 14.970 2404.780 15.290 ;
        RECT 2411.880 14.970 2412.140 15.290 ;
        RECT 2453.340 14.270 2453.480 16.330 ;
        RECT 2453.280 13.950 2453.540 14.270 ;
        RECT 2589.440 13.950 2589.700 14.270 ;
        RECT 2589.500 2.400 2589.640 13.950 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
      LAYER via2 ;
        RECT 2318.950 589.080 2319.230 589.360 ;
        RECT 2320.790 589.080 2321.070 589.360 ;
      LAYER met3 ;
        RECT 2318.925 589.370 2319.255 589.385 ;
        RECT 2320.765 589.370 2321.095 589.385 ;
        RECT 2318.925 589.070 2321.095 589.370 ;
        RECT 2318.925 589.055 2319.255 589.070 ;
        RECT 2320.765 589.055 2321.095 589.070 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 879.590 592.520 879.910 592.580 ;
        RECT 1092.110 592.520 1092.430 592.580 ;
        RECT 879.590 592.380 1092.430 592.520 ;
        RECT 879.590 592.320 879.910 592.380 ;
        RECT 1092.110 592.320 1092.430 592.380 ;
        RECT 823.470 19.620 823.790 19.680 ;
        RECT 879.590 19.620 879.910 19.680 ;
        RECT 823.470 19.480 879.910 19.620 ;
        RECT 823.470 19.420 823.790 19.480 ;
        RECT 879.590 19.420 879.910 19.480 ;
      LAYER via ;
        RECT 879.620 592.320 879.880 592.580 ;
        RECT 1092.140 592.320 1092.400 592.580 ;
        RECT 823.500 19.420 823.760 19.680 ;
        RECT 879.620 19.420 879.880 19.680 ;
      LAYER met2 ;
        RECT 1093.750 600.170 1094.030 604.000 ;
        RECT 1092.200 600.030 1094.030 600.170 ;
        RECT 1092.200 592.610 1092.340 600.030 ;
        RECT 1093.750 600.000 1094.030 600.030 ;
        RECT 879.620 592.290 879.880 592.610 ;
        RECT 1092.140 592.290 1092.400 592.610 ;
        RECT 879.680 19.710 879.820 592.290 ;
        RECT 823.500 19.390 823.760 19.710 ;
        RECT 879.620 19.390 879.880 19.710 ;
        RECT 823.560 2.400 823.700 19.390 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2014.410 19.620 2014.730 19.680 ;
        RECT 2607.350 19.620 2607.670 19.680 ;
        RECT 2014.410 19.480 2607.670 19.620 ;
        RECT 2014.410 19.420 2014.730 19.480 ;
        RECT 2607.350 19.420 2607.670 19.480 ;
      LAYER via ;
        RECT 2014.440 19.420 2014.700 19.680 ;
        RECT 2607.380 19.420 2607.640 19.680 ;
      LAYER met2 ;
        RECT 2011.910 600.170 2012.190 604.000 ;
        RECT 2011.910 600.030 2014.640 600.170 ;
        RECT 2011.910 600.000 2012.190 600.030 ;
        RECT 2014.500 19.710 2014.640 600.030 ;
        RECT 2014.440 19.390 2014.700 19.710 ;
        RECT 2607.380 19.390 2607.640 19.710 ;
        RECT 2607.440 2.400 2607.580 19.390 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2021.310 588.100 2021.630 588.160 ;
        RECT 2113.310 588.100 2113.630 588.160 ;
        RECT 2021.310 587.960 2113.630 588.100 ;
        RECT 2021.310 587.900 2021.630 587.960 ;
        RECT 2113.310 587.900 2113.630 587.960 ;
        RECT 2114.230 588.100 2114.550 588.160 ;
        RECT 2411.390 588.100 2411.710 588.160 ;
        RECT 2114.230 587.960 2411.710 588.100 ;
        RECT 2114.230 587.900 2114.550 587.960 ;
        RECT 2411.390 587.900 2411.710 587.960 ;
        RECT 2453.710 16.560 2454.030 16.620 ;
        RECT 2476.250 16.560 2476.570 16.620 ;
        RECT 2453.710 16.420 2476.570 16.560 ;
        RECT 2453.710 16.360 2454.030 16.420 ;
        RECT 2476.250 16.360 2476.570 16.420 ;
        RECT 2453.710 14.520 2454.030 14.580 ;
        RECT 2452.880 14.380 2454.030 14.520 ;
        RECT 2412.770 14.180 2413.090 14.240 ;
        RECT 2452.880 14.180 2453.020 14.380 ;
        RECT 2453.710 14.320 2454.030 14.380 ;
        RECT 2476.250 14.520 2476.570 14.580 ;
        RECT 2625.290 14.520 2625.610 14.580 ;
        RECT 2476.250 14.380 2625.610 14.520 ;
        RECT 2476.250 14.320 2476.570 14.380 ;
        RECT 2625.290 14.320 2625.610 14.380 ;
        RECT 2412.770 14.040 2453.020 14.180 ;
        RECT 2412.770 13.980 2413.090 14.040 ;
      LAYER via ;
        RECT 2021.340 587.900 2021.600 588.160 ;
        RECT 2113.340 587.900 2113.600 588.160 ;
        RECT 2114.260 587.900 2114.520 588.160 ;
        RECT 2411.420 587.900 2411.680 588.160 ;
        RECT 2453.740 16.360 2454.000 16.620 ;
        RECT 2476.280 16.360 2476.540 16.620 ;
        RECT 2412.800 13.980 2413.060 14.240 ;
        RECT 2453.740 14.320 2454.000 14.580 ;
        RECT 2476.280 14.320 2476.540 14.580 ;
        RECT 2625.320 14.320 2625.580 14.580 ;
      LAYER met2 ;
        RECT 2021.110 600.000 2021.390 604.000 ;
        RECT 2021.170 598.810 2021.310 600.000 ;
        RECT 2021.170 598.670 2021.540 598.810 ;
        RECT 2021.400 588.190 2021.540 598.670 ;
        RECT 2021.340 587.870 2021.600 588.190 ;
        RECT 2113.340 587.930 2113.600 588.190 ;
        RECT 2114.260 587.930 2114.520 588.190 ;
        RECT 2113.340 587.870 2114.520 587.930 ;
        RECT 2411.420 587.870 2411.680 588.190 ;
        RECT 2113.400 587.790 2114.460 587.870 ;
        RECT 2411.480 38.490 2411.620 587.870 ;
        RECT 2411.480 38.350 2413.000 38.490 ;
        RECT 2412.860 14.270 2413.000 38.350 ;
        RECT 2453.740 16.330 2454.000 16.650 ;
        RECT 2476.280 16.330 2476.540 16.650 ;
        RECT 2453.800 14.610 2453.940 16.330 ;
        RECT 2476.340 14.610 2476.480 16.330 ;
        RECT 2453.740 14.290 2454.000 14.610 ;
        RECT 2476.280 14.290 2476.540 14.610 ;
        RECT 2625.320 14.290 2625.580 14.610 ;
        RECT 2412.800 13.950 2413.060 14.270 ;
        RECT 2625.380 2.400 2625.520 14.290 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2031.890 586.740 2032.210 586.800 ;
        RECT 2035.110 586.740 2035.430 586.800 ;
        RECT 2031.890 586.600 2035.430 586.740 ;
        RECT 2031.890 586.540 2032.210 586.600 ;
        RECT 2035.110 586.540 2035.430 586.600 ;
        RECT 2035.110 19.280 2035.430 19.340 ;
        RECT 2643.230 19.280 2643.550 19.340 ;
        RECT 2035.110 19.140 2643.550 19.280 ;
        RECT 2035.110 19.080 2035.430 19.140 ;
        RECT 2643.230 19.080 2643.550 19.140 ;
      LAYER via ;
        RECT 2031.920 586.540 2032.180 586.800 ;
        RECT 2035.140 586.540 2035.400 586.800 ;
        RECT 2035.140 19.080 2035.400 19.340 ;
        RECT 2643.260 19.080 2643.520 19.340 ;
      LAYER met2 ;
        RECT 2030.310 600.170 2030.590 604.000 ;
        RECT 2030.310 600.030 2032.120 600.170 ;
        RECT 2030.310 600.000 2030.590 600.030 ;
        RECT 2031.980 586.830 2032.120 600.030 ;
        RECT 2031.920 586.510 2032.180 586.830 ;
        RECT 2035.140 586.510 2035.400 586.830 ;
        RECT 2035.200 19.370 2035.340 586.510 ;
        RECT 2035.140 19.050 2035.400 19.370 ;
        RECT 2643.260 19.050 2643.520 19.370 ;
        RECT 2643.320 2.400 2643.460 19.050 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2041.090 587.080 2041.410 587.140 ;
        RECT 2432.090 587.080 2432.410 587.140 ;
        RECT 2041.090 586.940 2432.410 587.080 ;
        RECT 2041.090 586.880 2041.410 586.940 ;
        RECT 2432.090 586.880 2432.410 586.940 ;
        RECT 2661.170 15.200 2661.490 15.260 ;
        RECT 2452.880 15.060 2661.490 15.200 ;
        RECT 2432.090 14.860 2432.410 14.920 ;
        RECT 2452.880 14.860 2453.020 15.060 ;
        RECT 2661.170 15.000 2661.490 15.060 ;
        RECT 2432.090 14.720 2453.020 14.860 ;
        RECT 2432.090 14.660 2432.410 14.720 ;
      LAYER via ;
        RECT 2041.120 586.880 2041.380 587.140 ;
        RECT 2432.120 586.880 2432.380 587.140 ;
        RECT 2432.120 14.660 2432.380 14.920 ;
        RECT 2661.200 15.000 2661.460 15.260 ;
      LAYER met2 ;
        RECT 2039.510 600.170 2039.790 604.000 ;
        RECT 2039.510 600.030 2041.320 600.170 ;
        RECT 2039.510 600.000 2039.790 600.030 ;
        RECT 2041.180 587.170 2041.320 600.030 ;
        RECT 2041.120 586.850 2041.380 587.170 ;
        RECT 2432.120 586.850 2432.380 587.170 ;
        RECT 2432.180 14.950 2432.320 586.850 ;
        RECT 2661.200 14.970 2661.460 15.290 ;
        RECT 2432.120 14.630 2432.380 14.950 ;
        RECT 2661.260 2.400 2661.400 14.970 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2047.530 46.140 2047.850 46.200 ;
        RECT 2048.910 46.140 2049.230 46.200 ;
        RECT 2047.530 46.000 2049.230 46.140 ;
        RECT 2047.530 45.940 2047.850 46.000 ;
        RECT 2048.910 45.940 2049.230 46.000 ;
        RECT 2047.530 18.940 2047.850 19.000 ;
        RECT 2678.650 18.940 2678.970 19.000 ;
        RECT 2047.530 18.800 2678.970 18.940 ;
        RECT 2047.530 18.740 2047.850 18.800 ;
        RECT 2678.650 18.740 2678.970 18.800 ;
      LAYER via ;
        RECT 2047.560 45.940 2047.820 46.200 ;
        RECT 2048.940 45.940 2049.200 46.200 ;
        RECT 2047.560 18.740 2047.820 19.000 ;
        RECT 2678.680 18.740 2678.940 19.000 ;
      LAYER met2 ;
        RECT 2048.710 600.000 2048.990 604.000 ;
        RECT 2048.770 598.810 2048.910 600.000 ;
        RECT 2048.770 598.670 2049.140 598.810 ;
        RECT 2049.000 46.230 2049.140 598.670 ;
        RECT 2047.560 45.910 2047.820 46.230 ;
        RECT 2048.940 45.910 2049.200 46.230 ;
        RECT 2047.620 19.030 2047.760 45.910 ;
        RECT 2047.560 18.710 2047.820 19.030 ;
        RECT 2678.680 18.710 2678.940 19.030 ;
        RECT 2678.740 2.400 2678.880 18.710 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2059.490 588.440 2059.810 588.500 ;
        RECT 2084.330 588.440 2084.650 588.500 ;
        RECT 2059.490 588.300 2084.650 588.440 ;
        RECT 2059.490 588.240 2059.810 588.300 ;
        RECT 2084.330 588.240 2084.650 588.300 ;
        RECT 2084.330 586.740 2084.650 586.800 ;
        RECT 2445.890 586.740 2446.210 586.800 ;
        RECT 2084.330 586.600 2446.210 586.740 ;
        RECT 2084.330 586.540 2084.650 586.600 ;
        RECT 2445.890 586.540 2446.210 586.600 ;
        RECT 2696.590 15.540 2696.910 15.600 ;
        RECT 2447.360 15.400 2696.910 15.540 ;
        RECT 2445.890 15.200 2446.210 15.260 ;
        RECT 2447.360 15.200 2447.500 15.400 ;
        RECT 2696.590 15.340 2696.910 15.400 ;
        RECT 2445.890 15.060 2447.500 15.200 ;
        RECT 2445.890 15.000 2446.210 15.060 ;
      LAYER via ;
        RECT 2059.520 588.240 2059.780 588.500 ;
        RECT 2084.360 588.240 2084.620 588.500 ;
        RECT 2084.360 586.540 2084.620 586.800 ;
        RECT 2445.920 586.540 2446.180 586.800 ;
        RECT 2445.920 15.000 2446.180 15.260 ;
        RECT 2696.620 15.340 2696.880 15.600 ;
      LAYER met2 ;
        RECT 2057.910 600.170 2058.190 604.000 ;
        RECT 2057.910 600.030 2059.720 600.170 ;
        RECT 2057.910 600.000 2058.190 600.030 ;
        RECT 2059.580 588.530 2059.720 600.030 ;
        RECT 2059.520 588.210 2059.780 588.530 ;
        RECT 2084.360 588.210 2084.620 588.530 ;
        RECT 2084.420 586.830 2084.560 588.210 ;
        RECT 2084.360 586.510 2084.620 586.830 ;
        RECT 2445.920 586.510 2446.180 586.830 ;
        RECT 2445.980 15.290 2446.120 586.510 ;
        RECT 2696.620 15.310 2696.880 15.630 ;
        RECT 2445.920 14.970 2446.180 15.290 ;
        RECT 2696.680 2.400 2696.820 15.310 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2068.690 587.420 2069.010 587.480 ;
        RECT 2080.190 587.420 2080.510 587.480 ;
        RECT 2068.690 587.280 2080.510 587.420 ;
        RECT 2068.690 587.220 2069.010 587.280 ;
        RECT 2080.190 587.220 2080.510 587.280 ;
        RECT 2114.690 18.600 2115.010 18.660 ;
        RECT 2714.530 18.600 2714.850 18.660 ;
        RECT 2114.690 18.460 2714.850 18.600 ;
        RECT 2114.690 18.400 2115.010 18.460 ;
        RECT 2714.530 18.400 2714.850 18.460 ;
        RECT 2080.190 14.860 2080.510 14.920 ;
        RECT 2114.690 14.860 2115.010 14.920 ;
        RECT 2080.190 14.720 2115.010 14.860 ;
        RECT 2080.190 14.660 2080.510 14.720 ;
        RECT 2114.690 14.660 2115.010 14.720 ;
      LAYER via ;
        RECT 2068.720 587.220 2068.980 587.480 ;
        RECT 2080.220 587.220 2080.480 587.480 ;
        RECT 2114.720 18.400 2114.980 18.660 ;
        RECT 2714.560 18.400 2714.820 18.660 ;
        RECT 2080.220 14.660 2080.480 14.920 ;
        RECT 2114.720 14.660 2114.980 14.920 ;
      LAYER met2 ;
        RECT 2067.110 600.170 2067.390 604.000 ;
        RECT 2067.110 600.030 2068.920 600.170 ;
        RECT 2067.110 600.000 2067.390 600.030 ;
        RECT 2068.780 587.510 2068.920 600.030 ;
        RECT 2068.720 587.190 2068.980 587.510 ;
        RECT 2080.220 587.190 2080.480 587.510 ;
        RECT 2080.280 14.950 2080.420 587.190 ;
        RECT 2114.720 18.370 2114.980 18.690 ;
        RECT 2714.560 18.370 2714.820 18.690 ;
        RECT 2114.780 14.950 2114.920 18.370 ;
        RECT 2080.220 14.630 2080.480 14.950 ;
        RECT 2114.720 14.630 2114.980 14.950 ;
        RECT 2714.620 2.400 2714.760 18.370 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2222.330 592.860 2222.650 592.920 ;
        RECT 2283.510 592.860 2283.830 592.920 ;
        RECT 2222.330 592.720 2283.830 592.860 ;
        RECT 2222.330 592.660 2222.650 592.720 ;
        RECT 2283.510 592.660 2283.830 592.720 ;
        RECT 2334.110 590.480 2334.430 590.540 ;
        RECT 2380.110 590.480 2380.430 590.540 ;
        RECT 2334.110 590.340 2380.430 590.480 ;
        RECT 2334.110 590.280 2334.430 590.340 ;
        RECT 2380.110 590.280 2380.430 590.340 ;
        RECT 2462.910 589.120 2463.230 589.180 ;
        RECT 2466.590 589.120 2466.910 589.180 ;
        RECT 2462.910 588.980 2466.910 589.120 ;
        RECT 2462.910 588.920 2463.230 588.980 ;
        RECT 2466.590 588.920 2466.910 588.980 ;
        RECT 2076.510 588.780 2076.830 588.840 ;
        RECT 2090.770 588.780 2091.090 588.840 ;
        RECT 2076.510 588.640 2091.090 588.780 ;
        RECT 2076.510 588.580 2076.830 588.640 ;
        RECT 2090.770 588.580 2091.090 588.640 ;
        RECT 2173.110 588.440 2173.430 588.500 ;
        RECT 2221.870 588.440 2222.190 588.500 ;
        RECT 2173.110 588.300 2222.190 588.440 ;
        RECT 2173.110 588.240 2173.430 588.300 ;
        RECT 2221.870 588.240 2222.190 588.300 ;
        RECT 2283.510 588.440 2283.830 588.500 ;
        RECT 2318.470 588.440 2318.790 588.500 ;
        RECT 2283.510 588.300 2318.790 588.440 ;
        RECT 2283.510 588.240 2283.830 588.300 ;
        RECT 2318.470 588.240 2318.790 588.300 ;
        RECT 2380.110 588.440 2380.430 588.500 ;
        RECT 2415.070 588.440 2415.390 588.500 ;
        RECT 2380.110 588.300 2415.390 588.440 ;
        RECT 2380.110 588.240 2380.430 588.300 ;
        RECT 2415.070 588.240 2415.390 588.300 ;
        RECT 2090.770 586.400 2091.090 586.460 ;
        RECT 2125.270 586.400 2125.590 586.460 ;
        RECT 2090.770 586.260 2125.590 586.400 ;
        RECT 2090.770 586.200 2091.090 586.260 ;
        RECT 2125.270 586.200 2125.590 586.260 ;
        RECT 2125.270 585.720 2125.590 585.780 ;
        RECT 2173.110 585.720 2173.430 585.780 ;
        RECT 2125.270 585.580 2173.430 585.720 ;
        RECT 2125.270 585.520 2125.590 585.580 ;
        RECT 2173.110 585.520 2173.430 585.580 ;
        RECT 2466.590 16.900 2466.910 16.960 ;
        RECT 2479.930 16.900 2480.250 16.960 ;
        RECT 2466.590 16.760 2480.250 16.900 ;
        RECT 2466.590 16.700 2466.910 16.760 ;
        RECT 2479.930 16.700 2480.250 16.760 ;
        RECT 2483.150 15.880 2483.470 15.940 ;
        RECT 2732.470 15.880 2732.790 15.940 ;
        RECT 2483.150 15.740 2732.790 15.880 ;
        RECT 2483.150 15.680 2483.470 15.740 ;
        RECT 2732.470 15.680 2732.790 15.740 ;
      LAYER via ;
        RECT 2222.360 592.660 2222.620 592.920 ;
        RECT 2283.540 592.660 2283.800 592.920 ;
        RECT 2334.140 590.280 2334.400 590.540 ;
        RECT 2380.140 590.280 2380.400 590.540 ;
        RECT 2462.940 588.920 2463.200 589.180 ;
        RECT 2466.620 588.920 2466.880 589.180 ;
        RECT 2076.540 588.580 2076.800 588.840 ;
        RECT 2090.800 588.580 2091.060 588.840 ;
        RECT 2173.140 588.240 2173.400 588.500 ;
        RECT 2221.900 588.240 2222.160 588.500 ;
        RECT 2283.540 588.240 2283.800 588.500 ;
        RECT 2318.500 588.240 2318.760 588.500 ;
        RECT 2380.140 588.240 2380.400 588.500 ;
        RECT 2415.100 588.240 2415.360 588.500 ;
        RECT 2090.800 586.200 2091.060 586.460 ;
        RECT 2125.300 586.200 2125.560 586.460 ;
        RECT 2125.300 585.520 2125.560 585.780 ;
        RECT 2173.140 585.520 2173.400 585.780 ;
        RECT 2466.620 16.700 2466.880 16.960 ;
        RECT 2479.960 16.700 2480.220 16.960 ;
        RECT 2483.180 15.680 2483.440 15.940 ;
        RECT 2732.500 15.680 2732.760 15.940 ;
      LAYER met2 ;
        RECT 2076.310 600.000 2076.590 604.000 ;
        RECT 2076.370 598.810 2076.510 600.000 ;
        RECT 2076.370 598.670 2076.740 598.810 ;
        RECT 2076.600 588.870 2076.740 598.670 ;
        RECT 2222.360 592.630 2222.620 592.950 ;
        RECT 2283.540 592.630 2283.800 592.950 ;
        RECT 2076.540 588.550 2076.800 588.870 ;
        RECT 2090.800 588.550 2091.060 588.870 ;
        RECT 2090.860 586.490 2091.000 588.550 ;
        RECT 2173.140 588.210 2173.400 588.530 ;
        RECT 2221.900 588.440 2222.160 588.530 ;
        RECT 2222.420 588.440 2222.560 592.630 ;
        RECT 2283.600 588.530 2283.740 592.630 ;
        RECT 2334.140 590.250 2334.400 590.570 ;
        RECT 2380.140 590.250 2380.400 590.570 ;
        RECT 2334.200 588.725 2334.340 590.250 ;
        RECT 2221.900 588.300 2222.560 588.440 ;
        RECT 2221.900 588.210 2222.160 588.300 ;
        RECT 2283.540 588.210 2283.800 588.530 ;
        RECT 2318.490 588.355 2318.770 588.725 ;
        RECT 2334.130 588.355 2334.410 588.725 ;
        RECT 2380.200 588.530 2380.340 590.250 ;
        RECT 2462.940 588.890 2463.200 589.210 ;
        RECT 2466.620 588.890 2466.880 589.210 ;
        RECT 2463.000 588.725 2463.140 588.890 ;
        RECT 2318.500 588.210 2318.760 588.355 ;
        RECT 2380.140 588.210 2380.400 588.530 ;
        RECT 2415.090 588.355 2415.370 588.725 ;
        RECT 2462.930 588.355 2463.210 588.725 ;
        RECT 2415.100 588.210 2415.360 588.355 ;
        RECT 2090.800 586.170 2091.060 586.490 ;
        RECT 2125.300 586.170 2125.560 586.490 ;
        RECT 2125.360 585.810 2125.500 586.170 ;
        RECT 2173.200 585.810 2173.340 588.210 ;
        RECT 2125.300 585.490 2125.560 585.810 ;
        RECT 2173.140 585.490 2173.400 585.810 ;
        RECT 2466.680 16.990 2466.820 588.890 ;
        RECT 2466.620 16.670 2466.880 16.990 ;
        RECT 2479.960 16.670 2480.220 16.990 ;
        RECT 2480.020 16.220 2480.160 16.670 ;
        RECT 2480.940 16.420 2483.380 16.560 ;
        RECT 2480.940 16.220 2481.080 16.420 ;
        RECT 2480.020 16.080 2481.080 16.220 ;
        RECT 2483.240 15.970 2483.380 16.420 ;
        RECT 2483.180 15.650 2483.440 15.970 ;
        RECT 2732.500 15.650 2732.760 15.970 ;
        RECT 2732.560 2.400 2732.700 15.650 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
      LAYER via2 ;
        RECT 2318.490 588.400 2318.770 588.680 ;
        RECT 2334.130 588.400 2334.410 588.680 ;
        RECT 2415.090 588.400 2415.370 588.680 ;
        RECT 2462.930 588.400 2463.210 588.680 ;
      LAYER met3 ;
        RECT 2318.465 588.690 2318.795 588.705 ;
        RECT 2334.105 588.690 2334.435 588.705 ;
        RECT 2318.465 588.390 2334.435 588.690 ;
        RECT 2318.465 588.375 2318.795 588.390 ;
        RECT 2334.105 588.375 2334.435 588.390 ;
        RECT 2415.065 588.690 2415.395 588.705 ;
        RECT 2462.905 588.690 2463.235 588.705 ;
        RECT 2415.065 588.390 2463.235 588.690 ;
        RECT 2415.065 588.375 2415.395 588.390 ;
        RECT 2462.905 588.375 2463.235 588.390 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2085.480 598.980 2085.800 599.040 ;
        RECT 2111.930 598.980 2112.250 599.040 ;
        RECT 2085.480 598.840 2112.250 598.980 ;
        RECT 2085.480 598.780 2085.800 598.840 ;
        RECT 2111.930 598.780 2112.250 598.840 ;
        RECT 2111.930 587.760 2112.250 587.820 ;
        RECT 2480.390 587.760 2480.710 587.820 ;
        RECT 2111.930 587.620 2480.710 587.760 ;
        RECT 2111.930 587.560 2112.250 587.620 ;
        RECT 2480.390 587.560 2480.710 587.620 ;
        RECT 2480.390 16.900 2480.710 16.960 ;
        RECT 2480.390 16.760 2521.560 16.900 ;
        RECT 2480.390 16.700 2480.710 16.760 ;
        RECT 2521.420 16.220 2521.560 16.760 ;
        RECT 2750.410 16.220 2750.730 16.280 ;
        RECT 2521.420 16.080 2750.730 16.220 ;
        RECT 2750.410 16.020 2750.730 16.080 ;
      LAYER via ;
        RECT 2085.510 598.780 2085.770 599.040 ;
        RECT 2111.960 598.780 2112.220 599.040 ;
        RECT 2111.960 587.560 2112.220 587.820 ;
        RECT 2480.420 587.560 2480.680 587.820 ;
        RECT 2480.420 16.700 2480.680 16.960 ;
        RECT 2750.440 16.020 2750.700 16.280 ;
      LAYER met2 ;
        RECT 2085.510 600.000 2085.790 604.000 ;
        RECT 2085.570 599.070 2085.710 600.000 ;
        RECT 2085.510 598.750 2085.770 599.070 ;
        RECT 2111.960 598.750 2112.220 599.070 ;
        RECT 2112.020 587.850 2112.160 598.750 ;
        RECT 2111.960 587.530 2112.220 587.850 ;
        RECT 2480.420 587.530 2480.680 587.850 ;
        RECT 2480.480 16.990 2480.620 587.530 ;
        RECT 2480.420 16.670 2480.680 16.990 ;
        RECT 2750.440 15.990 2750.700 16.310 ;
        RECT 2750.500 2.400 2750.640 15.990 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2096.290 587.760 2096.610 587.820 ;
        RECT 2100.890 587.760 2101.210 587.820 ;
        RECT 2096.290 587.620 2101.210 587.760 ;
        RECT 2096.290 587.560 2096.610 587.620 ;
        RECT 2100.890 587.560 2101.210 587.620 ;
        RECT 2100.890 18.600 2101.210 18.660 ;
        RECT 2100.890 18.460 2112.160 18.600 ;
        RECT 2100.890 18.400 2101.210 18.460 ;
        RECT 2112.020 18.260 2112.160 18.460 ;
        RECT 2767.890 18.260 2768.210 18.320 ;
        RECT 2112.020 18.120 2768.210 18.260 ;
        RECT 2767.890 18.060 2768.210 18.120 ;
      LAYER via ;
        RECT 2096.320 587.560 2096.580 587.820 ;
        RECT 2100.920 587.560 2101.180 587.820 ;
        RECT 2100.920 18.400 2101.180 18.660 ;
        RECT 2767.920 18.060 2768.180 18.320 ;
      LAYER met2 ;
        RECT 2094.710 600.170 2094.990 604.000 ;
        RECT 2094.710 600.030 2096.520 600.170 ;
        RECT 2094.710 600.000 2094.990 600.030 ;
        RECT 2096.380 587.850 2096.520 600.030 ;
        RECT 2096.320 587.530 2096.580 587.850 ;
        RECT 2100.920 587.530 2101.180 587.850 ;
        RECT 2100.980 18.690 2101.120 587.530 ;
        RECT 2100.920 18.370 2101.180 18.690 ;
        RECT 2767.920 18.030 2768.180 18.350 ;
        RECT 2767.980 2.400 2768.120 18.030 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 880.050 591.500 880.370 591.560 ;
        RECT 1101.310 591.500 1101.630 591.560 ;
        RECT 880.050 591.360 1101.630 591.500 ;
        RECT 880.050 591.300 880.370 591.360 ;
        RECT 1101.310 591.300 1101.630 591.360 ;
        RECT 840.950 19.960 841.270 20.020 ;
        RECT 880.050 19.960 880.370 20.020 ;
        RECT 840.950 19.820 880.370 19.960 ;
        RECT 840.950 19.760 841.270 19.820 ;
        RECT 880.050 19.760 880.370 19.820 ;
      LAYER via ;
        RECT 880.080 591.300 880.340 591.560 ;
        RECT 1101.340 591.300 1101.600 591.560 ;
        RECT 840.980 19.760 841.240 20.020 ;
        RECT 880.080 19.760 880.340 20.020 ;
      LAYER met2 ;
        RECT 1102.950 600.170 1103.230 604.000 ;
        RECT 1101.400 600.030 1103.230 600.170 ;
        RECT 1101.400 591.590 1101.540 600.030 ;
        RECT 1102.950 600.000 1103.230 600.030 ;
        RECT 880.080 591.270 880.340 591.590 ;
        RECT 1101.340 591.270 1101.600 591.590 ;
        RECT 880.140 20.050 880.280 591.270 ;
        RECT 840.980 19.730 841.240 20.050 ;
        RECT 880.080 19.730 880.340 20.050 ;
        RECT 841.040 2.400 841.180 19.730 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2104.110 589.460 2104.430 589.520 ;
        RECT 2501.090 589.460 2501.410 589.520 ;
        RECT 2104.110 589.320 2501.410 589.460 ;
        RECT 2104.110 589.260 2104.430 589.320 ;
        RECT 2501.090 589.260 2501.410 589.320 ;
        RECT 2501.090 20.640 2501.410 20.700 ;
        RECT 2522.710 20.640 2523.030 20.700 ;
        RECT 2501.090 20.500 2523.030 20.640 ;
        RECT 2501.090 20.440 2501.410 20.500 ;
        RECT 2522.710 20.440 2523.030 20.500 ;
        RECT 2522.710 16.560 2523.030 16.620 ;
        RECT 2785.830 16.560 2786.150 16.620 ;
        RECT 2522.710 16.420 2786.150 16.560 ;
        RECT 2522.710 16.360 2523.030 16.420 ;
        RECT 2785.830 16.360 2786.150 16.420 ;
      LAYER via ;
        RECT 2104.140 589.260 2104.400 589.520 ;
        RECT 2501.120 589.260 2501.380 589.520 ;
        RECT 2501.120 20.440 2501.380 20.700 ;
        RECT 2522.740 20.440 2523.000 20.700 ;
        RECT 2522.740 16.360 2523.000 16.620 ;
        RECT 2785.860 16.360 2786.120 16.620 ;
      LAYER met2 ;
        RECT 2103.910 600.000 2104.190 604.000 ;
        RECT 2103.970 598.810 2104.110 600.000 ;
        RECT 2103.970 598.670 2104.340 598.810 ;
        RECT 2104.200 589.550 2104.340 598.670 ;
        RECT 2104.140 589.230 2104.400 589.550 ;
        RECT 2501.120 589.230 2501.380 589.550 ;
        RECT 2501.180 20.730 2501.320 589.230 ;
        RECT 2501.120 20.410 2501.380 20.730 ;
        RECT 2522.740 20.410 2523.000 20.730 ;
        RECT 2522.800 16.650 2522.940 20.410 ;
        RECT 2522.740 16.330 2523.000 16.650 ;
        RECT 2785.860 16.330 2786.120 16.650 ;
        RECT 2785.920 2.400 2786.060 16.330 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2114.690 588.440 2115.010 588.500 ;
        RECT 2121.590 588.440 2121.910 588.500 ;
        RECT 2114.690 588.300 2121.910 588.440 ;
        RECT 2114.690 588.240 2115.010 588.300 ;
        RECT 2121.590 588.240 2121.910 588.300 ;
        RECT 2121.590 17.920 2121.910 17.980 ;
        RECT 2803.770 17.920 2804.090 17.980 ;
        RECT 2121.590 17.780 2804.090 17.920 ;
        RECT 2121.590 17.720 2121.910 17.780 ;
        RECT 2803.770 17.720 2804.090 17.780 ;
      LAYER via ;
        RECT 2114.720 588.240 2114.980 588.500 ;
        RECT 2121.620 588.240 2121.880 588.500 ;
        RECT 2121.620 17.720 2121.880 17.980 ;
        RECT 2803.800 17.720 2804.060 17.980 ;
      LAYER met2 ;
        RECT 2113.110 600.170 2113.390 604.000 ;
        RECT 2113.110 600.030 2114.920 600.170 ;
        RECT 2113.110 600.000 2113.390 600.030 ;
        RECT 2114.780 588.530 2114.920 600.030 ;
        RECT 2114.720 588.210 2114.980 588.530 ;
        RECT 2121.620 588.210 2121.880 588.530 ;
        RECT 2121.680 18.010 2121.820 588.210 ;
        RECT 2121.620 17.690 2121.880 18.010 ;
        RECT 2803.800 17.690 2804.060 18.010 ;
        RECT 2803.860 2.400 2804.000 17.690 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2123.890 593.540 2124.210 593.600 ;
        RECT 2123.890 593.400 2127.340 593.540 ;
        RECT 2123.890 593.340 2124.210 593.400 ;
        RECT 2127.200 593.200 2127.340 593.400 ;
        RECT 2131.340 593.400 2149.880 593.540 ;
        RECT 2131.340 593.200 2131.480 593.400 ;
        RECT 2127.200 593.060 2131.480 593.200 ;
        RECT 2149.740 593.200 2149.880 593.400 ;
        RECT 2157.930 593.200 2158.250 593.260 ;
        RECT 2149.740 593.060 2158.250 593.200 ;
        RECT 2157.930 593.000 2158.250 593.060 ;
        RECT 2163.450 588.780 2163.770 588.840 ;
        RECT 2428.410 588.780 2428.730 588.840 ;
        RECT 2163.450 588.640 2428.730 588.780 ;
        RECT 2163.450 588.580 2163.770 588.640 ;
        RECT 2428.410 588.580 2428.730 588.640 ;
        RECT 2429.330 588.780 2429.650 588.840 ;
        RECT 2514.890 588.780 2515.210 588.840 ;
        RECT 2429.330 588.640 2515.210 588.780 ;
        RECT 2429.330 588.580 2429.650 588.640 ;
        RECT 2514.890 588.580 2515.210 588.640 ;
        RECT 2157.930 587.420 2158.250 587.480 ;
        RECT 2163.450 587.420 2163.770 587.480 ;
        RECT 2157.930 587.280 2163.770 587.420 ;
        RECT 2157.930 587.220 2158.250 587.280 ;
        RECT 2163.450 587.220 2163.770 587.280 ;
        RECT 2521.790 16.900 2522.110 16.960 ;
        RECT 2821.710 16.900 2822.030 16.960 ;
        RECT 2521.790 16.760 2822.030 16.900 ;
        RECT 2521.790 16.700 2522.110 16.760 ;
        RECT 2821.710 16.700 2822.030 16.760 ;
        RECT 2514.890 16.560 2515.210 16.620 ;
        RECT 2520.870 16.560 2521.190 16.620 ;
        RECT 2514.890 16.420 2521.190 16.560 ;
        RECT 2514.890 16.360 2515.210 16.420 ;
        RECT 2520.870 16.360 2521.190 16.420 ;
      LAYER via ;
        RECT 2123.920 593.340 2124.180 593.600 ;
        RECT 2157.960 593.000 2158.220 593.260 ;
        RECT 2163.480 588.580 2163.740 588.840 ;
        RECT 2428.440 588.580 2428.700 588.840 ;
        RECT 2429.360 588.580 2429.620 588.840 ;
        RECT 2514.920 588.580 2515.180 588.840 ;
        RECT 2157.960 587.220 2158.220 587.480 ;
        RECT 2163.480 587.220 2163.740 587.480 ;
        RECT 2521.820 16.700 2522.080 16.960 ;
        RECT 2821.740 16.700 2822.000 16.960 ;
        RECT 2514.920 16.360 2515.180 16.620 ;
        RECT 2520.900 16.360 2521.160 16.620 ;
      LAYER met2 ;
        RECT 2122.310 600.170 2122.590 604.000 ;
        RECT 2122.310 600.030 2124.120 600.170 ;
        RECT 2122.310 600.000 2122.590 600.030 ;
        RECT 2123.980 593.630 2124.120 600.030 ;
        RECT 2123.920 593.310 2124.180 593.630 ;
        RECT 2157.960 592.970 2158.220 593.290 ;
        RECT 2158.020 587.510 2158.160 592.970 ;
        RECT 2163.480 588.550 2163.740 588.870 ;
        RECT 2428.440 588.610 2428.700 588.870 ;
        RECT 2429.360 588.610 2429.620 588.870 ;
        RECT 2428.440 588.550 2429.620 588.610 ;
        RECT 2514.920 588.550 2515.180 588.870 ;
        RECT 2163.540 587.510 2163.680 588.550 ;
        RECT 2428.500 588.470 2429.560 588.550 ;
        RECT 2157.960 587.190 2158.220 587.510 ;
        RECT 2163.480 587.190 2163.740 587.510 ;
        RECT 2514.980 16.650 2515.120 588.550 ;
        RECT 2521.820 16.730 2522.080 16.990 ;
        RECT 2520.960 16.670 2522.080 16.730 ;
        RECT 2821.740 16.670 2822.000 16.990 ;
        RECT 2520.960 16.650 2522.020 16.670 ;
        RECT 2514.920 16.330 2515.180 16.650 ;
        RECT 2520.900 16.590 2522.020 16.650 ;
        RECT 2520.900 16.330 2521.160 16.590 ;
        RECT 2821.800 2.400 2821.940 16.670 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2131.710 593.200 2132.030 593.260 ;
        RECT 2149.190 593.200 2149.510 593.260 ;
        RECT 2131.710 593.060 2149.510 593.200 ;
        RECT 2131.710 593.000 2132.030 593.060 ;
        RECT 2149.190 593.000 2149.510 593.060 ;
        RECT 2162.070 17.580 2162.390 17.640 ;
        RECT 2839.190 17.580 2839.510 17.640 ;
        RECT 2162.070 17.440 2839.510 17.580 ;
        RECT 2162.070 17.380 2162.390 17.440 ;
        RECT 2839.190 17.380 2839.510 17.440 ;
        RECT 2149.190 14.860 2149.510 14.920 ;
        RECT 2162.070 14.860 2162.390 14.920 ;
        RECT 2149.190 14.720 2162.390 14.860 ;
        RECT 2149.190 14.660 2149.510 14.720 ;
        RECT 2162.070 14.660 2162.390 14.720 ;
      LAYER via ;
        RECT 2131.740 593.000 2132.000 593.260 ;
        RECT 2149.220 593.000 2149.480 593.260 ;
        RECT 2162.100 17.380 2162.360 17.640 ;
        RECT 2839.220 17.380 2839.480 17.640 ;
        RECT 2149.220 14.660 2149.480 14.920 ;
        RECT 2162.100 14.660 2162.360 14.920 ;
      LAYER met2 ;
        RECT 2131.510 600.000 2131.790 604.000 ;
        RECT 2131.570 598.810 2131.710 600.000 ;
        RECT 2131.570 598.670 2131.940 598.810 ;
        RECT 2131.800 593.290 2131.940 598.670 ;
        RECT 2131.740 592.970 2132.000 593.290 ;
        RECT 2149.220 592.970 2149.480 593.290 ;
        RECT 2149.280 14.950 2149.420 592.970 ;
        RECT 2162.100 17.350 2162.360 17.670 ;
        RECT 2839.220 17.350 2839.480 17.670 ;
        RECT 2162.160 14.950 2162.300 17.350 ;
        RECT 2149.220 14.630 2149.480 14.950 ;
        RECT 2162.100 14.630 2162.360 14.950 ;
        RECT 2839.280 2.400 2839.420 17.350 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2142.290 587.420 2142.610 587.480 ;
        RECT 2151.030 587.420 2151.350 587.480 ;
        RECT 2142.290 587.280 2151.350 587.420 ;
        RECT 2142.290 587.220 2142.610 587.280 ;
        RECT 2151.030 587.220 2151.350 587.280 ;
        RECT 2166.670 587.420 2166.990 587.480 ;
        RECT 2535.590 587.420 2535.910 587.480 ;
        RECT 2166.670 587.280 2535.910 587.420 ;
        RECT 2166.670 587.220 2166.990 587.280 ;
        RECT 2535.590 587.220 2535.910 587.280 ;
        RECT 2151.030 586.400 2151.350 586.460 ;
        RECT 2166.670 586.400 2166.990 586.460 ;
        RECT 2151.030 586.260 2166.990 586.400 ;
        RECT 2151.030 586.200 2151.350 586.260 ;
        RECT 2166.670 586.200 2166.990 586.260 ;
        RECT 2535.590 20.640 2535.910 20.700 ;
        RECT 2857.130 20.640 2857.450 20.700 ;
        RECT 2535.590 20.500 2857.450 20.640 ;
        RECT 2535.590 20.440 2535.910 20.500 ;
        RECT 2857.130 20.440 2857.450 20.500 ;
      LAYER via ;
        RECT 2142.320 587.220 2142.580 587.480 ;
        RECT 2151.060 587.220 2151.320 587.480 ;
        RECT 2166.700 587.220 2166.960 587.480 ;
        RECT 2535.620 587.220 2535.880 587.480 ;
        RECT 2151.060 586.200 2151.320 586.460 ;
        RECT 2166.700 586.200 2166.960 586.460 ;
        RECT 2535.620 20.440 2535.880 20.700 ;
        RECT 2857.160 20.440 2857.420 20.700 ;
      LAYER met2 ;
        RECT 2140.710 600.170 2140.990 604.000 ;
        RECT 2140.710 600.030 2142.520 600.170 ;
        RECT 2140.710 600.000 2140.990 600.030 ;
        RECT 2142.380 587.510 2142.520 600.030 ;
        RECT 2142.320 587.190 2142.580 587.510 ;
        RECT 2151.060 587.190 2151.320 587.510 ;
        RECT 2166.700 587.190 2166.960 587.510 ;
        RECT 2535.620 587.190 2535.880 587.510 ;
        RECT 2151.120 586.490 2151.260 587.190 ;
        RECT 2166.760 586.490 2166.900 587.190 ;
        RECT 2151.060 586.170 2151.320 586.490 ;
        RECT 2166.700 586.170 2166.960 586.490 ;
        RECT 2535.680 20.730 2535.820 587.190 ;
        RECT 2535.620 20.410 2535.880 20.730 ;
        RECT 2857.160 20.410 2857.420 20.730 ;
        RECT 2857.220 2.400 2857.360 20.410 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2151.490 587.420 2151.810 587.480 ;
        RECT 2156.090 587.420 2156.410 587.480 ;
        RECT 2151.490 587.280 2156.410 587.420 ;
        RECT 2151.490 587.220 2151.810 587.280 ;
        RECT 2156.090 587.220 2156.410 587.280 ;
      LAYER via ;
        RECT 2151.520 587.220 2151.780 587.480 ;
        RECT 2156.120 587.220 2156.380 587.480 ;
      LAYER met2 ;
        RECT 2149.910 600.170 2150.190 604.000 ;
        RECT 2149.910 600.030 2151.720 600.170 ;
        RECT 2149.910 600.000 2150.190 600.030 ;
        RECT 2151.580 587.510 2151.720 600.030 ;
        RECT 2151.520 587.190 2151.780 587.510 ;
        RECT 2156.120 587.190 2156.380 587.510 ;
        RECT 2156.180 16.845 2156.320 587.190 ;
        RECT 2156.110 16.475 2156.390 16.845 ;
        RECT 2875.090 16.475 2875.370 16.845 ;
        RECT 2875.160 2.400 2875.300 16.475 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 2156.110 16.520 2156.390 16.800 ;
        RECT 2875.090 16.520 2875.370 16.800 ;
      LAYER met3 ;
        RECT 2156.085 16.810 2156.415 16.825 ;
        RECT 2875.065 16.810 2875.395 16.825 ;
        RECT 2156.085 16.510 2875.395 16.810 ;
        RECT 2156.085 16.495 2156.415 16.510 ;
        RECT 2875.065 16.495 2875.395 16.510 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2158.850 593.200 2159.170 593.260 ;
        RECT 2556.290 593.200 2556.610 593.260 ;
        RECT 2158.850 593.060 2556.610 593.200 ;
        RECT 2158.850 593.000 2159.170 593.060 ;
        RECT 2556.290 593.000 2556.610 593.060 ;
        RECT 2556.290 20.300 2556.610 20.360 ;
        RECT 2893.010 20.300 2893.330 20.360 ;
        RECT 2556.290 20.160 2893.330 20.300 ;
        RECT 2556.290 20.100 2556.610 20.160 ;
        RECT 2893.010 20.100 2893.330 20.160 ;
      LAYER via ;
        RECT 2158.880 593.000 2159.140 593.260 ;
        RECT 2556.320 593.000 2556.580 593.260 ;
        RECT 2556.320 20.100 2556.580 20.360 ;
        RECT 2893.040 20.100 2893.300 20.360 ;
      LAYER met2 ;
        RECT 2159.110 600.000 2159.390 604.000 ;
        RECT 2159.170 598.810 2159.310 600.000 ;
        RECT 2158.940 598.670 2159.310 598.810 ;
        RECT 2158.940 593.290 2159.080 598.670 ;
        RECT 2158.880 592.970 2159.140 593.290 ;
        RECT 2556.320 592.970 2556.580 593.290 ;
        RECT 2556.380 20.390 2556.520 592.970 ;
        RECT 2556.320 20.070 2556.580 20.390 ;
        RECT 2893.040 20.070 2893.300 20.390 ;
        RECT 2893.100 2.400 2893.240 20.070 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2211.290 17.240 2211.610 17.300 ;
        RECT 2910.950 17.240 2911.270 17.300 ;
        RECT 2211.290 17.100 2911.270 17.240 ;
        RECT 2211.290 17.040 2211.610 17.100 ;
        RECT 2910.950 17.040 2911.270 17.100 ;
      LAYER via ;
        RECT 2211.320 17.040 2211.580 17.300 ;
        RECT 2910.980 17.040 2911.240 17.300 ;
      LAYER met2 ;
        RECT 2168.310 600.170 2168.590 604.000 ;
        RECT 2168.310 600.030 2170.120 600.170 ;
        RECT 2168.310 600.000 2168.590 600.030 ;
        RECT 2169.980 590.085 2170.120 600.030 ;
        RECT 2169.910 589.715 2170.190 590.085 ;
        RECT 2211.310 589.715 2211.590 590.085 ;
        RECT 2211.380 17.330 2211.520 589.715 ;
        RECT 2211.320 17.010 2211.580 17.330 ;
        RECT 2910.980 17.010 2911.240 17.330 ;
        RECT 2911.040 2.400 2911.180 17.010 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 2169.910 589.760 2170.190 590.040 ;
        RECT 2211.310 589.760 2211.590 590.040 ;
      LAYER met3 ;
        RECT 2169.885 590.050 2170.215 590.065 ;
        RECT 2211.285 590.050 2211.615 590.065 ;
        RECT 2169.885 589.750 2211.615 590.050 ;
        RECT 2169.885 589.735 2170.215 589.750 ;
        RECT 2211.285 589.735 2211.615 589.750 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 872.690 589.800 873.010 589.860 ;
        RECT 1110.970 589.800 1111.290 589.860 ;
        RECT 872.690 589.660 1111.290 589.800 ;
        RECT 872.690 589.600 873.010 589.660 ;
        RECT 1110.970 589.600 1111.290 589.660 ;
        RECT 858.890 20.640 859.210 20.700 ;
        RECT 872.690 20.640 873.010 20.700 ;
        RECT 858.890 20.500 873.010 20.640 ;
        RECT 858.890 20.440 859.210 20.500 ;
        RECT 872.690 20.440 873.010 20.500 ;
      LAYER via ;
        RECT 872.720 589.600 872.980 589.860 ;
        RECT 1111.000 589.600 1111.260 589.860 ;
        RECT 858.920 20.440 859.180 20.700 ;
        RECT 872.720 20.440 872.980 20.700 ;
      LAYER met2 ;
        RECT 1112.150 600.170 1112.430 604.000 ;
        RECT 1111.060 600.030 1112.430 600.170 ;
        RECT 1111.060 589.890 1111.200 600.030 ;
        RECT 1112.150 600.000 1112.430 600.030 ;
        RECT 872.720 589.570 872.980 589.890 ;
        RECT 1111.000 589.570 1111.260 589.890 ;
        RECT 872.780 20.730 872.920 589.570 ;
        RECT 858.920 20.410 859.180 20.730 ;
        RECT 872.720 20.410 872.980 20.730 ;
        RECT 858.980 2.400 859.120 20.410 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 886.490 590.820 886.810 590.880 ;
        RECT 1119.710 590.820 1120.030 590.880 ;
        RECT 886.490 590.680 1120.030 590.820 ;
        RECT 886.490 590.620 886.810 590.680 ;
        RECT 1119.710 590.620 1120.030 590.680 ;
        RECT 876.830 17.580 877.150 17.640 ;
        RECT 886.490 17.580 886.810 17.640 ;
        RECT 876.830 17.440 886.810 17.580 ;
        RECT 876.830 17.380 877.150 17.440 ;
        RECT 886.490 17.380 886.810 17.440 ;
      LAYER via ;
        RECT 886.520 590.620 886.780 590.880 ;
        RECT 1119.740 590.620 1120.000 590.880 ;
        RECT 876.860 17.380 877.120 17.640 ;
        RECT 886.520 17.380 886.780 17.640 ;
      LAYER met2 ;
        RECT 1121.350 600.170 1121.630 604.000 ;
        RECT 1119.800 600.030 1121.630 600.170 ;
        RECT 1119.800 590.910 1119.940 600.030 ;
        RECT 1121.350 600.000 1121.630 600.030 ;
        RECT 886.520 590.590 886.780 590.910 ;
        RECT 1119.740 590.590 1120.000 590.910 ;
        RECT 886.580 17.670 886.720 590.590 ;
        RECT 876.860 17.350 877.120 17.670 ;
        RECT 886.520 17.350 886.780 17.670 ;
        RECT 876.920 2.400 877.060 17.350 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.610 591.160 896.930 591.220 ;
        RECT 1128.910 591.160 1129.230 591.220 ;
        RECT 896.610 591.020 1129.230 591.160 ;
        RECT 896.610 590.960 896.930 591.020 ;
        RECT 1128.910 590.960 1129.230 591.020 ;
        RECT 894.770 2.960 895.090 3.020 ;
        RECT 896.610 2.960 896.930 3.020 ;
        RECT 894.770 2.820 896.930 2.960 ;
        RECT 894.770 2.760 895.090 2.820 ;
        RECT 896.610 2.760 896.930 2.820 ;
      LAYER via ;
        RECT 896.640 590.960 896.900 591.220 ;
        RECT 1128.940 590.960 1129.200 591.220 ;
        RECT 894.800 2.760 895.060 3.020 ;
        RECT 896.640 2.760 896.900 3.020 ;
      LAYER met2 ;
        RECT 1130.550 600.170 1130.830 604.000 ;
        RECT 1129.000 600.030 1130.830 600.170 ;
        RECT 1129.000 591.250 1129.140 600.030 ;
        RECT 1130.550 600.000 1130.830 600.030 ;
        RECT 896.640 590.930 896.900 591.250 ;
        RECT 1128.940 590.930 1129.200 591.250 ;
        RECT 896.700 3.050 896.840 590.930 ;
        RECT 894.800 2.730 895.060 3.050 ;
        RECT 896.640 2.730 896.900 3.050 ;
        RECT 894.860 2.400 895.000 2.730 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 590.140 917.630 590.200 ;
        RECT 1138.570 590.140 1138.890 590.200 ;
        RECT 917.310 590.000 1138.890 590.140 ;
        RECT 917.310 589.940 917.630 590.000 ;
        RECT 1138.570 589.940 1138.890 590.000 ;
        RECT 912.710 16.560 913.030 16.620 ;
        RECT 917.310 16.560 917.630 16.620 ;
        RECT 912.710 16.420 917.630 16.560 ;
        RECT 912.710 16.360 913.030 16.420 ;
        RECT 917.310 16.360 917.630 16.420 ;
      LAYER via ;
        RECT 917.340 589.940 917.600 590.200 ;
        RECT 1138.600 589.940 1138.860 590.200 ;
        RECT 912.740 16.360 913.000 16.620 ;
        RECT 917.340 16.360 917.600 16.620 ;
      LAYER met2 ;
        RECT 1139.750 600.170 1140.030 604.000 ;
        RECT 1138.660 600.030 1140.030 600.170 ;
        RECT 1138.660 590.230 1138.800 600.030 ;
        RECT 1139.750 600.000 1140.030 600.030 ;
        RECT 917.340 589.910 917.600 590.230 ;
        RECT 1138.600 589.910 1138.860 590.230 ;
        RECT 917.400 16.650 917.540 589.910 ;
        RECT 912.740 16.330 913.000 16.650 ;
        RECT 917.340 16.330 917.600 16.650 ;
        RECT 912.800 2.400 912.940 16.330 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.110 591.840 931.430 591.900 ;
        RECT 1147.310 591.840 1147.630 591.900 ;
        RECT 931.110 591.700 1147.630 591.840 ;
        RECT 931.110 591.640 931.430 591.700 ;
        RECT 1147.310 591.640 1147.630 591.700 ;
        RECT 931.110 579.600 931.430 579.660 ;
        RECT 931.570 579.600 931.890 579.660 ;
        RECT 931.110 579.460 931.890 579.600 ;
        RECT 931.110 579.400 931.430 579.460 ;
        RECT 931.570 579.400 931.890 579.460 ;
        RECT 931.110 531.660 931.430 531.720 ;
        RECT 931.570 531.660 931.890 531.720 ;
        RECT 931.110 531.520 931.890 531.660 ;
        RECT 931.110 531.460 931.430 531.520 ;
        RECT 931.570 531.460 931.890 531.520 ;
        RECT 930.190 524.180 930.510 524.240 ;
        RECT 931.110 524.180 931.430 524.240 ;
        RECT 930.190 524.040 931.430 524.180 ;
        RECT 930.190 523.980 930.510 524.040 ;
        RECT 931.110 523.980 931.430 524.040 ;
        RECT 930.190 476.240 930.510 476.300 ;
        RECT 931.110 476.240 931.430 476.300 ;
        RECT 930.190 476.100 931.430 476.240 ;
        RECT 930.190 476.040 930.510 476.100 ;
        RECT 931.110 476.040 931.430 476.100 ;
        RECT 930.650 289.580 930.970 289.640 ;
        RECT 931.110 289.580 931.430 289.640 ;
        RECT 930.650 289.440 931.430 289.580 ;
        RECT 930.650 289.380 930.970 289.440 ;
        RECT 931.110 289.380 931.430 289.440 ;
        RECT 929.730 282.780 930.050 282.840 ;
        RECT 930.650 282.780 930.970 282.840 ;
        RECT 929.730 282.640 930.970 282.780 ;
        RECT 929.730 282.580 930.050 282.640 ;
        RECT 930.650 282.580 930.970 282.640 ;
        RECT 930.650 234.500 930.970 234.560 ;
        RECT 931.110 234.500 931.430 234.560 ;
        RECT 930.650 234.360 931.430 234.500 ;
        RECT 930.650 234.300 930.970 234.360 ;
        RECT 931.110 234.300 931.430 234.360 ;
        RECT 930.650 186.560 930.970 186.620 ;
        RECT 931.110 186.560 931.430 186.620 ;
        RECT 930.650 186.420 931.430 186.560 ;
        RECT 930.650 186.360 930.970 186.420 ;
        RECT 931.110 186.360 931.430 186.420 ;
        RECT 931.110 137.740 931.430 138.000 ;
        RECT 931.200 137.320 931.340 137.740 ;
        RECT 931.110 137.060 931.430 137.320 ;
        RECT 931.110 62.460 931.430 62.520 ;
        RECT 930.280 62.320 931.430 62.460 ;
        RECT 930.280 62.180 930.420 62.320 ;
        RECT 931.110 62.260 931.430 62.320 ;
        RECT 930.190 61.920 930.510 62.180 ;
      LAYER via ;
        RECT 931.140 591.640 931.400 591.900 ;
        RECT 1147.340 591.640 1147.600 591.900 ;
        RECT 931.140 579.400 931.400 579.660 ;
        RECT 931.600 579.400 931.860 579.660 ;
        RECT 931.140 531.460 931.400 531.720 ;
        RECT 931.600 531.460 931.860 531.720 ;
        RECT 930.220 523.980 930.480 524.240 ;
        RECT 931.140 523.980 931.400 524.240 ;
        RECT 930.220 476.040 930.480 476.300 ;
        RECT 931.140 476.040 931.400 476.300 ;
        RECT 930.680 289.380 930.940 289.640 ;
        RECT 931.140 289.380 931.400 289.640 ;
        RECT 929.760 282.580 930.020 282.840 ;
        RECT 930.680 282.580 930.940 282.840 ;
        RECT 930.680 234.300 930.940 234.560 ;
        RECT 931.140 234.300 931.400 234.560 ;
        RECT 930.680 186.360 930.940 186.620 ;
        RECT 931.140 186.360 931.400 186.620 ;
        RECT 931.140 137.740 931.400 138.000 ;
        RECT 931.140 137.060 931.400 137.320 ;
        RECT 931.140 62.260 931.400 62.520 ;
        RECT 930.220 61.920 930.480 62.180 ;
      LAYER met2 ;
        RECT 1148.950 600.170 1149.230 604.000 ;
        RECT 1147.400 600.030 1149.230 600.170 ;
        RECT 1147.400 591.930 1147.540 600.030 ;
        RECT 1148.950 600.000 1149.230 600.030 ;
        RECT 931.140 591.610 931.400 591.930 ;
        RECT 1147.340 591.610 1147.600 591.930 ;
        RECT 931.200 579.690 931.340 591.610 ;
        RECT 931.140 579.370 931.400 579.690 ;
        RECT 931.600 579.370 931.860 579.690 ;
        RECT 931.660 531.750 931.800 579.370 ;
        RECT 931.140 531.430 931.400 531.750 ;
        RECT 931.600 531.430 931.860 531.750 ;
        RECT 931.200 524.270 931.340 531.430 ;
        RECT 930.220 523.950 930.480 524.270 ;
        RECT 931.140 523.950 931.400 524.270 ;
        RECT 930.280 476.330 930.420 523.950 ;
        RECT 930.220 476.010 930.480 476.330 ;
        RECT 931.140 476.010 931.400 476.330 ;
        RECT 931.200 289.670 931.340 476.010 ;
        RECT 930.680 289.350 930.940 289.670 ;
        RECT 931.140 289.350 931.400 289.670 ;
        RECT 930.740 282.870 930.880 289.350 ;
        RECT 929.760 282.550 930.020 282.870 ;
        RECT 930.680 282.550 930.940 282.870 ;
        RECT 929.820 235.125 929.960 282.550 ;
        RECT 929.750 234.755 930.030 235.125 ;
        RECT 931.130 234.755 931.410 235.125 ;
        RECT 931.200 234.590 931.340 234.755 ;
        RECT 930.680 234.270 930.940 234.590 ;
        RECT 931.140 234.270 931.400 234.590 ;
        RECT 930.740 186.650 930.880 234.270 ;
        RECT 930.680 186.330 930.940 186.650 ;
        RECT 931.140 186.330 931.400 186.650 ;
        RECT 931.200 138.030 931.340 186.330 ;
        RECT 931.140 137.710 931.400 138.030 ;
        RECT 931.140 137.030 931.400 137.350 ;
        RECT 931.200 62.550 931.340 137.030 ;
        RECT 931.140 62.230 931.400 62.550 ;
        RECT 930.220 61.890 930.480 62.210 ;
        RECT 930.280 2.400 930.420 61.890 ;
        RECT 930.070 -4.800 930.630 2.400 ;
      LAYER via2 ;
        RECT 929.750 234.800 930.030 235.080 ;
        RECT 931.130 234.800 931.410 235.080 ;
      LAYER met3 ;
        RECT 929.725 235.090 930.055 235.105 ;
        RECT 931.105 235.090 931.435 235.105 ;
        RECT 929.725 234.790 931.435 235.090 ;
        RECT 929.725 234.775 930.055 234.790 ;
        RECT 931.105 234.775 931.435 234.790 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 592.860 952.130 592.920 ;
        RECT 1156.510 592.860 1156.830 592.920 ;
        RECT 951.810 592.720 1156.830 592.860 ;
        RECT 951.810 592.660 952.130 592.720 ;
        RECT 1156.510 592.660 1156.830 592.720 ;
        RECT 948.130 20.640 948.450 20.700 ;
        RECT 951.810 20.640 952.130 20.700 ;
        RECT 948.130 20.500 952.130 20.640 ;
        RECT 948.130 20.440 948.450 20.500 ;
        RECT 951.810 20.440 952.130 20.500 ;
      LAYER via ;
        RECT 951.840 592.660 952.100 592.920 ;
        RECT 1156.540 592.660 1156.800 592.920 ;
        RECT 948.160 20.440 948.420 20.700 ;
        RECT 951.840 20.440 952.100 20.700 ;
      LAYER met2 ;
        RECT 1158.150 600.170 1158.430 604.000 ;
        RECT 1156.600 600.030 1158.430 600.170 ;
        RECT 1156.600 592.950 1156.740 600.030 ;
        RECT 1158.150 600.000 1158.430 600.030 ;
        RECT 951.840 592.630 952.100 592.950 ;
        RECT 1156.540 592.630 1156.800 592.950 ;
        RECT 951.900 20.730 952.040 592.630 ;
        RECT 948.160 20.410 948.420 20.730 ;
        RECT 951.840 20.410 952.100 20.730 ;
        RECT 948.220 2.400 948.360 20.410 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.510 592.180 972.830 592.240 ;
        RECT 1166.170 592.180 1166.490 592.240 ;
        RECT 972.510 592.040 1166.490 592.180 ;
        RECT 972.510 591.980 972.830 592.040 ;
        RECT 1166.170 591.980 1166.490 592.040 ;
        RECT 966.070 16.560 966.390 16.620 ;
        RECT 972.510 16.560 972.830 16.620 ;
        RECT 966.070 16.420 972.830 16.560 ;
        RECT 966.070 16.360 966.390 16.420 ;
        RECT 972.510 16.360 972.830 16.420 ;
      LAYER via ;
        RECT 972.540 591.980 972.800 592.240 ;
        RECT 1166.200 591.980 1166.460 592.240 ;
        RECT 966.100 16.360 966.360 16.620 ;
        RECT 972.540 16.360 972.800 16.620 ;
      LAYER met2 ;
        RECT 1167.350 600.170 1167.630 604.000 ;
        RECT 1166.260 600.030 1167.630 600.170 ;
        RECT 1166.260 592.270 1166.400 600.030 ;
        RECT 1167.350 600.000 1167.630 600.030 ;
        RECT 972.540 591.950 972.800 592.270 ;
        RECT 1166.200 591.950 1166.460 592.270 ;
        RECT 972.600 16.650 972.740 591.950 ;
        RECT 966.100 16.330 966.360 16.650 ;
        RECT 972.540 16.330 972.800 16.650 ;
        RECT 966.160 2.400 966.300 16.330 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 986.310 588.440 986.630 588.500 ;
        RECT 1077.390 588.440 1077.710 588.500 ;
        RECT 986.310 588.300 1077.710 588.440 ;
        RECT 986.310 588.240 986.630 588.300 ;
        RECT 1077.390 588.240 1077.710 588.300 ;
        RECT 1100.390 588.100 1100.710 588.160 ;
        RECT 1152.370 588.100 1152.690 588.160 ;
        RECT 1100.390 587.960 1152.690 588.100 ;
        RECT 1100.390 587.900 1100.710 587.960 ;
        RECT 1152.370 587.900 1152.690 587.960 ;
        RECT 984.010 17.920 984.330 17.980 ;
        RECT 986.310 17.920 986.630 17.980 ;
        RECT 984.010 17.780 986.630 17.920 ;
        RECT 984.010 17.720 984.330 17.780 ;
        RECT 986.310 17.720 986.630 17.780 ;
      LAYER via ;
        RECT 986.340 588.240 986.600 588.500 ;
        RECT 1077.420 588.240 1077.680 588.500 ;
        RECT 1100.420 587.900 1100.680 588.160 ;
        RECT 1152.400 587.900 1152.660 588.160 ;
        RECT 984.040 17.720 984.300 17.980 ;
        RECT 986.340 17.720 986.600 17.980 ;
      LAYER met2 ;
        RECT 1176.550 600.170 1176.830 604.000 ;
        RECT 1175.000 600.030 1176.830 600.170 ;
        RECT 986.340 588.210 986.600 588.530 ;
        RECT 1077.410 588.355 1077.690 588.725 ;
        RECT 1100.410 588.355 1100.690 588.725 ;
        RECT 1077.420 588.210 1077.680 588.355 ;
        RECT 986.400 18.010 986.540 588.210 ;
        RECT 1100.480 588.190 1100.620 588.355 ;
        RECT 1100.420 587.870 1100.680 588.190 ;
        RECT 1152.400 588.045 1152.660 588.190 ;
        RECT 1175.000 588.045 1175.140 600.030 ;
        RECT 1176.550 600.000 1176.830 600.030 ;
        RECT 1152.390 587.675 1152.670 588.045 ;
        RECT 1174.930 587.675 1175.210 588.045 ;
        RECT 984.040 17.690 984.300 18.010 ;
        RECT 986.340 17.690 986.600 18.010 ;
        RECT 984.100 2.400 984.240 17.690 ;
        RECT 983.890 -4.800 984.450 2.400 ;
      LAYER via2 ;
        RECT 1077.410 588.400 1077.690 588.680 ;
        RECT 1100.410 588.400 1100.690 588.680 ;
        RECT 1152.390 587.720 1152.670 588.000 ;
        RECT 1174.930 587.720 1175.210 588.000 ;
      LAYER met3 ;
        RECT 1077.385 588.690 1077.715 588.705 ;
        RECT 1100.385 588.690 1100.715 588.705 ;
        RECT 1077.385 588.390 1100.715 588.690 ;
        RECT 1077.385 588.375 1077.715 588.390 ;
        RECT 1100.385 588.375 1100.715 588.390 ;
        RECT 1152.365 588.010 1152.695 588.025 ;
        RECT 1174.905 588.010 1175.235 588.025 ;
        RECT 1152.365 587.710 1175.235 588.010 ;
        RECT 1152.365 587.695 1152.695 587.710 ;
        RECT 1174.905 587.695 1175.235 587.710 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.470 583.000 1007.790 583.060 ;
        RECT 1009.310 583.000 1009.630 583.060 ;
        RECT 1007.470 582.860 1009.630 583.000 ;
        RECT 1007.470 582.800 1007.790 582.860 ;
        RECT 1009.310 582.800 1009.630 582.860 ;
        RECT 662.930 35.260 663.250 35.320 ;
        RECT 1007.470 35.260 1007.790 35.320 ;
        RECT 662.930 35.120 1007.790 35.260 ;
        RECT 662.930 35.060 663.250 35.120 ;
        RECT 1007.470 35.060 1007.790 35.120 ;
      LAYER via ;
        RECT 1007.500 582.800 1007.760 583.060 ;
        RECT 1009.340 582.800 1009.600 583.060 ;
        RECT 662.960 35.060 663.220 35.320 ;
        RECT 1007.500 35.060 1007.760 35.320 ;
      LAYER met2 ;
        RECT 1010.950 600.170 1011.230 604.000 ;
        RECT 1009.400 600.030 1011.230 600.170 ;
        RECT 1009.400 583.090 1009.540 600.030 ;
        RECT 1010.950 600.000 1011.230 600.030 ;
        RECT 1007.500 582.770 1007.760 583.090 ;
        RECT 1009.340 582.770 1009.600 583.090 ;
        RECT 1007.560 35.350 1007.700 582.770 ;
        RECT 662.960 35.030 663.220 35.350 ;
        RECT 1007.500 35.030 1007.760 35.350 ;
        RECT 663.020 2.400 663.160 35.030 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 587.760 1007.330 587.820 ;
        RECT 1184.110 587.760 1184.430 587.820 ;
        RECT 1007.010 587.620 1184.430 587.760 ;
        RECT 1007.010 587.560 1007.330 587.620 ;
        RECT 1184.110 587.560 1184.430 587.620 ;
        RECT 1001.950 17.920 1002.270 17.980 ;
        RECT 1007.010 17.920 1007.330 17.980 ;
        RECT 1001.950 17.780 1007.330 17.920 ;
        RECT 1001.950 17.720 1002.270 17.780 ;
        RECT 1007.010 17.720 1007.330 17.780 ;
      LAYER via ;
        RECT 1007.040 587.560 1007.300 587.820 ;
        RECT 1184.140 587.560 1184.400 587.820 ;
        RECT 1001.980 17.720 1002.240 17.980 ;
        RECT 1007.040 17.720 1007.300 17.980 ;
      LAYER met2 ;
        RECT 1185.750 600.170 1186.030 604.000 ;
        RECT 1184.200 600.030 1186.030 600.170 ;
        RECT 1184.200 587.850 1184.340 600.030 ;
        RECT 1185.750 600.000 1186.030 600.030 ;
        RECT 1007.040 587.530 1007.300 587.850 ;
        RECT 1184.140 587.530 1184.400 587.850 ;
        RECT 1007.100 18.010 1007.240 587.530 ;
        RECT 1001.980 17.690 1002.240 18.010 ;
        RECT 1007.040 17.690 1007.300 18.010 ;
        RECT 1002.040 2.400 1002.180 17.690 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1169.390 588.780 1169.710 588.840 ;
        RECT 1194.230 588.780 1194.550 588.840 ;
        RECT 1169.390 588.640 1194.550 588.780 ;
        RECT 1169.390 588.580 1169.710 588.640 ;
        RECT 1194.230 588.580 1194.550 588.640 ;
        RECT 1019.430 15.880 1019.750 15.940 ;
        RECT 1169.390 15.880 1169.710 15.940 ;
        RECT 1019.430 15.740 1169.710 15.880 ;
        RECT 1019.430 15.680 1019.750 15.740 ;
        RECT 1169.390 15.680 1169.710 15.740 ;
      LAYER via ;
        RECT 1169.420 588.580 1169.680 588.840 ;
        RECT 1194.260 588.580 1194.520 588.840 ;
        RECT 1019.460 15.680 1019.720 15.940 ;
        RECT 1169.420 15.680 1169.680 15.940 ;
      LAYER met2 ;
        RECT 1194.950 600.170 1195.230 604.000 ;
        RECT 1194.320 600.030 1195.230 600.170 ;
        RECT 1194.320 588.870 1194.460 600.030 ;
        RECT 1194.950 600.000 1195.230 600.030 ;
        RECT 1169.420 588.550 1169.680 588.870 ;
        RECT 1194.260 588.550 1194.520 588.870 ;
        RECT 1169.480 15.970 1169.620 588.550 ;
        RECT 1019.460 15.650 1019.720 15.970 ;
        RECT 1169.420 15.650 1169.680 15.970 ;
        RECT 1019.520 2.400 1019.660 15.650 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1187.790 588.100 1188.110 588.160 ;
        RECT 1202.050 588.100 1202.370 588.160 ;
        RECT 1187.790 587.960 1202.370 588.100 ;
        RECT 1187.790 587.900 1188.110 587.960 ;
        RECT 1202.050 587.900 1202.370 587.960 ;
        RECT 1041.510 587.420 1041.830 587.480 ;
        RECT 1041.510 587.280 1148.920 587.420 ;
        RECT 1041.510 587.220 1041.830 587.280 ;
        RECT 1148.780 586.740 1148.920 587.280 ;
        RECT 1187.790 586.740 1188.110 586.800 ;
        RECT 1148.780 586.600 1188.110 586.740 ;
        RECT 1187.790 586.540 1188.110 586.600 ;
        RECT 1037.370 18.600 1037.690 18.660 ;
        RECT 1041.510 18.600 1041.830 18.660 ;
        RECT 1037.370 18.460 1041.830 18.600 ;
        RECT 1037.370 18.400 1037.690 18.460 ;
        RECT 1041.510 18.400 1041.830 18.460 ;
      LAYER via ;
        RECT 1187.820 587.900 1188.080 588.160 ;
        RECT 1202.080 587.900 1202.340 588.160 ;
        RECT 1041.540 587.220 1041.800 587.480 ;
        RECT 1187.820 586.540 1188.080 586.800 ;
        RECT 1037.400 18.400 1037.660 18.660 ;
        RECT 1041.540 18.400 1041.800 18.660 ;
      LAYER met2 ;
        RECT 1203.690 600.170 1203.970 604.000 ;
        RECT 1202.140 600.030 1203.970 600.170 ;
        RECT 1202.140 588.190 1202.280 600.030 ;
        RECT 1203.690 600.000 1203.970 600.030 ;
        RECT 1187.820 587.870 1188.080 588.190 ;
        RECT 1202.080 587.870 1202.340 588.190 ;
        RECT 1041.540 587.190 1041.800 587.510 ;
        RECT 1041.600 18.690 1041.740 587.190 ;
        RECT 1187.880 586.830 1188.020 587.870 ;
        RECT 1187.820 586.510 1188.080 586.830 ;
        RECT 1037.400 18.370 1037.660 18.690 ;
        RECT 1041.540 18.370 1041.800 18.690 ;
        RECT 1037.460 2.400 1037.600 18.370 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1183.190 587.080 1183.510 587.140 ;
        RECT 1211.250 587.080 1211.570 587.140 ;
        RECT 1183.190 586.940 1211.570 587.080 ;
        RECT 1183.190 586.880 1183.510 586.940 ;
        RECT 1211.250 586.880 1211.570 586.940 ;
        RECT 1148.690 19.620 1149.010 19.680 ;
        RECT 1183.190 19.620 1183.510 19.680 ;
        RECT 1148.690 19.480 1183.510 19.620 ;
        RECT 1148.690 19.420 1149.010 19.480 ;
        RECT 1183.190 19.420 1183.510 19.480 ;
        RECT 1076.930 18.600 1077.250 18.660 ;
        RECT 1076.930 18.460 1099.700 18.600 ;
        RECT 1076.930 18.400 1077.250 18.460 ;
        RECT 1099.560 18.260 1099.700 18.460 ;
        RECT 1099.560 18.120 1119.020 18.260 ;
        RECT 1054.850 17.920 1055.170 17.980 ;
        RECT 1076.470 17.920 1076.790 17.980 ;
        RECT 1054.850 17.780 1076.790 17.920 ;
        RECT 1054.850 17.720 1055.170 17.780 ;
        RECT 1076.470 17.720 1076.790 17.780 ;
        RECT 1118.880 17.580 1119.020 18.120 ;
        RECT 1148.690 17.580 1149.010 17.640 ;
        RECT 1118.880 17.440 1149.010 17.580 ;
        RECT 1148.690 17.380 1149.010 17.440 ;
      LAYER via ;
        RECT 1183.220 586.880 1183.480 587.140 ;
        RECT 1211.280 586.880 1211.540 587.140 ;
        RECT 1148.720 19.420 1148.980 19.680 ;
        RECT 1183.220 19.420 1183.480 19.680 ;
        RECT 1076.960 18.400 1077.220 18.660 ;
        RECT 1054.880 17.720 1055.140 17.980 ;
        RECT 1076.500 17.720 1076.760 17.980 ;
        RECT 1148.720 17.380 1148.980 17.640 ;
      LAYER met2 ;
        RECT 1212.890 600.170 1213.170 604.000 ;
        RECT 1211.340 600.030 1213.170 600.170 ;
        RECT 1211.340 587.170 1211.480 600.030 ;
        RECT 1212.890 600.000 1213.170 600.030 ;
        RECT 1183.220 586.850 1183.480 587.170 ;
        RECT 1211.280 586.850 1211.540 587.170 ;
        RECT 1183.280 19.710 1183.420 586.850 ;
        RECT 1148.720 19.390 1148.980 19.710 ;
        RECT 1183.220 19.390 1183.480 19.710 ;
        RECT 1076.960 18.370 1077.220 18.690 ;
        RECT 1077.020 18.090 1077.160 18.370 ;
        RECT 1076.560 18.010 1077.160 18.090 ;
        RECT 1054.880 17.690 1055.140 18.010 ;
        RECT 1076.500 17.950 1077.160 18.010 ;
        RECT 1076.500 17.690 1076.760 17.950 ;
        RECT 1054.940 9.250 1055.080 17.690 ;
        RECT 1148.780 17.670 1148.920 19.390 ;
        RECT 1148.720 17.350 1148.980 17.670 ;
        RECT 1054.940 9.110 1055.540 9.250 ;
        RECT 1055.400 2.400 1055.540 9.110 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.990 586.740 1197.310 586.800 ;
        RECT 1221.370 586.740 1221.690 586.800 ;
        RECT 1196.990 586.600 1221.690 586.740 ;
        RECT 1196.990 586.540 1197.310 586.600 ;
        RECT 1221.370 586.540 1221.690 586.600 ;
        RECT 1073.250 14.520 1073.570 14.580 ;
        RECT 1196.990 14.520 1197.310 14.580 ;
        RECT 1073.250 14.380 1197.310 14.520 ;
        RECT 1073.250 14.320 1073.570 14.380 ;
        RECT 1196.990 14.320 1197.310 14.380 ;
      LAYER via ;
        RECT 1197.020 586.540 1197.280 586.800 ;
        RECT 1221.400 586.540 1221.660 586.800 ;
        RECT 1073.280 14.320 1073.540 14.580 ;
        RECT 1197.020 14.320 1197.280 14.580 ;
      LAYER met2 ;
        RECT 1222.090 600.170 1222.370 604.000 ;
        RECT 1221.460 600.030 1222.370 600.170 ;
        RECT 1221.460 586.830 1221.600 600.030 ;
        RECT 1222.090 600.000 1222.370 600.030 ;
        RECT 1197.020 586.510 1197.280 586.830 ;
        RECT 1221.400 586.510 1221.660 586.830 ;
        RECT 1197.080 14.610 1197.220 586.510 ;
        RECT 1073.280 14.290 1073.540 14.610 ;
        RECT 1197.020 14.290 1197.280 14.610 ;
        RECT 1073.340 2.400 1073.480 14.290 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.250 590.480 1096.570 590.540 ;
        RECT 1229.650 590.480 1229.970 590.540 ;
        RECT 1096.250 590.340 1229.970 590.480 ;
        RECT 1096.250 590.280 1096.570 590.340 ;
        RECT 1229.650 590.280 1229.970 590.340 ;
        RECT 1090.730 19.280 1091.050 19.340 ;
        RECT 1096.250 19.280 1096.570 19.340 ;
        RECT 1090.730 19.140 1096.570 19.280 ;
        RECT 1090.730 19.080 1091.050 19.140 ;
        RECT 1096.250 19.080 1096.570 19.140 ;
      LAYER via ;
        RECT 1096.280 590.280 1096.540 590.540 ;
        RECT 1229.680 590.280 1229.940 590.540 ;
        RECT 1090.760 19.080 1091.020 19.340 ;
        RECT 1096.280 19.080 1096.540 19.340 ;
      LAYER met2 ;
        RECT 1231.290 600.170 1231.570 604.000 ;
        RECT 1229.740 600.030 1231.570 600.170 ;
        RECT 1229.740 590.570 1229.880 600.030 ;
        RECT 1231.290 600.000 1231.570 600.030 ;
        RECT 1096.280 590.250 1096.540 590.570 ;
        RECT 1229.680 590.250 1229.940 590.570 ;
        RECT 1096.340 19.370 1096.480 590.250 ;
        RECT 1090.760 19.050 1091.020 19.370 ;
        RECT 1096.280 19.050 1096.540 19.370 ;
        RECT 1090.820 2.400 1090.960 19.050 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 592.520 1204.210 592.580 ;
        RECT 1238.850 592.520 1239.170 592.580 ;
        RECT 1203.890 592.380 1239.170 592.520 ;
        RECT 1203.890 592.320 1204.210 592.380 ;
        RECT 1238.850 592.320 1239.170 592.380 ;
        RECT 1108.670 18.600 1108.990 18.660 ;
        RECT 1203.430 18.600 1203.750 18.660 ;
        RECT 1108.670 18.460 1203.750 18.600 ;
        RECT 1108.670 18.400 1108.990 18.460 ;
        RECT 1203.430 18.400 1203.750 18.460 ;
      LAYER via ;
        RECT 1203.920 592.320 1204.180 592.580 ;
        RECT 1238.880 592.320 1239.140 592.580 ;
        RECT 1108.700 18.400 1108.960 18.660 ;
        RECT 1203.460 18.400 1203.720 18.660 ;
      LAYER met2 ;
        RECT 1240.490 600.170 1240.770 604.000 ;
        RECT 1238.940 600.030 1240.770 600.170 ;
        RECT 1238.940 592.610 1239.080 600.030 ;
        RECT 1240.490 600.000 1240.770 600.030 ;
        RECT 1203.920 592.290 1204.180 592.610 ;
        RECT 1238.880 592.290 1239.140 592.610 ;
        RECT 1203.980 21.490 1204.120 592.290 ;
        RECT 1203.520 21.350 1204.120 21.490 ;
        RECT 1203.520 18.690 1203.660 21.350 ;
        RECT 1108.700 18.370 1108.960 18.690 ;
        RECT 1203.460 18.370 1203.720 18.690 ;
        RECT 1108.760 2.400 1108.900 18.370 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 590.820 1131.530 590.880 ;
        RECT 1248.970 590.820 1249.290 590.880 ;
        RECT 1131.210 590.680 1249.290 590.820 ;
        RECT 1131.210 590.620 1131.530 590.680 ;
        RECT 1248.970 590.620 1249.290 590.680 ;
        RECT 1126.610 16.900 1126.930 16.960 ;
        RECT 1131.210 16.900 1131.530 16.960 ;
        RECT 1126.610 16.760 1131.530 16.900 ;
        RECT 1126.610 16.700 1126.930 16.760 ;
        RECT 1131.210 16.700 1131.530 16.760 ;
      LAYER via ;
        RECT 1131.240 590.620 1131.500 590.880 ;
        RECT 1249.000 590.620 1249.260 590.880 ;
        RECT 1126.640 16.700 1126.900 16.960 ;
        RECT 1131.240 16.700 1131.500 16.960 ;
      LAYER met2 ;
        RECT 1249.690 600.170 1249.970 604.000 ;
        RECT 1249.060 600.030 1249.970 600.170 ;
        RECT 1249.060 590.910 1249.200 600.030 ;
        RECT 1249.690 600.000 1249.970 600.030 ;
        RECT 1131.240 590.590 1131.500 590.910 ;
        RECT 1249.000 590.590 1249.260 590.910 ;
        RECT 1131.300 16.990 1131.440 590.590 ;
        RECT 1126.640 16.670 1126.900 16.990 ;
        RECT 1131.240 16.670 1131.500 16.990 ;
        RECT 1126.700 2.400 1126.840 16.670 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1238.390 587.080 1238.710 587.140 ;
        RECT 1257.250 587.080 1257.570 587.140 ;
        RECT 1238.390 586.940 1257.570 587.080 ;
        RECT 1238.390 586.880 1238.710 586.940 ;
        RECT 1257.250 586.880 1257.570 586.940 ;
        RECT 1144.550 18.260 1144.870 18.320 ;
        RECT 1238.390 18.260 1238.710 18.320 ;
        RECT 1144.550 18.120 1238.710 18.260 ;
        RECT 1144.550 18.060 1144.870 18.120 ;
        RECT 1238.390 18.060 1238.710 18.120 ;
      LAYER via ;
        RECT 1238.420 586.880 1238.680 587.140 ;
        RECT 1257.280 586.880 1257.540 587.140 ;
        RECT 1144.580 18.060 1144.840 18.320 ;
        RECT 1238.420 18.060 1238.680 18.320 ;
      LAYER met2 ;
        RECT 1258.890 600.170 1259.170 604.000 ;
        RECT 1257.340 600.030 1259.170 600.170 ;
        RECT 1257.340 587.170 1257.480 600.030 ;
        RECT 1258.890 600.000 1259.170 600.030 ;
        RECT 1238.420 586.850 1238.680 587.170 ;
        RECT 1257.280 586.850 1257.540 587.170 ;
        RECT 1238.480 18.350 1238.620 586.850 ;
        RECT 1144.580 18.030 1144.840 18.350 ;
        RECT 1238.420 18.030 1238.680 18.350 ;
        RECT 1144.640 2.400 1144.780 18.030 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1218.150 593.200 1218.470 593.260 ;
        RECT 1266.450 593.200 1266.770 593.260 ;
        RECT 1218.150 593.060 1266.770 593.200 ;
        RECT 1218.150 593.000 1218.470 593.060 ;
        RECT 1266.450 593.000 1266.770 593.060 ;
        RECT 1218.150 588.780 1218.470 588.840 ;
        RECT 1197.080 588.640 1218.470 588.780 ;
        RECT 1165.710 588.440 1166.030 588.500 ;
        RECT 1197.080 588.440 1197.220 588.640 ;
        RECT 1218.150 588.580 1218.470 588.640 ;
        RECT 1165.710 588.300 1197.220 588.440 ;
        RECT 1165.710 588.240 1166.030 588.300 ;
        RECT 1162.490 20.640 1162.810 20.700 ;
        RECT 1165.710 20.640 1166.030 20.700 ;
        RECT 1162.490 20.500 1166.030 20.640 ;
        RECT 1162.490 20.440 1162.810 20.500 ;
        RECT 1165.710 20.440 1166.030 20.500 ;
      LAYER via ;
        RECT 1218.180 593.000 1218.440 593.260 ;
        RECT 1266.480 593.000 1266.740 593.260 ;
        RECT 1165.740 588.240 1166.000 588.500 ;
        RECT 1218.180 588.580 1218.440 588.840 ;
        RECT 1162.520 20.440 1162.780 20.700 ;
        RECT 1165.740 20.440 1166.000 20.700 ;
      LAYER met2 ;
        RECT 1268.090 600.170 1268.370 604.000 ;
        RECT 1266.540 600.030 1268.370 600.170 ;
        RECT 1266.540 593.290 1266.680 600.030 ;
        RECT 1268.090 600.000 1268.370 600.030 ;
        RECT 1218.180 592.970 1218.440 593.290 ;
        RECT 1266.480 592.970 1266.740 593.290 ;
        RECT 1218.240 588.870 1218.380 592.970 ;
        RECT 1218.180 588.550 1218.440 588.870 ;
        RECT 1165.740 588.210 1166.000 588.530 ;
        RECT 1165.800 20.730 1165.940 588.210 ;
        RECT 1162.520 20.410 1162.780 20.730 ;
        RECT 1165.740 20.410 1166.000 20.730 ;
        RECT 1162.580 2.400 1162.720 20.410 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1014.830 583.000 1015.150 583.060 ;
        RECT 1018.510 583.000 1018.830 583.060 ;
        RECT 1014.830 582.860 1018.830 583.000 ;
        RECT 1014.830 582.800 1015.150 582.860 ;
        RECT 1018.510 582.800 1018.830 582.860 ;
        RECT 680.410 38.660 680.730 38.720 ;
        RECT 1014.830 38.660 1015.150 38.720 ;
        RECT 680.410 38.520 1015.150 38.660 ;
        RECT 680.410 38.460 680.730 38.520 ;
        RECT 1014.830 38.460 1015.150 38.520 ;
      LAYER via ;
        RECT 1014.860 582.800 1015.120 583.060 ;
        RECT 1018.540 582.800 1018.800 583.060 ;
        RECT 680.440 38.460 680.700 38.720 ;
        RECT 1014.860 38.460 1015.120 38.720 ;
      LAYER met2 ;
        RECT 1020.150 600.170 1020.430 604.000 ;
        RECT 1018.600 600.030 1020.430 600.170 ;
        RECT 1018.600 583.090 1018.740 600.030 ;
        RECT 1020.150 600.000 1020.430 600.030 ;
        RECT 1014.860 582.770 1015.120 583.090 ;
        RECT 1018.540 582.770 1018.800 583.090 ;
        RECT 1014.920 38.750 1015.060 582.770 ;
        RECT 680.440 38.430 680.700 38.750 ;
        RECT 1014.860 38.430 1015.120 38.750 ;
        RECT 680.500 2.400 680.640 38.430 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1208.950 592.860 1209.270 592.920 ;
        RECT 1276.570 592.860 1276.890 592.920 ;
        RECT 1208.950 592.720 1276.890 592.860 ;
        RECT 1208.950 592.660 1209.270 592.720 ;
        RECT 1276.570 592.660 1276.890 592.720 ;
        RECT 1208.950 588.100 1209.270 588.160 ;
        RECT 1202.600 587.960 1209.270 588.100 ;
        RECT 1197.450 587.760 1197.770 587.820 ;
        RECT 1202.600 587.760 1202.740 587.960 ;
        RECT 1208.950 587.900 1209.270 587.960 ;
        RECT 1197.450 587.620 1202.740 587.760 ;
        RECT 1197.450 587.560 1197.770 587.620 ;
        RECT 1196.530 586.740 1196.850 586.800 ;
        RECT 1188.340 586.600 1196.850 586.740 ;
        RECT 1185.950 586.400 1186.270 586.460 ;
        RECT 1188.340 586.400 1188.480 586.600 ;
        RECT 1196.530 586.540 1196.850 586.600 ;
        RECT 1185.950 586.260 1188.480 586.400 ;
        RECT 1185.950 586.200 1186.270 586.260 ;
        RECT 1185.950 62.260 1186.270 62.520 ;
        RECT 1186.040 61.840 1186.180 62.260 ;
        RECT 1185.950 61.580 1186.270 61.840 ;
        RECT 1179.970 22.680 1180.290 22.740 ;
        RECT 1185.950 22.680 1186.270 22.740 ;
        RECT 1179.970 22.540 1186.270 22.680 ;
        RECT 1179.970 22.480 1180.290 22.540 ;
        RECT 1185.950 22.480 1186.270 22.540 ;
      LAYER via ;
        RECT 1208.980 592.660 1209.240 592.920 ;
        RECT 1276.600 592.660 1276.860 592.920 ;
        RECT 1197.480 587.560 1197.740 587.820 ;
        RECT 1208.980 587.900 1209.240 588.160 ;
        RECT 1185.980 586.200 1186.240 586.460 ;
        RECT 1196.560 586.540 1196.820 586.800 ;
        RECT 1185.980 62.260 1186.240 62.520 ;
        RECT 1185.980 61.580 1186.240 61.840 ;
        RECT 1180.000 22.480 1180.260 22.740 ;
        RECT 1185.980 22.480 1186.240 22.740 ;
      LAYER met2 ;
        RECT 1277.290 600.170 1277.570 604.000 ;
        RECT 1276.660 600.030 1277.570 600.170 ;
        RECT 1276.660 592.950 1276.800 600.030 ;
        RECT 1277.290 600.000 1277.570 600.030 ;
        RECT 1208.980 592.630 1209.240 592.950 ;
        RECT 1276.600 592.630 1276.860 592.950 ;
        RECT 1209.040 588.190 1209.180 592.630 ;
        RECT 1208.980 587.870 1209.240 588.190 ;
        RECT 1197.480 587.530 1197.740 587.850 ;
        RECT 1197.540 587.250 1197.680 587.530 ;
        RECT 1196.620 587.110 1197.680 587.250 ;
        RECT 1196.620 586.830 1196.760 587.110 ;
        RECT 1196.560 586.510 1196.820 586.830 ;
        RECT 1185.980 586.170 1186.240 586.490 ;
        RECT 1186.040 62.550 1186.180 586.170 ;
        RECT 1185.980 62.230 1186.240 62.550 ;
        RECT 1185.980 61.550 1186.240 61.870 ;
        RECT 1186.040 22.770 1186.180 61.550 ;
        RECT 1180.000 22.450 1180.260 22.770 ;
        RECT 1185.980 22.450 1186.240 22.770 ;
        RECT 1180.060 2.400 1180.200 22.450 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 588.440 1200.530 588.500 ;
        RECT 1284.850 588.440 1285.170 588.500 ;
        RECT 1200.210 588.300 1285.170 588.440 ;
        RECT 1200.210 588.240 1200.530 588.300 ;
        RECT 1284.850 588.240 1285.170 588.300 ;
        RECT 1197.910 20.640 1198.230 20.700 ;
        RECT 1200.210 20.640 1200.530 20.700 ;
        RECT 1197.910 20.500 1200.530 20.640 ;
        RECT 1197.910 20.440 1198.230 20.500 ;
        RECT 1200.210 20.440 1200.530 20.500 ;
      LAYER via ;
        RECT 1200.240 588.240 1200.500 588.500 ;
        RECT 1284.880 588.240 1285.140 588.500 ;
        RECT 1197.940 20.440 1198.200 20.700 ;
        RECT 1200.240 20.440 1200.500 20.700 ;
      LAYER met2 ;
        RECT 1286.490 600.170 1286.770 604.000 ;
        RECT 1284.940 600.030 1286.770 600.170 ;
        RECT 1284.940 588.530 1285.080 600.030 ;
        RECT 1286.490 600.000 1286.770 600.030 ;
        RECT 1200.240 588.210 1200.500 588.530 ;
        RECT 1284.880 588.210 1285.140 588.530 ;
        RECT 1200.300 20.730 1200.440 588.210 ;
        RECT 1197.940 20.410 1198.200 20.730 ;
        RECT 1200.240 20.410 1200.500 20.730 ;
        RECT 1198.000 2.400 1198.140 20.410 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 588.100 1221.230 588.160 ;
        RECT 1294.050 588.100 1294.370 588.160 ;
        RECT 1220.910 587.960 1294.370 588.100 ;
        RECT 1220.910 587.900 1221.230 587.960 ;
        RECT 1294.050 587.900 1294.370 587.960 ;
        RECT 1215.850 20.640 1216.170 20.700 ;
        RECT 1220.910 20.640 1221.230 20.700 ;
        RECT 1215.850 20.500 1221.230 20.640 ;
        RECT 1215.850 20.440 1216.170 20.500 ;
        RECT 1220.910 20.440 1221.230 20.500 ;
      LAYER via ;
        RECT 1220.940 587.900 1221.200 588.160 ;
        RECT 1294.080 587.900 1294.340 588.160 ;
        RECT 1215.880 20.440 1216.140 20.700 ;
        RECT 1220.940 20.440 1221.200 20.700 ;
      LAYER met2 ;
        RECT 1295.690 600.170 1295.970 604.000 ;
        RECT 1294.140 600.030 1295.970 600.170 ;
        RECT 1294.140 588.190 1294.280 600.030 ;
        RECT 1295.690 600.000 1295.970 600.030 ;
        RECT 1220.940 587.870 1221.200 588.190 ;
        RECT 1294.080 587.870 1294.340 588.190 ;
        RECT 1221.000 20.730 1221.140 587.870 ;
        RECT 1215.880 20.410 1216.140 20.730 ;
        RECT 1220.940 20.410 1221.200 20.730 ;
        RECT 1215.940 2.400 1216.080 20.410 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1252.650 591.500 1252.970 591.560 ;
        RECT 1304.170 591.500 1304.490 591.560 ;
        RECT 1252.650 591.360 1304.490 591.500 ;
        RECT 1252.650 591.300 1252.970 591.360 ;
        RECT 1304.170 591.300 1304.490 591.360 ;
        RECT 1233.790 16.220 1234.110 16.280 ;
        RECT 1252.650 16.220 1252.970 16.280 ;
        RECT 1233.790 16.080 1252.970 16.220 ;
        RECT 1233.790 16.020 1234.110 16.080 ;
        RECT 1252.650 16.020 1252.970 16.080 ;
      LAYER via ;
        RECT 1252.680 591.300 1252.940 591.560 ;
        RECT 1304.200 591.300 1304.460 591.560 ;
        RECT 1233.820 16.020 1234.080 16.280 ;
        RECT 1252.680 16.020 1252.940 16.280 ;
      LAYER met2 ;
        RECT 1304.890 600.170 1305.170 604.000 ;
        RECT 1304.260 600.030 1305.170 600.170 ;
        RECT 1304.260 591.590 1304.400 600.030 ;
        RECT 1304.890 600.000 1305.170 600.030 ;
        RECT 1252.680 591.270 1252.940 591.590 ;
        RECT 1304.200 591.270 1304.460 591.590 ;
        RECT 1252.740 16.310 1252.880 591.270 ;
        RECT 1233.820 15.990 1234.080 16.310 ;
        RECT 1252.680 15.990 1252.940 16.310 ;
        RECT 1233.880 2.400 1234.020 15.990 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 590.820 1255.730 590.880 ;
        RECT 1312.450 590.820 1312.770 590.880 ;
        RECT 1255.410 590.680 1312.770 590.820 ;
        RECT 1255.410 590.620 1255.730 590.680 ;
        RECT 1312.450 590.620 1312.770 590.680 ;
        RECT 1251.730 16.900 1252.050 16.960 ;
        RECT 1255.410 16.900 1255.730 16.960 ;
        RECT 1251.730 16.760 1255.730 16.900 ;
        RECT 1251.730 16.700 1252.050 16.760 ;
        RECT 1255.410 16.700 1255.730 16.760 ;
      LAYER via ;
        RECT 1255.440 590.620 1255.700 590.880 ;
        RECT 1312.480 590.620 1312.740 590.880 ;
        RECT 1251.760 16.700 1252.020 16.960 ;
        RECT 1255.440 16.700 1255.700 16.960 ;
      LAYER met2 ;
        RECT 1314.090 600.170 1314.370 604.000 ;
        RECT 1312.540 600.030 1314.370 600.170 ;
        RECT 1312.540 590.910 1312.680 600.030 ;
        RECT 1314.090 600.000 1314.370 600.030 ;
        RECT 1255.440 590.590 1255.700 590.910 ;
        RECT 1312.480 590.590 1312.740 590.910 ;
        RECT 1255.500 16.990 1255.640 590.590 ;
        RECT 1251.760 16.670 1252.020 16.990 ;
        RECT 1255.440 16.670 1255.700 16.990 ;
        RECT 1251.820 2.400 1251.960 16.670 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1286.690 592.860 1287.010 592.920 ;
        RECT 1321.650 592.860 1321.970 592.920 ;
        RECT 1286.690 592.720 1321.970 592.860 ;
        RECT 1286.690 592.660 1287.010 592.720 ;
        RECT 1321.650 592.660 1321.970 592.720 ;
        RECT 1269.210 16.560 1269.530 16.620 ;
        RECT 1286.690 16.560 1287.010 16.620 ;
        RECT 1269.210 16.420 1287.010 16.560 ;
        RECT 1269.210 16.360 1269.530 16.420 ;
        RECT 1286.690 16.360 1287.010 16.420 ;
      LAYER via ;
        RECT 1286.720 592.660 1286.980 592.920 ;
        RECT 1321.680 592.660 1321.940 592.920 ;
        RECT 1269.240 16.360 1269.500 16.620 ;
        RECT 1286.720 16.360 1286.980 16.620 ;
      LAYER met2 ;
        RECT 1323.290 600.170 1323.570 604.000 ;
        RECT 1321.740 600.030 1323.570 600.170 ;
        RECT 1321.740 592.950 1321.880 600.030 ;
        RECT 1323.290 600.000 1323.570 600.030 ;
        RECT 1286.720 592.630 1286.980 592.950 ;
        RECT 1321.680 592.630 1321.940 592.950 ;
        RECT 1286.780 16.650 1286.920 592.630 ;
        RECT 1269.240 16.330 1269.500 16.650 ;
        RECT 1286.720 16.330 1286.980 16.650 ;
        RECT 1269.300 2.400 1269.440 16.330 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 591.840 1290.230 591.900 ;
        RECT 1331.770 591.840 1332.090 591.900 ;
        RECT 1289.910 591.700 1332.090 591.840 ;
        RECT 1289.910 591.640 1290.230 591.700 ;
        RECT 1331.770 591.640 1332.090 591.700 ;
        RECT 1287.150 17.580 1287.470 17.640 ;
        RECT 1289.910 17.580 1290.230 17.640 ;
        RECT 1287.150 17.440 1290.230 17.580 ;
        RECT 1287.150 17.380 1287.470 17.440 ;
        RECT 1289.910 17.380 1290.230 17.440 ;
      LAYER via ;
        RECT 1289.940 591.640 1290.200 591.900 ;
        RECT 1331.800 591.640 1332.060 591.900 ;
        RECT 1287.180 17.380 1287.440 17.640 ;
        RECT 1289.940 17.380 1290.200 17.640 ;
      LAYER met2 ;
        RECT 1332.490 600.170 1332.770 604.000 ;
        RECT 1331.860 600.030 1332.770 600.170 ;
        RECT 1331.860 591.930 1332.000 600.030 ;
        RECT 1332.490 600.000 1332.770 600.030 ;
        RECT 1289.940 591.610 1290.200 591.930 ;
        RECT 1331.800 591.610 1332.060 591.930 ;
        RECT 1290.000 17.670 1290.140 591.610 ;
        RECT 1287.180 17.350 1287.440 17.670 ;
        RECT 1289.940 17.350 1290.200 17.670 ;
        RECT 1287.240 2.400 1287.380 17.350 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 590.140 1310.930 590.200 ;
        RECT 1340.050 590.140 1340.370 590.200 ;
        RECT 1310.610 590.000 1340.370 590.140 ;
        RECT 1310.610 589.940 1310.930 590.000 ;
        RECT 1340.050 589.940 1340.370 590.000 ;
        RECT 1305.090 16.220 1305.410 16.280 ;
        RECT 1310.610 16.220 1310.930 16.280 ;
        RECT 1305.090 16.080 1310.930 16.220 ;
        RECT 1305.090 16.020 1305.410 16.080 ;
        RECT 1310.610 16.020 1310.930 16.080 ;
      LAYER via ;
        RECT 1310.640 589.940 1310.900 590.200 ;
        RECT 1340.080 589.940 1340.340 590.200 ;
        RECT 1305.120 16.020 1305.380 16.280 ;
        RECT 1310.640 16.020 1310.900 16.280 ;
      LAYER met2 ;
        RECT 1341.690 600.170 1341.970 604.000 ;
        RECT 1340.140 600.030 1341.970 600.170 ;
        RECT 1340.140 590.230 1340.280 600.030 ;
        RECT 1341.690 600.000 1341.970 600.030 ;
        RECT 1310.640 589.910 1310.900 590.230 ;
        RECT 1340.080 589.910 1340.340 590.230 ;
        RECT 1310.700 16.310 1310.840 589.910 ;
        RECT 1305.120 15.990 1305.380 16.310 ;
        RECT 1310.640 15.990 1310.900 16.310 ;
        RECT 1305.180 2.400 1305.320 15.990 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1341.890 586.740 1342.210 586.800 ;
        RECT 1349.250 586.740 1349.570 586.800 ;
        RECT 1341.890 586.600 1349.570 586.740 ;
        RECT 1341.890 586.540 1342.210 586.600 ;
        RECT 1349.250 586.540 1349.570 586.600 ;
        RECT 1323.030 15.540 1323.350 15.600 ;
        RECT 1341.890 15.540 1342.210 15.600 ;
        RECT 1323.030 15.400 1342.210 15.540 ;
        RECT 1323.030 15.340 1323.350 15.400 ;
        RECT 1341.890 15.340 1342.210 15.400 ;
      LAYER via ;
        RECT 1341.920 586.540 1342.180 586.800 ;
        RECT 1349.280 586.540 1349.540 586.800 ;
        RECT 1323.060 15.340 1323.320 15.600 ;
        RECT 1341.920 15.340 1342.180 15.600 ;
      LAYER met2 ;
        RECT 1350.890 600.170 1351.170 604.000 ;
        RECT 1349.340 600.030 1351.170 600.170 ;
        RECT 1349.340 586.830 1349.480 600.030 ;
        RECT 1350.890 600.000 1351.170 600.030 ;
        RECT 1341.920 586.510 1342.180 586.830 ;
        RECT 1349.280 586.510 1349.540 586.830 ;
        RECT 1341.980 15.630 1342.120 586.510 ;
        RECT 1323.060 15.310 1323.320 15.630 ;
        RECT 1341.920 15.310 1342.180 15.630 ;
        RECT 1323.120 2.400 1323.260 15.310 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1348.790 587.080 1349.110 587.140 ;
        RECT 1359.370 587.080 1359.690 587.140 ;
        RECT 1348.790 586.940 1359.690 587.080 ;
        RECT 1348.790 586.880 1349.110 586.940 ;
        RECT 1359.370 586.880 1359.690 586.940 ;
        RECT 1340.510 20.640 1340.830 20.700 ;
        RECT 1348.790 20.640 1349.110 20.700 ;
        RECT 1340.510 20.500 1349.110 20.640 ;
        RECT 1340.510 20.440 1340.830 20.500 ;
        RECT 1348.790 20.440 1349.110 20.500 ;
      LAYER via ;
        RECT 1348.820 586.880 1349.080 587.140 ;
        RECT 1359.400 586.880 1359.660 587.140 ;
        RECT 1340.540 20.440 1340.800 20.700 ;
        RECT 1348.820 20.440 1349.080 20.700 ;
      LAYER met2 ;
        RECT 1360.090 600.170 1360.370 604.000 ;
        RECT 1359.460 600.030 1360.370 600.170 ;
        RECT 1359.460 587.170 1359.600 600.030 ;
        RECT 1360.090 600.000 1360.370 600.030 ;
        RECT 1348.820 586.850 1349.080 587.170 ;
        RECT 1359.400 586.850 1359.660 587.170 ;
        RECT 1348.880 20.730 1349.020 586.850 ;
        RECT 1340.540 20.410 1340.800 20.730 ;
        RECT 1348.820 20.410 1349.080 20.730 ;
        RECT 1340.600 2.400 1340.740 20.410 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 698.350 39.000 698.670 39.060 ;
        RECT 1028.630 39.000 1028.950 39.060 ;
        RECT 698.350 38.860 1028.950 39.000 ;
        RECT 698.350 38.800 698.670 38.860 ;
        RECT 1028.630 38.800 1028.950 38.860 ;
      LAYER via ;
        RECT 698.380 38.800 698.640 39.060 ;
        RECT 1028.660 38.800 1028.920 39.060 ;
      LAYER met2 ;
        RECT 1029.350 600.170 1029.630 604.000 ;
        RECT 1028.720 600.030 1029.630 600.170 ;
        RECT 1028.720 39.090 1028.860 600.030 ;
        RECT 1029.350 600.000 1029.630 600.030 ;
        RECT 698.380 38.770 698.640 39.090 ;
        RECT 1028.660 38.770 1028.920 39.090 ;
        RECT 698.440 2.400 698.580 38.770 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1362.590 587.080 1362.910 587.140 ;
        RECT 1367.650 587.080 1367.970 587.140 ;
        RECT 1362.590 586.940 1367.970 587.080 ;
        RECT 1362.590 586.880 1362.910 586.940 ;
        RECT 1367.650 586.880 1367.970 586.940 ;
        RECT 1358.450 20.640 1358.770 20.700 ;
        RECT 1362.590 20.640 1362.910 20.700 ;
        RECT 1358.450 20.500 1362.910 20.640 ;
        RECT 1358.450 20.440 1358.770 20.500 ;
        RECT 1362.590 20.440 1362.910 20.500 ;
      LAYER via ;
        RECT 1362.620 586.880 1362.880 587.140 ;
        RECT 1367.680 586.880 1367.940 587.140 ;
        RECT 1358.480 20.440 1358.740 20.700 ;
        RECT 1362.620 20.440 1362.880 20.700 ;
      LAYER met2 ;
        RECT 1369.290 600.170 1369.570 604.000 ;
        RECT 1367.740 600.030 1369.570 600.170 ;
        RECT 1367.740 587.170 1367.880 600.030 ;
        RECT 1369.290 600.000 1369.570 600.030 ;
        RECT 1362.620 586.850 1362.880 587.170 ;
        RECT 1367.680 586.850 1367.940 587.170 ;
        RECT 1362.680 20.730 1362.820 586.850 ;
        RECT 1358.480 20.410 1358.740 20.730 ;
        RECT 1362.620 20.410 1362.880 20.730 ;
        RECT 1358.540 2.400 1358.680 20.410 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1374.550 524.520 1374.870 524.580 ;
        RECT 1376.850 524.520 1377.170 524.580 ;
        RECT 1374.550 524.380 1377.170 524.520 ;
        RECT 1374.550 524.320 1374.870 524.380 ;
        RECT 1376.850 524.320 1377.170 524.380 ;
        RECT 1374.090 62.260 1374.410 62.520 ;
        RECT 1374.180 61.780 1374.320 62.260 ;
        RECT 1376.390 61.780 1376.710 61.840 ;
        RECT 1374.180 61.640 1376.710 61.780 ;
        RECT 1376.390 61.580 1376.710 61.640 ;
      LAYER via ;
        RECT 1374.580 524.320 1374.840 524.580 ;
        RECT 1376.880 524.320 1377.140 524.580 ;
        RECT 1374.120 62.260 1374.380 62.520 ;
        RECT 1376.420 61.580 1376.680 61.840 ;
      LAYER met2 ;
        RECT 1378.490 600.170 1378.770 604.000 ;
        RECT 1376.940 600.030 1378.770 600.170 ;
        RECT 1376.940 524.610 1377.080 600.030 ;
        RECT 1378.490 600.000 1378.770 600.030 ;
        RECT 1374.580 524.290 1374.840 524.610 ;
        RECT 1376.880 524.290 1377.140 524.610 ;
        RECT 1374.640 524.125 1374.780 524.290 ;
        RECT 1373.650 523.755 1373.930 524.125 ;
        RECT 1374.570 523.755 1374.850 524.125 ;
        RECT 1373.720 447.170 1373.860 523.755 ;
        RECT 1373.720 447.030 1374.320 447.170 ;
        RECT 1374.180 62.550 1374.320 447.030 ;
        RECT 1374.120 62.230 1374.380 62.550 ;
        RECT 1376.420 61.550 1376.680 61.870 ;
        RECT 1376.480 2.400 1376.620 61.550 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
      LAYER via2 ;
        RECT 1373.650 523.800 1373.930 524.080 ;
        RECT 1374.570 523.800 1374.850 524.080 ;
      LAYER met3 ;
        RECT 1373.625 524.090 1373.955 524.105 ;
        RECT 1374.545 524.090 1374.875 524.105 ;
        RECT 1373.625 523.790 1374.875 524.090 ;
        RECT 1373.625 523.775 1373.955 523.790 ;
        RECT 1374.545 523.775 1374.875 523.790 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1389.270 586.740 1389.590 586.800 ;
        RECT 1394.330 586.740 1394.650 586.800 ;
        RECT 1389.270 586.600 1394.650 586.740 ;
        RECT 1389.270 586.540 1389.590 586.600 ;
        RECT 1394.330 586.540 1394.650 586.600 ;
      LAYER via ;
        RECT 1389.300 586.540 1389.560 586.800 ;
        RECT 1394.360 586.540 1394.620 586.800 ;
      LAYER met2 ;
        RECT 1387.690 600.170 1387.970 604.000 ;
        RECT 1387.690 600.030 1389.500 600.170 ;
        RECT 1387.690 600.000 1387.970 600.030 ;
        RECT 1389.360 586.830 1389.500 600.030 ;
        RECT 1389.300 586.510 1389.560 586.830 ;
        RECT 1394.360 586.510 1394.620 586.830 ;
        RECT 1394.420 2.400 1394.560 586.510 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1398.470 524.180 1398.790 524.240 ;
        RECT 1398.930 524.180 1399.250 524.240 ;
        RECT 1398.470 524.040 1399.250 524.180 ;
        RECT 1398.470 523.980 1398.790 524.040 ;
        RECT 1398.930 523.980 1399.250 524.040 ;
        RECT 1398.470 496.980 1398.790 497.040 ;
        RECT 1398.470 496.840 1399.160 496.980 ;
        RECT 1398.470 496.780 1398.790 496.840 ;
        RECT 1399.020 496.700 1399.160 496.840 ;
        RECT 1398.930 496.440 1399.250 496.700 ;
        RECT 1398.470 435.100 1398.790 435.160 ;
        RECT 1398.930 435.100 1399.250 435.160 ;
        RECT 1398.470 434.960 1399.250 435.100 ;
        RECT 1398.470 434.900 1398.790 434.960 ;
        RECT 1398.930 434.900 1399.250 434.960 ;
        RECT 1397.550 379.340 1397.870 379.400 ;
        RECT 1398.470 379.340 1398.790 379.400 ;
        RECT 1397.550 379.200 1398.790 379.340 ;
        RECT 1397.550 379.140 1397.870 379.200 ;
        RECT 1398.470 379.140 1398.790 379.200 ;
        RECT 1397.550 331.400 1397.870 331.460 ;
        RECT 1398.930 331.400 1399.250 331.460 ;
        RECT 1397.550 331.260 1399.250 331.400 ;
        RECT 1397.550 331.200 1397.870 331.260 ;
        RECT 1398.930 331.200 1399.250 331.260 ;
        RECT 1399.390 303.520 1399.710 303.580 ;
        RECT 1400.310 303.520 1400.630 303.580 ;
        RECT 1399.390 303.380 1400.630 303.520 ;
        RECT 1399.390 303.320 1399.710 303.380 ;
        RECT 1400.310 303.320 1400.630 303.380 ;
        RECT 1399.390 289.580 1399.710 289.640 ;
        RECT 1400.310 289.580 1400.630 289.640 ;
        RECT 1399.390 289.440 1400.630 289.580 ;
        RECT 1399.390 289.380 1399.710 289.440 ;
        RECT 1400.310 289.380 1400.630 289.440 ;
        RECT 1399.390 241.640 1399.710 241.700 ;
        RECT 1400.310 241.640 1400.630 241.700 ;
        RECT 1399.390 241.500 1400.630 241.640 ;
        RECT 1399.390 241.440 1399.710 241.500 ;
        RECT 1400.310 241.440 1400.630 241.500 ;
        RECT 1399.390 193.360 1399.710 193.420 ;
        RECT 1400.310 193.360 1400.630 193.420 ;
        RECT 1399.390 193.220 1400.630 193.360 ;
        RECT 1399.390 193.160 1399.710 193.220 ;
        RECT 1400.310 193.160 1400.630 193.220 ;
        RECT 1399.390 158.680 1399.710 158.740 ;
        RECT 1400.310 158.680 1400.630 158.740 ;
        RECT 1399.390 158.540 1400.630 158.680 ;
        RECT 1399.390 158.480 1399.710 158.540 ;
        RECT 1400.310 158.480 1400.630 158.540 ;
        RECT 1398.930 144.740 1399.250 144.800 ;
        RECT 1400.310 144.740 1400.630 144.800 ;
        RECT 1398.930 144.600 1400.630 144.740 ;
        RECT 1398.930 144.540 1399.250 144.600 ;
        RECT 1400.310 144.540 1400.630 144.600 ;
        RECT 1398.930 96.800 1399.250 96.860 ;
        RECT 1399.850 96.800 1400.170 96.860 ;
        RECT 1398.930 96.660 1400.170 96.800 ;
        RECT 1398.930 96.600 1399.250 96.660 ;
        RECT 1399.850 96.600 1400.170 96.660 ;
        RECT 1400.310 20.640 1400.630 20.700 ;
        RECT 1412.270 20.640 1412.590 20.700 ;
        RECT 1400.310 20.500 1412.590 20.640 ;
        RECT 1400.310 20.440 1400.630 20.500 ;
        RECT 1412.270 20.440 1412.590 20.500 ;
      LAYER via ;
        RECT 1398.500 523.980 1398.760 524.240 ;
        RECT 1398.960 523.980 1399.220 524.240 ;
        RECT 1398.500 496.780 1398.760 497.040 ;
        RECT 1398.960 496.440 1399.220 496.700 ;
        RECT 1398.500 434.900 1398.760 435.160 ;
        RECT 1398.960 434.900 1399.220 435.160 ;
        RECT 1397.580 379.140 1397.840 379.400 ;
        RECT 1398.500 379.140 1398.760 379.400 ;
        RECT 1397.580 331.200 1397.840 331.460 ;
        RECT 1398.960 331.200 1399.220 331.460 ;
        RECT 1399.420 303.320 1399.680 303.580 ;
        RECT 1400.340 303.320 1400.600 303.580 ;
        RECT 1399.420 289.380 1399.680 289.640 ;
        RECT 1400.340 289.380 1400.600 289.640 ;
        RECT 1399.420 241.440 1399.680 241.700 ;
        RECT 1400.340 241.440 1400.600 241.700 ;
        RECT 1399.420 193.160 1399.680 193.420 ;
        RECT 1400.340 193.160 1400.600 193.420 ;
        RECT 1399.420 158.480 1399.680 158.740 ;
        RECT 1400.340 158.480 1400.600 158.740 ;
        RECT 1398.960 144.540 1399.220 144.800 ;
        RECT 1400.340 144.540 1400.600 144.800 ;
        RECT 1398.960 96.600 1399.220 96.860 ;
        RECT 1399.880 96.600 1400.140 96.860 ;
        RECT 1400.340 20.440 1400.600 20.700 ;
        RECT 1412.300 20.440 1412.560 20.700 ;
      LAYER met2 ;
        RECT 1396.890 600.170 1397.170 604.000 ;
        RECT 1396.890 600.030 1398.700 600.170 ;
        RECT 1396.890 600.000 1397.170 600.030 ;
        RECT 1398.560 596.770 1398.700 600.030 ;
        RECT 1398.560 596.630 1400.080 596.770 ;
        RECT 1399.940 545.090 1400.080 596.630 ;
        RECT 1399.020 544.950 1400.080 545.090 ;
        RECT 1399.020 524.270 1399.160 544.950 ;
        RECT 1398.500 523.950 1398.760 524.270 ;
        RECT 1398.960 523.950 1399.220 524.270 ;
        RECT 1398.560 497.070 1398.700 523.950 ;
        RECT 1398.500 496.750 1398.760 497.070 ;
        RECT 1398.960 496.410 1399.220 496.730 ;
        RECT 1399.020 435.190 1399.160 496.410 ;
        RECT 1398.500 434.870 1398.760 435.190 ;
        RECT 1398.960 434.870 1399.220 435.190 ;
        RECT 1398.560 379.430 1398.700 434.870 ;
        RECT 1397.580 379.110 1397.840 379.430 ;
        RECT 1398.500 379.110 1398.760 379.430 ;
        RECT 1397.640 331.490 1397.780 379.110 ;
        RECT 1397.580 331.170 1397.840 331.490 ;
        RECT 1398.960 331.170 1399.220 331.490 ;
        RECT 1399.020 303.690 1399.160 331.170 ;
        RECT 1399.020 303.610 1399.620 303.690 ;
        RECT 1399.020 303.550 1399.680 303.610 ;
        RECT 1399.420 303.290 1399.680 303.550 ;
        RECT 1400.340 303.290 1400.600 303.610 ;
        RECT 1400.400 289.670 1400.540 303.290 ;
        RECT 1399.420 289.350 1399.680 289.670 ;
        RECT 1400.340 289.350 1400.600 289.670 ;
        RECT 1399.480 241.730 1399.620 289.350 ;
        RECT 1399.420 241.410 1399.680 241.730 ;
        RECT 1400.340 241.410 1400.600 241.730 ;
        RECT 1400.400 193.450 1400.540 241.410 ;
        RECT 1399.420 193.130 1399.680 193.450 ;
        RECT 1400.340 193.130 1400.600 193.450 ;
        RECT 1399.480 158.770 1399.620 193.130 ;
        RECT 1399.420 158.450 1399.680 158.770 ;
        RECT 1400.340 158.450 1400.600 158.770 ;
        RECT 1400.400 144.830 1400.540 158.450 ;
        RECT 1398.960 144.510 1399.220 144.830 ;
        RECT 1400.340 144.510 1400.600 144.830 ;
        RECT 1399.020 96.890 1399.160 144.510 ;
        RECT 1398.960 96.570 1399.220 96.890 ;
        RECT 1399.880 96.570 1400.140 96.890 ;
        RECT 1399.940 62.290 1400.080 96.570 ;
        RECT 1399.940 62.150 1400.540 62.290 ;
        RECT 1400.400 20.730 1400.540 62.150 ;
        RECT 1400.340 20.410 1400.600 20.730 ;
        RECT 1412.300 20.410 1412.560 20.730 ;
        RECT 1412.360 2.400 1412.500 20.410 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1407.210 16.220 1407.530 16.280 ;
        RECT 1429.750 16.220 1430.070 16.280 ;
        RECT 1407.210 16.080 1430.070 16.220 ;
        RECT 1407.210 16.020 1407.530 16.080 ;
        RECT 1429.750 16.020 1430.070 16.080 ;
      LAYER via ;
        RECT 1407.240 16.020 1407.500 16.280 ;
        RECT 1429.780 16.020 1430.040 16.280 ;
      LAYER met2 ;
        RECT 1406.090 600.170 1406.370 604.000 ;
        RECT 1406.090 600.030 1407.440 600.170 ;
        RECT 1406.090 600.000 1406.370 600.030 ;
        RECT 1407.300 16.310 1407.440 600.030 ;
        RECT 1407.240 15.990 1407.500 16.310 ;
        RECT 1429.780 15.990 1430.040 16.310 ;
        RECT 1429.840 2.400 1429.980 15.990 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1416.870 586.740 1417.190 586.800 ;
        RECT 1421.010 586.740 1421.330 586.800 ;
        RECT 1416.870 586.600 1421.330 586.740 ;
        RECT 1416.870 586.540 1417.190 586.600 ;
        RECT 1421.010 586.540 1421.330 586.600 ;
        RECT 1421.010 18.260 1421.330 18.320 ;
        RECT 1447.690 18.260 1448.010 18.320 ;
        RECT 1421.010 18.120 1448.010 18.260 ;
        RECT 1421.010 18.060 1421.330 18.120 ;
        RECT 1447.690 18.060 1448.010 18.120 ;
      LAYER via ;
        RECT 1416.900 586.540 1417.160 586.800 ;
        RECT 1421.040 586.540 1421.300 586.800 ;
        RECT 1421.040 18.060 1421.300 18.320 ;
        RECT 1447.720 18.060 1447.980 18.320 ;
      LAYER met2 ;
        RECT 1415.290 600.170 1415.570 604.000 ;
        RECT 1415.290 600.030 1417.100 600.170 ;
        RECT 1415.290 600.000 1415.570 600.030 ;
        RECT 1416.960 586.830 1417.100 600.030 ;
        RECT 1416.900 586.510 1417.160 586.830 ;
        RECT 1421.040 586.510 1421.300 586.830 ;
        RECT 1421.100 18.350 1421.240 586.510 ;
        RECT 1421.040 18.030 1421.300 18.350 ;
        RECT 1447.720 18.030 1447.980 18.350 ;
        RECT 1447.780 2.400 1447.920 18.030 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1426.070 586.740 1426.390 586.800 ;
        RECT 1427.910 586.740 1428.230 586.800 ;
        RECT 1426.070 586.600 1428.230 586.740 ;
        RECT 1426.070 586.540 1426.390 586.600 ;
        RECT 1427.910 586.540 1428.230 586.600 ;
        RECT 1465.630 19.960 1465.950 20.020 ;
        RECT 1436.740 19.820 1465.950 19.960 ;
        RECT 1427.910 19.620 1428.230 19.680 ;
        RECT 1436.740 19.620 1436.880 19.820 ;
        RECT 1465.630 19.760 1465.950 19.820 ;
        RECT 1427.910 19.480 1436.880 19.620 ;
        RECT 1427.910 19.420 1428.230 19.480 ;
      LAYER via ;
        RECT 1426.100 586.540 1426.360 586.800 ;
        RECT 1427.940 586.540 1428.200 586.800 ;
        RECT 1427.940 19.420 1428.200 19.680 ;
        RECT 1465.660 19.760 1465.920 20.020 ;
      LAYER met2 ;
        RECT 1424.490 600.170 1424.770 604.000 ;
        RECT 1424.490 600.030 1426.300 600.170 ;
        RECT 1424.490 600.000 1424.770 600.030 ;
        RECT 1426.160 586.830 1426.300 600.030 ;
        RECT 1426.100 586.510 1426.360 586.830 ;
        RECT 1427.940 586.510 1428.200 586.830 ;
        RECT 1428.000 19.710 1428.140 586.510 ;
        RECT 1465.660 19.730 1465.920 20.050 ;
        RECT 1427.940 19.390 1428.200 19.710 ;
        RECT 1465.720 2.400 1465.860 19.730 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.350 18.600 1434.670 18.660 ;
        RECT 1483.570 18.600 1483.890 18.660 ;
        RECT 1434.350 18.460 1483.890 18.600 ;
        RECT 1434.350 18.400 1434.670 18.460 ;
        RECT 1483.570 18.400 1483.890 18.460 ;
      LAYER via ;
        RECT 1434.380 18.400 1434.640 18.660 ;
        RECT 1483.600 18.400 1483.860 18.660 ;
      LAYER met2 ;
        RECT 1433.690 600.170 1433.970 604.000 ;
        RECT 1433.690 600.030 1434.580 600.170 ;
        RECT 1433.690 600.000 1433.970 600.030 ;
        RECT 1434.440 18.690 1434.580 600.030 ;
        RECT 1434.380 18.370 1434.640 18.690 ;
        RECT 1483.600 18.370 1483.860 18.690 ;
        RECT 1483.660 2.400 1483.800 18.370 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1444.470 589.460 1444.790 589.520 ;
        RECT 1444.470 589.320 1465.400 589.460 ;
        RECT 1444.470 589.260 1444.790 589.320 ;
        RECT 1465.260 589.120 1465.400 589.320 ;
        RECT 1486.790 589.120 1487.110 589.180 ;
        RECT 1465.260 588.980 1487.110 589.120 ;
        RECT 1486.790 588.920 1487.110 588.980 ;
        RECT 1486.790 15.880 1487.110 15.940 ;
        RECT 1501.510 15.880 1501.830 15.940 ;
        RECT 1486.790 15.740 1501.830 15.880 ;
        RECT 1486.790 15.680 1487.110 15.740 ;
        RECT 1501.510 15.680 1501.830 15.740 ;
      LAYER via ;
        RECT 1444.500 589.260 1444.760 589.520 ;
        RECT 1486.820 588.920 1487.080 589.180 ;
        RECT 1486.820 15.680 1487.080 15.940 ;
        RECT 1501.540 15.680 1501.800 15.940 ;
      LAYER met2 ;
        RECT 1442.890 600.170 1443.170 604.000 ;
        RECT 1442.890 600.030 1444.700 600.170 ;
        RECT 1442.890 600.000 1443.170 600.030 ;
        RECT 1444.560 589.550 1444.700 600.030 ;
        RECT 1444.500 589.230 1444.760 589.550 ;
        RECT 1486.820 588.890 1487.080 589.210 ;
        RECT 1486.880 15.970 1487.020 588.890 ;
        RECT 1486.820 15.650 1487.080 15.970 ;
        RECT 1501.540 15.650 1501.800 15.970 ;
        RECT 1501.600 2.400 1501.740 15.650 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1453.210 497.320 1453.530 497.380 ;
        RECT 1452.840 497.180 1453.530 497.320 ;
        RECT 1452.840 496.700 1452.980 497.180 ;
        RECT 1453.210 497.120 1453.530 497.180 ;
        RECT 1452.750 496.440 1453.070 496.700 ;
        RECT 1451.370 483.040 1451.690 483.100 ;
        RECT 1452.750 483.040 1453.070 483.100 ;
        RECT 1451.370 482.900 1453.070 483.040 ;
        RECT 1451.370 482.840 1451.690 482.900 ;
        RECT 1452.750 482.840 1453.070 482.900 ;
        RECT 1451.370 324.260 1451.690 324.320 ;
        RECT 1452.290 324.260 1452.610 324.320 ;
        RECT 1451.370 324.120 1452.610 324.260 ;
        RECT 1451.370 324.060 1451.690 324.120 ;
        RECT 1452.290 324.060 1452.610 324.120 ;
        RECT 1451.370 276.320 1451.690 276.380 ;
        RECT 1452.750 276.320 1453.070 276.380 ;
        RECT 1451.370 276.180 1453.070 276.320 ;
        RECT 1451.370 276.120 1451.690 276.180 ;
        RECT 1452.750 276.120 1453.070 276.180 ;
        RECT 1453.210 193.160 1453.530 193.420 ;
        RECT 1453.300 192.740 1453.440 193.160 ;
        RECT 1453.210 192.480 1453.530 192.740 ;
        RECT 1453.210 158.820 1453.530 159.080 ;
        RECT 1453.300 158.400 1453.440 158.820 ;
        RECT 1453.210 158.140 1453.530 158.400 ;
        RECT 1453.670 110.400 1453.990 110.460 ;
        RECT 1454.590 110.400 1454.910 110.460 ;
        RECT 1453.670 110.260 1454.910 110.400 ;
        RECT 1453.670 110.200 1453.990 110.260 ;
        RECT 1454.590 110.200 1454.910 110.260 ;
        RECT 1453.670 96.460 1453.990 96.520 ;
        RECT 1454.590 96.460 1454.910 96.520 ;
        RECT 1453.670 96.320 1454.910 96.460 ;
        RECT 1453.670 96.260 1453.990 96.320 ;
        RECT 1454.590 96.260 1454.910 96.320 ;
        RECT 1453.670 62.120 1453.990 62.180 ;
        RECT 1454.590 62.120 1454.910 62.180 ;
        RECT 1453.670 61.980 1454.910 62.120 ;
        RECT 1453.670 61.920 1453.990 61.980 ;
        RECT 1454.590 61.920 1454.910 61.980 ;
        RECT 1454.590 18.260 1454.910 18.320 ;
        RECT 1518.990 18.260 1519.310 18.320 ;
        RECT 1454.590 18.120 1519.310 18.260 ;
        RECT 1454.590 18.060 1454.910 18.120 ;
        RECT 1518.990 18.060 1519.310 18.120 ;
      LAYER via ;
        RECT 1453.240 497.120 1453.500 497.380 ;
        RECT 1452.780 496.440 1453.040 496.700 ;
        RECT 1451.400 482.840 1451.660 483.100 ;
        RECT 1452.780 482.840 1453.040 483.100 ;
        RECT 1451.400 324.060 1451.660 324.320 ;
        RECT 1452.320 324.060 1452.580 324.320 ;
        RECT 1451.400 276.120 1451.660 276.380 ;
        RECT 1452.780 276.120 1453.040 276.380 ;
        RECT 1453.240 193.160 1453.500 193.420 ;
        RECT 1453.240 192.480 1453.500 192.740 ;
        RECT 1453.240 158.820 1453.500 159.080 ;
        RECT 1453.240 158.140 1453.500 158.400 ;
        RECT 1453.700 110.200 1453.960 110.460 ;
        RECT 1454.620 110.200 1454.880 110.460 ;
        RECT 1453.700 96.260 1453.960 96.520 ;
        RECT 1454.620 96.260 1454.880 96.520 ;
        RECT 1453.700 61.920 1453.960 62.180 ;
        RECT 1454.620 61.920 1454.880 62.180 ;
        RECT 1454.620 18.060 1454.880 18.320 ;
        RECT 1519.020 18.060 1519.280 18.320 ;
      LAYER met2 ;
        RECT 1452.090 600.170 1452.370 604.000 ;
        RECT 1452.090 600.030 1453.900 600.170 ;
        RECT 1452.090 600.000 1452.370 600.030 ;
        RECT 1453.760 583.170 1453.900 600.030 ;
        RECT 1453.760 583.030 1454.820 583.170 ;
        RECT 1454.680 565.490 1454.820 583.030 ;
        RECT 1454.220 565.350 1454.820 565.490 ;
        RECT 1454.220 545.090 1454.360 565.350 ;
        RECT 1453.300 544.950 1454.360 545.090 ;
        RECT 1453.300 497.410 1453.440 544.950 ;
        RECT 1453.240 497.090 1453.500 497.410 ;
        RECT 1452.780 496.410 1453.040 496.730 ;
        RECT 1452.840 483.130 1452.980 496.410 ;
        RECT 1451.400 482.810 1451.660 483.130 ;
        RECT 1452.780 482.810 1453.040 483.130 ;
        RECT 1451.460 435.045 1451.600 482.810 ;
        RECT 1451.390 434.675 1451.670 435.045 ;
        RECT 1452.310 434.675 1452.590 435.045 ;
        RECT 1452.380 399.570 1452.520 434.675 ;
        RECT 1452.380 399.430 1452.980 399.570 ;
        RECT 1452.840 338.485 1452.980 399.430 ;
        RECT 1452.770 338.115 1453.050 338.485 ;
        RECT 1452.310 331.315 1452.590 331.685 ;
        RECT 1452.380 324.350 1452.520 331.315 ;
        RECT 1451.400 324.030 1451.660 324.350 ;
        RECT 1452.320 324.030 1452.580 324.350 ;
        RECT 1451.460 276.410 1451.600 324.030 ;
        RECT 1451.400 276.090 1451.660 276.410 ;
        RECT 1452.780 276.090 1453.040 276.410 ;
        RECT 1452.840 234.330 1452.980 276.090 ;
        RECT 1452.840 234.190 1453.440 234.330 ;
        RECT 1453.300 193.450 1453.440 234.190 ;
        RECT 1453.240 193.130 1453.500 193.450 ;
        RECT 1453.240 192.450 1453.500 192.770 ;
        RECT 1453.300 159.110 1453.440 192.450 ;
        RECT 1453.240 158.790 1453.500 159.110 ;
        RECT 1453.240 158.110 1453.500 158.430 ;
        RECT 1453.300 110.570 1453.440 158.110 ;
        RECT 1453.300 110.490 1453.900 110.570 ;
        RECT 1453.300 110.430 1453.960 110.490 ;
        RECT 1453.700 110.170 1453.960 110.430 ;
        RECT 1454.620 110.170 1454.880 110.490 ;
        RECT 1454.680 96.550 1454.820 110.170 ;
        RECT 1453.700 96.230 1453.960 96.550 ;
        RECT 1454.620 96.230 1454.880 96.550 ;
        RECT 1453.760 62.210 1453.900 96.230 ;
        RECT 1453.700 61.890 1453.960 62.210 ;
        RECT 1454.620 61.890 1454.880 62.210 ;
        RECT 1454.680 18.350 1454.820 61.890 ;
        RECT 1454.620 18.030 1454.880 18.350 ;
        RECT 1519.020 18.030 1519.280 18.350 ;
        RECT 1519.080 2.400 1519.220 18.030 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
      LAYER via2 ;
        RECT 1451.390 434.720 1451.670 435.000 ;
        RECT 1452.310 434.720 1452.590 435.000 ;
        RECT 1452.770 338.160 1453.050 338.440 ;
        RECT 1452.310 331.360 1452.590 331.640 ;
      LAYER met3 ;
        RECT 1451.365 435.010 1451.695 435.025 ;
        RECT 1452.285 435.010 1452.615 435.025 ;
        RECT 1451.365 434.710 1452.615 435.010 ;
        RECT 1451.365 434.695 1451.695 434.710 ;
        RECT 1452.285 434.695 1452.615 434.710 ;
        RECT 1452.030 338.450 1452.410 338.460 ;
        RECT 1452.745 338.450 1453.075 338.465 ;
        RECT 1452.030 338.150 1453.075 338.450 ;
        RECT 1452.030 338.140 1452.410 338.150 ;
        RECT 1452.745 338.135 1453.075 338.150 ;
        RECT 1452.285 331.660 1452.615 331.665 ;
        RECT 1452.030 331.650 1452.615 331.660 ;
        RECT 1452.030 331.350 1452.840 331.650 ;
        RECT 1452.030 331.340 1452.615 331.350 ;
        RECT 1452.285 331.335 1452.615 331.340 ;
      LAYER via3 ;
        RECT 1452.060 338.140 1452.380 338.460 ;
        RECT 1452.060 331.340 1452.380 331.660 ;
      LAYER met4 ;
        RECT 1452.055 338.135 1452.385 338.465 ;
        RECT 1452.070 331.665 1452.370 338.135 ;
        RECT 1452.055 331.335 1452.385 331.665 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1037.370 579.600 1037.690 579.660 ;
        RECT 1037.830 579.600 1038.150 579.660 ;
        RECT 1037.370 579.460 1038.150 579.600 ;
        RECT 1037.370 579.400 1037.690 579.460 ;
        RECT 1037.830 579.400 1038.150 579.460 ;
        RECT 1035.990 496.980 1036.310 497.040 ;
        RECT 1036.910 496.980 1037.230 497.040 ;
        RECT 1035.990 496.840 1037.230 496.980 ;
        RECT 1035.990 496.780 1036.310 496.840 ;
        RECT 1036.910 496.780 1037.230 496.840 ;
        RECT 1035.990 483.040 1036.310 483.100 ;
        RECT 1036.450 483.040 1036.770 483.100 ;
        RECT 1035.990 482.900 1036.770 483.040 ;
        RECT 1035.990 482.840 1036.310 482.900 ;
        RECT 1036.450 482.840 1036.770 482.900 ;
        RECT 1036.450 448.700 1036.770 448.760 ;
        RECT 1036.080 448.560 1036.770 448.700 ;
        RECT 1036.080 448.420 1036.220 448.560 ;
        RECT 1036.450 448.500 1036.770 448.560 ;
        RECT 1035.990 448.160 1036.310 448.420 ;
        RECT 1034.610 410.620 1034.930 410.680 ;
        RECT 1036.450 410.620 1036.770 410.680 ;
        RECT 1034.610 410.480 1036.770 410.620 ;
        RECT 1034.610 410.420 1034.930 410.480 ;
        RECT 1036.450 410.420 1036.770 410.480 ;
        RECT 1034.610 386.480 1034.930 386.540 ;
        RECT 1035.530 386.480 1035.850 386.540 ;
        RECT 1034.610 386.340 1035.850 386.480 ;
        RECT 1034.610 386.280 1034.930 386.340 ;
        RECT 1035.530 386.280 1035.850 386.340 ;
        RECT 1034.610 355.540 1034.930 355.600 ;
        RECT 1035.530 355.540 1035.850 355.600 ;
        RECT 1034.610 355.400 1035.850 355.540 ;
        RECT 1034.610 355.340 1034.930 355.400 ;
        RECT 1035.530 355.340 1035.850 355.400 ;
        RECT 1034.610 331.400 1034.930 331.460 ;
        RECT 1035.990 331.400 1036.310 331.460 ;
        RECT 1034.610 331.260 1036.310 331.400 ;
        RECT 1034.610 331.200 1034.930 331.260 ;
        RECT 1035.990 331.200 1036.310 331.260 ;
        RECT 1035.530 289.720 1035.850 289.980 ;
        RECT 1034.610 289.240 1034.930 289.300 ;
        RECT 1035.620 289.240 1035.760 289.720 ;
        RECT 1034.610 289.100 1035.760 289.240 ;
        RECT 1034.610 289.040 1034.930 289.100 ;
        RECT 1034.610 241.980 1034.930 242.040 ;
        RECT 1037.370 241.980 1037.690 242.040 ;
        RECT 1034.610 241.840 1037.690 241.980 ;
        RECT 1034.610 241.780 1034.930 241.840 ;
        RECT 1037.370 241.780 1037.690 241.840 ;
        RECT 1036.450 234.500 1036.770 234.560 ;
        RECT 1037.370 234.500 1037.690 234.560 ;
        RECT 1036.450 234.360 1037.690 234.500 ;
        RECT 1036.450 234.300 1036.770 234.360 ;
        RECT 1037.370 234.300 1037.690 234.360 ;
        RECT 1036.450 186.560 1036.770 186.620 ;
        RECT 1037.370 186.560 1037.690 186.620 ;
        RECT 1036.450 186.420 1037.690 186.560 ;
        RECT 1036.450 186.360 1036.770 186.420 ;
        RECT 1037.370 186.360 1037.690 186.420 ;
        RECT 1037.370 145.080 1037.690 145.140 ;
        RECT 1037.370 144.940 1038.060 145.080 ;
        RECT 1037.370 144.880 1037.690 144.940 ;
        RECT 1037.920 144.800 1038.060 144.940 ;
        RECT 1037.830 144.540 1038.150 144.800 ;
        RECT 1037.370 138.280 1037.690 138.340 ;
        RECT 1037.830 138.280 1038.150 138.340 ;
        RECT 1037.370 138.140 1038.150 138.280 ;
        RECT 1037.370 138.080 1037.690 138.140 ;
        RECT 1037.830 138.080 1038.150 138.140 ;
        RECT 1035.530 90.000 1035.850 90.060 ;
        RECT 1036.910 90.000 1037.230 90.060 ;
        RECT 1035.530 89.860 1037.230 90.000 ;
        RECT 1035.530 89.800 1035.850 89.860 ;
        RECT 1036.910 89.800 1037.230 89.860 ;
        RECT 1010.230 54.980 1010.550 55.040 ;
        RECT 1035.990 54.980 1036.310 55.040 ;
        RECT 1010.230 54.840 1036.310 54.980 ;
        RECT 1010.230 54.780 1010.550 54.840 ;
        RECT 1035.990 54.780 1036.310 54.840 ;
        RECT 716.290 44.780 716.610 44.840 ;
        RECT 1010.230 44.780 1010.550 44.840 ;
        RECT 716.290 44.640 1010.550 44.780 ;
        RECT 716.290 44.580 716.610 44.640 ;
        RECT 1010.230 44.580 1010.550 44.640 ;
      LAYER via ;
        RECT 1037.400 579.400 1037.660 579.660 ;
        RECT 1037.860 579.400 1038.120 579.660 ;
        RECT 1036.020 496.780 1036.280 497.040 ;
        RECT 1036.940 496.780 1037.200 497.040 ;
        RECT 1036.020 482.840 1036.280 483.100 ;
        RECT 1036.480 482.840 1036.740 483.100 ;
        RECT 1036.480 448.500 1036.740 448.760 ;
        RECT 1036.020 448.160 1036.280 448.420 ;
        RECT 1034.640 410.420 1034.900 410.680 ;
        RECT 1036.480 410.420 1036.740 410.680 ;
        RECT 1034.640 386.280 1034.900 386.540 ;
        RECT 1035.560 386.280 1035.820 386.540 ;
        RECT 1034.640 355.340 1034.900 355.600 ;
        RECT 1035.560 355.340 1035.820 355.600 ;
        RECT 1034.640 331.200 1034.900 331.460 ;
        RECT 1036.020 331.200 1036.280 331.460 ;
        RECT 1035.560 289.720 1035.820 289.980 ;
        RECT 1034.640 289.040 1034.900 289.300 ;
        RECT 1034.640 241.780 1034.900 242.040 ;
        RECT 1037.400 241.780 1037.660 242.040 ;
        RECT 1036.480 234.300 1036.740 234.560 ;
        RECT 1037.400 234.300 1037.660 234.560 ;
        RECT 1036.480 186.360 1036.740 186.620 ;
        RECT 1037.400 186.360 1037.660 186.620 ;
        RECT 1037.400 144.880 1037.660 145.140 ;
        RECT 1037.860 144.540 1038.120 144.800 ;
        RECT 1037.400 138.080 1037.660 138.340 ;
        RECT 1037.860 138.080 1038.120 138.340 ;
        RECT 1035.560 89.800 1035.820 90.060 ;
        RECT 1036.940 89.800 1037.200 90.060 ;
        RECT 1010.260 54.780 1010.520 55.040 ;
        RECT 1036.020 54.780 1036.280 55.040 ;
        RECT 716.320 44.580 716.580 44.840 ;
        RECT 1010.260 44.580 1010.520 44.840 ;
      LAYER met2 ;
        RECT 1038.550 600.850 1038.830 604.000 ;
        RECT 1037.920 600.710 1038.830 600.850 ;
        RECT 1037.920 579.690 1038.060 600.710 ;
        RECT 1038.550 600.000 1038.830 600.710 ;
        RECT 1037.400 579.370 1037.660 579.690 ;
        RECT 1037.860 579.370 1038.120 579.690 ;
        RECT 1037.460 531.490 1037.600 579.370 ;
        RECT 1037.000 531.350 1037.600 531.490 ;
        RECT 1037.000 497.070 1037.140 531.350 ;
        RECT 1036.020 496.750 1036.280 497.070 ;
        RECT 1036.940 496.750 1037.200 497.070 ;
        RECT 1036.080 483.130 1036.220 496.750 ;
        RECT 1036.020 482.810 1036.280 483.130 ;
        RECT 1036.480 482.810 1036.740 483.130 ;
        RECT 1036.540 448.790 1036.680 482.810 ;
        RECT 1036.480 448.470 1036.740 448.790 ;
        RECT 1036.020 448.130 1036.280 448.450 ;
        RECT 1036.080 434.930 1036.220 448.130 ;
        RECT 1036.080 434.790 1036.680 434.930 ;
        RECT 1036.540 410.710 1036.680 434.790 ;
        RECT 1034.640 410.390 1034.900 410.710 ;
        RECT 1036.480 410.390 1036.740 410.710 ;
        RECT 1034.700 386.570 1034.840 410.390 ;
        RECT 1034.640 386.250 1034.900 386.570 ;
        RECT 1035.560 386.250 1035.820 386.570 ;
        RECT 1035.620 355.630 1035.760 386.250 ;
        RECT 1034.640 355.310 1034.900 355.630 ;
        RECT 1035.560 355.310 1035.820 355.630 ;
        RECT 1034.700 331.490 1034.840 355.310 ;
        RECT 1034.640 331.170 1034.900 331.490 ;
        RECT 1036.020 331.170 1036.280 331.490 ;
        RECT 1036.080 330.890 1036.220 331.170 ;
        RECT 1035.620 330.750 1036.220 330.890 ;
        RECT 1035.620 290.010 1035.760 330.750 ;
        RECT 1035.560 289.690 1035.820 290.010 ;
        RECT 1034.640 289.010 1034.900 289.330 ;
        RECT 1034.700 242.070 1034.840 289.010 ;
        RECT 1034.640 241.750 1034.900 242.070 ;
        RECT 1037.400 241.750 1037.660 242.070 ;
        RECT 1037.460 234.590 1037.600 241.750 ;
        RECT 1036.480 234.270 1036.740 234.590 ;
        RECT 1037.400 234.270 1037.660 234.590 ;
        RECT 1036.540 186.650 1036.680 234.270 ;
        RECT 1036.480 186.330 1036.740 186.650 ;
        RECT 1037.400 186.330 1037.660 186.650 ;
        RECT 1037.460 145.170 1037.600 186.330 ;
        RECT 1037.400 144.850 1037.660 145.170 ;
        RECT 1037.860 144.510 1038.120 144.830 ;
        RECT 1037.920 138.370 1038.060 144.510 ;
        RECT 1037.400 138.050 1037.660 138.370 ;
        RECT 1037.860 138.050 1038.120 138.370 ;
        RECT 1037.460 137.770 1037.600 138.050 ;
        RECT 1037.000 137.630 1037.600 137.770 ;
        RECT 1037.000 90.090 1037.140 137.630 ;
        RECT 1035.560 89.770 1035.820 90.090 ;
        RECT 1036.940 89.770 1037.200 90.090 ;
        RECT 1035.620 89.490 1035.760 89.770 ;
        RECT 1035.620 89.350 1036.220 89.490 ;
        RECT 1036.080 55.070 1036.220 89.350 ;
        RECT 1010.260 54.750 1010.520 55.070 ;
        RECT 1036.020 54.750 1036.280 55.070 ;
        RECT 1010.320 44.870 1010.460 54.750 ;
        RECT 716.320 44.550 716.580 44.870 ;
        RECT 1010.260 44.550 1010.520 44.870 ;
        RECT 716.380 2.400 716.520 44.550 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1461.950 20.640 1462.270 20.700 ;
        RECT 1536.930 20.640 1537.250 20.700 ;
        RECT 1461.950 20.500 1537.250 20.640 ;
        RECT 1461.950 20.440 1462.270 20.500 ;
        RECT 1536.930 20.440 1537.250 20.500 ;
      LAYER via ;
        RECT 1461.980 20.440 1462.240 20.700 ;
        RECT 1536.960 20.440 1537.220 20.700 ;
      LAYER met2 ;
        RECT 1461.290 600.170 1461.570 604.000 ;
        RECT 1461.290 600.030 1462.180 600.170 ;
        RECT 1461.290 600.000 1461.570 600.030 ;
        RECT 1462.040 20.730 1462.180 600.030 ;
        RECT 1461.980 20.410 1462.240 20.730 ;
        RECT 1536.960 20.410 1537.220 20.730 ;
        RECT 1537.020 2.400 1537.160 20.410 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1471.610 589.800 1471.930 589.860 ;
        RECT 1476.210 589.800 1476.530 589.860 ;
        RECT 1471.610 589.660 1476.530 589.800 ;
        RECT 1471.610 589.600 1471.930 589.660 ;
        RECT 1476.210 589.600 1476.530 589.660 ;
        RECT 1476.210 17.240 1476.530 17.300 ;
        RECT 1554.870 17.240 1555.190 17.300 ;
        RECT 1476.210 17.100 1555.190 17.240 ;
        RECT 1476.210 17.040 1476.530 17.100 ;
        RECT 1554.870 17.040 1555.190 17.100 ;
      LAYER via ;
        RECT 1471.640 589.600 1471.900 589.860 ;
        RECT 1476.240 589.600 1476.500 589.860 ;
        RECT 1476.240 17.040 1476.500 17.300 ;
        RECT 1554.900 17.040 1555.160 17.300 ;
      LAYER met2 ;
        RECT 1470.030 600.170 1470.310 604.000 ;
        RECT 1470.030 600.030 1471.840 600.170 ;
        RECT 1470.030 600.000 1470.310 600.030 ;
        RECT 1471.700 589.890 1471.840 600.030 ;
        RECT 1471.640 589.570 1471.900 589.890 ;
        RECT 1476.240 589.570 1476.500 589.890 ;
        RECT 1476.300 17.330 1476.440 589.570 ;
        RECT 1476.240 17.010 1476.500 17.330 ;
        RECT 1554.900 17.010 1555.160 17.330 ;
        RECT 1554.960 2.400 1555.100 17.010 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1480.810 591.500 1481.130 591.560 ;
        RECT 1528.190 591.500 1528.510 591.560 ;
        RECT 1480.810 591.360 1528.510 591.500 ;
        RECT 1480.810 591.300 1481.130 591.360 ;
        RECT 1528.190 591.300 1528.510 591.360 ;
        RECT 1528.190 17.580 1528.510 17.640 ;
        RECT 1531.410 17.580 1531.730 17.640 ;
        RECT 1528.190 17.440 1531.730 17.580 ;
        RECT 1528.190 17.380 1528.510 17.440 ;
        RECT 1531.410 17.380 1531.730 17.440 ;
        RECT 1531.410 16.560 1531.730 16.620 ;
        RECT 1572.810 16.560 1573.130 16.620 ;
        RECT 1531.410 16.420 1573.130 16.560 ;
        RECT 1531.410 16.360 1531.730 16.420 ;
        RECT 1572.810 16.360 1573.130 16.420 ;
      LAYER via ;
        RECT 1480.840 591.300 1481.100 591.560 ;
        RECT 1528.220 591.300 1528.480 591.560 ;
        RECT 1528.220 17.380 1528.480 17.640 ;
        RECT 1531.440 17.380 1531.700 17.640 ;
        RECT 1531.440 16.360 1531.700 16.620 ;
        RECT 1572.840 16.360 1573.100 16.620 ;
      LAYER met2 ;
        RECT 1479.230 600.170 1479.510 604.000 ;
        RECT 1479.230 600.030 1481.040 600.170 ;
        RECT 1479.230 600.000 1479.510 600.030 ;
        RECT 1480.900 591.590 1481.040 600.030 ;
        RECT 1480.840 591.270 1481.100 591.590 ;
        RECT 1528.220 591.270 1528.480 591.590 ;
        RECT 1528.280 17.670 1528.420 591.270 ;
        RECT 1528.220 17.350 1528.480 17.670 ;
        RECT 1531.440 17.350 1531.700 17.670 ;
        RECT 1531.500 16.650 1531.640 17.350 ;
        RECT 1531.440 16.330 1531.700 16.650 ;
        RECT 1572.840 16.330 1573.100 16.650 ;
        RECT 1572.900 2.400 1573.040 16.330 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1489.550 20.100 1489.870 20.360 ;
        RECT 1489.640 19.960 1489.780 20.100 ;
        RECT 1590.290 19.960 1590.610 20.020 ;
        RECT 1489.640 19.820 1590.610 19.960 ;
        RECT 1590.290 19.760 1590.610 19.820 ;
      LAYER via ;
        RECT 1489.580 20.100 1489.840 20.360 ;
        RECT 1590.320 19.760 1590.580 20.020 ;
      LAYER met2 ;
        RECT 1488.430 600.170 1488.710 604.000 ;
        RECT 1488.430 600.030 1489.780 600.170 ;
        RECT 1488.430 600.000 1488.710 600.030 ;
        RECT 1489.640 20.390 1489.780 600.030 ;
        RECT 1489.580 20.070 1489.840 20.390 ;
        RECT 1590.320 19.730 1590.580 20.050 ;
        RECT 1590.380 2.400 1590.520 19.730 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1499.210 587.760 1499.530 587.820 ;
        RECT 1576.490 587.760 1576.810 587.820 ;
        RECT 1499.210 587.620 1576.810 587.760 ;
        RECT 1499.210 587.560 1499.530 587.620 ;
        RECT 1576.490 587.560 1576.810 587.620 ;
        RECT 1576.490 20.640 1576.810 20.700 ;
        RECT 1579.250 20.640 1579.570 20.700 ;
        RECT 1576.490 20.500 1579.570 20.640 ;
        RECT 1576.490 20.440 1576.810 20.500 ;
        RECT 1579.250 20.440 1579.570 20.500 ;
        RECT 1579.250 16.220 1579.570 16.280 ;
        RECT 1608.230 16.220 1608.550 16.280 ;
        RECT 1579.250 16.080 1608.550 16.220 ;
        RECT 1579.250 16.020 1579.570 16.080 ;
        RECT 1608.230 16.020 1608.550 16.080 ;
      LAYER via ;
        RECT 1499.240 587.560 1499.500 587.820 ;
        RECT 1576.520 587.560 1576.780 587.820 ;
        RECT 1576.520 20.440 1576.780 20.700 ;
        RECT 1579.280 20.440 1579.540 20.700 ;
        RECT 1579.280 16.020 1579.540 16.280 ;
        RECT 1608.260 16.020 1608.520 16.280 ;
      LAYER met2 ;
        RECT 1497.630 600.170 1497.910 604.000 ;
        RECT 1497.630 600.030 1499.440 600.170 ;
        RECT 1497.630 600.000 1497.910 600.030 ;
        RECT 1499.300 587.850 1499.440 600.030 ;
        RECT 1499.240 587.530 1499.500 587.850 ;
        RECT 1576.520 587.530 1576.780 587.850 ;
        RECT 1576.580 20.730 1576.720 587.530 ;
        RECT 1576.520 20.410 1576.780 20.730 ;
        RECT 1579.280 20.410 1579.540 20.730 ;
        RECT 1579.340 16.310 1579.480 20.410 ;
        RECT 1579.280 15.990 1579.540 16.310 ;
        RECT 1608.260 15.990 1608.520 16.310 ;
        RECT 1608.320 2.400 1608.460 15.990 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1508.410 579.600 1508.730 579.660 ;
        RECT 1509.790 579.600 1510.110 579.660 ;
        RECT 1508.410 579.460 1510.110 579.600 ;
        RECT 1508.410 579.400 1508.730 579.460 ;
        RECT 1509.790 579.400 1510.110 579.460 ;
        RECT 1509.790 531.320 1510.110 531.380 ;
        RECT 1510.250 531.320 1510.570 531.380 ;
        RECT 1509.790 531.180 1510.570 531.320 ;
        RECT 1509.790 531.120 1510.110 531.180 ;
        RECT 1510.250 531.120 1510.570 531.180 ;
        RECT 1510.250 496.980 1510.570 497.040 ;
        RECT 1509.880 496.840 1510.570 496.980 ;
        RECT 1509.880 496.700 1510.020 496.840 ;
        RECT 1510.250 496.780 1510.570 496.840 ;
        RECT 1509.790 496.440 1510.110 496.700 ;
        RECT 1509.330 386.820 1509.650 386.880 ;
        RECT 1510.250 386.820 1510.570 386.880 ;
        RECT 1509.330 386.680 1510.570 386.820 ;
        RECT 1509.330 386.620 1509.650 386.680 ;
        RECT 1510.250 386.620 1510.570 386.680 ;
        RECT 1509.790 338.200 1510.110 338.260 ;
        RECT 1511.630 338.200 1511.950 338.260 ;
        RECT 1509.790 338.060 1511.950 338.200 ;
        RECT 1509.790 338.000 1510.110 338.060 ;
        RECT 1511.630 338.000 1511.950 338.060 ;
        RECT 1508.870 289.920 1509.190 289.980 ;
        RECT 1510.250 289.920 1510.570 289.980 ;
        RECT 1508.870 289.780 1510.570 289.920 ;
        RECT 1508.870 289.720 1509.190 289.780 ;
        RECT 1510.250 289.720 1510.570 289.780 ;
        RECT 1507.490 241.640 1507.810 241.700 ;
        RECT 1509.330 241.640 1509.650 241.700 ;
        RECT 1507.490 241.500 1509.650 241.640 ;
        RECT 1507.490 241.440 1507.810 241.500 ;
        RECT 1509.330 241.440 1509.650 241.500 ;
        RECT 1509.790 169.220 1510.110 169.280 ;
        RECT 1511.170 169.220 1511.490 169.280 ;
        RECT 1509.790 169.080 1511.490 169.220 ;
        RECT 1509.790 169.020 1510.110 169.080 ;
        RECT 1511.170 169.020 1511.490 169.080 ;
        RECT 1508.410 137.940 1508.730 138.000 ;
        RECT 1509.790 137.940 1510.110 138.000 ;
        RECT 1508.410 137.800 1510.110 137.940 ;
        RECT 1508.410 137.740 1508.730 137.800 ;
        RECT 1509.790 137.740 1510.110 137.800 ;
        RECT 1508.410 90.000 1508.730 90.060 ;
        RECT 1509.330 90.000 1509.650 90.060 ;
        RECT 1508.410 89.860 1509.650 90.000 ;
        RECT 1508.410 89.800 1508.730 89.860 ;
        RECT 1509.330 89.800 1509.650 89.860 ;
        RECT 1509.330 48.520 1509.650 48.580 ;
        RECT 1510.250 48.520 1510.570 48.580 ;
        RECT 1509.330 48.380 1510.570 48.520 ;
        RECT 1509.330 48.320 1509.650 48.380 ;
        RECT 1510.250 48.320 1510.570 48.380 ;
        RECT 1510.250 18.940 1510.570 19.000 ;
        RECT 1626.170 18.940 1626.490 19.000 ;
        RECT 1510.250 18.800 1626.490 18.940 ;
        RECT 1510.250 18.740 1510.570 18.800 ;
        RECT 1626.170 18.740 1626.490 18.800 ;
      LAYER via ;
        RECT 1508.440 579.400 1508.700 579.660 ;
        RECT 1509.820 579.400 1510.080 579.660 ;
        RECT 1509.820 531.120 1510.080 531.380 ;
        RECT 1510.280 531.120 1510.540 531.380 ;
        RECT 1510.280 496.780 1510.540 497.040 ;
        RECT 1509.820 496.440 1510.080 496.700 ;
        RECT 1509.360 386.620 1509.620 386.880 ;
        RECT 1510.280 386.620 1510.540 386.880 ;
        RECT 1509.820 338.000 1510.080 338.260 ;
        RECT 1511.660 338.000 1511.920 338.260 ;
        RECT 1508.900 289.720 1509.160 289.980 ;
        RECT 1510.280 289.720 1510.540 289.980 ;
        RECT 1507.520 241.440 1507.780 241.700 ;
        RECT 1509.360 241.440 1509.620 241.700 ;
        RECT 1509.820 169.020 1510.080 169.280 ;
        RECT 1511.200 169.020 1511.460 169.280 ;
        RECT 1508.440 137.740 1508.700 138.000 ;
        RECT 1509.820 137.740 1510.080 138.000 ;
        RECT 1508.440 89.800 1508.700 90.060 ;
        RECT 1509.360 89.800 1509.620 90.060 ;
        RECT 1509.360 48.320 1509.620 48.580 ;
        RECT 1510.280 48.320 1510.540 48.580 ;
        RECT 1510.280 18.740 1510.540 19.000 ;
        RECT 1626.200 18.740 1626.460 19.000 ;
      LAYER met2 ;
        RECT 1506.830 600.000 1507.110 604.000 ;
        RECT 1506.890 598.810 1507.030 600.000 ;
        RECT 1506.890 598.670 1507.260 598.810 ;
        RECT 1507.120 580.565 1507.260 598.670 ;
        RECT 1507.050 580.195 1507.330 580.565 ;
        RECT 1508.890 579.770 1509.170 579.885 ;
        RECT 1508.500 579.690 1509.170 579.770 ;
        RECT 1508.440 579.630 1509.170 579.690 ;
        RECT 1508.440 579.370 1508.700 579.630 ;
        RECT 1508.890 579.515 1509.170 579.630 ;
        RECT 1509.820 579.370 1510.080 579.690 ;
        RECT 1508.500 579.215 1508.640 579.370 ;
        RECT 1509.880 531.410 1510.020 579.370 ;
        RECT 1509.820 531.090 1510.080 531.410 ;
        RECT 1510.280 531.090 1510.540 531.410 ;
        RECT 1510.340 497.070 1510.480 531.090 ;
        RECT 1510.280 496.750 1510.540 497.070 ;
        RECT 1509.820 496.410 1510.080 496.730 ;
        RECT 1509.880 483.210 1510.020 496.410 ;
        RECT 1509.880 483.070 1510.480 483.210 ;
        RECT 1510.340 448.530 1510.480 483.070 ;
        RECT 1509.420 448.390 1510.480 448.530 ;
        RECT 1509.420 386.910 1509.560 448.390 ;
        RECT 1509.360 386.590 1509.620 386.910 ;
        RECT 1510.280 386.590 1510.540 386.910 ;
        RECT 1510.340 386.085 1510.480 386.590 ;
        RECT 1510.270 385.715 1510.550 386.085 ;
        RECT 1511.650 385.715 1511.930 386.085 ;
        RECT 1511.720 338.290 1511.860 385.715 ;
        RECT 1509.820 337.970 1510.080 338.290 ;
        RECT 1511.660 337.970 1511.920 338.290 ;
        RECT 1509.880 304.370 1510.020 337.970 ;
        RECT 1509.880 304.230 1510.480 304.370 ;
        RECT 1510.340 290.010 1510.480 304.230 ;
        RECT 1508.900 289.690 1509.160 290.010 ;
        RECT 1510.280 289.690 1510.540 290.010 ;
        RECT 1508.960 289.525 1509.100 289.690 ;
        RECT 1507.510 289.155 1507.790 289.525 ;
        RECT 1508.890 289.155 1509.170 289.525 ;
        RECT 1507.580 241.730 1507.720 289.155 ;
        RECT 1507.520 241.410 1507.780 241.730 ;
        RECT 1509.360 241.410 1509.620 241.730 ;
        RECT 1509.420 207.130 1509.560 241.410 ;
        RECT 1509.420 206.990 1510.020 207.130 ;
        RECT 1509.880 169.310 1510.020 206.990 ;
        RECT 1509.820 168.990 1510.080 169.310 ;
        RECT 1511.200 168.990 1511.460 169.310 ;
        RECT 1511.260 145.365 1511.400 168.990 ;
        RECT 1510.270 145.250 1510.550 145.365 ;
        RECT 1509.880 145.110 1510.550 145.250 ;
        RECT 1509.880 138.030 1510.020 145.110 ;
        RECT 1510.270 144.995 1510.550 145.110 ;
        RECT 1511.190 144.995 1511.470 145.365 ;
        RECT 1508.440 137.710 1508.700 138.030 ;
        RECT 1509.820 137.710 1510.080 138.030 ;
        RECT 1508.500 90.090 1508.640 137.710 ;
        RECT 1508.440 89.770 1508.700 90.090 ;
        RECT 1509.360 89.770 1509.620 90.090 ;
        RECT 1509.420 48.610 1509.560 89.770 ;
        RECT 1509.360 48.290 1509.620 48.610 ;
        RECT 1510.280 48.290 1510.540 48.610 ;
        RECT 1510.340 19.030 1510.480 48.290 ;
        RECT 1510.280 18.710 1510.540 19.030 ;
        RECT 1626.200 18.710 1626.460 19.030 ;
        RECT 1626.260 2.400 1626.400 18.710 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
      LAYER via2 ;
        RECT 1507.050 580.240 1507.330 580.520 ;
        RECT 1508.890 579.560 1509.170 579.840 ;
        RECT 1510.270 385.760 1510.550 386.040 ;
        RECT 1511.650 385.760 1511.930 386.040 ;
        RECT 1507.510 289.200 1507.790 289.480 ;
        RECT 1508.890 289.200 1509.170 289.480 ;
        RECT 1510.270 145.040 1510.550 145.320 ;
        RECT 1511.190 145.040 1511.470 145.320 ;
      LAYER met3 ;
        RECT 1507.025 580.530 1507.355 580.545 ;
        RECT 1507.025 580.230 1509.410 580.530 ;
        RECT 1507.025 580.215 1507.355 580.230 ;
        RECT 1509.110 579.865 1509.410 580.230 ;
        RECT 1508.865 579.550 1509.410 579.865 ;
        RECT 1508.865 579.535 1509.195 579.550 ;
        RECT 1510.245 386.050 1510.575 386.065 ;
        RECT 1511.625 386.050 1511.955 386.065 ;
        RECT 1510.245 385.750 1511.955 386.050 ;
        RECT 1510.245 385.735 1510.575 385.750 ;
        RECT 1511.625 385.735 1511.955 385.750 ;
        RECT 1507.485 289.490 1507.815 289.505 ;
        RECT 1508.865 289.490 1509.195 289.505 ;
        RECT 1507.485 289.190 1509.195 289.490 ;
        RECT 1507.485 289.175 1507.815 289.190 ;
        RECT 1508.865 289.175 1509.195 289.190 ;
        RECT 1510.245 145.330 1510.575 145.345 ;
        RECT 1511.165 145.330 1511.495 145.345 ;
        RECT 1510.245 145.030 1511.495 145.330 ;
        RECT 1510.245 145.015 1510.575 145.030 ;
        RECT 1511.165 145.015 1511.495 145.030 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.150 17.920 1517.470 17.980 ;
        RECT 1644.110 17.920 1644.430 17.980 ;
        RECT 1517.150 17.780 1644.430 17.920 ;
        RECT 1517.150 17.720 1517.470 17.780 ;
        RECT 1644.110 17.720 1644.430 17.780 ;
      LAYER via ;
        RECT 1517.180 17.720 1517.440 17.980 ;
        RECT 1644.140 17.720 1644.400 17.980 ;
      LAYER met2 ;
        RECT 1516.030 600.170 1516.310 604.000 ;
        RECT 1516.030 600.030 1517.380 600.170 ;
        RECT 1516.030 600.000 1516.310 600.030 ;
        RECT 1517.240 18.010 1517.380 600.030 ;
        RECT 1517.180 17.690 1517.440 18.010 ;
        RECT 1644.140 17.690 1644.400 18.010 ;
        RECT 1644.200 2.400 1644.340 17.690 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1526.810 586.740 1527.130 586.800 ;
        RECT 1531.410 586.740 1531.730 586.800 ;
        RECT 1526.810 586.600 1531.730 586.740 ;
        RECT 1526.810 586.540 1527.130 586.600 ;
        RECT 1531.410 586.540 1531.730 586.600 ;
        RECT 1531.410 18.260 1531.730 18.320 ;
        RECT 1662.050 18.260 1662.370 18.320 ;
        RECT 1531.410 18.120 1662.370 18.260 ;
        RECT 1531.410 18.060 1531.730 18.120 ;
        RECT 1662.050 18.060 1662.370 18.120 ;
      LAYER via ;
        RECT 1526.840 586.540 1527.100 586.800 ;
        RECT 1531.440 586.540 1531.700 586.800 ;
        RECT 1531.440 18.060 1531.700 18.320 ;
        RECT 1662.080 18.060 1662.340 18.320 ;
      LAYER met2 ;
        RECT 1525.230 600.170 1525.510 604.000 ;
        RECT 1525.230 600.030 1527.040 600.170 ;
        RECT 1525.230 600.000 1525.510 600.030 ;
        RECT 1526.900 586.830 1527.040 600.030 ;
        RECT 1526.840 586.510 1527.100 586.830 ;
        RECT 1531.440 586.510 1531.700 586.830 ;
        RECT 1531.500 18.350 1531.640 586.510 ;
        RECT 1531.440 18.030 1531.700 18.350 ;
        RECT 1662.080 18.030 1662.340 18.350 ;
        RECT 1662.140 2.400 1662.280 18.030 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1536.010 591.500 1536.330 591.560 ;
        RECT 1673.090 591.500 1673.410 591.560 ;
        RECT 1536.010 591.360 1673.410 591.500 ;
        RECT 1536.010 591.300 1536.330 591.360 ;
        RECT 1673.090 591.300 1673.410 591.360 ;
        RECT 1673.090 25.060 1673.410 25.120 ;
        RECT 1679.530 25.060 1679.850 25.120 ;
        RECT 1673.090 24.920 1679.850 25.060 ;
        RECT 1673.090 24.860 1673.410 24.920 ;
        RECT 1679.530 24.860 1679.850 24.920 ;
      LAYER via ;
        RECT 1536.040 591.300 1536.300 591.560 ;
        RECT 1673.120 591.300 1673.380 591.560 ;
        RECT 1673.120 24.860 1673.380 25.120 ;
        RECT 1679.560 24.860 1679.820 25.120 ;
      LAYER met2 ;
        RECT 1534.430 600.170 1534.710 604.000 ;
        RECT 1534.430 600.030 1536.240 600.170 ;
        RECT 1534.430 600.000 1534.710 600.030 ;
        RECT 1536.100 591.590 1536.240 600.030 ;
        RECT 1536.040 591.270 1536.300 591.590 ;
        RECT 1673.120 591.270 1673.380 591.590 ;
        RECT 1673.180 25.150 1673.320 591.270 ;
        RECT 1673.120 24.830 1673.380 25.150 ;
        RECT 1679.560 24.830 1679.820 25.150 ;
        RECT 1679.620 2.400 1679.760 24.830 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 17.580 1545.530 17.640 ;
        RECT 1697.470 17.580 1697.790 17.640 ;
        RECT 1545.210 17.440 1697.790 17.580 ;
        RECT 1545.210 17.380 1545.530 17.440 ;
        RECT 1697.470 17.380 1697.790 17.440 ;
      LAYER via ;
        RECT 1545.240 17.380 1545.500 17.640 ;
        RECT 1697.500 17.380 1697.760 17.640 ;
      LAYER met2 ;
        RECT 1543.630 600.170 1543.910 604.000 ;
        RECT 1543.630 600.030 1545.440 600.170 ;
        RECT 1543.630 600.000 1543.910 600.030 ;
        RECT 1545.300 17.670 1545.440 600.030 ;
        RECT 1545.240 17.350 1545.500 17.670 ;
        RECT 1697.500 17.350 1697.760 17.670 ;
        RECT 1697.560 2.400 1697.700 17.350 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1042.430 569.400 1042.750 569.460 ;
        RECT 1046.110 569.400 1046.430 569.460 ;
        RECT 1042.430 569.260 1046.430 569.400 ;
        RECT 1042.430 569.200 1042.750 569.260 ;
        RECT 1046.110 569.200 1046.430 569.260 ;
        RECT 841.410 21.320 841.730 21.380 ;
        RECT 1042.430 21.320 1042.750 21.380 ;
        RECT 841.410 21.180 1042.750 21.320 ;
        RECT 841.410 21.120 841.730 21.180 ;
        RECT 1042.430 21.120 1042.750 21.180 ;
        RECT 734.230 18.600 734.550 18.660 ;
        RECT 841.410 18.600 841.730 18.660 ;
        RECT 734.230 18.460 841.730 18.600 ;
        RECT 734.230 18.400 734.550 18.460 ;
        RECT 841.410 18.400 841.730 18.460 ;
      LAYER via ;
        RECT 1042.460 569.200 1042.720 569.460 ;
        RECT 1046.140 569.200 1046.400 569.460 ;
        RECT 841.440 21.120 841.700 21.380 ;
        RECT 1042.460 21.120 1042.720 21.380 ;
        RECT 734.260 18.400 734.520 18.660 ;
        RECT 841.440 18.400 841.700 18.660 ;
      LAYER met2 ;
        RECT 1047.750 600.170 1048.030 604.000 ;
        RECT 1046.200 600.030 1048.030 600.170 ;
        RECT 1046.200 569.490 1046.340 600.030 ;
        RECT 1047.750 600.000 1048.030 600.030 ;
        RECT 1042.460 569.170 1042.720 569.490 ;
        RECT 1046.140 569.170 1046.400 569.490 ;
        RECT 1042.520 21.410 1042.660 569.170 ;
        RECT 841.440 21.090 841.700 21.410 ;
        RECT 1042.460 21.090 1042.720 21.410 ;
        RECT 841.500 18.690 841.640 21.090 ;
        RECT 734.260 18.370 734.520 18.690 ;
        RECT 841.440 18.370 841.700 18.690 ;
        RECT 734.320 2.400 734.460 18.370 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1554.410 592.520 1554.730 592.580 ;
        RECT 1706.210 592.520 1706.530 592.580 ;
        RECT 1554.410 592.380 1706.530 592.520 ;
        RECT 1554.410 592.320 1554.730 592.380 ;
        RECT 1706.210 592.320 1706.530 592.380 ;
        RECT 1704.830 579.600 1705.150 579.660 ;
        RECT 1706.210 579.600 1706.530 579.660 ;
        RECT 1704.830 579.460 1706.530 579.600 ;
        RECT 1704.830 579.400 1705.150 579.460 ;
        RECT 1706.210 579.400 1706.530 579.460 ;
        RECT 1704.830 531.660 1705.150 531.720 ;
        RECT 1705.750 531.660 1706.070 531.720 ;
        RECT 1704.830 531.520 1706.070 531.660 ;
        RECT 1704.830 531.460 1705.150 531.520 ;
        RECT 1705.750 531.460 1706.070 531.520 ;
        RECT 1705.750 496.780 1706.070 497.040 ;
        RECT 1705.840 496.640 1705.980 496.780 ;
        RECT 1706.670 496.640 1706.990 496.700 ;
        RECT 1705.840 496.500 1706.990 496.640 ;
        RECT 1706.670 496.440 1706.990 496.500 ;
        RECT 1705.290 483.040 1705.610 483.100 ;
        RECT 1706.670 483.040 1706.990 483.100 ;
        RECT 1705.290 482.900 1706.990 483.040 ;
        RECT 1705.290 482.840 1705.610 482.900 ;
        RECT 1706.670 482.840 1706.990 482.900 ;
        RECT 1706.670 385.800 1706.990 385.860 ;
        RECT 1708.050 385.800 1708.370 385.860 ;
        RECT 1706.670 385.660 1708.370 385.800 ;
        RECT 1706.670 385.600 1706.990 385.660 ;
        RECT 1708.050 385.600 1708.370 385.660 ;
        RECT 1707.130 338.200 1707.450 338.260 ;
        RECT 1708.050 338.200 1708.370 338.260 ;
        RECT 1707.130 338.060 1708.370 338.200 ;
        RECT 1707.130 338.000 1707.450 338.060 ;
        RECT 1708.050 338.000 1708.370 338.060 ;
        RECT 1707.590 265.780 1707.910 265.840 ;
        RECT 1708.970 265.780 1709.290 265.840 ;
        RECT 1707.590 265.640 1709.290 265.780 ;
        RECT 1707.590 265.580 1707.910 265.640 ;
        RECT 1708.970 265.580 1709.290 265.640 ;
        RECT 1706.210 234.500 1706.530 234.560 ;
        RECT 1707.590 234.500 1707.910 234.560 ;
        RECT 1706.210 234.360 1707.910 234.500 ;
        RECT 1706.210 234.300 1706.530 234.360 ;
        RECT 1707.590 234.300 1707.910 234.360 ;
        RECT 1706.210 186.560 1706.530 186.620 ;
        RECT 1707.130 186.560 1707.450 186.620 ;
        RECT 1706.210 186.420 1707.450 186.560 ;
        RECT 1706.210 186.360 1706.530 186.420 ;
        RECT 1707.130 186.360 1707.450 186.420 ;
        RECT 1708.050 17.920 1708.370 17.980 ;
        RECT 1715.410 17.920 1715.730 17.980 ;
        RECT 1708.050 17.780 1715.730 17.920 ;
        RECT 1708.050 17.720 1708.370 17.780 ;
        RECT 1715.410 17.720 1715.730 17.780 ;
      LAYER via ;
        RECT 1554.440 592.320 1554.700 592.580 ;
        RECT 1706.240 592.320 1706.500 592.580 ;
        RECT 1704.860 579.400 1705.120 579.660 ;
        RECT 1706.240 579.400 1706.500 579.660 ;
        RECT 1704.860 531.460 1705.120 531.720 ;
        RECT 1705.780 531.460 1706.040 531.720 ;
        RECT 1705.780 496.780 1706.040 497.040 ;
        RECT 1706.700 496.440 1706.960 496.700 ;
        RECT 1705.320 482.840 1705.580 483.100 ;
        RECT 1706.700 482.840 1706.960 483.100 ;
        RECT 1706.700 385.600 1706.960 385.860 ;
        RECT 1708.080 385.600 1708.340 385.860 ;
        RECT 1707.160 338.000 1707.420 338.260 ;
        RECT 1708.080 338.000 1708.340 338.260 ;
        RECT 1707.620 265.580 1707.880 265.840 ;
        RECT 1709.000 265.580 1709.260 265.840 ;
        RECT 1706.240 234.300 1706.500 234.560 ;
        RECT 1707.620 234.300 1707.880 234.560 ;
        RECT 1706.240 186.360 1706.500 186.620 ;
        RECT 1707.160 186.360 1707.420 186.620 ;
        RECT 1708.080 17.720 1708.340 17.980 ;
        RECT 1715.440 17.720 1715.700 17.980 ;
      LAYER met2 ;
        RECT 1552.830 600.170 1553.110 604.000 ;
        RECT 1552.830 600.030 1554.640 600.170 ;
        RECT 1552.830 600.000 1553.110 600.030 ;
        RECT 1554.500 592.610 1554.640 600.030 ;
        RECT 1554.440 592.290 1554.700 592.610 ;
        RECT 1706.240 592.290 1706.500 592.610 ;
        RECT 1706.300 579.690 1706.440 592.290 ;
        RECT 1704.860 579.370 1705.120 579.690 ;
        RECT 1706.240 579.370 1706.500 579.690 ;
        RECT 1704.920 531.750 1705.060 579.370 ;
        RECT 1704.860 531.430 1705.120 531.750 ;
        RECT 1705.780 531.430 1706.040 531.750 ;
        RECT 1705.840 497.070 1705.980 531.430 ;
        RECT 1705.780 496.750 1706.040 497.070 ;
        RECT 1706.700 496.410 1706.960 496.730 ;
        RECT 1706.760 483.130 1706.900 496.410 ;
        RECT 1705.320 482.810 1705.580 483.130 ;
        RECT 1706.700 482.810 1706.960 483.130 ;
        RECT 1705.380 435.045 1705.520 482.810 ;
        RECT 1705.310 434.675 1705.590 435.045 ;
        RECT 1706.230 434.675 1706.510 435.045 ;
        RECT 1706.300 399.570 1706.440 434.675 ;
        RECT 1706.300 399.430 1706.900 399.570 ;
        RECT 1706.760 385.890 1706.900 399.430 ;
        RECT 1706.700 385.570 1706.960 385.890 ;
        RECT 1708.080 385.570 1708.340 385.890 ;
        RECT 1708.140 338.290 1708.280 385.570 ;
        RECT 1707.160 337.970 1707.420 338.290 ;
        RECT 1708.080 337.970 1708.340 338.290 ;
        RECT 1707.220 303.690 1707.360 337.970 ;
        RECT 1707.220 303.550 1707.820 303.690 ;
        RECT 1707.680 265.870 1707.820 303.550 ;
        RECT 1707.620 265.550 1707.880 265.870 ;
        RECT 1709.000 265.550 1709.260 265.870 ;
        RECT 1709.060 241.925 1709.200 265.550 ;
        RECT 1708.070 241.810 1708.350 241.925 ;
        RECT 1707.680 241.670 1708.350 241.810 ;
        RECT 1707.680 234.590 1707.820 241.670 ;
        RECT 1708.070 241.555 1708.350 241.670 ;
        RECT 1708.990 241.555 1709.270 241.925 ;
        RECT 1706.240 234.270 1706.500 234.590 ;
        RECT 1707.620 234.270 1707.880 234.590 ;
        RECT 1706.300 186.650 1706.440 234.270 ;
        RECT 1706.240 186.330 1706.500 186.650 ;
        RECT 1707.160 186.330 1707.420 186.650 ;
        RECT 1707.220 158.170 1707.360 186.330 ;
        RECT 1707.220 158.030 1707.820 158.170 ;
        RECT 1707.680 62.290 1707.820 158.030 ;
        RECT 1707.680 62.150 1708.280 62.290 ;
        RECT 1708.140 18.010 1708.280 62.150 ;
        RECT 1708.080 17.690 1708.340 18.010 ;
        RECT 1715.440 17.690 1715.700 18.010 ;
        RECT 1715.500 2.400 1715.640 17.690 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
      LAYER via2 ;
        RECT 1705.310 434.720 1705.590 435.000 ;
        RECT 1706.230 434.720 1706.510 435.000 ;
        RECT 1708.070 241.600 1708.350 241.880 ;
        RECT 1708.990 241.600 1709.270 241.880 ;
      LAYER met3 ;
        RECT 1705.285 435.010 1705.615 435.025 ;
        RECT 1706.205 435.010 1706.535 435.025 ;
        RECT 1705.285 434.710 1706.535 435.010 ;
        RECT 1705.285 434.695 1705.615 434.710 ;
        RECT 1706.205 434.695 1706.535 434.710 ;
        RECT 1708.045 241.890 1708.375 241.905 ;
        RECT 1708.965 241.890 1709.295 241.905 ;
        RECT 1708.045 241.590 1709.295 241.890 ;
        RECT 1708.045 241.575 1708.375 241.590 ;
        RECT 1708.965 241.575 1709.295 241.590 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1563.610 586.740 1563.930 586.800 ;
        RECT 1565.910 586.740 1566.230 586.800 ;
        RECT 1563.610 586.600 1566.230 586.740 ;
        RECT 1563.610 586.540 1563.930 586.600 ;
        RECT 1565.910 586.540 1566.230 586.600 ;
        RECT 1565.910 17.240 1566.230 17.300 ;
        RECT 1733.350 17.240 1733.670 17.300 ;
        RECT 1565.910 17.100 1733.670 17.240 ;
        RECT 1565.910 17.040 1566.230 17.100 ;
        RECT 1733.350 17.040 1733.670 17.100 ;
      LAYER via ;
        RECT 1563.640 586.540 1563.900 586.800 ;
        RECT 1565.940 586.540 1566.200 586.800 ;
        RECT 1565.940 17.040 1566.200 17.300 ;
        RECT 1733.380 17.040 1733.640 17.300 ;
      LAYER met2 ;
        RECT 1562.030 600.170 1562.310 604.000 ;
        RECT 1562.030 600.030 1563.840 600.170 ;
        RECT 1562.030 600.000 1562.310 600.030 ;
        RECT 1563.700 586.830 1563.840 600.030 ;
        RECT 1563.640 586.510 1563.900 586.830 ;
        RECT 1565.940 586.510 1566.200 586.830 ;
        RECT 1566.000 17.330 1566.140 586.510 ;
        RECT 1565.940 17.010 1566.200 17.330 ;
        RECT 1733.380 17.010 1733.640 17.330 ;
        RECT 1733.440 2.400 1733.580 17.010 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.810 588.100 1573.130 588.160 ;
        RECT 1604.090 588.100 1604.410 588.160 ;
        RECT 1572.810 587.960 1604.410 588.100 ;
        RECT 1572.810 587.900 1573.130 587.960 ;
        RECT 1604.090 587.900 1604.410 587.960 ;
        RECT 1604.090 15.880 1604.410 15.940 ;
        RECT 1751.290 15.880 1751.610 15.940 ;
        RECT 1604.090 15.740 1751.610 15.880 ;
        RECT 1604.090 15.680 1604.410 15.740 ;
        RECT 1751.290 15.680 1751.610 15.740 ;
      LAYER via ;
        RECT 1572.840 587.900 1573.100 588.160 ;
        RECT 1604.120 587.900 1604.380 588.160 ;
        RECT 1604.120 15.680 1604.380 15.940 ;
        RECT 1751.320 15.680 1751.580 15.940 ;
      LAYER met2 ;
        RECT 1571.230 600.170 1571.510 604.000 ;
        RECT 1571.230 600.030 1573.040 600.170 ;
        RECT 1571.230 600.000 1571.510 600.030 ;
        RECT 1572.900 588.190 1573.040 600.030 ;
        RECT 1572.840 587.870 1573.100 588.190 ;
        RECT 1604.120 587.870 1604.380 588.190 ;
        RECT 1604.180 15.970 1604.320 587.870 ;
        RECT 1604.120 15.650 1604.380 15.970 ;
        RECT 1751.320 15.650 1751.580 15.970 ;
        RECT 1751.380 2.400 1751.520 15.650 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1582.010 586.740 1582.330 586.800 ;
        RECT 1586.610 586.740 1586.930 586.800 ;
        RECT 1582.010 586.600 1586.930 586.740 ;
        RECT 1582.010 586.540 1582.330 586.600 ;
        RECT 1586.610 586.540 1586.930 586.600 ;
        RECT 1586.610 16.560 1586.930 16.620 ;
        RECT 1768.770 16.560 1769.090 16.620 ;
        RECT 1586.610 16.420 1769.090 16.560 ;
        RECT 1586.610 16.360 1586.930 16.420 ;
        RECT 1768.770 16.360 1769.090 16.420 ;
      LAYER via ;
        RECT 1582.040 586.540 1582.300 586.800 ;
        RECT 1586.640 586.540 1586.900 586.800 ;
        RECT 1586.640 16.360 1586.900 16.620 ;
        RECT 1768.800 16.360 1769.060 16.620 ;
      LAYER met2 ;
        RECT 1580.430 600.170 1580.710 604.000 ;
        RECT 1580.430 600.030 1582.240 600.170 ;
        RECT 1580.430 600.000 1580.710 600.030 ;
        RECT 1582.100 586.830 1582.240 600.030 ;
        RECT 1582.040 586.510 1582.300 586.830 ;
        RECT 1586.640 586.510 1586.900 586.830 ;
        RECT 1586.700 16.650 1586.840 586.510 ;
        RECT 1586.640 16.330 1586.900 16.650 ;
        RECT 1768.800 16.330 1769.060 16.650 ;
        RECT 1768.860 2.400 1769.000 16.330 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1591.210 587.080 1591.530 587.140 ;
        RECT 1610.990 587.080 1611.310 587.140 ;
        RECT 1591.210 586.940 1611.310 587.080 ;
        RECT 1591.210 586.880 1591.530 586.940 ;
        RECT 1610.990 586.880 1611.310 586.940 ;
        RECT 1610.990 16.220 1611.310 16.280 ;
        RECT 1786.710 16.220 1787.030 16.280 ;
        RECT 1610.990 16.080 1787.030 16.220 ;
        RECT 1610.990 16.020 1611.310 16.080 ;
        RECT 1786.710 16.020 1787.030 16.080 ;
      LAYER via ;
        RECT 1591.240 586.880 1591.500 587.140 ;
        RECT 1611.020 586.880 1611.280 587.140 ;
        RECT 1611.020 16.020 1611.280 16.280 ;
        RECT 1786.740 16.020 1787.000 16.280 ;
      LAYER met2 ;
        RECT 1589.630 600.170 1589.910 604.000 ;
        RECT 1589.630 600.030 1591.440 600.170 ;
        RECT 1589.630 600.000 1589.910 600.030 ;
        RECT 1591.300 587.170 1591.440 600.030 ;
        RECT 1591.240 586.850 1591.500 587.170 ;
        RECT 1611.020 586.850 1611.280 587.170 ;
        RECT 1611.080 16.310 1611.220 586.850 ;
        RECT 1611.020 15.990 1611.280 16.310 ;
        RECT 1786.740 15.990 1787.000 16.310 ;
        RECT 1786.800 2.400 1786.940 15.990 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1666.190 590.480 1666.510 590.540 ;
        RECT 1762.790 590.480 1763.110 590.540 ;
        RECT 1666.190 590.340 1763.110 590.480 ;
        RECT 1666.190 590.280 1666.510 590.340 ;
        RECT 1762.790 590.280 1763.110 590.340 ;
        RECT 1600.410 590.140 1600.730 590.200 ;
        RECT 1600.410 590.000 1609.380 590.140 ;
        RECT 1600.410 589.940 1600.730 590.000 ;
        RECT 1609.240 589.800 1609.380 590.000 ;
        RECT 1666.190 589.800 1666.510 589.860 ;
        RECT 1609.240 589.660 1666.510 589.800 ;
        RECT 1666.190 589.600 1666.510 589.660 ;
        RECT 1762.790 587.080 1763.110 587.140 ;
        RECT 1790.390 587.080 1790.710 587.140 ;
        RECT 1762.790 586.940 1790.710 587.080 ;
        RECT 1762.790 586.880 1763.110 586.940 ;
        RECT 1790.390 586.880 1790.710 586.940 ;
        RECT 1790.390 20.640 1790.710 20.700 ;
        RECT 1804.650 20.640 1804.970 20.700 ;
        RECT 1790.390 20.500 1804.970 20.640 ;
        RECT 1790.390 20.440 1790.710 20.500 ;
        RECT 1804.650 20.440 1804.970 20.500 ;
      LAYER via ;
        RECT 1666.220 590.280 1666.480 590.540 ;
        RECT 1762.820 590.280 1763.080 590.540 ;
        RECT 1600.440 589.940 1600.700 590.200 ;
        RECT 1666.220 589.600 1666.480 589.860 ;
        RECT 1762.820 586.880 1763.080 587.140 ;
        RECT 1790.420 586.880 1790.680 587.140 ;
        RECT 1790.420 20.440 1790.680 20.700 ;
        RECT 1804.680 20.440 1804.940 20.700 ;
      LAYER met2 ;
        RECT 1598.830 600.170 1599.110 604.000 ;
        RECT 1598.830 600.030 1600.640 600.170 ;
        RECT 1598.830 600.000 1599.110 600.030 ;
        RECT 1600.500 590.230 1600.640 600.030 ;
        RECT 1666.220 590.250 1666.480 590.570 ;
        RECT 1762.820 590.250 1763.080 590.570 ;
        RECT 1600.440 589.910 1600.700 590.230 ;
        RECT 1666.280 589.890 1666.420 590.250 ;
        RECT 1666.220 589.570 1666.480 589.890 ;
        RECT 1762.880 587.170 1763.020 590.250 ;
        RECT 1762.820 586.850 1763.080 587.170 ;
        RECT 1790.420 586.850 1790.680 587.170 ;
        RECT 1790.480 20.730 1790.620 586.850 ;
        RECT 1790.420 20.410 1790.680 20.730 ;
        RECT 1804.680 20.410 1804.940 20.730 ;
        RECT 1804.740 2.400 1804.880 20.410 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1609.610 590.140 1609.930 590.200 ;
        RECT 1789.930 590.140 1790.250 590.200 ;
        RECT 1609.610 590.000 1790.250 590.140 ;
        RECT 1609.610 589.940 1609.930 590.000 ;
        RECT 1789.930 589.940 1790.250 590.000 ;
        RECT 1789.930 584.700 1790.250 584.760 ;
        RECT 1817.990 584.700 1818.310 584.760 ;
        RECT 1789.930 584.560 1818.310 584.700 ;
        RECT 1789.930 584.500 1790.250 584.560 ;
        RECT 1817.990 584.500 1818.310 584.560 ;
        RECT 1817.990 20.640 1818.310 20.700 ;
        RECT 1822.590 20.640 1822.910 20.700 ;
        RECT 1817.990 20.500 1822.910 20.640 ;
        RECT 1817.990 20.440 1818.310 20.500 ;
        RECT 1822.590 20.440 1822.910 20.500 ;
      LAYER via ;
        RECT 1609.640 589.940 1609.900 590.200 ;
        RECT 1789.960 589.940 1790.220 590.200 ;
        RECT 1789.960 584.500 1790.220 584.760 ;
        RECT 1818.020 584.500 1818.280 584.760 ;
        RECT 1818.020 20.440 1818.280 20.700 ;
        RECT 1822.620 20.440 1822.880 20.700 ;
      LAYER met2 ;
        RECT 1608.030 600.170 1608.310 604.000 ;
        RECT 1608.030 600.030 1609.840 600.170 ;
        RECT 1608.030 600.000 1608.310 600.030 ;
        RECT 1609.700 590.230 1609.840 600.030 ;
        RECT 1609.640 589.910 1609.900 590.230 ;
        RECT 1789.960 589.910 1790.220 590.230 ;
        RECT 1790.020 584.790 1790.160 589.910 ;
        RECT 1789.960 584.470 1790.220 584.790 ;
        RECT 1818.020 584.470 1818.280 584.790 ;
        RECT 1818.080 20.730 1818.220 584.470 ;
        RECT 1818.020 20.410 1818.280 20.730 ;
        RECT 1822.620 20.410 1822.880 20.730 ;
        RECT 1822.680 2.400 1822.820 20.410 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1618.810 586.740 1619.130 586.800 ;
        RECT 1621.110 586.740 1621.430 586.800 ;
        RECT 1618.810 586.600 1621.430 586.740 ;
        RECT 1618.810 586.540 1619.130 586.600 ;
        RECT 1621.110 586.540 1621.430 586.600 ;
        RECT 1770.240 20.500 1777.280 20.640 ;
        RECT 1621.110 20.300 1621.430 20.360 ;
        RECT 1770.240 20.300 1770.380 20.500 ;
        RECT 1621.110 20.160 1770.380 20.300 ;
        RECT 1777.140 20.300 1777.280 20.500 ;
        RECT 1840.070 20.300 1840.390 20.360 ;
        RECT 1777.140 20.160 1840.390 20.300 ;
        RECT 1621.110 20.100 1621.430 20.160 ;
        RECT 1840.070 20.100 1840.390 20.160 ;
      LAYER via ;
        RECT 1618.840 586.540 1619.100 586.800 ;
        RECT 1621.140 586.540 1621.400 586.800 ;
        RECT 1621.140 20.100 1621.400 20.360 ;
        RECT 1840.100 20.100 1840.360 20.360 ;
      LAYER met2 ;
        RECT 1617.230 600.170 1617.510 604.000 ;
        RECT 1617.230 600.030 1619.040 600.170 ;
        RECT 1617.230 600.000 1617.510 600.030 ;
        RECT 1618.900 586.830 1619.040 600.030 ;
        RECT 1618.840 586.510 1619.100 586.830 ;
        RECT 1621.140 586.510 1621.400 586.830 ;
        RECT 1621.200 20.390 1621.340 586.510 ;
        RECT 1621.140 20.070 1621.400 20.390 ;
        RECT 1840.100 20.070 1840.360 20.390 ;
        RECT 1840.160 2.400 1840.300 20.070 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1818.910 590.480 1819.230 590.540 ;
        RECT 1845.590 590.480 1845.910 590.540 ;
        RECT 1818.910 590.340 1845.910 590.480 ;
        RECT 1818.910 590.280 1819.230 590.340 ;
        RECT 1845.590 590.280 1845.910 590.340 ;
        RECT 1787.170 589.800 1787.490 589.860 ;
        RECT 1762.880 589.660 1787.490 589.800 ;
        RECT 1656.990 589.460 1657.310 589.520 ;
        RECT 1752.210 589.460 1752.530 589.520 ;
        RECT 1656.990 589.320 1752.530 589.460 ;
        RECT 1656.990 589.260 1657.310 589.320 ;
        RECT 1752.210 589.260 1752.530 589.320 ;
        RECT 1752.670 589.460 1752.990 589.520 ;
        RECT 1762.880 589.460 1763.020 589.660 ;
        RECT 1787.170 589.600 1787.490 589.660 ;
        RECT 1752.670 589.320 1763.020 589.460 ;
        RECT 1752.670 589.260 1752.990 589.320 ;
        RECT 1627.090 589.120 1627.410 589.180 ;
        RECT 1642.270 589.120 1642.590 589.180 ;
        RECT 1627.090 588.980 1642.590 589.120 ;
        RECT 1627.090 588.920 1627.410 588.980 ;
        RECT 1642.270 588.920 1642.590 588.980 ;
        RECT 1845.590 14.860 1845.910 14.920 ;
        RECT 1858.010 14.860 1858.330 14.920 ;
        RECT 1845.590 14.720 1858.330 14.860 ;
        RECT 1845.590 14.660 1845.910 14.720 ;
        RECT 1858.010 14.660 1858.330 14.720 ;
      LAYER via ;
        RECT 1818.940 590.280 1819.200 590.540 ;
        RECT 1845.620 590.280 1845.880 590.540 ;
        RECT 1657.020 589.260 1657.280 589.520 ;
        RECT 1752.240 589.260 1752.500 589.520 ;
        RECT 1752.700 589.260 1752.960 589.520 ;
        RECT 1787.200 589.600 1787.460 589.860 ;
        RECT 1627.120 588.920 1627.380 589.180 ;
        RECT 1642.300 588.920 1642.560 589.180 ;
        RECT 1845.620 14.660 1845.880 14.920 ;
        RECT 1858.040 14.660 1858.300 14.920 ;
      LAYER met2 ;
        RECT 1626.430 600.170 1626.710 604.000 ;
        RECT 1626.430 600.030 1627.320 600.170 ;
        RECT 1626.430 600.000 1626.710 600.030 ;
        RECT 1627.180 589.210 1627.320 600.030 ;
        RECT 1818.940 590.250 1819.200 590.570 ;
        RECT 1845.620 590.250 1845.880 590.570 ;
        RECT 1819.000 590.085 1819.140 590.250 ;
        RECT 1787.190 589.715 1787.470 590.085 ;
        RECT 1818.930 589.715 1819.210 590.085 ;
        RECT 1787.200 589.570 1787.460 589.715 ;
        RECT 1657.020 589.230 1657.280 589.550 ;
        RECT 1752.240 589.460 1752.500 589.550 ;
        RECT 1752.700 589.460 1752.960 589.550 ;
        RECT 1752.240 589.320 1752.960 589.460 ;
        RECT 1752.240 589.230 1752.500 589.320 ;
        RECT 1752.700 589.230 1752.960 589.320 ;
        RECT 1627.120 588.890 1627.380 589.210 ;
        RECT 1642.300 588.890 1642.560 589.210 ;
        RECT 1642.360 588.725 1642.500 588.890 ;
        RECT 1657.080 588.725 1657.220 589.230 ;
        RECT 1642.290 588.355 1642.570 588.725 ;
        RECT 1657.010 588.355 1657.290 588.725 ;
        RECT 1845.680 14.950 1845.820 590.250 ;
        RECT 1845.620 14.630 1845.880 14.950 ;
        RECT 1858.040 14.630 1858.300 14.950 ;
        RECT 1858.100 2.400 1858.240 14.630 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
      LAYER via2 ;
        RECT 1787.190 589.760 1787.470 590.040 ;
        RECT 1818.930 589.760 1819.210 590.040 ;
        RECT 1642.290 588.400 1642.570 588.680 ;
        RECT 1657.010 588.400 1657.290 588.680 ;
      LAYER met3 ;
        RECT 1787.165 590.050 1787.495 590.065 ;
        RECT 1818.905 590.050 1819.235 590.065 ;
        RECT 1787.165 589.750 1819.235 590.050 ;
        RECT 1787.165 589.735 1787.495 589.750 ;
        RECT 1818.905 589.735 1819.235 589.750 ;
        RECT 1642.265 588.690 1642.595 588.705 ;
        RECT 1656.985 588.690 1657.315 588.705 ;
        RECT 1642.265 588.390 1657.315 588.690 ;
        RECT 1642.265 588.375 1642.595 588.390 ;
        RECT 1656.985 588.375 1657.315 588.390 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1637.210 586.740 1637.530 586.800 ;
        RECT 1641.810 586.740 1642.130 586.800 ;
        RECT 1637.210 586.600 1642.130 586.740 ;
        RECT 1637.210 586.540 1637.530 586.600 ;
        RECT 1641.810 586.540 1642.130 586.600 ;
        RECT 1641.810 19.280 1642.130 19.340 ;
        RECT 1875.950 19.280 1876.270 19.340 ;
        RECT 1641.810 19.140 1876.270 19.280 ;
        RECT 1641.810 19.080 1642.130 19.140 ;
        RECT 1875.950 19.080 1876.270 19.140 ;
      LAYER via ;
        RECT 1637.240 586.540 1637.500 586.800 ;
        RECT 1641.840 586.540 1642.100 586.800 ;
        RECT 1641.840 19.080 1642.100 19.340 ;
        RECT 1875.980 19.080 1876.240 19.340 ;
      LAYER met2 ;
        RECT 1635.630 600.170 1635.910 604.000 ;
        RECT 1635.630 600.030 1637.440 600.170 ;
        RECT 1635.630 600.000 1635.910 600.030 ;
        RECT 1637.300 586.830 1637.440 600.030 ;
        RECT 1637.240 586.510 1637.500 586.830 ;
        RECT 1641.840 586.510 1642.100 586.830 ;
        RECT 1641.900 19.370 1642.040 586.510 ;
        RECT 1641.840 19.050 1642.100 19.370 ;
        RECT 1875.980 19.050 1876.240 19.370 ;
        RECT 1876.040 2.400 1876.180 19.050 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 752.170 27.780 752.490 27.840 ;
        RECT 1056.230 27.780 1056.550 27.840 ;
        RECT 752.170 27.640 1056.550 27.780 ;
        RECT 752.170 27.580 752.490 27.640 ;
        RECT 1056.230 27.580 1056.550 27.640 ;
      LAYER via ;
        RECT 752.200 27.580 752.460 27.840 ;
        RECT 1056.260 27.580 1056.520 27.840 ;
      LAYER met2 ;
        RECT 1056.950 600.170 1057.230 604.000 ;
        RECT 1056.320 600.030 1057.230 600.170 ;
        RECT 1056.320 27.870 1056.460 600.030 ;
        RECT 1056.950 600.000 1057.230 600.030 ;
        RECT 752.200 27.550 752.460 27.870 ;
        RECT 1056.260 27.550 1056.520 27.870 ;
        RECT 752.260 2.400 752.400 27.550 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1644.800 598.980 1645.120 599.040 ;
        RECT 1670.330 598.980 1670.650 599.040 ;
        RECT 1644.800 598.840 1670.650 598.980 ;
        RECT 1644.800 598.780 1645.120 598.840 ;
        RECT 1670.330 598.780 1670.650 598.840 ;
        RECT 1670.330 588.780 1670.650 588.840 ;
        RECT 1670.330 588.640 1763.020 588.780 ;
        RECT 1670.330 588.580 1670.650 588.640 ;
        RECT 1762.880 588.440 1763.020 588.640 ;
        RECT 1790.850 588.440 1791.170 588.500 ;
        RECT 1762.880 588.300 1791.170 588.440 ;
        RECT 1790.850 588.240 1791.170 588.300 ;
        RECT 1790.850 16.560 1791.170 16.620 ;
        RECT 1893.890 16.560 1894.210 16.620 ;
        RECT 1790.850 16.420 1894.210 16.560 ;
        RECT 1790.850 16.360 1791.170 16.420 ;
        RECT 1893.890 16.360 1894.210 16.420 ;
      LAYER via ;
        RECT 1644.830 598.780 1645.090 599.040 ;
        RECT 1670.360 598.780 1670.620 599.040 ;
        RECT 1670.360 588.580 1670.620 588.840 ;
        RECT 1790.880 588.240 1791.140 588.500 ;
        RECT 1790.880 16.360 1791.140 16.620 ;
        RECT 1893.920 16.360 1894.180 16.620 ;
      LAYER met2 ;
        RECT 1644.830 600.000 1645.110 604.000 ;
        RECT 1644.890 599.070 1645.030 600.000 ;
        RECT 1644.830 598.750 1645.090 599.070 ;
        RECT 1670.360 598.750 1670.620 599.070 ;
        RECT 1670.420 588.870 1670.560 598.750 ;
        RECT 1670.360 588.550 1670.620 588.870 ;
        RECT 1790.880 588.210 1791.140 588.530 ;
        RECT 1790.940 16.650 1791.080 588.210 ;
        RECT 1790.880 16.330 1791.140 16.650 ;
        RECT 1893.920 16.330 1894.180 16.650 ;
        RECT 1893.980 2.400 1894.120 16.330 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1680.450 18.600 1680.770 18.660 ;
        RECT 1911.830 18.600 1912.150 18.660 ;
        RECT 1680.450 18.460 1912.150 18.600 ;
        RECT 1680.450 18.400 1680.770 18.460 ;
        RECT 1911.830 18.400 1912.150 18.460 ;
        RECT 1655.610 17.920 1655.930 17.980 ;
        RECT 1656.070 17.920 1656.390 17.980 ;
        RECT 1655.610 17.780 1656.390 17.920 ;
        RECT 1655.610 17.720 1655.930 17.780 ;
        RECT 1656.070 17.720 1656.390 17.780 ;
        RECT 1656.070 15.540 1656.390 15.600 ;
        RECT 1680.450 15.540 1680.770 15.600 ;
        RECT 1656.070 15.400 1680.770 15.540 ;
        RECT 1656.070 15.340 1656.390 15.400 ;
        RECT 1680.450 15.340 1680.770 15.400 ;
      LAYER via ;
        RECT 1680.480 18.400 1680.740 18.660 ;
        RECT 1911.860 18.400 1912.120 18.660 ;
        RECT 1655.640 17.720 1655.900 17.980 ;
        RECT 1656.100 17.720 1656.360 17.980 ;
        RECT 1656.100 15.340 1656.360 15.600 ;
        RECT 1680.480 15.340 1680.740 15.600 ;
      LAYER met2 ;
        RECT 1654.030 600.170 1654.310 604.000 ;
        RECT 1654.030 600.030 1655.840 600.170 ;
        RECT 1654.030 600.000 1654.310 600.030 ;
        RECT 1655.700 18.010 1655.840 600.030 ;
        RECT 1680.480 18.370 1680.740 18.690 ;
        RECT 1911.860 18.370 1912.120 18.690 ;
        RECT 1655.640 17.690 1655.900 18.010 ;
        RECT 1656.100 17.690 1656.360 18.010 ;
        RECT 1656.160 15.630 1656.300 17.690 ;
        RECT 1680.540 15.630 1680.680 18.370 ;
        RECT 1656.100 15.310 1656.360 15.630 ;
        RECT 1680.480 15.310 1680.740 15.630 ;
        RECT 1911.920 2.400 1912.060 18.370 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1664.810 587.080 1665.130 587.140 ;
        RECT 1669.410 587.080 1669.730 587.140 ;
        RECT 1664.810 586.940 1669.730 587.080 ;
        RECT 1664.810 586.880 1665.130 586.940 ;
        RECT 1669.410 586.880 1669.730 586.940 ;
        RECT 1929.310 18.940 1929.630 19.000 ;
        RECT 1680.080 18.800 1929.630 18.940 ;
        RECT 1669.410 18.600 1669.730 18.660 ;
        RECT 1680.080 18.600 1680.220 18.800 ;
        RECT 1929.310 18.740 1929.630 18.800 ;
        RECT 1669.410 18.460 1680.220 18.600 ;
        RECT 1669.410 18.400 1669.730 18.460 ;
      LAYER via ;
        RECT 1664.840 586.880 1665.100 587.140 ;
        RECT 1669.440 586.880 1669.700 587.140 ;
        RECT 1669.440 18.400 1669.700 18.660 ;
        RECT 1929.340 18.740 1929.600 19.000 ;
      LAYER met2 ;
        RECT 1663.230 600.170 1663.510 604.000 ;
        RECT 1663.230 600.030 1665.040 600.170 ;
        RECT 1663.230 600.000 1663.510 600.030 ;
        RECT 1664.900 587.170 1665.040 600.030 ;
        RECT 1664.840 586.850 1665.100 587.170 ;
        RECT 1669.440 586.850 1669.700 587.170 ;
        RECT 1669.500 18.690 1669.640 586.850 ;
        RECT 1929.340 18.710 1929.600 19.030 ;
        RECT 1669.440 18.370 1669.700 18.690 ;
        RECT 1929.400 2.400 1929.540 18.710 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1674.010 586.740 1674.330 586.800 ;
        RECT 1676.310 586.740 1676.630 586.800 ;
        RECT 1674.010 586.600 1676.630 586.740 ;
        RECT 1674.010 586.540 1674.330 586.600 ;
        RECT 1676.310 586.540 1676.630 586.600 ;
        RECT 1676.310 18.260 1676.630 18.320 ;
        RECT 1947.250 18.260 1947.570 18.320 ;
        RECT 1676.310 18.120 1947.570 18.260 ;
        RECT 1676.310 18.060 1676.630 18.120 ;
        RECT 1947.250 18.060 1947.570 18.120 ;
      LAYER via ;
        RECT 1674.040 586.540 1674.300 586.800 ;
        RECT 1676.340 586.540 1676.600 586.800 ;
        RECT 1676.340 18.060 1676.600 18.320 ;
        RECT 1947.280 18.060 1947.540 18.320 ;
      LAYER met2 ;
        RECT 1672.430 600.170 1672.710 604.000 ;
        RECT 1672.430 600.030 1674.240 600.170 ;
        RECT 1672.430 600.000 1672.710 600.030 ;
        RECT 1674.100 586.830 1674.240 600.030 ;
        RECT 1674.040 586.510 1674.300 586.830 ;
        RECT 1676.340 586.510 1676.600 586.830 ;
        RECT 1676.400 18.350 1676.540 586.510 ;
        RECT 1676.340 18.030 1676.600 18.350 ;
        RECT 1947.280 18.030 1947.540 18.350 ;
        RECT 1947.340 2.400 1947.480 18.030 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.210 591.500 1683.530 591.560 ;
        RECT 1873.190 591.500 1873.510 591.560 ;
        RECT 1683.210 591.360 1873.510 591.500 ;
        RECT 1683.210 591.300 1683.530 591.360 ;
        RECT 1873.190 591.300 1873.510 591.360 ;
        RECT 1873.190 19.620 1873.510 19.680 ;
        RECT 1873.190 19.480 1877.100 19.620 ;
        RECT 1873.190 19.420 1873.510 19.480 ;
        RECT 1876.960 19.280 1877.100 19.480 ;
        RECT 1965.190 19.280 1965.510 19.340 ;
        RECT 1876.960 19.140 1965.510 19.280 ;
        RECT 1965.190 19.080 1965.510 19.140 ;
      LAYER via ;
        RECT 1683.240 591.300 1683.500 591.560 ;
        RECT 1873.220 591.300 1873.480 591.560 ;
        RECT 1873.220 19.420 1873.480 19.680 ;
        RECT 1965.220 19.080 1965.480 19.340 ;
      LAYER met2 ;
        RECT 1681.630 600.170 1681.910 604.000 ;
        RECT 1681.630 600.030 1683.440 600.170 ;
        RECT 1681.630 600.000 1681.910 600.030 ;
        RECT 1683.300 591.590 1683.440 600.030 ;
        RECT 1683.240 591.270 1683.500 591.590 ;
        RECT 1873.220 591.270 1873.480 591.590 ;
        RECT 1873.280 19.710 1873.420 591.270 ;
        RECT 1873.220 19.390 1873.480 19.710 ;
        RECT 1965.220 19.050 1965.480 19.370 ;
        RECT 1965.280 2.400 1965.420 19.050 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1692.410 591.160 1692.730 591.220 ;
        RECT 1921.030 591.160 1921.350 591.220 ;
        RECT 1692.410 591.020 1921.350 591.160 ;
        RECT 1692.410 590.960 1692.730 591.020 ;
        RECT 1921.030 590.960 1921.350 591.020 ;
        RECT 1921.490 18.600 1921.810 18.660 ;
        RECT 1983.130 18.600 1983.450 18.660 ;
        RECT 1921.490 18.460 1983.450 18.600 ;
        RECT 1921.490 18.400 1921.810 18.460 ;
        RECT 1983.130 18.400 1983.450 18.460 ;
      LAYER via ;
        RECT 1692.440 590.960 1692.700 591.220 ;
        RECT 1921.060 590.960 1921.320 591.220 ;
        RECT 1921.520 18.400 1921.780 18.660 ;
        RECT 1983.160 18.400 1983.420 18.660 ;
      LAYER met2 ;
        RECT 1690.830 600.170 1691.110 604.000 ;
        RECT 1690.830 600.030 1692.640 600.170 ;
        RECT 1690.830 600.000 1691.110 600.030 ;
        RECT 1692.500 591.250 1692.640 600.030 ;
        RECT 1692.440 590.930 1692.700 591.250 ;
        RECT 1921.060 590.930 1921.320 591.250 ;
        RECT 1921.120 589.290 1921.260 590.930 ;
        RECT 1921.120 589.150 1921.720 589.290 ;
        RECT 1921.580 18.690 1921.720 589.150 ;
        RECT 1921.520 18.370 1921.780 18.690 ;
        RECT 1983.160 18.370 1983.420 18.690 ;
        RECT 1983.220 2.400 1983.360 18.370 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1701.610 586.740 1701.930 586.800 ;
        RECT 1703.910 586.740 1704.230 586.800 ;
        RECT 1701.610 586.600 1704.230 586.740 ;
        RECT 1701.610 586.540 1701.930 586.600 ;
        RECT 1703.910 586.540 1704.230 586.600 ;
        RECT 1703.910 14.180 1704.230 14.240 ;
        RECT 2001.070 14.180 2001.390 14.240 ;
        RECT 1703.910 14.040 2001.390 14.180 ;
        RECT 1703.910 13.980 1704.230 14.040 ;
        RECT 2001.070 13.980 2001.390 14.040 ;
      LAYER via ;
        RECT 1701.640 586.540 1701.900 586.800 ;
        RECT 1703.940 586.540 1704.200 586.800 ;
        RECT 1703.940 13.980 1704.200 14.240 ;
        RECT 2001.100 13.980 2001.360 14.240 ;
      LAYER met2 ;
        RECT 1700.030 600.170 1700.310 604.000 ;
        RECT 1700.030 600.030 1701.840 600.170 ;
        RECT 1700.030 600.000 1700.310 600.030 ;
        RECT 1701.700 586.830 1701.840 600.030 ;
        RECT 1701.640 586.510 1701.900 586.830 ;
        RECT 1703.940 586.510 1704.200 586.830 ;
        RECT 1704.000 14.270 1704.140 586.510 ;
        RECT 1703.940 13.950 1704.200 14.270 ;
        RECT 2001.100 13.950 2001.360 14.270 ;
        RECT 2001.160 2.400 2001.300 13.950 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 592.180 1711.130 592.240 ;
        RECT 1949.090 592.180 1949.410 592.240 ;
        RECT 1710.810 592.040 1949.410 592.180 ;
        RECT 1710.810 591.980 1711.130 592.040 ;
        RECT 1949.090 591.980 1949.410 592.040 ;
        RECT 1949.090 18.940 1949.410 19.000 ;
        RECT 2018.550 18.940 2018.870 19.000 ;
        RECT 1949.090 18.800 2018.870 18.940 ;
        RECT 1949.090 18.740 1949.410 18.800 ;
        RECT 2018.550 18.740 2018.870 18.800 ;
      LAYER via ;
        RECT 1710.840 591.980 1711.100 592.240 ;
        RECT 1949.120 591.980 1949.380 592.240 ;
        RECT 1949.120 18.740 1949.380 19.000 ;
        RECT 2018.580 18.740 2018.840 19.000 ;
      LAYER met2 ;
        RECT 1709.230 600.170 1709.510 604.000 ;
        RECT 1709.230 600.030 1711.040 600.170 ;
        RECT 1709.230 600.000 1709.510 600.030 ;
        RECT 1710.900 592.270 1711.040 600.030 ;
        RECT 1710.840 591.950 1711.100 592.270 ;
        RECT 1949.120 591.950 1949.380 592.270 ;
        RECT 1949.180 19.030 1949.320 591.950 ;
        RECT 1949.120 18.710 1949.380 19.030 ;
        RECT 2018.580 18.710 2018.840 19.030 ;
        RECT 2018.640 2.400 2018.780 18.710 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1720.010 589.120 1720.330 589.180 ;
        RECT 1724.610 589.120 1724.930 589.180 ;
        RECT 1720.010 588.980 1724.930 589.120 ;
        RECT 1720.010 588.920 1720.330 588.980 ;
        RECT 1724.610 588.920 1724.930 588.980 ;
        RECT 1724.610 17.580 1724.930 17.640 ;
        RECT 2036.490 17.580 2036.810 17.640 ;
        RECT 1724.610 17.440 2036.810 17.580 ;
        RECT 1724.610 17.380 1724.930 17.440 ;
        RECT 2036.490 17.380 2036.810 17.440 ;
      LAYER via ;
        RECT 1720.040 588.920 1720.300 589.180 ;
        RECT 1724.640 588.920 1724.900 589.180 ;
        RECT 1724.640 17.380 1724.900 17.640 ;
        RECT 2036.520 17.380 2036.780 17.640 ;
      LAYER met2 ;
        RECT 1718.430 600.170 1718.710 604.000 ;
        RECT 1718.430 600.030 1720.240 600.170 ;
        RECT 1718.430 600.000 1718.710 600.030 ;
        RECT 1720.100 589.210 1720.240 600.030 ;
        RECT 1720.040 588.890 1720.300 589.210 ;
        RECT 1724.640 588.890 1724.900 589.210 ;
        RECT 1724.700 17.670 1724.840 588.890 ;
        RECT 1724.640 17.350 1724.900 17.670 ;
        RECT 2036.520 17.350 2036.780 17.670 ;
        RECT 2036.580 2.400 2036.720 17.350 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1729.210 589.120 1729.530 589.180 ;
        RECT 1983.590 589.120 1983.910 589.180 ;
        RECT 1729.210 588.980 1983.910 589.120 ;
        RECT 1729.210 588.920 1729.530 588.980 ;
        RECT 1983.590 588.920 1983.910 588.980 ;
        RECT 1983.590 18.600 1983.910 18.660 ;
        RECT 2054.430 18.600 2054.750 18.660 ;
        RECT 1983.590 18.460 2054.750 18.600 ;
        RECT 1983.590 18.400 1983.910 18.460 ;
        RECT 2054.430 18.400 2054.750 18.460 ;
      LAYER via ;
        RECT 1729.240 588.920 1729.500 589.180 ;
        RECT 1983.620 588.920 1983.880 589.180 ;
        RECT 1983.620 18.400 1983.880 18.660 ;
        RECT 2054.460 18.400 2054.720 18.660 ;
      LAYER met2 ;
        RECT 1727.630 600.170 1727.910 604.000 ;
        RECT 1727.630 600.030 1729.440 600.170 ;
        RECT 1727.630 600.000 1727.910 600.030 ;
        RECT 1729.300 589.210 1729.440 600.030 ;
        RECT 1729.240 588.890 1729.500 589.210 ;
        RECT 1983.620 588.890 1983.880 589.210 ;
        RECT 1983.680 18.690 1983.820 588.890 ;
        RECT 1983.620 18.370 1983.880 18.690 ;
        RECT 2054.460 18.370 2054.720 18.690 ;
        RECT 2054.520 2.400 2054.660 18.370 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 858.890 586.740 859.210 586.800 ;
        RECT 1064.510 586.740 1064.830 586.800 ;
        RECT 858.890 586.600 1064.830 586.740 ;
        RECT 858.890 586.540 859.210 586.600 ;
        RECT 1064.510 586.540 1064.830 586.600 ;
        RECT 769.650 19.280 769.970 19.340 ;
        RECT 857.510 19.280 857.830 19.340 ;
        RECT 769.650 19.140 857.830 19.280 ;
        RECT 769.650 19.080 769.970 19.140 ;
        RECT 857.510 19.080 857.830 19.140 ;
      LAYER via ;
        RECT 858.920 586.540 859.180 586.800 ;
        RECT 1064.540 586.540 1064.800 586.800 ;
        RECT 769.680 19.080 769.940 19.340 ;
        RECT 857.540 19.080 857.800 19.340 ;
      LAYER met2 ;
        RECT 1066.150 600.170 1066.430 604.000 ;
        RECT 1064.600 600.030 1066.430 600.170 ;
        RECT 1064.600 586.830 1064.740 600.030 ;
        RECT 1066.150 600.000 1066.430 600.030 ;
        RECT 858.920 586.510 859.180 586.830 ;
        RECT 1064.540 586.510 1064.800 586.830 ;
        RECT 858.980 28.290 859.120 586.510 ;
        RECT 857.600 28.150 859.120 28.290 ;
        RECT 857.600 19.370 857.740 28.150 ;
        RECT 769.680 19.050 769.940 19.370 ;
        RECT 857.540 19.050 857.800 19.370 ;
        RECT 769.740 2.400 769.880 19.050 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1737.950 592.520 1738.270 592.580 ;
        RECT 1880.090 592.520 1880.410 592.580 ;
        RECT 1737.950 592.380 1880.410 592.520 ;
        RECT 1737.950 592.320 1738.270 592.380 ;
        RECT 1880.090 592.320 1880.410 592.380 ;
        RECT 1880.090 14.860 1880.410 14.920 ;
        RECT 2072.370 14.860 2072.690 14.920 ;
        RECT 1880.090 14.720 2072.690 14.860 ;
        RECT 1880.090 14.660 1880.410 14.720 ;
        RECT 2072.370 14.660 2072.690 14.720 ;
      LAYER via ;
        RECT 1737.980 592.320 1738.240 592.580 ;
        RECT 1880.120 592.320 1880.380 592.580 ;
        RECT 1880.120 14.660 1880.380 14.920 ;
        RECT 2072.400 14.660 2072.660 14.920 ;
      LAYER met2 ;
        RECT 1736.370 600.170 1736.650 604.000 ;
        RECT 1736.370 600.030 1738.180 600.170 ;
        RECT 1736.370 600.000 1736.650 600.030 ;
        RECT 1738.040 592.610 1738.180 600.030 ;
        RECT 1737.980 592.290 1738.240 592.610 ;
        RECT 1880.120 592.290 1880.380 592.610 ;
        RECT 1880.180 14.950 1880.320 592.290 ;
        RECT 1880.120 14.630 1880.380 14.950 ;
        RECT 2072.400 14.630 2072.660 14.950 ;
        RECT 2072.460 2.400 2072.600 14.630 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.710 589.460 1787.030 589.520 ;
        RECT 2083.870 589.460 2084.190 589.520 ;
        RECT 1786.710 589.320 2084.190 589.460 ;
        RECT 1786.710 589.260 1787.030 589.320 ;
        RECT 2083.870 589.260 2084.190 589.320 ;
        RECT 2083.870 37.980 2084.190 38.040 ;
        RECT 2089.850 37.980 2090.170 38.040 ;
        RECT 2083.870 37.840 2090.170 37.980 ;
        RECT 2083.870 37.780 2084.190 37.840 ;
        RECT 2089.850 37.780 2090.170 37.840 ;
      LAYER via ;
        RECT 1786.740 589.260 1787.000 589.520 ;
        RECT 2083.900 589.260 2084.160 589.520 ;
        RECT 2083.900 37.780 2084.160 38.040 ;
        RECT 2089.880 37.780 2090.140 38.040 ;
      LAYER met2 ;
        RECT 1745.570 600.170 1745.850 604.000 ;
        RECT 1745.570 600.030 1747.380 600.170 ;
        RECT 1745.570 600.000 1745.850 600.030 ;
        RECT 1747.240 589.405 1747.380 600.030 ;
        RECT 1786.740 589.405 1787.000 589.550 ;
        RECT 1747.170 589.035 1747.450 589.405 ;
        RECT 1786.730 589.035 1787.010 589.405 ;
        RECT 2083.900 589.230 2084.160 589.550 ;
        RECT 2083.960 38.070 2084.100 589.230 ;
        RECT 2083.900 37.750 2084.160 38.070 ;
        RECT 2089.880 37.750 2090.140 38.070 ;
        RECT 2089.940 2.400 2090.080 37.750 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
      LAYER via2 ;
        RECT 1747.170 589.080 1747.450 589.360 ;
        RECT 1786.730 589.080 1787.010 589.360 ;
      LAYER met3 ;
        RECT 1747.145 589.370 1747.475 589.385 ;
        RECT 1786.705 589.370 1787.035 589.385 ;
        RECT 1747.145 589.070 1787.035 589.370 ;
        RECT 1747.145 589.055 1747.475 589.070 ;
        RECT 1786.705 589.055 1787.035 589.070 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1756.350 586.740 1756.670 586.800 ;
        RECT 1759.110 586.740 1759.430 586.800 ;
        RECT 1756.350 586.600 1759.430 586.740 ;
        RECT 1756.350 586.540 1756.670 586.600 ;
        RECT 1759.110 586.540 1759.430 586.600 ;
        RECT 2107.790 17.580 2108.110 17.640 ;
        RECT 2091.320 17.440 2108.110 17.580 ;
        RECT 1759.110 17.240 1759.430 17.300 ;
        RECT 2091.320 17.240 2091.460 17.440 ;
        RECT 2107.790 17.380 2108.110 17.440 ;
        RECT 1759.110 17.100 2091.460 17.240 ;
        RECT 1759.110 17.040 1759.430 17.100 ;
      LAYER via ;
        RECT 1756.380 586.540 1756.640 586.800 ;
        RECT 1759.140 586.540 1759.400 586.800 ;
        RECT 1759.140 17.040 1759.400 17.300 ;
        RECT 2107.820 17.380 2108.080 17.640 ;
      LAYER met2 ;
        RECT 1754.770 600.170 1755.050 604.000 ;
        RECT 1754.770 600.030 1756.580 600.170 ;
        RECT 1754.770 600.000 1755.050 600.030 ;
        RECT 1756.440 586.830 1756.580 600.030 ;
        RECT 1756.380 586.510 1756.640 586.830 ;
        RECT 1759.140 586.510 1759.400 586.830 ;
        RECT 1759.200 17.330 1759.340 586.510 ;
        RECT 2107.820 17.350 2108.080 17.670 ;
        RECT 1759.140 17.010 1759.400 17.330 ;
        RECT 2107.880 2.400 2108.020 17.350 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1765.550 593.200 1765.870 593.260 ;
        RECT 2126.650 593.200 2126.970 593.260 ;
        RECT 1765.550 593.060 2126.970 593.200 ;
        RECT 1765.550 593.000 1765.870 593.060 ;
        RECT 2126.650 593.000 2126.970 593.060 ;
        RECT 2125.730 2.960 2126.050 3.020 ;
        RECT 2126.650 2.960 2126.970 3.020 ;
        RECT 2125.730 2.820 2126.970 2.960 ;
        RECT 2125.730 2.760 2126.050 2.820 ;
        RECT 2126.650 2.760 2126.970 2.820 ;
      LAYER via ;
        RECT 1765.580 593.000 1765.840 593.260 ;
        RECT 2126.680 593.000 2126.940 593.260 ;
        RECT 2125.760 2.760 2126.020 3.020 ;
        RECT 2126.680 2.760 2126.940 3.020 ;
      LAYER met2 ;
        RECT 1763.970 600.170 1764.250 604.000 ;
        RECT 1763.970 600.030 1765.780 600.170 ;
        RECT 1763.970 600.000 1764.250 600.030 ;
        RECT 1765.640 593.290 1765.780 600.030 ;
        RECT 1765.580 592.970 1765.840 593.290 ;
        RECT 2126.680 592.970 2126.940 593.290 ;
        RECT 2126.740 3.050 2126.880 592.970 ;
        RECT 2125.760 2.730 2126.020 3.050 ;
        RECT 2126.680 2.730 2126.940 3.050 ;
        RECT 2125.820 2.400 2125.960 2.730 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1774.750 588.100 1775.070 588.160 ;
        RECT 1774.750 587.960 1793.840 588.100 ;
        RECT 1774.750 587.900 1775.070 587.960 ;
        RECT 1793.700 587.760 1793.840 587.960 ;
        RECT 1846.050 587.760 1846.370 587.820 ;
        RECT 1793.700 587.620 1846.370 587.760 ;
        RECT 1846.050 587.560 1846.370 587.620 ;
        RECT 1846.970 14.520 1847.290 14.580 ;
        RECT 2143.670 14.520 2143.990 14.580 ;
        RECT 1846.970 14.380 2143.990 14.520 ;
        RECT 1846.970 14.320 1847.290 14.380 ;
        RECT 2143.670 14.320 2143.990 14.380 ;
      LAYER via ;
        RECT 1774.780 587.900 1775.040 588.160 ;
        RECT 1846.080 587.560 1846.340 587.820 ;
        RECT 1847.000 14.320 1847.260 14.580 ;
        RECT 2143.700 14.320 2143.960 14.580 ;
      LAYER met2 ;
        RECT 1773.170 600.170 1773.450 604.000 ;
        RECT 1773.170 600.030 1774.980 600.170 ;
        RECT 1773.170 600.000 1773.450 600.030 ;
        RECT 1774.840 588.190 1774.980 600.030 ;
        RECT 1774.780 587.870 1775.040 588.190 ;
        RECT 1846.080 587.530 1846.340 587.850 ;
        RECT 1846.140 24.210 1846.280 587.530 ;
        RECT 1846.140 24.070 1847.200 24.210 ;
        RECT 1847.060 14.610 1847.200 24.070 ;
        RECT 1847.000 14.290 1847.260 14.610 ;
        RECT 2143.700 14.290 2143.960 14.610 ;
        RECT 2143.760 2.400 2143.900 14.290 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1846.600 587.620 1921.720 587.760 ;
        RECT 1783.950 587.420 1784.270 587.480 ;
        RECT 1846.600 587.420 1846.740 587.620 ;
        RECT 1783.950 587.280 1846.740 587.420 ;
        RECT 1921.580 587.420 1921.720 587.620 ;
        RECT 1969.790 587.420 1970.110 587.480 ;
        RECT 1921.580 587.280 1970.110 587.420 ;
        RECT 1783.950 587.220 1784.270 587.280 ;
        RECT 1969.790 587.220 1970.110 587.280 ;
        RECT 1994.170 19.280 1994.490 19.340 ;
        RECT 1994.170 19.140 2019.240 19.280 ;
        RECT 1994.170 19.080 1994.490 19.140 ;
        RECT 2019.100 18.940 2019.240 19.140 ;
        RECT 2036.950 18.940 2037.270 19.000 ;
        RECT 2019.100 18.800 2037.270 18.940 ;
        RECT 2036.950 18.740 2037.270 18.800 ;
        RECT 1969.790 18.260 1970.110 18.320 ;
        RECT 1994.170 18.260 1994.490 18.320 ;
        RECT 1969.790 18.120 1994.490 18.260 ;
        RECT 1969.790 18.060 1970.110 18.120 ;
        RECT 1994.170 18.060 1994.490 18.120 ;
        RECT 2036.950 17.580 2037.270 17.640 ;
        RECT 2089.390 17.580 2089.710 17.640 ;
        RECT 2161.610 17.580 2161.930 17.640 ;
        RECT 2036.950 17.440 2089.710 17.580 ;
        RECT 2036.950 17.380 2037.270 17.440 ;
        RECT 2089.390 17.380 2089.710 17.440 ;
        RECT 2139.160 17.440 2161.930 17.580 ;
        RECT 2091.690 17.240 2092.010 17.300 ;
        RECT 2139.160 17.240 2139.300 17.440 ;
        RECT 2161.610 17.380 2161.930 17.440 ;
        RECT 2091.690 17.100 2139.300 17.240 ;
        RECT 2091.690 17.040 2092.010 17.100 ;
      LAYER via ;
        RECT 1783.980 587.220 1784.240 587.480 ;
        RECT 1969.820 587.220 1970.080 587.480 ;
        RECT 1994.200 19.080 1994.460 19.340 ;
        RECT 2036.980 18.740 2037.240 19.000 ;
        RECT 1969.820 18.060 1970.080 18.320 ;
        RECT 1994.200 18.060 1994.460 18.320 ;
        RECT 2036.980 17.380 2037.240 17.640 ;
        RECT 2089.420 17.380 2089.680 17.640 ;
        RECT 2091.720 17.040 2091.980 17.300 ;
        RECT 2161.640 17.380 2161.900 17.640 ;
      LAYER met2 ;
        RECT 1782.370 600.170 1782.650 604.000 ;
        RECT 1782.370 600.030 1784.180 600.170 ;
        RECT 1782.370 600.000 1782.650 600.030 ;
        RECT 1784.040 587.510 1784.180 600.030 ;
        RECT 1783.980 587.190 1784.240 587.510 ;
        RECT 1969.820 587.190 1970.080 587.510 ;
        RECT 1969.880 18.350 1970.020 587.190 ;
        RECT 1994.200 19.050 1994.460 19.370 ;
        RECT 1994.260 18.350 1994.400 19.050 ;
        RECT 2036.980 18.710 2037.240 19.030 ;
        RECT 1969.820 18.030 1970.080 18.350 ;
        RECT 1994.200 18.030 1994.460 18.350 ;
        RECT 2037.040 17.670 2037.180 18.710 ;
        RECT 2089.410 17.835 2089.690 18.205 ;
        RECT 2091.710 17.835 2091.990 18.205 ;
        RECT 2089.480 17.670 2089.620 17.835 ;
        RECT 2036.980 17.350 2037.240 17.670 ;
        RECT 2089.420 17.350 2089.680 17.670 ;
        RECT 2091.780 17.330 2091.920 17.835 ;
        RECT 2161.640 17.350 2161.900 17.670 ;
        RECT 2091.720 17.010 2091.980 17.330 ;
        RECT 2161.700 2.400 2161.840 17.350 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
      LAYER via2 ;
        RECT 2089.410 17.880 2089.690 18.160 ;
        RECT 2091.710 17.880 2091.990 18.160 ;
      LAYER met3 ;
        RECT 2089.385 18.170 2089.715 18.185 ;
        RECT 2091.685 18.170 2092.015 18.185 ;
        RECT 2089.385 17.870 2092.015 18.170 ;
        RECT 2089.385 17.855 2089.715 17.870 ;
        RECT 2091.685 17.855 2092.015 17.870 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 35.600 1793.930 35.660 ;
        RECT 2179.090 35.600 2179.410 35.660 ;
        RECT 1793.610 35.460 2179.410 35.600 ;
        RECT 1793.610 35.400 1793.930 35.460 ;
        RECT 2179.090 35.400 2179.410 35.460 ;
      LAYER via ;
        RECT 1793.640 35.400 1793.900 35.660 ;
        RECT 2179.120 35.400 2179.380 35.660 ;
      LAYER met2 ;
        RECT 1791.570 600.170 1791.850 604.000 ;
        RECT 1791.570 600.030 1793.840 600.170 ;
        RECT 1791.570 600.000 1791.850 600.030 ;
        RECT 1793.700 35.690 1793.840 600.030 ;
        RECT 1793.640 35.370 1793.900 35.690 ;
        RECT 2179.120 35.370 2179.380 35.690 ;
        RECT 2179.180 2.400 2179.320 35.370 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1802.350 588.440 1802.670 588.500 ;
        RECT 1990.490 588.440 1990.810 588.500 ;
        RECT 1802.350 588.300 1990.810 588.440 ;
        RECT 1802.350 588.240 1802.670 588.300 ;
        RECT 1990.490 588.240 1990.810 588.300 ;
        RECT 1990.490 17.920 1990.810 17.980 ;
        RECT 2041.550 17.920 2041.870 17.980 ;
        RECT 1990.490 17.780 2041.870 17.920 ;
        RECT 1990.490 17.720 1990.810 17.780 ;
        RECT 2041.550 17.720 2041.870 17.780 ;
        RECT 2042.470 17.920 2042.790 17.980 ;
        RECT 2042.470 17.780 2114.920 17.920 ;
        RECT 2042.470 17.720 2042.790 17.780 ;
        RECT 2114.780 17.580 2114.920 17.780 ;
        RECT 2138.610 17.580 2138.930 17.640 ;
        RECT 2114.780 17.440 2138.930 17.580 ;
        RECT 2138.610 17.380 2138.930 17.440 ;
        RECT 2139.530 17.240 2139.850 17.300 ;
        RECT 2197.030 17.240 2197.350 17.300 ;
        RECT 2139.530 17.100 2197.350 17.240 ;
        RECT 2139.530 17.040 2139.850 17.100 ;
        RECT 2197.030 17.040 2197.350 17.100 ;
      LAYER via ;
        RECT 1802.380 588.240 1802.640 588.500 ;
        RECT 1990.520 588.240 1990.780 588.500 ;
        RECT 1990.520 17.720 1990.780 17.980 ;
        RECT 2041.580 17.720 2041.840 17.980 ;
        RECT 2042.500 17.720 2042.760 17.980 ;
        RECT 2138.640 17.380 2138.900 17.640 ;
        RECT 2139.560 17.040 2139.820 17.300 ;
        RECT 2197.060 17.040 2197.320 17.300 ;
      LAYER met2 ;
        RECT 1800.770 600.170 1801.050 604.000 ;
        RECT 1800.770 600.030 1802.580 600.170 ;
        RECT 1800.770 600.000 1801.050 600.030 ;
        RECT 1802.440 588.530 1802.580 600.030 ;
        RECT 1802.380 588.210 1802.640 588.530 ;
        RECT 1990.520 588.210 1990.780 588.530 ;
        RECT 1990.580 18.010 1990.720 588.210 ;
        RECT 1990.520 17.690 1990.780 18.010 ;
        RECT 2041.570 17.835 2041.850 18.205 ;
        RECT 2042.490 17.835 2042.770 18.205 ;
        RECT 2041.580 17.690 2041.840 17.835 ;
        RECT 2042.500 17.690 2042.760 17.835 ;
        RECT 2138.640 17.525 2138.900 17.670 ;
        RECT 2138.630 17.155 2138.910 17.525 ;
        RECT 2139.550 17.155 2139.830 17.525 ;
        RECT 2139.560 17.010 2139.820 17.155 ;
        RECT 2197.060 17.010 2197.320 17.330 ;
        RECT 2197.120 2.400 2197.260 17.010 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
      LAYER via2 ;
        RECT 2041.570 17.880 2041.850 18.160 ;
        RECT 2042.490 17.880 2042.770 18.160 ;
        RECT 2138.630 17.200 2138.910 17.480 ;
        RECT 2139.550 17.200 2139.830 17.480 ;
      LAYER met3 ;
        RECT 2041.545 18.170 2041.875 18.185 ;
        RECT 2042.465 18.170 2042.795 18.185 ;
        RECT 2041.545 17.870 2042.795 18.170 ;
        RECT 2041.545 17.855 2041.875 17.870 ;
        RECT 2042.465 17.855 2042.795 17.870 ;
        RECT 2138.605 17.490 2138.935 17.505 ;
        RECT 2139.525 17.490 2139.855 17.505 ;
        RECT 2138.605 17.190 2139.855 17.490 ;
        RECT 2138.605 17.175 2138.935 17.190 ;
        RECT 2139.525 17.175 2139.855 17.190 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1811.550 592.860 1811.870 592.920 ;
        RECT 2214.970 592.860 2215.290 592.920 ;
        RECT 1811.550 592.720 2215.290 592.860 ;
        RECT 1811.550 592.660 1811.870 592.720 ;
        RECT 2214.970 592.660 2215.290 592.720 ;
      LAYER via ;
        RECT 1811.580 592.660 1811.840 592.920 ;
        RECT 2215.000 592.660 2215.260 592.920 ;
      LAYER met2 ;
        RECT 1809.970 600.170 1810.250 604.000 ;
        RECT 1809.970 600.030 1811.780 600.170 ;
        RECT 1809.970 600.000 1810.250 600.030 ;
        RECT 1811.640 592.950 1811.780 600.030 ;
        RECT 1811.580 592.630 1811.840 592.950 ;
        RECT 2215.000 592.630 2215.260 592.950 ;
        RECT 2215.060 2.400 2215.200 592.630 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1820.290 588.780 1820.610 588.840 ;
        RECT 1941.730 588.780 1942.050 588.840 ;
        RECT 1820.290 588.640 1942.050 588.780 ;
        RECT 1820.290 588.580 1820.610 588.640 ;
        RECT 1941.730 588.580 1942.050 588.640 ;
        RECT 1941.730 587.080 1942.050 587.140 ;
        RECT 1980.370 587.080 1980.690 587.140 ;
        RECT 1941.730 586.940 1980.690 587.080 ;
        RECT 1941.730 586.880 1942.050 586.940 ;
        RECT 1980.370 586.880 1980.690 586.940 ;
        RECT 1980.370 584.700 1980.690 584.760 ;
        RECT 2011.190 584.700 2011.510 584.760 ;
        RECT 1980.370 584.560 2011.510 584.700 ;
        RECT 1980.370 584.500 1980.690 584.560 ;
        RECT 2011.190 584.500 2011.510 584.560 ;
        RECT 2185.990 14.860 2186.310 14.920 ;
        RECT 2163.080 14.720 2186.310 14.860 ;
        RECT 2011.190 14.180 2011.510 14.240 ;
        RECT 2163.080 14.180 2163.220 14.720 ;
        RECT 2185.990 14.660 2186.310 14.720 ;
        RECT 2232.910 14.180 2233.230 14.240 ;
        RECT 2011.190 14.040 2163.220 14.180 ;
        RECT 2221.500 14.040 2233.230 14.180 ;
        RECT 2011.190 13.980 2011.510 14.040 ;
        RECT 2185.990 13.840 2186.310 13.900 ;
        RECT 2221.500 13.840 2221.640 14.040 ;
        RECT 2232.910 13.980 2233.230 14.040 ;
        RECT 2185.990 13.700 2221.640 13.840 ;
        RECT 2185.990 13.640 2186.310 13.700 ;
      LAYER via ;
        RECT 1820.320 588.580 1820.580 588.840 ;
        RECT 1941.760 588.580 1942.020 588.840 ;
        RECT 1941.760 586.880 1942.020 587.140 ;
        RECT 1980.400 586.880 1980.660 587.140 ;
        RECT 1980.400 584.500 1980.660 584.760 ;
        RECT 2011.220 584.500 2011.480 584.760 ;
        RECT 2011.220 13.980 2011.480 14.240 ;
        RECT 2186.020 14.660 2186.280 14.920 ;
        RECT 2186.020 13.640 2186.280 13.900 ;
        RECT 2232.940 13.980 2233.200 14.240 ;
      LAYER met2 ;
        RECT 1819.170 600.170 1819.450 604.000 ;
        RECT 1819.170 600.030 1820.520 600.170 ;
        RECT 1819.170 600.000 1819.450 600.030 ;
        RECT 1820.380 588.870 1820.520 600.030 ;
        RECT 1820.320 588.550 1820.580 588.870 ;
        RECT 1941.760 588.550 1942.020 588.870 ;
        RECT 1941.820 587.170 1941.960 588.550 ;
        RECT 1941.760 586.850 1942.020 587.170 ;
        RECT 1980.400 586.850 1980.660 587.170 ;
        RECT 1980.460 584.790 1980.600 586.850 ;
        RECT 1980.400 584.470 1980.660 584.790 ;
        RECT 2011.220 584.470 2011.480 584.790 ;
        RECT 2011.280 14.270 2011.420 584.470 ;
        RECT 2186.020 14.630 2186.280 14.950 ;
        RECT 2011.220 13.950 2011.480 14.270 ;
        RECT 2186.080 13.930 2186.220 14.630 ;
        RECT 2232.940 13.950 2233.200 14.270 ;
        RECT 2186.020 13.610 2186.280 13.930 ;
        RECT 2233.000 2.400 2233.140 13.950 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 787.590 30.840 787.910 30.900 ;
        RECT 1070.490 30.840 1070.810 30.900 ;
        RECT 787.590 30.700 1070.810 30.840 ;
        RECT 787.590 30.640 787.910 30.700 ;
        RECT 1070.490 30.640 1070.810 30.700 ;
      LAYER via ;
        RECT 787.620 30.640 787.880 30.900 ;
        RECT 1070.520 30.640 1070.780 30.900 ;
      LAYER met2 ;
        RECT 1075.350 600.170 1075.630 604.000 ;
        RECT 1072.880 600.030 1075.630 600.170 ;
        RECT 1072.880 587.250 1073.020 600.030 ;
        RECT 1075.350 600.000 1075.630 600.030 ;
        RECT 1070.580 587.110 1073.020 587.250 ;
        RECT 1070.580 30.930 1070.720 587.110 ;
        RECT 787.620 30.610 787.880 30.930 ;
        RECT 1070.520 30.610 1070.780 30.930 ;
        RECT 787.680 2.400 787.820 30.610 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1829.950 591.840 1830.270 591.900 ;
        RECT 2249.470 591.840 2249.790 591.900 ;
        RECT 1829.950 591.700 2249.790 591.840 ;
        RECT 1829.950 591.640 1830.270 591.700 ;
        RECT 2249.470 591.640 2249.790 591.700 ;
      LAYER via ;
        RECT 1829.980 591.640 1830.240 591.900 ;
        RECT 2249.500 591.640 2249.760 591.900 ;
      LAYER met2 ;
        RECT 1828.370 600.170 1828.650 604.000 ;
        RECT 1828.370 600.030 1830.180 600.170 ;
        RECT 1828.370 600.000 1828.650 600.030 ;
        RECT 1830.040 591.930 1830.180 600.030 ;
        RECT 1829.980 591.610 1830.240 591.930 ;
        RECT 2249.500 591.610 2249.760 591.930 ;
        RECT 2249.560 3.130 2249.700 591.610 ;
        RECT 2249.560 2.990 2251.080 3.130 ;
        RECT 2250.940 2.400 2251.080 2.990 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1839.150 590.140 1839.470 590.200 ;
        RECT 1853.410 590.140 1853.730 590.200 ;
        RECT 1839.150 590.000 1853.730 590.140 ;
        RECT 1839.150 589.940 1839.470 590.000 ;
        RECT 1853.410 589.940 1853.730 590.000 ;
        RECT 1853.410 587.420 1853.730 587.480 ;
        RECT 1886.990 587.420 1887.310 587.480 ;
        RECT 1853.410 587.280 1887.310 587.420 ;
        RECT 1853.410 587.220 1853.730 587.280 ;
        RECT 1886.990 587.220 1887.310 587.280 ;
        RECT 1886.990 15.200 1887.310 15.260 ;
        RECT 2268.330 15.200 2268.650 15.260 ;
        RECT 1886.990 15.060 2268.650 15.200 ;
        RECT 1886.990 15.000 1887.310 15.060 ;
        RECT 2268.330 15.000 2268.650 15.060 ;
      LAYER via ;
        RECT 1839.180 589.940 1839.440 590.200 ;
        RECT 1853.440 589.940 1853.700 590.200 ;
        RECT 1853.440 587.220 1853.700 587.480 ;
        RECT 1887.020 587.220 1887.280 587.480 ;
        RECT 1887.020 15.000 1887.280 15.260 ;
        RECT 2268.360 15.000 2268.620 15.260 ;
      LAYER met2 ;
        RECT 1837.570 600.170 1837.850 604.000 ;
        RECT 1837.570 600.030 1839.380 600.170 ;
        RECT 1837.570 600.000 1837.850 600.030 ;
        RECT 1839.240 590.230 1839.380 600.030 ;
        RECT 1839.180 589.910 1839.440 590.230 ;
        RECT 1853.440 589.910 1853.700 590.230 ;
        RECT 1853.500 587.510 1853.640 589.910 ;
        RECT 1853.440 587.190 1853.700 587.510 ;
        RECT 1887.020 587.190 1887.280 587.510 ;
        RECT 1887.080 15.290 1887.220 587.190 ;
        RECT 1887.020 14.970 1887.280 15.290 ;
        RECT 2268.360 14.970 2268.620 15.290 ;
        RECT 2268.420 2.400 2268.560 14.970 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.350 590.820 1848.670 590.880 ;
        RECT 2283.970 590.820 2284.290 590.880 ;
        RECT 1848.350 590.680 2284.290 590.820 ;
        RECT 1848.350 590.620 1848.670 590.680 ;
        RECT 2283.970 590.620 2284.290 590.680 ;
        RECT 2283.970 2.960 2284.290 3.020 ;
        RECT 2286.270 2.960 2286.590 3.020 ;
        RECT 2283.970 2.820 2286.590 2.960 ;
        RECT 2283.970 2.760 2284.290 2.820 ;
        RECT 2286.270 2.760 2286.590 2.820 ;
      LAYER via ;
        RECT 1848.380 590.620 1848.640 590.880 ;
        RECT 2284.000 590.620 2284.260 590.880 ;
        RECT 2284.000 2.760 2284.260 3.020 ;
        RECT 2286.300 2.760 2286.560 3.020 ;
      LAYER met2 ;
        RECT 1846.770 600.170 1847.050 604.000 ;
        RECT 1846.770 600.030 1848.580 600.170 ;
        RECT 1846.770 600.000 1847.050 600.030 ;
        RECT 1848.440 590.910 1848.580 600.030 ;
        RECT 1848.380 590.590 1848.640 590.910 ;
        RECT 2284.000 590.590 2284.260 590.910 ;
        RECT 2284.060 3.050 2284.200 590.590 ;
        RECT 2284.000 2.730 2284.260 3.050 ;
        RECT 2286.300 2.730 2286.560 3.050 ;
        RECT 2286.360 2.400 2286.500 2.730 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1857.550 587.080 1857.870 587.140 ;
        RECT 1862.610 587.080 1862.930 587.140 ;
        RECT 1857.550 586.940 1862.930 587.080 ;
        RECT 1857.550 586.880 1857.870 586.940 ;
        RECT 1862.610 586.880 1862.930 586.940 ;
        RECT 1862.610 15.540 1862.930 15.600 ;
        RECT 2304.210 15.540 2304.530 15.600 ;
        RECT 1862.610 15.400 2304.530 15.540 ;
        RECT 1862.610 15.340 1862.930 15.400 ;
        RECT 2304.210 15.340 2304.530 15.400 ;
      LAYER via ;
        RECT 1857.580 586.880 1857.840 587.140 ;
        RECT 1862.640 586.880 1862.900 587.140 ;
        RECT 1862.640 15.340 1862.900 15.600 ;
        RECT 2304.240 15.340 2304.500 15.600 ;
      LAYER met2 ;
        RECT 1855.970 600.170 1856.250 604.000 ;
        RECT 1855.970 600.030 1857.780 600.170 ;
        RECT 1855.970 600.000 1856.250 600.030 ;
        RECT 1857.640 587.170 1857.780 600.030 ;
        RECT 1857.580 586.850 1857.840 587.170 ;
        RECT 1862.640 586.850 1862.900 587.170 ;
        RECT 1862.700 15.630 1862.840 586.850 ;
        RECT 1862.640 15.310 1862.900 15.630 ;
        RECT 2304.240 15.310 2304.500 15.630 ;
        RECT 2304.300 2.400 2304.440 15.310 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1866.750 590.480 1867.070 590.540 ;
        RECT 2319.850 590.480 2320.170 590.540 ;
        RECT 1866.750 590.340 2320.170 590.480 ;
        RECT 1866.750 590.280 1867.070 590.340 ;
        RECT 2319.850 590.280 2320.170 590.340 ;
        RECT 2318.470 585.040 2318.790 585.100 ;
        RECT 2321.230 585.040 2321.550 585.100 ;
        RECT 2318.470 584.900 2321.550 585.040 ;
        RECT 2318.470 584.840 2318.790 584.900 ;
        RECT 2321.230 584.840 2321.550 584.900 ;
        RECT 2318.470 62.120 2318.790 62.180 ;
        RECT 2321.690 62.120 2322.010 62.180 ;
        RECT 2318.470 61.980 2322.010 62.120 ;
        RECT 2318.470 61.920 2318.790 61.980 ;
        RECT 2321.690 61.920 2322.010 61.980 ;
      LAYER via ;
        RECT 1866.780 590.280 1867.040 590.540 ;
        RECT 2319.880 590.280 2320.140 590.540 ;
        RECT 2318.500 584.840 2318.760 585.100 ;
        RECT 2321.260 584.840 2321.520 585.100 ;
        RECT 2318.500 61.920 2318.760 62.180 ;
        RECT 2321.720 61.920 2321.980 62.180 ;
      LAYER met2 ;
        RECT 1865.170 600.170 1865.450 604.000 ;
        RECT 1865.170 600.030 1866.980 600.170 ;
        RECT 1865.170 600.000 1865.450 600.030 ;
        RECT 1866.840 590.570 1866.980 600.030 ;
        RECT 2319.940 591.020 2321.460 591.160 ;
        RECT 2319.940 590.570 2320.080 591.020 ;
        RECT 1866.780 590.250 1867.040 590.570 ;
        RECT 2319.880 590.250 2320.140 590.570 ;
        RECT 2321.320 585.130 2321.460 591.020 ;
        RECT 2318.500 584.810 2318.760 585.130 ;
        RECT 2321.260 584.810 2321.520 585.130 ;
        RECT 2318.560 62.210 2318.700 584.810 ;
        RECT 2318.500 61.890 2318.760 62.210 ;
        RECT 2321.720 61.890 2321.980 62.210 ;
        RECT 2321.780 61.610 2321.920 61.890 ;
        RECT 2321.780 61.470 2322.380 61.610 ;
        RECT 2322.240 2.400 2322.380 61.470 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.410 15.880 1876.730 15.940 ;
        RECT 2339.630 15.880 2339.950 15.940 ;
        RECT 1876.410 15.740 2339.950 15.880 ;
        RECT 1876.410 15.680 1876.730 15.740 ;
        RECT 2339.630 15.680 2339.950 15.740 ;
      LAYER via ;
        RECT 1876.440 15.680 1876.700 15.940 ;
        RECT 2339.660 15.680 2339.920 15.940 ;
      LAYER met2 ;
        RECT 1874.370 600.170 1874.650 604.000 ;
        RECT 1874.370 600.030 1876.640 600.170 ;
        RECT 1874.370 600.000 1874.650 600.030 ;
        RECT 1876.500 15.970 1876.640 600.030 ;
        RECT 1876.440 15.650 1876.700 15.970 ;
        RECT 2339.660 15.650 2339.920 15.970 ;
        RECT 2339.720 2.400 2339.860 15.650 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1885.150 591.500 1885.470 591.560 ;
        RECT 1921.490 591.500 1921.810 591.560 ;
        RECT 1885.150 591.360 1921.810 591.500 ;
        RECT 1885.150 591.300 1885.470 591.360 ;
        RECT 1921.490 591.300 1921.810 591.360 ;
        RECT 1921.490 590.140 1921.810 590.200 ;
        RECT 2352.970 590.140 2353.290 590.200 ;
        RECT 1921.490 590.000 2353.290 590.140 ;
        RECT 1921.490 589.940 1921.810 590.000 ;
        RECT 2352.970 589.940 2353.290 590.000 ;
        RECT 2352.970 2.960 2353.290 3.020 ;
        RECT 2357.570 2.960 2357.890 3.020 ;
        RECT 2352.970 2.820 2357.890 2.960 ;
        RECT 2352.970 2.760 2353.290 2.820 ;
        RECT 2357.570 2.760 2357.890 2.820 ;
      LAYER via ;
        RECT 1885.180 591.300 1885.440 591.560 ;
        RECT 1921.520 591.300 1921.780 591.560 ;
        RECT 1921.520 589.940 1921.780 590.200 ;
        RECT 2353.000 589.940 2353.260 590.200 ;
        RECT 2353.000 2.760 2353.260 3.020 ;
        RECT 2357.600 2.760 2357.860 3.020 ;
      LAYER met2 ;
        RECT 1883.570 600.170 1883.850 604.000 ;
        RECT 1883.570 600.030 1885.380 600.170 ;
        RECT 1883.570 600.000 1883.850 600.030 ;
        RECT 1885.240 591.590 1885.380 600.030 ;
        RECT 1885.180 591.270 1885.440 591.590 ;
        RECT 1921.520 591.270 1921.780 591.590 ;
        RECT 1921.580 590.230 1921.720 591.270 ;
        RECT 1921.520 589.910 1921.780 590.230 ;
        RECT 2353.000 589.910 2353.260 590.230 ;
        RECT 2353.060 3.050 2353.200 589.910 ;
        RECT 2353.000 2.730 2353.260 3.050 ;
        RECT 2357.600 2.730 2357.860 3.050 ;
        RECT 2357.660 2.400 2357.800 2.730 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1894.350 586.740 1894.670 586.800 ;
        RECT 1897.110 586.740 1897.430 586.800 ;
        RECT 1894.350 586.600 1897.430 586.740 ;
        RECT 1894.350 586.540 1894.670 586.600 ;
        RECT 1897.110 586.540 1897.430 586.600 ;
        RECT 1897.110 16.220 1897.430 16.280 ;
        RECT 2375.510 16.220 2375.830 16.280 ;
        RECT 1897.110 16.080 2375.830 16.220 ;
        RECT 1897.110 16.020 1897.430 16.080 ;
        RECT 2375.510 16.020 2375.830 16.080 ;
      LAYER via ;
        RECT 1894.380 586.540 1894.640 586.800 ;
        RECT 1897.140 586.540 1897.400 586.800 ;
        RECT 1897.140 16.020 1897.400 16.280 ;
        RECT 2375.540 16.020 2375.800 16.280 ;
      LAYER met2 ;
        RECT 1892.770 600.170 1893.050 604.000 ;
        RECT 1892.770 600.030 1894.580 600.170 ;
        RECT 1892.770 600.000 1893.050 600.030 ;
        RECT 1894.440 586.830 1894.580 600.030 ;
        RECT 1894.380 586.510 1894.640 586.830 ;
        RECT 1897.140 586.510 1897.400 586.830 ;
        RECT 1897.200 16.310 1897.340 586.510 ;
        RECT 1897.140 15.990 1897.400 16.310 ;
        RECT 2375.540 15.990 2375.800 16.310 ;
        RECT 2375.600 2.400 2375.740 15.990 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1903.550 589.800 1903.870 589.860 ;
        RECT 2387.470 589.800 2387.790 589.860 ;
        RECT 1903.550 589.660 2387.790 589.800 ;
        RECT 1903.550 589.600 1903.870 589.660 ;
        RECT 2387.470 589.600 2387.790 589.660 ;
        RECT 2387.470 37.640 2387.790 37.700 ;
        RECT 2393.450 37.640 2393.770 37.700 ;
        RECT 2387.470 37.500 2393.770 37.640 ;
        RECT 2387.470 37.440 2387.790 37.500 ;
        RECT 2393.450 37.440 2393.770 37.500 ;
      LAYER via ;
        RECT 1903.580 589.600 1903.840 589.860 ;
        RECT 2387.500 589.600 2387.760 589.860 ;
        RECT 2387.500 37.440 2387.760 37.700 ;
        RECT 2393.480 37.440 2393.740 37.700 ;
      LAYER met2 ;
        RECT 1901.970 600.170 1902.250 604.000 ;
        RECT 1901.970 600.030 1903.780 600.170 ;
        RECT 1901.970 600.000 1902.250 600.030 ;
        RECT 1903.640 589.890 1903.780 600.030 ;
        RECT 1903.580 589.570 1903.840 589.890 ;
        RECT 2387.500 589.570 2387.760 589.890 ;
        RECT 2387.560 37.730 2387.700 589.570 ;
        RECT 2387.500 37.410 2387.760 37.730 ;
        RECT 2393.480 37.410 2393.740 37.730 ;
        RECT 2393.540 2.400 2393.680 37.410 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1912.750 586.740 1913.070 586.800 ;
        RECT 1917.810 586.740 1918.130 586.800 ;
        RECT 1912.750 586.600 1918.130 586.740 ;
        RECT 1912.750 586.540 1913.070 586.600 ;
        RECT 1917.810 586.540 1918.130 586.600 ;
        RECT 1917.350 16.560 1917.670 16.620 ;
        RECT 2411.390 16.560 2411.710 16.620 ;
        RECT 1917.350 16.420 2411.710 16.560 ;
        RECT 1917.350 16.360 1917.670 16.420 ;
        RECT 2411.390 16.360 2411.710 16.420 ;
      LAYER via ;
        RECT 1912.780 586.540 1913.040 586.800 ;
        RECT 1917.840 586.540 1918.100 586.800 ;
        RECT 1917.380 16.360 1917.640 16.620 ;
        RECT 2411.420 16.360 2411.680 16.620 ;
      LAYER met2 ;
        RECT 1911.170 600.170 1911.450 604.000 ;
        RECT 1911.170 600.030 1912.980 600.170 ;
        RECT 1911.170 600.000 1911.450 600.030 ;
        RECT 1912.840 586.830 1912.980 600.030 ;
        RECT 1912.780 586.510 1913.040 586.830 ;
        RECT 1917.840 586.510 1918.100 586.830 ;
        RECT 1917.900 29.140 1918.040 586.510 ;
        RECT 1917.440 29.000 1918.040 29.140 ;
        RECT 1917.440 16.650 1917.580 29.000 ;
        RECT 1917.380 16.330 1917.640 16.650 ;
        RECT 2411.420 16.330 2411.680 16.650 ;
        RECT 2411.480 2.400 2411.620 16.330 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.990 590.480 852.310 590.540 ;
        RECT 1083.370 590.480 1083.690 590.540 ;
        RECT 851.990 590.340 1083.690 590.480 ;
        RECT 851.990 590.280 852.310 590.340 ;
        RECT 1083.370 590.280 1083.690 590.340 ;
        RECT 851.990 20.300 852.310 20.360 ;
        RECT 840.580 20.160 852.310 20.300 ;
        RECT 805.530 19.960 805.850 20.020 ;
        RECT 840.580 19.960 840.720 20.160 ;
        RECT 851.990 20.100 852.310 20.160 ;
        RECT 805.530 19.820 840.720 19.960 ;
        RECT 805.530 19.760 805.850 19.820 ;
      LAYER via ;
        RECT 852.020 590.280 852.280 590.540 ;
        RECT 1083.400 590.280 1083.660 590.540 ;
        RECT 805.560 19.760 805.820 20.020 ;
        RECT 852.020 20.100 852.280 20.360 ;
      LAYER met2 ;
        RECT 1084.550 600.170 1084.830 604.000 ;
        RECT 1083.460 600.030 1084.830 600.170 ;
        RECT 1083.460 590.570 1083.600 600.030 ;
        RECT 1084.550 600.000 1084.830 600.030 ;
        RECT 852.020 590.250 852.280 590.570 ;
        RECT 1083.400 590.250 1083.660 590.570 ;
        RECT 852.080 20.390 852.220 590.250 ;
        RECT 852.020 20.070 852.280 20.390 ;
        RECT 805.560 19.730 805.820 20.050 ;
        RECT 805.620 2.400 805.760 19.730 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 37.980 3.150 38.040 ;
        RECT 669.370 37.980 669.690 38.040 ;
        RECT 2.830 37.840 669.690 37.980 ;
        RECT 2.830 37.780 3.150 37.840 ;
        RECT 669.370 37.780 669.690 37.840 ;
      LAYER via ;
        RECT 2.860 37.780 3.120 38.040 ;
        RECT 669.400 37.780 669.660 38.040 ;
      LAYER met2 ;
        RECT 671.470 600.170 671.750 604.000 ;
        RECT 669.460 600.030 671.750 600.170 ;
        RECT 669.460 38.070 669.600 600.030 ;
        RECT 671.470 600.000 671.750 600.030 ;
        RECT 2.860 37.750 3.120 38.070 ;
        RECT 669.400 37.750 669.660 38.070 ;
        RECT 2.920 2.400 3.060 37.750 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 670.290 596.940 670.610 597.000 ;
        RECT 673.050 596.940 673.370 597.000 ;
        RECT 670.290 596.800 673.370 596.940 ;
        RECT 670.290 596.740 670.610 596.800 ;
        RECT 673.050 596.740 673.370 596.800 ;
        RECT 670.290 572.460 670.610 572.520 ;
        RECT 671.210 572.460 671.530 572.520 ;
        RECT 670.290 572.320 671.530 572.460 ;
        RECT 670.290 572.260 670.610 572.320 ;
        RECT 671.210 572.260 671.530 572.320 ;
        RECT 669.830 524.520 670.150 524.580 ;
        RECT 671.210 524.520 671.530 524.580 ;
        RECT 669.830 524.380 671.530 524.520 ;
        RECT 669.830 524.320 670.150 524.380 ;
        RECT 671.210 524.320 671.530 524.380 ;
        RECT 8.350 38.660 8.670 38.720 ;
        RECT 670.290 38.660 670.610 38.720 ;
        RECT 8.350 38.520 670.610 38.660 ;
        RECT 8.350 38.460 8.670 38.520 ;
        RECT 670.290 38.460 670.610 38.520 ;
      LAYER via ;
        RECT 670.320 596.740 670.580 597.000 ;
        RECT 673.080 596.740 673.340 597.000 ;
        RECT 670.320 572.260 670.580 572.520 ;
        RECT 671.240 572.260 671.500 572.520 ;
        RECT 669.860 524.320 670.120 524.580 ;
        RECT 671.240 524.320 671.500 524.580 ;
        RECT 8.380 38.460 8.640 38.720 ;
        RECT 670.320 38.460 670.580 38.720 ;
      LAYER met2 ;
        RECT 674.230 600.170 674.510 604.000 ;
        RECT 673.140 600.030 674.510 600.170 ;
        RECT 673.140 597.030 673.280 600.030 ;
        RECT 674.230 600.000 674.510 600.030 ;
        RECT 670.320 596.710 670.580 597.030 ;
        RECT 673.080 596.710 673.340 597.030 ;
        RECT 670.380 572.550 670.520 596.710 ;
        RECT 670.320 572.230 670.580 572.550 ;
        RECT 671.240 572.230 671.500 572.550 ;
        RECT 671.300 524.610 671.440 572.230 ;
        RECT 669.860 524.290 670.120 524.610 ;
        RECT 671.240 524.290 671.500 524.610 ;
        RECT 669.920 458.730 670.060 524.290 ;
        RECT 669.920 458.590 670.520 458.730 ;
        RECT 670.380 303.690 670.520 458.590 ;
        RECT 669.920 303.550 670.520 303.690 ;
        RECT 669.920 303.010 670.060 303.550 ;
        RECT 669.920 302.870 670.520 303.010 ;
        RECT 670.380 207.130 670.520 302.870 ;
        RECT 669.920 206.990 670.520 207.130 ;
        RECT 669.920 206.450 670.060 206.990 ;
        RECT 669.920 206.310 670.520 206.450 ;
        RECT 670.380 110.570 670.520 206.310 ;
        RECT 669.920 110.430 670.520 110.570 ;
        RECT 669.920 109.890 670.060 110.430 ;
        RECT 669.920 109.750 670.520 109.890 ;
        RECT 670.380 38.750 670.520 109.750 ;
        RECT 8.380 38.430 8.640 38.750 ;
        RECT 670.320 38.430 670.580 38.750 ;
        RECT 8.440 2.400 8.580 38.430 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 38.320 14.650 38.380 ;
        RECT 676.730 38.320 677.050 38.380 ;
        RECT 14.330 38.180 677.050 38.320 ;
        RECT 14.330 38.120 14.650 38.180 ;
        RECT 676.730 38.120 677.050 38.180 ;
      LAYER via ;
        RECT 14.360 38.120 14.620 38.380 ;
        RECT 676.760 38.120 677.020 38.380 ;
      LAYER met2 ;
        RECT 677.450 600.170 677.730 604.000 ;
        RECT 676.820 600.030 677.730 600.170 ;
        RECT 676.820 38.410 676.960 600.030 ;
        RECT 677.450 600.000 677.730 600.030 ;
        RECT 14.360 38.090 14.620 38.410 ;
        RECT 676.760 38.090 677.020 38.410 ;
        RECT 14.420 2.400 14.560 38.090 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 683.630 554.440 683.950 554.500 ;
        RECT 687.770 554.440 688.090 554.500 ;
        RECT 683.630 554.300 688.090 554.440 ;
        RECT 683.630 554.240 683.950 554.300 ;
        RECT 687.770 554.240 688.090 554.300 ;
        RECT 38.250 39.340 38.570 39.400 ;
        RECT 683.630 39.340 683.950 39.400 ;
        RECT 38.250 39.200 683.950 39.340 ;
        RECT 38.250 39.140 38.570 39.200 ;
        RECT 683.630 39.140 683.950 39.200 ;
      LAYER via ;
        RECT 683.660 554.240 683.920 554.500 ;
        RECT 687.800 554.240 688.060 554.500 ;
        RECT 38.280 39.140 38.540 39.400 ;
        RECT 683.660 39.140 683.920 39.400 ;
      LAYER met2 ;
        RECT 689.410 600.170 689.690 604.000 ;
        RECT 687.860 600.030 689.690 600.170 ;
        RECT 687.860 554.530 688.000 600.030 ;
        RECT 689.410 600.000 689.690 600.030 ;
        RECT 683.660 554.210 683.920 554.530 ;
        RECT 687.800 554.210 688.060 554.530 ;
        RECT 683.720 39.430 683.860 554.210 ;
        RECT 38.280 39.110 38.540 39.430 ;
        RECT 683.660 39.110 683.920 39.430 ;
        RECT 38.340 2.400 38.480 39.110 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 240.650 40.020 240.970 40.080 ;
        RECT 794.030 40.020 794.350 40.080 ;
        RECT 240.650 39.880 794.350 40.020 ;
        RECT 240.650 39.820 240.970 39.880 ;
        RECT 794.030 39.820 794.350 39.880 ;
      LAYER via ;
        RECT 240.680 39.820 240.940 40.080 ;
        RECT 794.060 39.820 794.320 40.080 ;
      LAYER met2 ;
        RECT 793.830 600.000 794.110 604.000 ;
        RECT 793.890 598.810 794.030 600.000 ;
        RECT 793.890 598.670 794.260 598.810 ;
        RECT 794.120 40.110 794.260 598.670 ;
        RECT 240.680 39.790 240.940 40.110 ;
        RECT 794.060 39.790 794.320 40.110 ;
        RECT 240.740 2.400 240.880 39.790 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 47.160 258.450 47.220 ;
        RECT 800.930 47.160 801.250 47.220 ;
        RECT 258.130 47.020 801.250 47.160 ;
        RECT 258.130 46.960 258.450 47.020 ;
        RECT 800.930 46.960 801.250 47.020 ;
      LAYER via ;
        RECT 258.160 46.960 258.420 47.220 ;
        RECT 800.960 46.960 801.220 47.220 ;
      LAYER met2 ;
        RECT 803.030 600.170 803.310 604.000 ;
        RECT 801.020 600.030 803.310 600.170 ;
        RECT 801.020 47.250 801.160 600.030 ;
        RECT 803.030 600.000 803.310 600.030 ;
        RECT 258.160 46.930 258.420 47.250 ;
        RECT 800.960 46.930 801.220 47.250 ;
        RECT 258.220 2.400 258.360 46.930 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 808.750 524.180 809.070 524.240 ;
        RECT 809.670 524.180 809.990 524.240 ;
        RECT 808.750 524.040 809.990 524.180 ;
        RECT 808.750 523.980 809.070 524.040 ;
        RECT 809.670 523.980 809.990 524.040 ;
        RECT 807.830 476.240 808.150 476.300 ;
        RECT 809.670 476.240 809.990 476.300 ;
        RECT 807.830 476.100 809.990 476.240 ;
        RECT 807.830 476.040 808.150 476.100 ;
        RECT 809.670 476.040 809.990 476.100 ;
        RECT 807.830 448.500 808.150 448.760 ;
        RECT 807.920 448.020 808.060 448.500 ;
        RECT 808.290 448.020 808.610 448.080 ;
        RECT 807.920 447.880 808.610 448.020 ;
        RECT 808.290 447.820 808.610 447.880 ;
        RECT 808.290 420.820 808.610 420.880 ;
        RECT 809.670 420.820 809.990 420.880 ;
        RECT 808.290 420.680 809.990 420.820 ;
        RECT 808.290 420.620 808.610 420.680 ;
        RECT 809.670 420.620 809.990 420.680 ;
        RECT 808.750 372.880 809.070 372.940 ;
        RECT 809.670 372.880 809.990 372.940 ;
        RECT 808.750 372.740 809.990 372.880 ;
        RECT 808.750 372.680 809.070 372.740 ;
        RECT 809.670 372.680 809.990 372.740 ;
        RECT 807.830 303.520 808.150 303.580 ;
        RECT 808.750 303.520 809.070 303.580 ;
        RECT 807.830 303.380 809.070 303.520 ;
        RECT 807.830 303.320 808.150 303.380 ;
        RECT 808.750 303.320 809.070 303.380 ;
        RECT 807.830 282.780 808.150 282.840 ;
        RECT 808.750 282.780 809.070 282.840 ;
        RECT 807.830 282.640 809.070 282.780 ;
        RECT 807.830 282.580 808.150 282.640 ;
        RECT 808.750 282.580 809.070 282.640 ;
        RECT 807.830 234.840 808.150 234.900 ;
        RECT 808.750 234.840 809.070 234.900 ;
        RECT 807.830 234.700 809.070 234.840 ;
        RECT 807.830 234.640 808.150 234.700 ;
        RECT 808.750 234.640 809.070 234.700 ;
        RECT 808.750 111.420 809.070 111.480 ;
        RECT 807.920 111.280 809.070 111.420 ;
        RECT 807.920 110.460 808.060 111.280 ;
        RECT 808.750 111.220 809.070 111.280 ;
        RECT 807.830 110.200 808.150 110.460 ;
        RECT 276.070 47.500 276.390 47.560 ;
        RECT 808.750 47.500 809.070 47.560 ;
        RECT 276.070 47.360 809.070 47.500 ;
        RECT 276.070 47.300 276.390 47.360 ;
        RECT 808.750 47.300 809.070 47.360 ;
      LAYER via ;
        RECT 808.780 523.980 809.040 524.240 ;
        RECT 809.700 523.980 809.960 524.240 ;
        RECT 807.860 476.040 808.120 476.300 ;
        RECT 809.700 476.040 809.960 476.300 ;
        RECT 807.860 448.500 808.120 448.760 ;
        RECT 808.320 447.820 808.580 448.080 ;
        RECT 808.320 420.620 808.580 420.880 ;
        RECT 809.700 420.620 809.960 420.880 ;
        RECT 808.780 372.680 809.040 372.940 ;
        RECT 809.700 372.680 809.960 372.940 ;
        RECT 807.860 303.320 808.120 303.580 ;
        RECT 808.780 303.320 809.040 303.580 ;
        RECT 807.860 282.580 808.120 282.840 ;
        RECT 808.780 282.580 809.040 282.840 ;
        RECT 807.860 234.640 808.120 234.900 ;
        RECT 808.780 234.640 809.040 234.900 ;
        RECT 808.780 111.220 809.040 111.480 ;
        RECT 807.860 110.200 808.120 110.460 ;
        RECT 276.100 47.300 276.360 47.560 ;
        RECT 808.780 47.300 809.040 47.560 ;
      LAYER met2 ;
        RECT 812.230 600.170 812.510 604.000 ;
        RECT 810.680 600.030 812.510 600.170 ;
        RECT 810.680 579.885 810.820 600.030 ;
        RECT 812.230 600.000 812.510 600.030 ;
        RECT 808.770 579.515 809.050 579.885 ;
        RECT 810.610 579.515 810.890 579.885 ;
        RECT 808.840 524.270 808.980 579.515 ;
        RECT 808.780 523.950 809.040 524.270 ;
        RECT 809.700 523.950 809.960 524.270 ;
        RECT 809.760 476.330 809.900 523.950 ;
        RECT 807.860 476.010 808.120 476.330 ;
        RECT 809.700 476.010 809.960 476.330 ;
        RECT 807.920 448.790 808.060 476.010 ;
        RECT 807.860 448.470 808.120 448.790 ;
        RECT 808.320 447.790 808.580 448.110 ;
        RECT 808.380 420.910 808.520 447.790 ;
        RECT 808.320 420.590 808.580 420.910 ;
        RECT 809.700 420.590 809.960 420.910 ;
        RECT 809.760 372.970 809.900 420.590 ;
        RECT 808.780 372.650 809.040 372.970 ;
        RECT 809.700 372.650 809.960 372.970 ;
        RECT 808.840 304.370 808.980 372.650 ;
        RECT 808.380 304.230 808.980 304.370 ;
        RECT 808.380 303.690 808.520 304.230 ;
        RECT 807.920 303.610 808.520 303.690 ;
        RECT 807.860 303.550 808.520 303.610 ;
        RECT 807.860 303.290 808.120 303.550 ;
        RECT 808.780 303.290 809.040 303.610 ;
        RECT 808.840 282.870 808.980 303.290 ;
        RECT 807.860 282.550 808.120 282.870 ;
        RECT 808.780 282.550 809.040 282.870 ;
        RECT 807.920 234.930 808.060 282.550 ;
        RECT 807.860 234.610 808.120 234.930 ;
        RECT 808.780 234.610 809.040 234.930 ;
        RECT 808.840 111.510 808.980 234.610 ;
        RECT 808.780 111.190 809.040 111.510 ;
        RECT 807.860 110.170 808.120 110.490 ;
        RECT 807.920 58.890 808.060 110.170 ;
        RECT 807.920 58.750 808.980 58.890 ;
        RECT 808.840 47.590 808.980 58.750 ;
        RECT 276.100 47.270 276.360 47.590 ;
        RECT 808.780 47.270 809.040 47.590 ;
        RECT 276.160 2.400 276.300 47.270 ;
        RECT 275.950 -4.800 276.510 2.400 ;
      LAYER via2 ;
        RECT 808.770 579.560 809.050 579.840 ;
        RECT 810.610 579.560 810.890 579.840 ;
      LAYER met3 ;
        RECT 808.745 579.850 809.075 579.865 ;
        RECT 810.585 579.850 810.915 579.865 ;
        RECT 808.745 579.550 810.915 579.850 ;
        RECT 808.745 579.535 809.075 579.550 ;
        RECT 810.585 579.535 810.915 579.550 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 47.840 294.330 47.900 ;
        RECT 821.630 47.840 821.950 47.900 ;
        RECT 294.010 47.700 821.950 47.840 ;
        RECT 294.010 47.640 294.330 47.700 ;
        RECT 821.630 47.640 821.950 47.700 ;
      LAYER via ;
        RECT 294.040 47.640 294.300 47.900 ;
        RECT 821.660 47.640 821.920 47.900 ;
      LAYER met2 ;
        RECT 821.430 600.000 821.710 604.000 ;
        RECT 821.490 598.810 821.630 600.000 ;
        RECT 821.490 598.670 821.860 598.810 ;
        RECT 821.720 47.930 821.860 598.670 ;
        RECT 294.040 47.610 294.300 47.930 ;
        RECT 821.660 47.610 821.920 47.930 ;
        RECT 294.100 2.400 294.240 47.610 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 26.420 312.270 26.480 ;
        RECT 828.530 26.420 828.850 26.480 ;
        RECT 311.950 26.280 828.850 26.420 ;
        RECT 311.950 26.220 312.270 26.280 ;
        RECT 828.530 26.220 828.850 26.280 ;
      LAYER via ;
        RECT 311.980 26.220 312.240 26.480 ;
        RECT 828.560 26.220 828.820 26.480 ;
      LAYER met2 ;
        RECT 830.630 600.170 830.910 604.000 ;
        RECT 828.620 600.030 830.910 600.170 ;
        RECT 828.620 26.510 828.760 600.030 ;
        RECT 830.630 600.000 830.910 600.030 ;
        RECT 311.980 26.190 312.240 26.510 ;
        RECT 828.560 26.190 828.820 26.510 ;
        RECT 312.040 2.400 312.180 26.190 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.970 569.400 835.290 569.460 ;
        RECT 838.190 569.400 838.510 569.460 ;
        RECT 834.970 569.260 838.510 569.400 ;
        RECT 834.970 569.200 835.290 569.260 ;
        RECT 838.190 569.200 838.510 569.260 ;
        RECT 329.890 26.760 330.210 26.820 ;
        RECT 834.970 26.760 835.290 26.820 ;
        RECT 329.890 26.620 835.290 26.760 ;
        RECT 329.890 26.560 330.210 26.620 ;
        RECT 834.970 26.560 835.290 26.620 ;
      LAYER via ;
        RECT 835.000 569.200 835.260 569.460 ;
        RECT 838.220 569.200 838.480 569.460 ;
        RECT 329.920 26.560 330.180 26.820 ;
        RECT 835.000 26.560 835.260 26.820 ;
      LAYER met2 ;
        RECT 839.830 600.170 840.110 604.000 ;
        RECT 838.280 600.030 840.110 600.170 ;
        RECT 838.280 569.490 838.420 600.030 ;
        RECT 839.830 600.000 840.110 600.030 ;
        RECT 835.000 569.170 835.260 569.490 ;
        RECT 838.220 569.170 838.480 569.490 ;
        RECT 835.060 26.850 835.200 569.170 ;
        RECT 329.920 26.530 330.180 26.850 ;
        RECT 835.000 26.530 835.260 26.850 ;
        RECT 329.980 2.400 330.120 26.530 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 27.100 347.690 27.160 ;
        RECT 849.690 27.100 850.010 27.160 ;
        RECT 347.370 26.960 850.010 27.100 ;
        RECT 347.370 26.900 347.690 26.960 ;
        RECT 849.690 26.900 850.010 26.960 ;
      LAYER via ;
        RECT 347.400 26.900 347.660 27.160 ;
        RECT 849.720 26.900 849.980 27.160 ;
      LAYER met2 ;
        RECT 848.570 600.170 848.850 604.000 ;
        RECT 848.570 600.030 849.920 600.170 ;
        RECT 848.570 600.000 848.850 600.030 ;
        RECT 849.780 27.190 849.920 600.030 ;
        RECT 347.400 26.870 347.660 27.190 ;
        RECT 849.720 26.870 849.980 27.190 ;
        RECT 347.460 2.400 347.600 26.870 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 27.440 365.630 27.500 ;
        RECT 856.130 27.440 856.450 27.500 ;
        RECT 365.310 27.300 856.450 27.440 ;
        RECT 365.310 27.240 365.630 27.300 ;
        RECT 856.130 27.240 856.450 27.300 ;
      LAYER via ;
        RECT 365.340 27.240 365.600 27.500 ;
        RECT 856.160 27.240 856.420 27.500 ;
      LAYER met2 ;
        RECT 857.770 600.170 858.050 604.000 ;
        RECT 856.220 600.030 858.050 600.170 ;
        RECT 856.220 27.530 856.360 600.030 ;
        RECT 857.770 600.000 858.050 600.030 ;
        RECT 365.340 27.210 365.600 27.530 ;
        RECT 856.160 27.210 856.420 27.530 ;
        RECT 365.400 2.400 365.540 27.210 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.570 569.400 862.890 569.460 ;
        RECT 865.330 569.400 865.650 569.460 ;
        RECT 862.570 569.260 865.650 569.400 ;
        RECT 862.570 569.200 862.890 569.260 ;
        RECT 865.330 569.200 865.650 569.260 ;
        RECT 383.250 23.700 383.570 23.760 ;
        RECT 862.570 23.700 862.890 23.760 ;
        RECT 383.250 23.560 862.890 23.700 ;
        RECT 383.250 23.500 383.570 23.560 ;
        RECT 862.570 23.500 862.890 23.560 ;
      LAYER via ;
        RECT 862.600 569.200 862.860 569.460 ;
        RECT 865.360 569.200 865.620 569.460 ;
        RECT 383.280 23.500 383.540 23.760 ;
        RECT 862.600 23.500 862.860 23.760 ;
      LAYER met2 ;
        RECT 866.970 600.170 867.250 604.000 ;
        RECT 865.420 600.030 867.250 600.170 ;
        RECT 865.420 569.490 865.560 600.030 ;
        RECT 866.970 600.000 867.250 600.030 ;
        RECT 862.600 569.170 862.860 569.490 ;
        RECT 865.360 569.170 865.620 569.490 ;
        RECT 862.660 23.790 862.800 569.170 ;
        RECT 383.280 23.470 383.540 23.790 ;
        RECT 862.600 23.470 862.860 23.790 ;
        RECT 383.340 2.400 383.480 23.470 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 23.360 401.510 23.420 ;
        RECT 877.750 23.360 878.070 23.420 ;
        RECT 401.190 23.220 878.070 23.360 ;
        RECT 401.190 23.160 401.510 23.220 ;
        RECT 877.750 23.160 878.070 23.220 ;
      LAYER via ;
        RECT 401.220 23.160 401.480 23.420 ;
        RECT 877.780 23.160 878.040 23.420 ;
      LAYER met2 ;
        RECT 876.170 600.170 876.450 604.000 ;
        RECT 876.170 600.030 877.980 600.170 ;
        RECT 876.170 600.000 876.450 600.030 ;
        RECT 877.840 23.450 877.980 600.030 ;
        RECT 401.220 23.130 401.480 23.450 ;
        RECT 877.780 23.130 878.040 23.450 ;
        RECT 401.280 2.400 401.420 23.130 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 696.970 569.400 697.290 569.460 ;
        RECT 700.190 569.400 700.510 569.460 ;
        RECT 696.970 569.260 700.510 569.400 ;
        RECT 696.970 569.200 697.290 569.260 ;
        RECT 700.190 569.200 700.510 569.260 ;
        RECT 62.170 24.380 62.490 24.440 ;
        RECT 696.970 24.380 697.290 24.440 ;
        RECT 62.170 24.240 697.290 24.380 ;
        RECT 62.170 24.180 62.490 24.240 ;
        RECT 696.970 24.180 697.290 24.240 ;
      LAYER via ;
        RECT 697.000 569.200 697.260 569.460 ;
        RECT 700.220 569.200 700.480 569.460 ;
        RECT 62.200 24.180 62.460 24.440 ;
        RECT 697.000 24.180 697.260 24.440 ;
      LAYER met2 ;
        RECT 701.830 600.170 702.110 604.000 ;
        RECT 700.280 600.030 702.110 600.170 ;
        RECT 700.280 569.490 700.420 600.030 ;
        RECT 701.830 600.000 702.110 600.030 ;
        RECT 697.000 569.170 697.260 569.490 ;
        RECT 700.220 569.170 700.480 569.490 ;
        RECT 697.060 24.470 697.200 569.170 ;
        RECT 62.200 24.150 62.460 24.470 ;
        RECT 697.000 24.150 697.260 24.470 ;
        RECT 62.260 2.400 62.400 24.150 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 23.020 419.450 23.080 ;
        RECT 883.730 23.020 884.050 23.080 ;
        RECT 419.130 22.880 884.050 23.020 ;
        RECT 419.130 22.820 419.450 22.880 ;
        RECT 883.730 22.820 884.050 22.880 ;
      LAYER via ;
        RECT 419.160 22.820 419.420 23.080 ;
        RECT 883.760 22.820 884.020 23.080 ;
      LAYER met2 ;
        RECT 885.370 600.170 885.650 604.000 ;
        RECT 883.820 600.030 885.650 600.170 ;
        RECT 883.820 23.110 883.960 600.030 ;
        RECT 885.370 600.000 885.650 600.030 ;
        RECT 419.160 22.790 419.420 23.110 ;
        RECT 883.760 22.790 884.020 23.110 ;
        RECT 419.220 2.400 419.360 22.790 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 890.170 569.400 890.490 569.460 ;
        RECT 892.930 569.400 893.250 569.460 ;
        RECT 890.170 569.260 893.250 569.400 ;
        RECT 890.170 569.200 890.490 569.260 ;
        RECT 892.930 569.200 893.250 569.260 ;
        RECT 436.610 22.680 436.930 22.740 ;
        RECT 890.170 22.680 890.490 22.740 ;
        RECT 436.610 22.540 890.490 22.680 ;
        RECT 436.610 22.480 436.930 22.540 ;
        RECT 890.170 22.480 890.490 22.540 ;
      LAYER via ;
        RECT 890.200 569.200 890.460 569.460 ;
        RECT 892.960 569.200 893.220 569.460 ;
        RECT 436.640 22.480 436.900 22.740 ;
        RECT 890.200 22.480 890.460 22.740 ;
      LAYER met2 ;
        RECT 894.570 600.170 894.850 604.000 ;
        RECT 893.020 600.030 894.850 600.170 ;
        RECT 893.020 569.490 893.160 600.030 ;
        RECT 894.570 600.000 894.850 600.030 ;
        RECT 890.200 569.170 890.460 569.490 ;
        RECT 892.960 569.170 893.220 569.490 ;
        RECT 890.260 22.770 890.400 569.170 ;
        RECT 436.640 22.450 436.900 22.770 ;
        RECT 890.200 22.450 890.460 22.770 ;
        RECT 436.700 2.400 436.840 22.450 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 33.560 454.870 33.620 ;
        RECT 904.430 33.560 904.750 33.620 ;
        RECT 454.550 33.420 904.750 33.560 ;
        RECT 454.550 33.360 454.870 33.420 ;
        RECT 904.430 33.360 904.750 33.420 ;
      LAYER via ;
        RECT 454.580 33.360 454.840 33.620 ;
        RECT 904.460 33.360 904.720 33.620 ;
      LAYER met2 ;
        RECT 903.770 600.170 904.050 604.000 ;
        RECT 903.770 600.030 904.660 600.170 ;
        RECT 903.770 600.000 904.050 600.030 ;
        RECT 904.520 33.650 904.660 600.030 ;
        RECT 454.580 33.330 454.840 33.650 ;
        RECT 904.460 33.330 904.720 33.650 ;
        RECT 454.640 2.400 454.780 33.330 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 34.240 472.810 34.300 ;
        RECT 911.330 34.240 911.650 34.300 ;
        RECT 472.490 34.100 911.650 34.240 ;
        RECT 472.490 34.040 472.810 34.100 ;
        RECT 911.330 34.040 911.650 34.100 ;
      LAYER via ;
        RECT 472.520 34.040 472.780 34.300 ;
        RECT 911.360 34.040 911.620 34.300 ;
      LAYER met2 ;
        RECT 912.970 600.170 913.250 604.000 ;
        RECT 911.420 600.030 913.250 600.170 ;
        RECT 911.420 34.330 911.560 600.030 ;
        RECT 912.970 600.000 913.250 600.030 ;
        RECT 472.520 34.010 472.780 34.330 ;
        RECT 911.360 34.010 911.620 34.330 ;
        RECT 472.580 2.400 472.720 34.010 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 918.690 572.800 919.010 572.860 ;
        RECT 920.530 572.800 920.850 572.860 ;
        RECT 918.690 572.660 920.850 572.800 ;
        RECT 918.690 572.600 919.010 572.660 ;
        RECT 920.530 572.600 920.850 572.660 ;
        RECT 918.230 531.660 918.550 531.720 ;
        RECT 918.690 531.660 919.010 531.720 ;
        RECT 918.230 531.520 919.010 531.660 ;
        RECT 918.230 531.460 918.550 531.520 ;
        RECT 918.690 531.460 919.010 531.520 ;
        RECT 918.690 524.180 919.010 524.240 ;
        RECT 919.150 524.180 919.470 524.240 ;
        RECT 918.690 524.040 919.470 524.180 ;
        RECT 918.690 523.980 919.010 524.040 ;
        RECT 919.150 523.980 919.470 524.040 ;
        RECT 918.690 380.160 919.010 380.420 ;
        RECT 918.780 379.740 918.920 380.160 ;
        RECT 918.690 379.480 919.010 379.740 ;
        RECT 918.690 351.940 919.010 352.200 ;
        RECT 918.780 351.800 918.920 351.940 ;
        RECT 919.150 351.800 919.470 351.860 ;
        RECT 918.780 351.660 919.470 351.800 ;
        RECT 919.150 351.600 919.470 351.660 ;
        RECT 918.690 331.400 919.010 331.460 ;
        RECT 919.150 331.400 919.470 331.460 ;
        RECT 918.690 331.260 919.470 331.400 ;
        RECT 918.690 331.200 919.010 331.260 ;
        RECT 919.150 331.200 919.470 331.260 ;
        RECT 918.230 303.520 918.550 303.580 ;
        RECT 919.150 303.520 919.470 303.580 ;
        RECT 918.230 303.380 919.470 303.520 ;
        RECT 918.230 303.320 918.550 303.380 ;
        RECT 919.150 303.320 919.470 303.380 ;
        RECT 918.690 137.740 919.010 138.000 ;
        RECT 918.780 137.320 918.920 137.740 ;
        RECT 918.690 137.060 919.010 137.320 ;
        RECT 918.230 90.000 918.550 90.060 ;
        RECT 918.690 90.000 919.010 90.060 ;
        RECT 918.230 89.860 919.010 90.000 ;
        RECT 918.230 89.800 918.550 89.860 ;
        RECT 918.690 89.800 919.010 89.860 ;
        RECT 490.430 30.160 490.750 30.220 ;
        RECT 919.150 30.160 919.470 30.220 ;
        RECT 490.430 30.020 919.470 30.160 ;
        RECT 490.430 29.960 490.750 30.020 ;
        RECT 919.150 29.960 919.470 30.020 ;
      LAYER via ;
        RECT 918.720 572.600 918.980 572.860 ;
        RECT 920.560 572.600 920.820 572.860 ;
        RECT 918.260 531.460 918.520 531.720 ;
        RECT 918.720 531.460 918.980 531.720 ;
        RECT 918.720 523.980 918.980 524.240 ;
        RECT 919.180 523.980 919.440 524.240 ;
        RECT 918.720 380.160 918.980 380.420 ;
        RECT 918.720 379.480 918.980 379.740 ;
        RECT 918.720 351.940 918.980 352.200 ;
        RECT 919.180 351.600 919.440 351.860 ;
        RECT 918.720 331.200 918.980 331.460 ;
        RECT 919.180 331.200 919.440 331.460 ;
        RECT 918.260 303.320 918.520 303.580 ;
        RECT 919.180 303.320 919.440 303.580 ;
        RECT 918.720 137.740 918.980 138.000 ;
        RECT 918.720 137.060 918.980 137.320 ;
        RECT 918.260 89.800 918.520 90.060 ;
        RECT 918.720 89.800 918.980 90.060 ;
        RECT 490.460 29.960 490.720 30.220 ;
        RECT 919.180 29.960 919.440 30.220 ;
      LAYER met2 ;
        RECT 922.170 600.170 922.450 604.000 ;
        RECT 920.620 600.030 922.450 600.170 ;
        RECT 920.620 572.890 920.760 600.030 ;
        RECT 922.170 600.000 922.450 600.030 ;
        RECT 918.720 572.570 918.980 572.890 ;
        RECT 920.560 572.570 920.820 572.890 ;
        RECT 918.780 555.970 918.920 572.570 ;
        RECT 918.320 555.830 918.920 555.970 ;
        RECT 918.320 531.750 918.460 555.830 ;
        RECT 918.260 531.430 918.520 531.750 ;
        RECT 918.720 531.430 918.980 531.750 ;
        RECT 918.780 524.270 918.920 531.430 ;
        RECT 918.720 523.950 918.980 524.270 ;
        RECT 919.180 523.950 919.440 524.270 ;
        RECT 919.240 447.170 919.380 523.950 ;
        RECT 918.780 447.030 919.380 447.170 ;
        RECT 918.780 380.450 918.920 447.030 ;
        RECT 918.720 380.130 918.980 380.450 ;
        RECT 918.720 379.450 918.980 379.770 ;
        RECT 918.780 352.230 918.920 379.450 ;
        RECT 918.720 351.910 918.980 352.230 ;
        RECT 919.180 351.570 919.440 351.890 ;
        RECT 919.240 331.490 919.380 351.570 ;
        RECT 918.720 331.170 918.980 331.490 ;
        RECT 919.180 331.170 919.440 331.490 ;
        RECT 918.780 303.690 918.920 331.170 ;
        RECT 918.320 303.610 918.920 303.690 ;
        RECT 918.260 303.550 918.920 303.610 ;
        RECT 918.260 303.290 918.520 303.550 ;
        RECT 919.180 303.290 919.440 303.610 ;
        RECT 919.240 211.210 919.380 303.290 ;
        RECT 918.780 211.070 919.380 211.210 ;
        RECT 918.780 158.850 918.920 211.070 ;
        RECT 918.320 158.710 918.920 158.850 ;
        RECT 918.320 158.170 918.460 158.710 ;
        RECT 918.320 158.030 918.920 158.170 ;
        RECT 918.780 138.030 918.920 158.030 ;
        RECT 918.720 137.710 918.980 138.030 ;
        RECT 918.720 137.030 918.980 137.350 ;
        RECT 918.780 90.090 918.920 137.030 ;
        RECT 918.260 89.770 918.520 90.090 ;
        RECT 918.720 89.770 918.980 90.090 ;
        RECT 918.320 58.890 918.460 89.770 ;
        RECT 918.320 58.750 919.380 58.890 ;
        RECT 919.240 30.250 919.380 58.750 ;
        RECT 490.460 29.930 490.720 30.250 ;
        RECT 919.180 29.930 919.440 30.250 ;
        RECT 490.520 2.400 490.660 29.930 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 30.500 508.230 30.560 ;
        RECT 932.490 30.500 932.810 30.560 ;
        RECT 507.910 30.360 932.810 30.500 ;
        RECT 507.910 30.300 508.230 30.360 ;
        RECT 932.490 30.300 932.810 30.360 ;
      LAYER via ;
        RECT 507.940 30.300 508.200 30.560 ;
        RECT 932.520 30.300 932.780 30.560 ;
      LAYER met2 ;
        RECT 931.370 600.170 931.650 604.000 ;
        RECT 931.370 600.030 932.720 600.170 ;
        RECT 931.370 600.000 931.650 600.030 ;
        RECT 932.580 30.590 932.720 600.030 ;
        RECT 507.940 30.270 508.200 30.590 ;
        RECT 932.520 30.270 932.780 30.590 ;
        RECT 508.000 2.400 508.140 30.270 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 32.540 526.170 32.600 ;
        RECT 938.470 32.540 938.790 32.600 ;
        RECT 525.850 32.400 938.790 32.540 ;
        RECT 525.850 32.340 526.170 32.400 ;
        RECT 938.470 32.340 938.790 32.400 ;
      LAYER via ;
        RECT 525.880 32.340 526.140 32.600 ;
        RECT 938.500 32.340 938.760 32.600 ;
      LAYER met2 ;
        RECT 940.570 600.170 940.850 604.000 ;
        RECT 938.560 600.030 940.850 600.170 ;
        RECT 938.560 32.630 938.700 600.030 ;
        RECT 940.570 600.000 940.850 600.030 ;
        RECT 525.880 32.310 526.140 32.630 ;
        RECT 938.500 32.310 938.760 32.630 ;
        RECT 525.940 2.400 526.080 32.310 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 945.370 557.840 945.690 557.900 ;
        RECT 948.130 557.840 948.450 557.900 ;
        RECT 945.370 557.700 948.450 557.840 ;
        RECT 945.370 557.640 945.690 557.700 ;
        RECT 948.130 557.640 948.450 557.700 ;
        RECT 543.790 29.820 544.110 29.880 ;
        RECT 945.370 29.820 945.690 29.880 ;
        RECT 543.790 29.680 945.690 29.820 ;
        RECT 543.790 29.620 544.110 29.680 ;
        RECT 945.370 29.620 945.690 29.680 ;
      LAYER via ;
        RECT 945.400 557.640 945.660 557.900 ;
        RECT 948.160 557.640 948.420 557.900 ;
        RECT 543.820 29.620 544.080 29.880 ;
        RECT 945.400 29.620 945.660 29.880 ;
      LAYER met2 ;
        RECT 949.770 600.170 950.050 604.000 ;
        RECT 948.220 600.030 950.050 600.170 ;
        RECT 948.220 557.930 948.360 600.030 ;
        RECT 949.770 600.000 950.050 600.030 ;
        RECT 945.400 557.610 945.660 557.930 ;
        RECT 948.160 557.610 948.420 557.930 ;
        RECT 945.460 29.910 945.600 557.610 ;
        RECT 543.820 29.590 544.080 29.910 ;
        RECT 945.400 29.590 945.660 29.910 ;
        RECT 543.880 2.400 544.020 29.590 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 29.480 562.050 29.540 ;
        RECT 959.170 29.480 959.490 29.540 ;
        RECT 561.730 29.340 959.490 29.480 ;
        RECT 561.730 29.280 562.050 29.340 ;
        RECT 959.170 29.280 959.490 29.340 ;
      LAYER via ;
        RECT 561.760 29.280 562.020 29.540 ;
        RECT 959.200 29.280 959.460 29.540 ;
      LAYER met2 ;
        RECT 958.970 600.000 959.250 604.000 ;
        RECT 959.030 598.810 959.170 600.000 ;
        RECT 959.030 598.670 959.400 598.810 ;
        RECT 959.260 29.570 959.400 598.670 ;
        RECT 561.760 29.250 562.020 29.570 ;
        RECT 959.200 29.250 959.460 29.570 ;
        RECT 561.820 2.400 561.960 29.250 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 28.800 579.990 28.860 ;
        RECT 966.070 28.800 966.390 28.860 ;
        RECT 579.670 28.660 966.390 28.800 ;
        RECT 579.670 28.600 579.990 28.660 ;
        RECT 966.070 28.600 966.390 28.660 ;
      LAYER via ;
        RECT 579.700 28.600 579.960 28.860 ;
        RECT 966.100 28.600 966.360 28.860 ;
      LAYER met2 ;
        RECT 968.170 600.170 968.450 604.000 ;
        RECT 966.160 600.030 968.450 600.170 ;
        RECT 966.160 28.890 966.300 600.030 ;
        RECT 968.170 600.000 968.450 600.030 ;
        RECT 579.700 28.570 579.960 28.890 ;
        RECT 966.100 28.570 966.360 28.890 ;
        RECT 579.760 2.400 579.900 28.570 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 654.650 594.560 654.970 594.620 ;
        RECT 711.230 594.560 711.550 594.620 ;
        RECT 712.610 594.560 712.930 594.620 ;
        RECT 654.650 594.420 712.930 594.560 ;
        RECT 654.650 594.360 654.970 594.420 ;
        RECT 711.230 594.360 711.550 594.420 ;
        RECT 712.610 594.360 712.930 594.420 ;
        RECT 86.090 24.040 86.410 24.100 ;
        RECT 711.230 24.040 711.550 24.100 ;
        RECT 86.090 23.900 711.550 24.040 ;
        RECT 86.090 23.840 86.410 23.900 ;
        RECT 711.230 23.840 711.550 23.900 ;
      LAYER via ;
        RECT 654.680 594.360 654.940 594.620 ;
        RECT 711.260 594.360 711.520 594.620 ;
        RECT 712.640 594.360 712.900 594.620 ;
        RECT 86.120 23.840 86.380 24.100 ;
        RECT 711.260 23.840 711.520 24.100 ;
      LAYER met2 ;
        RECT 654.670 2500.515 654.950 2500.885 ;
        RECT 654.740 594.650 654.880 2500.515 ;
        RECT 714.250 600.170 714.530 604.000 ;
        RECT 712.700 600.030 714.530 600.170 ;
        RECT 712.700 594.650 712.840 600.030 ;
        RECT 714.250 600.000 714.530 600.030 ;
        RECT 654.680 594.330 654.940 594.650 ;
        RECT 711.260 594.330 711.520 594.650 ;
        RECT 712.640 594.330 712.900 594.650 ;
        RECT 711.320 24.130 711.460 594.330 ;
        RECT 86.120 23.810 86.380 24.130 ;
        RECT 711.260 23.810 711.520 24.130 ;
        RECT 86.180 2.400 86.320 23.810 ;
        RECT 85.970 -4.800 86.530 2.400 ;
      LAYER via2 ;
        RECT 654.670 2500.560 654.950 2500.840 ;
      LAYER met3 ;
        RECT 1885.335 2707.080 1889.335 2707.360 ;
        RECT 1885.335 2706.760 1889.370 2707.080 ;
        RECT 1889.070 2705.530 1889.370 2706.760 ;
        RECT 1898.230 2705.530 1898.610 2705.540 ;
        RECT 1889.070 2705.230 1898.610 2705.530 ;
        RECT 1898.230 2705.220 1898.610 2705.230 ;
        RECT 654.645 2500.850 654.975 2500.865 ;
        RECT 1898.230 2500.850 1898.610 2500.860 ;
        RECT 654.645 2500.550 1898.610 2500.850 ;
        RECT 654.645 2500.535 654.975 2500.550 ;
        RECT 1898.230 2500.540 1898.610 2500.550 ;
      LAYER via3 ;
        RECT 1898.260 2705.220 1898.580 2705.540 ;
        RECT 1898.260 2500.540 1898.580 2500.860 ;
      LAYER met4 ;
        RECT 1898.255 2705.215 1898.585 2705.545 ;
        RECT 1898.270 2500.865 1898.570 2705.215 ;
        RECT 1898.255 2500.535 1898.585 2500.865 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 973.430 569.400 973.750 569.460 ;
        RECT 975.730 569.400 976.050 569.460 ;
        RECT 973.430 569.260 976.050 569.400 ;
        RECT 973.430 569.200 973.750 569.260 ;
        RECT 975.730 569.200 976.050 569.260 ;
        RECT 597.150 28.460 597.470 28.520 ;
        RECT 973.430 28.460 973.750 28.520 ;
        RECT 597.150 28.320 973.750 28.460 ;
        RECT 597.150 28.260 597.470 28.320 ;
        RECT 973.430 28.260 973.750 28.320 ;
      LAYER via ;
        RECT 973.460 569.200 973.720 569.460 ;
        RECT 975.760 569.200 976.020 569.460 ;
        RECT 597.180 28.260 597.440 28.520 ;
        RECT 973.460 28.260 973.720 28.520 ;
      LAYER met2 ;
        RECT 977.370 600.170 977.650 604.000 ;
        RECT 975.820 600.030 977.650 600.170 ;
        RECT 975.820 569.490 975.960 600.030 ;
        RECT 977.370 600.000 977.650 600.030 ;
        RECT 973.460 569.170 973.720 569.490 ;
        RECT 975.760 569.170 976.020 569.490 ;
        RECT 973.520 28.550 973.660 569.170 ;
        RECT 597.180 28.230 597.440 28.550 ;
        RECT 973.460 28.230 973.720 28.550 ;
        RECT 597.240 2.400 597.380 28.230 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 28.120 615.410 28.180 ;
        RECT 986.770 28.120 987.090 28.180 ;
        RECT 615.090 27.980 987.090 28.120 ;
        RECT 615.090 27.920 615.410 27.980 ;
        RECT 986.770 27.920 987.090 27.980 ;
      LAYER via ;
        RECT 615.120 27.920 615.380 28.180 ;
        RECT 986.800 27.920 987.060 28.180 ;
      LAYER met2 ;
        RECT 986.570 600.000 986.850 604.000 ;
        RECT 986.630 598.810 986.770 600.000 ;
        RECT 986.630 598.670 987.000 598.810 ;
        RECT 986.860 28.210 987.000 598.670 ;
        RECT 615.120 27.890 615.380 28.210 ;
        RECT 986.800 27.890 987.060 28.210 ;
        RECT 615.180 2.400 615.320 27.890 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 647.750 2815.440 648.070 2815.500 ;
        RECT 1483.570 2815.440 1483.890 2815.500 ;
        RECT 647.750 2815.300 1483.890 2815.440 ;
        RECT 647.750 2815.240 648.070 2815.300 ;
        RECT 1483.570 2815.240 1483.890 2815.300 ;
        RECT 647.750 594.220 648.070 594.280 ;
        RECT 724.570 594.220 724.890 594.280 ;
        RECT 647.750 594.080 724.890 594.220 ;
        RECT 647.750 594.020 648.070 594.080 ;
        RECT 724.570 594.020 724.890 594.080 ;
        RECT 724.570 572.460 724.890 572.520 ;
        RECT 725.490 572.460 725.810 572.520 ;
        RECT 724.570 572.320 725.810 572.460 ;
        RECT 724.570 572.260 724.890 572.320 ;
        RECT 725.490 572.260 725.810 572.320 ;
        RECT 725.030 338.200 725.350 338.260 ;
        RECT 725.490 338.200 725.810 338.260 ;
        RECT 725.030 338.060 725.810 338.200 ;
        RECT 725.030 338.000 725.350 338.060 ;
        RECT 725.490 338.000 725.810 338.060 ;
        RECT 723.650 324.260 723.970 324.320 ;
        RECT 725.030 324.260 725.350 324.320 ;
        RECT 723.650 324.120 725.350 324.260 ;
        RECT 723.650 324.060 723.970 324.120 ;
        RECT 725.030 324.060 725.350 324.120 ;
        RECT 723.650 276.320 723.970 276.380 ;
        RECT 724.570 276.320 724.890 276.380 ;
        RECT 723.650 276.180 724.890 276.320 ;
        RECT 723.650 276.120 723.970 276.180 ;
        RECT 724.570 276.120 724.890 276.180 ;
        RECT 724.110 234.500 724.430 234.560 ;
        RECT 725.030 234.500 725.350 234.560 ;
        RECT 724.110 234.360 725.350 234.500 ;
        RECT 724.110 234.300 724.430 234.360 ;
        RECT 725.030 234.300 725.350 234.360 ;
        RECT 722.730 227.700 723.050 227.760 ;
        RECT 724.110 227.700 724.430 227.760 ;
        RECT 722.730 227.560 724.430 227.700 ;
        RECT 722.730 227.500 723.050 227.560 ;
        RECT 724.110 227.500 724.430 227.560 ;
        RECT 722.730 179.760 723.050 179.820 ;
        RECT 723.650 179.760 723.970 179.820 ;
        RECT 722.730 179.620 723.970 179.760 ;
        RECT 722.730 179.560 723.050 179.620 ;
        RECT 723.650 179.560 723.970 179.620 ;
        RECT 723.650 138.280 723.970 138.340 ;
        RECT 724.570 138.280 724.890 138.340 ;
        RECT 723.650 138.140 724.890 138.280 ;
        RECT 723.650 138.080 723.970 138.140 ;
        RECT 724.570 138.080 724.890 138.140 ;
        RECT 724.570 110.400 724.890 110.460 ;
        RECT 725.490 110.400 725.810 110.460 ;
        RECT 724.570 110.260 725.810 110.400 ;
        RECT 724.570 110.200 724.890 110.260 ;
        RECT 725.490 110.200 725.810 110.260 ;
        RECT 109.550 24.720 109.870 24.780 ;
        RECT 725.490 24.720 725.810 24.780 ;
        RECT 109.550 24.580 725.810 24.720 ;
        RECT 109.550 24.520 109.870 24.580 ;
        RECT 725.490 24.520 725.810 24.580 ;
      LAYER via ;
        RECT 647.780 2815.240 648.040 2815.500 ;
        RECT 1483.600 2815.240 1483.860 2815.500 ;
        RECT 647.780 594.020 648.040 594.280 ;
        RECT 724.600 594.020 724.860 594.280 ;
        RECT 724.600 572.260 724.860 572.520 ;
        RECT 725.520 572.260 725.780 572.520 ;
        RECT 725.060 338.000 725.320 338.260 ;
        RECT 725.520 338.000 725.780 338.260 ;
        RECT 723.680 324.060 723.940 324.320 ;
        RECT 725.060 324.060 725.320 324.320 ;
        RECT 723.680 276.120 723.940 276.380 ;
        RECT 724.600 276.120 724.860 276.380 ;
        RECT 724.140 234.300 724.400 234.560 ;
        RECT 725.060 234.300 725.320 234.560 ;
        RECT 722.760 227.500 723.020 227.760 ;
        RECT 724.140 227.500 724.400 227.760 ;
        RECT 722.760 179.560 723.020 179.820 ;
        RECT 723.680 179.560 723.940 179.820 ;
        RECT 723.680 138.080 723.940 138.340 ;
        RECT 724.600 138.080 724.860 138.340 ;
        RECT 724.600 110.200 724.860 110.460 ;
        RECT 725.520 110.200 725.780 110.460 ;
        RECT 109.580 24.520 109.840 24.780 ;
        RECT 725.520 24.520 725.780 24.780 ;
      LAYER met2 ;
        RECT 1483.590 2816.035 1483.870 2816.405 ;
        RECT 1483.660 2815.530 1483.800 2816.035 ;
        RECT 647.780 2815.210 648.040 2815.530 ;
        RECT 1483.600 2815.210 1483.860 2815.530 ;
        RECT 647.840 594.310 647.980 2815.210 ;
        RECT 726.210 600.850 726.490 604.000 ;
        RECT 724.660 600.710 726.490 600.850 ;
        RECT 724.660 594.310 724.800 600.710 ;
        RECT 726.210 600.000 726.490 600.710 ;
        RECT 647.780 593.990 648.040 594.310 ;
        RECT 724.600 593.990 724.860 594.310 ;
        RECT 724.660 572.550 724.800 593.990 ;
        RECT 724.600 572.230 724.860 572.550 ;
        RECT 725.520 572.230 725.780 572.550 ;
        RECT 725.580 500.210 725.720 572.230 ;
        RECT 725.120 500.070 725.720 500.210 ;
        RECT 725.120 448.530 725.260 500.070 ;
        RECT 725.120 448.390 725.720 448.530 ;
        RECT 725.580 338.290 725.720 448.390 ;
        RECT 725.060 337.970 725.320 338.290 ;
        RECT 725.520 337.970 725.780 338.290 ;
        RECT 725.120 324.350 725.260 337.970 ;
        RECT 723.680 324.030 723.940 324.350 ;
        RECT 725.060 324.030 725.320 324.350 ;
        RECT 723.740 276.410 723.880 324.030 ;
        RECT 723.680 276.090 723.940 276.410 ;
        RECT 724.600 276.090 724.860 276.410 ;
        RECT 724.660 235.010 724.800 276.090 ;
        RECT 724.660 234.870 725.260 235.010 ;
        RECT 725.120 234.590 725.260 234.870 ;
        RECT 724.140 234.270 724.400 234.590 ;
        RECT 725.060 234.270 725.320 234.590 ;
        RECT 724.200 227.790 724.340 234.270 ;
        RECT 722.760 227.470 723.020 227.790 ;
        RECT 724.140 227.470 724.400 227.790 ;
        RECT 722.820 179.850 722.960 227.470 ;
        RECT 722.760 179.530 723.020 179.850 ;
        RECT 723.680 179.530 723.940 179.850 ;
        RECT 723.740 138.370 723.880 179.530 ;
        RECT 723.680 138.050 723.940 138.370 ;
        RECT 724.600 138.050 724.860 138.370 ;
        RECT 724.660 110.490 724.800 138.050 ;
        RECT 724.600 110.170 724.860 110.490 ;
        RECT 725.520 110.170 725.780 110.490 ;
        RECT 725.580 24.810 725.720 110.170 ;
        RECT 109.580 24.490 109.840 24.810 ;
        RECT 725.520 24.490 725.780 24.810 ;
        RECT 109.640 2.400 109.780 24.490 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 1483.590 2816.080 1483.870 2816.360 ;
      LAYER met3 ;
        RECT 1500.000 2818.600 1504.000 2818.880 ;
        RECT 1499.910 2818.280 1504.000 2818.600 ;
        RECT 1483.565 2816.370 1483.895 2816.385 ;
        RECT 1499.910 2816.370 1500.210 2818.280 ;
        RECT 1483.565 2816.070 1500.210 2816.370 ;
        RECT 1483.565 2816.055 1483.895 2816.070 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 593.540 648.530 593.600 ;
        RECT 738.830 593.540 739.150 593.600 ;
        RECT 648.210 593.400 739.150 593.540 ;
        RECT 648.210 593.340 648.530 593.400 ;
        RECT 738.830 593.340 739.150 593.400 ;
        RECT 133.470 25.060 133.790 25.120 ;
        RECT 738.830 25.060 739.150 25.120 ;
        RECT 133.470 24.920 739.150 25.060 ;
        RECT 133.470 24.860 133.790 24.920 ;
        RECT 738.830 24.860 739.150 24.920 ;
      LAYER via ;
        RECT 648.240 593.340 648.500 593.600 ;
        RECT 738.860 593.340 739.120 593.600 ;
        RECT 133.500 24.860 133.760 25.120 ;
        RECT 738.860 24.860 739.120 25.120 ;
      LAYER met2 ;
        RECT 648.230 2911.915 648.510 2912.285 ;
        RECT 1747.630 2911.915 1747.910 2912.285 ;
        RECT 648.300 593.630 648.440 2911.915 ;
        RECT 1747.700 2900.055 1747.840 2911.915 ;
        RECT 1747.570 2896.055 1747.850 2900.055 ;
        RECT 738.630 600.000 738.910 604.000 ;
        RECT 738.690 598.810 738.830 600.000 ;
        RECT 738.690 598.670 739.060 598.810 ;
        RECT 738.920 593.630 739.060 598.670 ;
        RECT 648.240 593.310 648.500 593.630 ;
        RECT 738.860 593.310 739.120 593.630 ;
        RECT 738.920 25.150 739.060 593.310 ;
        RECT 133.500 24.830 133.760 25.150 ;
        RECT 738.860 24.830 739.120 25.150 ;
        RECT 133.560 2.400 133.700 24.830 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 648.230 2911.960 648.510 2912.240 ;
        RECT 1747.630 2911.960 1747.910 2912.240 ;
      LAYER met3 ;
        RECT 648.205 2912.250 648.535 2912.265 ;
        RECT 1747.605 2912.250 1747.935 2912.265 ;
        RECT 648.205 2911.950 1747.935 2912.250 ;
        RECT 648.205 2911.935 648.535 2911.950 ;
        RECT 1747.605 2911.935 1747.935 2911.950 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 655.110 593.880 655.430 593.940 ;
        RECT 745.270 593.880 745.590 593.940 ;
        RECT 655.110 593.740 745.590 593.880 ;
        RECT 655.110 593.680 655.430 593.740 ;
        RECT 745.270 593.680 745.590 593.740 ;
      LAYER via ;
        RECT 655.140 593.680 655.400 593.940 ;
        RECT 745.300 593.680 745.560 593.940 ;
      LAYER met2 ;
        RECT 655.130 2501.195 655.410 2501.565 ;
        RECT 655.200 593.970 655.340 2501.195 ;
        RECT 747.830 600.170 748.110 604.000 ;
        RECT 745.360 600.030 748.110 600.170 ;
        RECT 745.360 593.970 745.500 600.030 ;
        RECT 747.830 600.000 748.110 600.030 ;
        RECT 655.140 593.650 655.400 593.970 ;
        RECT 745.300 593.650 745.560 593.970 ;
        RECT 745.360 24.325 745.500 593.650 ;
        RECT 151.430 23.955 151.710 24.325 ;
        RECT 745.290 23.955 745.570 24.325 ;
        RECT 151.500 2.400 151.640 23.955 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 655.130 2501.240 655.410 2501.520 ;
        RECT 151.430 24.000 151.710 24.280 ;
        RECT 745.290 24.000 745.570 24.280 ;
      LAYER met3 ;
        RECT 1885.335 2863.480 1889.335 2863.760 ;
        RECT 1885.335 2863.160 1889.370 2863.480 ;
        RECT 1889.070 2860.570 1889.370 2863.160 ;
        RECT 1897.310 2860.570 1897.690 2860.580 ;
        RECT 1889.070 2860.270 1897.690 2860.570 ;
        RECT 1897.310 2860.260 1897.690 2860.270 ;
        RECT 655.105 2501.530 655.435 2501.545 ;
        RECT 1897.310 2501.530 1897.690 2501.540 ;
        RECT 655.105 2501.230 1897.690 2501.530 ;
        RECT 655.105 2501.215 655.435 2501.230 ;
        RECT 1897.310 2501.220 1897.690 2501.230 ;
        RECT 151.405 24.290 151.735 24.305 ;
        RECT 745.265 24.290 745.595 24.305 ;
        RECT 151.405 23.990 745.595 24.290 ;
        RECT 151.405 23.975 151.735 23.990 ;
        RECT 745.265 23.975 745.595 23.990 ;
      LAYER via3 ;
        RECT 1897.340 2860.260 1897.660 2860.580 ;
        RECT 1897.340 2501.220 1897.660 2501.540 ;
      LAYER met4 ;
        RECT 1897.335 2860.255 1897.665 2860.585 ;
        RECT 1897.350 2501.545 1897.650 2860.255 ;
        RECT 1897.335 2501.215 1897.665 2501.545 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 753.550 476.580 753.870 476.640 ;
        RECT 753.180 476.440 753.870 476.580 ;
        RECT 753.180 476.300 753.320 476.440 ;
        RECT 753.550 476.380 753.870 476.440 ;
        RECT 753.090 476.040 753.410 476.300 ;
        RECT 753.550 448.700 753.870 448.760 ;
        RECT 753.180 448.560 753.870 448.700 ;
        RECT 753.180 448.420 753.320 448.560 ;
        RECT 753.550 448.500 753.870 448.560 ;
        RECT 753.090 448.160 753.410 448.420 ;
        RECT 752.630 427.960 752.950 428.020 ;
        RECT 753.090 427.960 753.410 428.020 ;
        RECT 752.630 427.820 753.410 427.960 ;
        RECT 752.630 427.760 752.950 427.820 ;
        RECT 753.090 427.760 753.410 427.820 ;
        RECT 752.630 379.680 752.950 379.740 ;
        RECT 753.550 379.680 753.870 379.740 ;
        RECT 752.630 379.540 753.870 379.680 ;
        RECT 752.630 379.480 752.950 379.540 ;
        RECT 753.550 379.480 753.870 379.540 ;
        RECT 753.550 352.480 753.870 352.540 ;
        RECT 753.180 352.340 753.870 352.480 ;
        RECT 753.180 351.860 753.320 352.340 ;
        RECT 753.550 352.280 753.870 352.340 ;
        RECT 753.090 351.600 753.410 351.860 ;
        RECT 752.630 303.520 752.950 303.580 ;
        RECT 753.550 303.520 753.870 303.580 ;
        RECT 752.630 303.380 753.870 303.520 ;
        RECT 752.630 303.320 752.950 303.380 ;
        RECT 753.550 303.320 753.870 303.380 ;
        RECT 753.090 234.500 753.410 234.560 ;
        RECT 754.010 234.500 754.330 234.560 ;
        RECT 753.090 234.360 754.330 234.500 ;
        RECT 753.090 234.300 753.410 234.360 ;
        RECT 754.010 234.300 754.330 234.360 ;
        RECT 169.350 25.740 169.670 25.800 ;
        RECT 753.550 25.740 753.870 25.800 ;
        RECT 169.350 25.600 753.870 25.740 ;
        RECT 169.350 25.540 169.670 25.600 ;
        RECT 753.550 25.540 753.870 25.600 ;
      LAYER via ;
        RECT 753.580 476.380 753.840 476.640 ;
        RECT 753.120 476.040 753.380 476.300 ;
        RECT 753.580 448.500 753.840 448.760 ;
        RECT 753.120 448.160 753.380 448.420 ;
        RECT 752.660 427.760 752.920 428.020 ;
        RECT 753.120 427.760 753.380 428.020 ;
        RECT 752.660 379.480 752.920 379.740 ;
        RECT 753.580 379.480 753.840 379.740 ;
        RECT 753.580 352.280 753.840 352.540 ;
        RECT 753.120 351.600 753.380 351.860 ;
        RECT 752.660 303.320 752.920 303.580 ;
        RECT 753.580 303.320 753.840 303.580 ;
        RECT 753.120 234.300 753.380 234.560 ;
        RECT 754.040 234.300 754.300 234.560 ;
        RECT 169.380 25.540 169.640 25.800 ;
        RECT 753.580 25.540 753.840 25.800 ;
      LAYER met2 ;
        RECT 757.030 601.530 757.310 604.000 ;
        RECT 755.480 601.390 757.310 601.530 ;
        RECT 755.480 545.090 755.620 601.390 ;
        RECT 757.030 600.000 757.310 601.390 ;
        RECT 753.640 544.950 755.620 545.090 ;
        RECT 753.640 476.670 753.780 544.950 ;
        RECT 753.580 476.350 753.840 476.670 ;
        RECT 753.120 476.010 753.380 476.330 ;
        RECT 753.180 475.730 753.320 476.010 ;
        RECT 753.180 475.590 753.780 475.730 ;
        RECT 753.640 448.790 753.780 475.590 ;
        RECT 753.580 448.470 753.840 448.790 ;
        RECT 753.120 448.130 753.380 448.450 ;
        RECT 753.180 428.050 753.320 448.130 ;
        RECT 752.660 427.730 752.920 428.050 ;
        RECT 753.120 427.730 753.380 428.050 ;
        RECT 752.720 379.770 752.860 427.730 ;
        RECT 752.660 379.450 752.920 379.770 ;
        RECT 753.580 379.450 753.840 379.770 ;
        RECT 753.640 352.570 753.780 379.450 ;
        RECT 753.580 352.250 753.840 352.570 ;
        RECT 753.120 351.570 753.380 351.890 ;
        RECT 753.180 303.690 753.320 351.570 ;
        RECT 752.720 303.610 753.320 303.690 ;
        RECT 752.660 303.550 753.320 303.610 ;
        RECT 752.660 303.290 752.920 303.550 ;
        RECT 753.580 303.290 753.840 303.610 ;
        RECT 753.640 258.810 753.780 303.290 ;
        RECT 753.180 258.670 753.780 258.810 ;
        RECT 753.180 254.730 753.320 258.670 ;
        RECT 753.180 254.590 754.240 254.730 ;
        RECT 754.100 234.590 754.240 254.590 ;
        RECT 753.120 234.270 753.380 234.590 ;
        RECT 754.040 234.270 754.300 234.590 ;
        RECT 753.180 62.290 753.320 234.270 ;
        RECT 753.180 62.150 753.780 62.290 ;
        RECT 753.640 25.830 753.780 62.150 ;
        RECT 169.380 25.510 169.640 25.830 ;
        RECT 753.580 25.510 753.840 25.830 ;
        RECT 169.440 2.400 169.580 25.510 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 26.080 187.150 26.140 ;
        RECT 766.430 26.080 766.750 26.140 ;
        RECT 186.830 25.940 766.750 26.080 ;
        RECT 186.830 25.880 187.150 25.940 ;
        RECT 766.430 25.880 766.750 25.940 ;
      LAYER via ;
        RECT 186.860 25.880 187.120 26.140 ;
        RECT 766.460 25.880 766.720 26.140 ;
      LAYER met2 ;
        RECT 766.230 600.000 766.510 604.000 ;
        RECT 766.290 598.810 766.430 600.000 ;
        RECT 766.290 598.670 766.660 598.810 ;
        RECT 766.520 26.170 766.660 598.670 ;
        RECT 186.860 25.850 187.120 26.170 ;
        RECT 766.460 25.850 766.720 26.170 ;
        RECT 186.920 2.400 187.060 25.850 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 46.480 205.090 46.540 ;
        RECT 773.330 46.480 773.650 46.540 ;
        RECT 204.770 46.340 773.650 46.480 ;
        RECT 204.770 46.280 205.090 46.340 ;
        RECT 773.330 46.280 773.650 46.340 ;
      LAYER via ;
        RECT 204.800 46.280 205.060 46.540 ;
        RECT 773.360 46.280 773.620 46.540 ;
      LAYER met2 ;
        RECT 775.430 600.170 775.710 604.000 ;
        RECT 773.420 600.030 775.710 600.170 ;
        RECT 773.420 46.570 773.560 600.030 ;
        RECT 775.430 600.000 775.710 600.030 ;
        RECT 204.800 46.250 205.060 46.570 ;
        RECT 773.360 46.250 773.620 46.570 ;
        RECT 204.860 2.400 205.000 46.250 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.770 569.400 780.090 569.460 ;
        RECT 782.990 569.400 783.310 569.460 ;
        RECT 779.770 569.260 783.310 569.400 ;
        RECT 779.770 569.200 780.090 569.260 ;
        RECT 782.990 569.200 783.310 569.260 ;
        RECT 222.710 30.840 223.030 30.900 ;
        RECT 779.770 30.840 780.090 30.900 ;
        RECT 222.710 30.700 780.090 30.840 ;
        RECT 222.710 30.640 223.030 30.700 ;
        RECT 779.770 30.640 780.090 30.700 ;
      LAYER via ;
        RECT 779.800 569.200 780.060 569.460 ;
        RECT 783.020 569.200 783.280 569.460 ;
        RECT 222.740 30.640 223.000 30.900 ;
        RECT 779.800 30.640 780.060 30.900 ;
      LAYER met2 ;
        RECT 784.630 600.170 784.910 604.000 ;
        RECT 783.080 600.030 784.910 600.170 ;
        RECT 783.080 569.490 783.220 600.030 ;
        RECT 784.630 600.000 784.910 600.030 ;
        RECT 779.800 569.170 780.060 569.490 ;
        RECT 783.020 569.170 783.280 569.490 ;
        RECT 779.860 30.930 780.000 569.170 ;
        RECT 222.740 30.610 223.000 30.930 ;
        RECT 779.800 30.610 780.060 30.930 ;
        RECT 222.800 2.400 222.940 30.610 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 676.270 569.400 676.590 569.460 ;
        RECT 678.570 569.400 678.890 569.460 ;
        RECT 676.270 569.260 678.890 569.400 ;
        RECT 676.270 569.200 676.590 569.260 ;
        RECT 678.570 569.200 678.890 569.260 ;
        RECT 20.310 39.000 20.630 39.060 ;
        RECT 676.270 39.000 676.590 39.060 ;
        RECT 20.310 38.860 676.590 39.000 ;
        RECT 20.310 38.800 20.630 38.860 ;
        RECT 676.270 38.800 676.590 38.860 ;
      LAYER via ;
        RECT 676.300 569.200 676.560 569.460 ;
        RECT 678.600 569.200 678.860 569.460 ;
        RECT 20.340 38.800 20.600 39.060 ;
        RECT 676.300 38.800 676.560 39.060 ;
      LAYER met2 ;
        RECT 680.210 600.170 680.490 604.000 ;
        RECT 678.660 600.030 680.490 600.170 ;
        RECT 678.660 569.490 678.800 600.030 ;
        RECT 680.210 600.000 680.490 600.030 ;
        RECT 676.300 569.170 676.560 569.490 ;
        RECT 678.600 569.170 678.860 569.490 ;
        RECT 676.360 39.090 676.500 569.170 ;
        RECT 20.340 38.770 20.600 39.090 ;
        RECT 676.300 38.770 676.560 39.090 ;
        RECT 20.400 2.400 20.540 38.770 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.570 2504.340 517.890 2504.400 ;
        RECT 524.010 2504.340 524.330 2504.400 ;
        RECT 1904.470 2504.340 1904.790 2504.400 ;
        RECT 517.570 2504.200 1904.790 2504.340 ;
        RECT 517.570 2504.140 517.890 2504.200 ;
        RECT 524.010 2504.140 524.330 2504.200 ;
        RECT 1904.470 2504.140 1904.790 2504.200 ;
        RECT 350.590 2039.220 350.910 2039.280 ;
        RECT 524.010 2039.220 524.330 2039.280 ;
        RECT 2084.790 2039.220 2085.110 2039.280 ;
        RECT 350.590 2039.080 2085.110 2039.220 ;
        RECT 350.590 2039.020 350.910 2039.080 ;
        RECT 524.010 2039.020 524.330 2039.080 ;
        RECT 2084.790 2039.020 2085.110 2039.080 ;
        RECT 44.230 32.540 44.550 32.600 ;
        RECT 517.570 32.540 517.890 32.600 ;
        RECT 44.230 32.400 517.890 32.540 ;
        RECT 44.230 32.340 44.550 32.400 ;
        RECT 517.570 32.340 517.890 32.400 ;
      LAYER via ;
        RECT 517.600 2504.140 517.860 2504.400 ;
        RECT 524.040 2504.140 524.300 2504.400 ;
        RECT 1904.500 2504.140 1904.760 2504.400 ;
        RECT 350.620 2039.020 350.880 2039.280 ;
        RECT 524.040 2039.020 524.300 2039.280 ;
        RECT 2084.820 2039.020 2085.080 2039.280 ;
        RECT 44.260 32.340 44.520 32.600 ;
        RECT 517.600 32.340 517.860 32.600 ;
      LAYER met2 ;
        RECT 519.330 2600.730 519.610 2604.000 ;
        RECT 517.660 2600.590 519.610 2600.730 ;
        RECT 517.660 2504.430 517.800 2600.590 ;
        RECT 519.330 2600.000 519.610 2600.590 ;
        RECT 1903.570 2595.715 1903.850 2596.085 ;
        RECT 1903.640 2515.730 1903.780 2595.715 ;
        RECT 1903.640 2515.590 1904.700 2515.730 ;
        RECT 1904.560 2504.430 1904.700 2515.590 ;
        RECT 517.600 2504.110 517.860 2504.430 ;
        RECT 524.040 2504.110 524.300 2504.430 ;
        RECT 1904.500 2504.110 1904.760 2504.430 ;
        RECT 524.100 2039.310 524.240 2504.110 ;
        RECT 350.620 2038.990 350.880 2039.310 ;
        RECT 524.040 2038.990 524.300 2039.310 ;
        RECT 2084.820 2038.990 2085.080 2039.310 ;
        RECT 350.680 1851.485 350.820 2038.990 ;
        RECT 2084.880 1873.245 2085.020 2038.990 ;
        RECT 2084.810 1872.875 2085.090 1873.245 ;
        RECT 350.610 1851.115 350.890 1851.485 ;
        RECT 357.970 1851.115 358.250 1851.485 ;
        RECT 358.040 589.405 358.180 1851.115 ;
        RECT 692.630 600.170 692.910 604.000 ;
        RECT 691.080 600.030 692.910 600.170 ;
        RECT 458.710 591.075 458.990 591.445 ;
        RECT 458.780 590.085 458.920 591.075 ;
        RECT 458.710 589.715 458.990 590.085 ;
        RECT 517.130 589.970 517.410 590.085 ;
        RECT 517.130 589.830 517.800 589.970 ;
        RECT 517.130 589.715 517.410 589.830 ;
        RECT 357.970 589.035 358.250 589.405 ;
        RECT 517.660 588.045 517.800 589.830 ;
        RECT 691.080 589.405 691.220 600.030 ;
        RECT 692.630 600.000 692.910 600.030 ;
        RECT 619.710 589.035 619.990 589.405 ;
        RECT 675.830 589.035 676.110 589.405 ;
        RECT 691.010 589.035 691.290 589.405 ;
        RECT 619.780 588.045 619.920 589.035 ;
        RECT 517.590 587.675 517.870 588.045 ;
        RECT 619.710 587.675 619.990 588.045 ;
        RECT 517.660 32.630 517.800 587.675 ;
        RECT 675.900 587.365 676.040 589.035 ;
        RECT 675.830 586.995 676.110 587.365 ;
        RECT 44.260 32.310 44.520 32.630 ;
        RECT 517.600 32.310 517.860 32.630 ;
        RECT 44.320 2.400 44.460 32.310 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 1903.570 2595.760 1903.850 2596.040 ;
        RECT 2084.810 1872.920 2085.090 1873.200 ;
        RECT 350.610 1851.160 350.890 1851.440 ;
        RECT 357.970 1851.160 358.250 1851.440 ;
        RECT 458.710 591.120 458.990 591.400 ;
        RECT 458.710 589.760 458.990 590.040 ;
        RECT 517.130 589.760 517.410 590.040 ;
        RECT 357.970 589.080 358.250 589.360 ;
        RECT 619.710 589.080 619.990 589.360 ;
        RECT 675.830 589.080 676.110 589.360 ;
        RECT 691.010 589.080 691.290 589.360 ;
        RECT 517.590 587.720 517.870 588.000 ;
        RECT 619.710 587.720 619.990 588.000 ;
        RECT 675.830 587.040 676.110 587.320 ;
      LAYER met3 ;
        RECT 1885.335 2596.920 1889.335 2597.200 ;
        RECT 1885.335 2596.600 1889.370 2596.920 ;
        RECT 1889.070 2596.050 1889.370 2596.600 ;
        RECT 1903.545 2596.050 1903.875 2596.065 ;
        RECT 1889.070 2595.750 1903.875 2596.050 ;
        RECT 1903.545 2595.735 1903.875 2595.750 ;
        RECT 2084.785 1873.210 2085.115 1873.225 ;
        RECT 2075.830 1872.910 2085.115 1873.210 ;
        RECT 2075.830 1870.320 2076.130 1872.910 ;
        RECT 2084.785 1872.895 2085.115 1872.910 ;
        RECT 2072.375 1869.720 2076.375 1870.320 ;
        RECT 350.585 1851.450 350.915 1851.465 ;
        RECT 357.945 1851.450 358.275 1851.465 ;
        RECT 360.000 1851.450 364.000 1851.600 ;
        RECT 350.585 1851.150 364.000 1851.450 ;
        RECT 350.585 1851.135 350.915 1851.150 ;
        RECT 357.945 1851.135 358.275 1851.150 ;
        RECT 360.000 1851.000 364.000 1851.150 ;
        RECT 434.510 591.410 434.890 591.420 ;
        RECT 458.685 591.410 459.015 591.425 ;
        RECT 434.510 591.110 459.015 591.410 ;
        RECT 434.510 591.100 434.890 591.110 ;
        RECT 458.685 591.095 459.015 591.110 ;
        RECT 399.590 590.050 400.810 590.220 ;
        RECT 434.510 590.050 434.890 590.060 ;
        RECT 399.590 589.920 434.890 590.050 ;
        RECT 357.945 589.370 358.275 589.385 ;
        RECT 399.590 589.370 399.890 589.920 ;
        RECT 400.510 589.750 434.890 589.920 ;
        RECT 434.510 589.740 434.890 589.750 ;
        RECT 458.685 590.050 459.015 590.065 ;
        RECT 517.105 590.050 517.435 590.065 ;
        RECT 458.685 589.750 482.690 590.050 ;
        RECT 458.685 589.735 459.015 589.750 ;
        RECT 357.945 589.070 399.890 589.370 ;
        RECT 482.390 589.370 482.690 589.750 ;
        RECT 483.310 589.750 517.435 590.050 ;
        RECT 483.310 589.370 483.610 589.750 ;
        RECT 517.105 589.735 517.435 589.750 ;
        RECT 482.390 589.070 483.610 589.370 ;
        RECT 619.685 589.370 620.015 589.385 ;
        RECT 627.710 589.370 628.090 589.380 ;
        RECT 619.685 589.070 628.090 589.370 ;
        RECT 357.945 589.055 358.275 589.070 ;
        RECT 619.685 589.055 620.015 589.070 ;
        RECT 627.710 589.060 628.090 589.070 ;
        RECT 675.805 589.370 676.135 589.385 ;
        RECT 690.985 589.370 691.315 589.385 ;
        RECT 675.805 589.070 691.315 589.370 ;
        RECT 675.805 589.055 676.135 589.070 ;
        RECT 690.985 589.055 691.315 589.070 ;
        RECT 517.565 588.010 517.895 588.025 ;
        RECT 531.110 588.010 531.490 588.020 ;
        RECT 517.565 587.710 531.490 588.010 ;
        RECT 517.565 587.695 517.895 587.710 ;
        RECT 531.110 587.700 531.490 587.710 ;
        RECT 572.510 588.010 572.890 588.020 ;
        RECT 619.685 588.010 620.015 588.025 ;
        RECT 572.510 587.710 620.015 588.010 ;
        RECT 572.510 587.700 572.890 587.710 ;
        RECT 619.685 587.695 620.015 587.710 ;
        RECT 627.710 587.330 628.090 587.340 ;
        RECT 675.805 587.330 676.135 587.345 ;
        RECT 627.710 587.030 676.135 587.330 ;
        RECT 627.710 587.020 628.090 587.030 ;
        RECT 675.805 587.015 676.135 587.030 ;
        RECT 531.110 586.650 531.490 586.660 ;
        RECT 572.510 586.650 572.890 586.660 ;
        RECT 531.110 586.350 572.890 586.650 ;
        RECT 531.110 586.340 531.490 586.350 ;
        RECT 572.510 586.340 572.890 586.350 ;
      LAYER via3 ;
        RECT 434.540 591.100 434.860 591.420 ;
        RECT 434.540 589.740 434.860 590.060 ;
        RECT 627.740 589.060 628.060 589.380 ;
        RECT 531.140 587.700 531.460 588.020 ;
        RECT 572.540 587.700 572.860 588.020 ;
        RECT 627.740 587.020 628.060 587.340 ;
        RECT 531.140 586.340 531.460 586.660 ;
        RECT 572.540 586.340 572.860 586.660 ;
      LAYER met4 ;
        RECT 434.535 591.095 434.865 591.425 ;
        RECT 434.550 590.065 434.850 591.095 ;
        RECT 434.535 589.735 434.865 590.065 ;
        RECT 627.735 589.055 628.065 589.385 ;
        RECT 531.135 587.695 531.465 588.025 ;
        RECT 572.535 587.695 572.865 588.025 ;
        RECT 531.150 586.665 531.450 587.695 ;
        RECT 572.550 586.665 572.850 587.695 ;
        RECT 627.750 587.345 628.050 589.055 ;
        RECT 627.735 587.015 628.065 587.345 ;
        RECT 531.135 586.335 531.465 586.665 ;
        RECT 572.535 586.335 572.865 586.665 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1554.870 2898.060 1555.190 2898.120 ;
        RECT 1528.280 2897.920 1555.190 2898.060 ;
        RECT 945.370 2895.680 945.690 2895.740 ;
        RECT 980.330 2895.680 980.650 2895.740 ;
        RECT 945.370 2895.540 980.650 2895.680 ;
        RECT 945.370 2895.480 945.690 2895.540 ;
        RECT 980.330 2895.480 980.650 2895.540 ;
        RECT 1495.530 2895.680 1495.850 2895.740 ;
        RECT 1495.530 2895.540 1503.120 2895.680 ;
        RECT 1495.530 2895.480 1495.850 2895.540 ;
        RECT 1502.980 2895.340 1503.120 2895.540 ;
        RECT 1528.280 2895.340 1528.420 2897.920 ;
        RECT 1554.870 2897.860 1555.190 2897.920 ;
        RECT 1502.980 2895.200 1528.420 2895.340 ;
        RECT 881.890 2895.000 882.210 2895.060 ;
        RECT 945.370 2895.000 945.690 2895.060 ;
        RECT 881.890 2894.860 945.690 2895.000 ;
        RECT 881.890 2894.800 882.210 2894.860 ;
        RECT 945.370 2894.800 945.690 2894.860 ;
        RECT 1186.870 2894.660 1187.190 2894.720 ;
        RECT 1234.710 2894.660 1235.030 2894.720 ;
        RECT 1186.870 2894.520 1235.030 2894.660 ;
        RECT 1186.870 2894.460 1187.190 2894.520 ;
        RECT 1234.710 2894.460 1235.030 2894.520 ;
        RECT 651.890 2894.320 652.210 2894.380 ;
        RECT 786.670 2894.320 786.990 2894.380 ;
        RECT 1249.430 2894.320 1249.750 2894.380 ;
        RECT 651.890 2894.180 691.220 2894.320 ;
        RECT 651.890 2894.120 652.210 2894.180 ;
        RECT 691.080 2893.980 691.220 2894.180 ;
        RECT 786.670 2894.180 834.740 2894.320 ;
        RECT 786.670 2894.120 786.990 2894.180 ;
        RECT 834.600 2893.980 834.740 2894.180 ;
        RECT 1249.430 2894.180 1317.740 2894.320 ;
        RECT 1249.430 2894.120 1249.750 2894.180 ;
        RECT 980.330 2893.980 980.650 2894.040 ;
        RECT 1000.570 2893.980 1000.890 2894.040 ;
        RECT 1076.930 2893.980 1077.250 2894.040 ;
        RECT 1097.170 2893.980 1097.490 2894.040 ;
        RECT 1173.530 2893.980 1173.850 2894.040 ;
        RECT 1186.870 2893.980 1187.190 2894.040 ;
        RECT 691.080 2893.840 762.520 2893.980 ;
        RECT 834.600 2893.840 836.120 2893.980 ;
        RECT 762.380 2893.640 762.520 2893.840 ;
        RECT 835.980 2893.640 836.120 2893.840 ;
        RECT 980.330 2893.840 993.900 2893.980 ;
        RECT 980.330 2893.780 980.650 2893.840 ;
        RECT 881.890 2893.640 882.210 2893.700 ;
        RECT 762.380 2893.500 786.440 2893.640 ;
        RECT 835.980 2893.500 882.210 2893.640 ;
        RECT 993.760 2893.640 993.900 2893.840 ;
        RECT 1000.570 2893.840 1028.860 2893.980 ;
        RECT 1000.570 2893.780 1000.890 2893.840 ;
        RECT 1000.110 2893.640 1000.430 2893.700 ;
        RECT 993.760 2893.500 1000.430 2893.640 ;
        RECT 1028.720 2893.640 1028.860 2893.840 ;
        RECT 1076.930 2893.840 1090.500 2893.980 ;
        RECT 1076.930 2893.780 1077.250 2893.840 ;
        RECT 1090.360 2893.640 1090.500 2893.840 ;
        RECT 1097.170 2893.840 1125.460 2893.980 ;
        RECT 1097.170 2893.780 1097.490 2893.840 ;
        RECT 1096.710 2893.640 1097.030 2893.700 ;
        RECT 1028.720 2893.500 1076.240 2893.640 ;
        RECT 1090.360 2893.500 1097.030 2893.640 ;
        RECT 1125.320 2893.640 1125.460 2893.840 ;
        RECT 1173.530 2893.840 1187.190 2893.980 ;
        RECT 1317.600 2893.980 1317.740 2894.180 ;
        RECT 1317.600 2893.840 1319.120 2893.980 ;
        RECT 1173.530 2893.780 1173.850 2893.840 ;
        RECT 1186.870 2893.780 1187.190 2893.840 ;
        RECT 1318.980 2893.640 1319.120 2893.840 ;
        RECT 1439.870 2893.640 1440.190 2893.700 ;
        RECT 1495.530 2893.640 1495.850 2893.700 ;
        RECT 1125.320 2893.500 1172.840 2893.640 ;
        RECT 1318.980 2893.500 1366.040 2893.640 ;
        RECT 786.300 2893.300 786.440 2893.500 ;
        RECT 881.890 2893.440 882.210 2893.500 ;
        RECT 1000.110 2893.440 1000.430 2893.500 ;
        RECT 1076.100 2893.360 1076.240 2893.500 ;
        RECT 1096.710 2893.440 1097.030 2893.500 ;
        RECT 1172.700 2893.360 1172.840 2893.500 ;
        RECT 786.670 2893.300 786.990 2893.360 ;
        RECT 786.300 2893.160 786.990 2893.300 ;
        RECT 786.670 2893.100 786.990 2893.160 ;
        RECT 1076.010 2893.100 1076.330 2893.360 ;
        RECT 1172.610 2893.100 1172.930 2893.360 ;
        RECT 1234.710 2893.300 1235.030 2893.360 ;
        RECT 1249.430 2893.300 1249.750 2893.360 ;
        RECT 1234.710 2893.160 1249.750 2893.300 ;
        RECT 1365.900 2893.300 1366.040 2893.500 ;
        RECT 1439.870 2893.500 1495.850 2893.640 ;
        RECT 1439.870 2893.440 1440.190 2893.500 ;
        RECT 1495.530 2893.440 1495.850 2893.500 ;
        RECT 1400.770 2893.300 1401.090 2893.360 ;
        RECT 1365.900 2893.160 1401.090 2893.300 ;
        RECT 1234.710 2893.100 1235.030 2893.160 ;
        RECT 1249.430 2893.100 1249.750 2893.160 ;
        RECT 1400.770 2893.100 1401.090 2893.160 ;
        RECT 446.730 2594.440 447.050 2594.500 ;
        RECT 649.130 2594.440 649.450 2594.500 ;
        RECT 651.890 2594.440 652.210 2594.500 ;
        RECT 446.730 2594.300 652.210 2594.440 ;
        RECT 446.730 2594.240 447.050 2594.300 ;
        RECT 649.130 2594.240 649.450 2594.300 ;
        RECT 651.890 2594.240 652.210 2594.300 ;
        RECT 644.990 1756.000 645.310 1756.060 ;
        RECT 649.130 1756.000 649.450 1756.060 ;
        RECT 651.890 1756.000 652.210 1756.060 ;
        RECT 644.990 1755.860 652.210 1756.000 ;
        RECT 644.990 1755.800 645.310 1755.860 ;
        RECT 649.130 1755.800 649.450 1755.860 ;
        RECT 651.890 1755.800 652.210 1755.860 ;
        RECT 651.890 1703.300 652.210 1703.360 ;
        RECT 1908.150 1703.300 1908.470 1703.360 ;
        RECT 651.890 1703.160 1908.470 1703.300 ;
        RECT 651.890 1703.100 652.210 1703.160 ;
        RECT 1908.150 1703.100 1908.470 1703.160 ;
        RECT 651.890 1642.440 652.210 1642.500 ;
        RECT 654.190 1642.440 654.510 1642.500 ;
        RECT 651.890 1642.300 654.510 1642.440 ;
        RECT 651.890 1642.240 652.210 1642.300 ;
        RECT 654.190 1642.240 654.510 1642.300 ;
        RECT 652.810 1607.760 653.130 1607.820 ;
        RECT 654.190 1607.760 654.510 1607.820 ;
        RECT 652.810 1607.620 654.510 1607.760 ;
        RECT 652.810 1607.560 653.130 1607.620 ;
        RECT 654.190 1607.560 654.510 1607.620 ;
        RECT 652.810 1559.480 653.130 1559.540 ;
        RECT 654.190 1559.480 654.510 1559.540 ;
        RECT 652.810 1559.340 654.510 1559.480 ;
        RECT 652.810 1559.280 653.130 1559.340 ;
        RECT 654.190 1559.280 654.510 1559.340 ;
        RECT 652.810 1510.860 653.130 1510.920 ;
        RECT 654.190 1510.860 654.510 1510.920 ;
        RECT 652.810 1510.720 654.510 1510.860 ;
        RECT 652.810 1510.660 653.130 1510.720 ;
        RECT 654.190 1510.660 654.510 1510.720 ;
        RECT 652.350 1497.260 652.670 1497.320 ;
        RECT 652.810 1497.260 653.130 1497.320 ;
        RECT 652.350 1497.120 653.130 1497.260 ;
        RECT 652.350 1497.060 652.670 1497.120 ;
        RECT 652.810 1497.060 653.130 1497.120 ;
        RECT 652.350 1449.320 652.670 1449.380 ;
        RECT 654.190 1449.320 654.510 1449.380 ;
        RECT 652.350 1449.180 654.510 1449.320 ;
        RECT 652.350 1449.120 652.670 1449.180 ;
        RECT 654.190 1449.120 654.510 1449.180 ;
        RECT 652.810 1414.300 653.130 1414.360 ;
        RECT 654.190 1414.300 654.510 1414.360 ;
        RECT 652.810 1414.160 654.510 1414.300 ;
        RECT 652.810 1414.100 653.130 1414.160 ;
        RECT 654.190 1414.100 654.510 1414.160 ;
        RECT 652.350 1400.700 652.670 1400.760 ;
        RECT 652.810 1400.700 653.130 1400.760 ;
        RECT 652.350 1400.560 653.130 1400.700 ;
        RECT 652.350 1400.500 652.670 1400.560 ;
        RECT 652.810 1400.500 653.130 1400.560 ;
        RECT 652.350 1352.760 652.670 1352.820 ;
        RECT 654.190 1352.760 654.510 1352.820 ;
        RECT 652.350 1352.620 654.510 1352.760 ;
        RECT 652.350 1352.560 652.670 1352.620 ;
        RECT 654.190 1352.560 654.510 1352.620 ;
        RECT 652.810 1317.740 653.130 1317.800 ;
        RECT 654.190 1317.740 654.510 1317.800 ;
        RECT 652.810 1317.600 654.510 1317.740 ;
        RECT 652.810 1317.540 653.130 1317.600 ;
        RECT 654.190 1317.540 654.510 1317.600 ;
        RECT 652.350 1304.140 652.670 1304.200 ;
        RECT 652.810 1304.140 653.130 1304.200 ;
        RECT 652.350 1304.000 653.130 1304.140 ;
        RECT 652.350 1303.940 652.670 1304.000 ;
        RECT 652.810 1303.940 653.130 1304.000 ;
        RECT 652.810 1221.180 653.130 1221.240 ;
        RECT 654.190 1221.180 654.510 1221.240 ;
        RECT 652.810 1221.040 654.510 1221.180 ;
        RECT 652.810 1220.980 653.130 1221.040 ;
        RECT 654.190 1220.980 654.510 1221.040 ;
        RECT 652.810 1159.300 653.130 1159.360 ;
        RECT 654.190 1159.300 654.510 1159.360 ;
        RECT 652.810 1159.160 654.510 1159.300 ;
        RECT 652.810 1159.100 653.130 1159.160 ;
        RECT 654.190 1159.100 654.510 1159.160 ;
        RECT 652.810 1124.620 653.130 1124.680 ;
        RECT 654.190 1124.620 654.510 1124.680 ;
        RECT 652.810 1124.480 654.510 1124.620 ;
        RECT 652.810 1124.420 653.130 1124.480 ;
        RECT 654.190 1124.420 654.510 1124.480 ;
        RECT 652.810 1062.740 653.130 1062.800 ;
        RECT 654.190 1062.740 654.510 1062.800 ;
        RECT 652.810 1062.600 654.510 1062.740 ;
        RECT 652.810 1062.540 653.130 1062.600 ;
        RECT 654.190 1062.540 654.510 1062.600 ;
        RECT 652.350 1028.060 652.670 1028.120 ;
        RECT 654.190 1028.060 654.510 1028.120 ;
        RECT 652.350 1027.920 654.510 1028.060 ;
        RECT 652.350 1027.860 652.670 1027.920 ;
        RECT 654.190 1027.860 654.510 1027.920 ;
        RECT 652.350 966.180 652.670 966.240 ;
        RECT 654.190 966.180 654.510 966.240 ;
        RECT 652.350 966.040 654.510 966.180 ;
        RECT 652.350 965.980 652.670 966.040 ;
        RECT 654.190 965.980 654.510 966.040 ;
        RECT 654.190 931.500 654.510 931.560 ;
        RECT 652.900 931.360 654.510 931.500 ;
        RECT 651.890 931.160 652.210 931.220 ;
        RECT 652.900 931.160 653.040 931.360 ;
        RECT 654.190 931.300 654.510 931.360 ;
        RECT 651.890 931.020 653.040 931.160 ;
        RECT 651.890 930.960 652.210 931.020 ;
        RECT 651.890 869.620 652.210 869.680 ;
        RECT 654.190 869.620 654.510 869.680 ;
        RECT 651.890 869.480 654.510 869.620 ;
        RECT 651.890 869.420 652.210 869.480 ;
        RECT 654.190 869.420 654.510 869.480 ;
        RECT 652.350 834.940 652.670 835.000 ;
        RECT 654.190 834.940 654.510 835.000 ;
        RECT 652.350 834.800 654.510 834.940 ;
        RECT 652.350 834.740 652.670 834.800 ;
        RECT 654.190 834.740 654.510 834.800 ;
        RECT 652.350 737.700 652.670 737.760 ;
        RECT 654.190 737.700 654.510 737.760 ;
        RECT 652.350 737.560 654.510 737.700 ;
        RECT 652.350 737.500 652.670 737.560 ;
        RECT 654.190 737.500 654.510 737.560 ;
        RECT 653.270 641.480 653.590 641.540 ;
        RECT 654.190 641.480 654.510 641.540 ;
        RECT 653.270 641.340 654.510 641.480 ;
        RECT 653.270 641.280 653.590 641.340 ;
        RECT 654.190 641.280 654.510 641.340 ;
        RECT 651.890 627.880 652.210 627.940 ;
        RECT 653.270 627.880 653.590 627.940 ;
        RECT 651.890 627.740 653.590 627.880 ;
        RECT 651.890 627.680 652.210 627.740 ;
        RECT 653.270 627.680 653.590 627.740 ;
        RECT 651.890 588.100 652.210 588.160 ;
        RECT 678.110 588.100 678.430 588.160 ;
        RECT 651.890 587.960 678.430 588.100 ;
        RECT 651.890 587.900 652.210 587.960 ;
        RECT 678.110 587.900 678.430 587.960 ;
        RECT 679.490 588.100 679.810 588.160 ;
        RECT 794.950 588.100 795.270 588.160 ;
        RECT 679.490 587.960 795.270 588.100 ;
        RECT 679.490 587.900 679.810 587.960 ;
        RECT 794.950 587.900 795.270 587.960 ;
        RECT 246.630 22.340 246.950 22.400 ;
        RECT 651.890 22.340 652.210 22.400 ;
        RECT 246.630 22.200 652.210 22.340 ;
        RECT 246.630 22.140 246.950 22.200 ;
        RECT 651.890 22.140 652.210 22.200 ;
      LAYER via ;
        RECT 945.400 2895.480 945.660 2895.740 ;
        RECT 980.360 2895.480 980.620 2895.740 ;
        RECT 1495.560 2895.480 1495.820 2895.740 ;
        RECT 1554.900 2897.860 1555.160 2898.120 ;
        RECT 881.920 2894.800 882.180 2895.060 ;
        RECT 945.400 2894.800 945.660 2895.060 ;
        RECT 1186.900 2894.460 1187.160 2894.720 ;
        RECT 1234.740 2894.460 1235.000 2894.720 ;
        RECT 651.920 2894.120 652.180 2894.380 ;
        RECT 786.700 2894.120 786.960 2894.380 ;
        RECT 1249.460 2894.120 1249.720 2894.380 ;
        RECT 980.360 2893.780 980.620 2894.040 ;
        RECT 881.920 2893.440 882.180 2893.700 ;
        RECT 1000.600 2893.780 1000.860 2894.040 ;
        RECT 1000.140 2893.440 1000.400 2893.700 ;
        RECT 1076.960 2893.780 1077.220 2894.040 ;
        RECT 1097.200 2893.780 1097.460 2894.040 ;
        RECT 1096.740 2893.440 1097.000 2893.700 ;
        RECT 1173.560 2893.780 1173.820 2894.040 ;
        RECT 1186.900 2893.780 1187.160 2894.040 ;
        RECT 786.700 2893.100 786.960 2893.360 ;
        RECT 1076.040 2893.100 1076.300 2893.360 ;
        RECT 1172.640 2893.100 1172.900 2893.360 ;
        RECT 1234.740 2893.100 1235.000 2893.360 ;
        RECT 1249.460 2893.100 1249.720 2893.360 ;
        RECT 1439.900 2893.440 1440.160 2893.700 ;
        RECT 1495.560 2893.440 1495.820 2893.700 ;
        RECT 1400.800 2893.100 1401.060 2893.360 ;
        RECT 446.760 2594.240 447.020 2594.500 ;
        RECT 649.160 2594.240 649.420 2594.500 ;
        RECT 651.920 2594.240 652.180 2594.500 ;
        RECT 645.020 1755.800 645.280 1756.060 ;
        RECT 649.160 1755.800 649.420 1756.060 ;
        RECT 651.920 1755.800 652.180 1756.060 ;
        RECT 651.920 1703.100 652.180 1703.360 ;
        RECT 1908.180 1703.100 1908.440 1703.360 ;
        RECT 651.920 1642.240 652.180 1642.500 ;
        RECT 654.220 1642.240 654.480 1642.500 ;
        RECT 652.840 1607.560 653.100 1607.820 ;
        RECT 654.220 1607.560 654.480 1607.820 ;
        RECT 652.840 1559.280 653.100 1559.540 ;
        RECT 654.220 1559.280 654.480 1559.540 ;
        RECT 652.840 1510.660 653.100 1510.920 ;
        RECT 654.220 1510.660 654.480 1510.920 ;
        RECT 652.380 1497.060 652.640 1497.320 ;
        RECT 652.840 1497.060 653.100 1497.320 ;
        RECT 652.380 1449.120 652.640 1449.380 ;
        RECT 654.220 1449.120 654.480 1449.380 ;
        RECT 652.840 1414.100 653.100 1414.360 ;
        RECT 654.220 1414.100 654.480 1414.360 ;
        RECT 652.380 1400.500 652.640 1400.760 ;
        RECT 652.840 1400.500 653.100 1400.760 ;
        RECT 652.380 1352.560 652.640 1352.820 ;
        RECT 654.220 1352.560 654.480 1352.820 ;
        RECT 652.840 1317.540 653.100 1317.800 ;
        RECT 654.220 1317.540 654.480 1317.800 ;
        RECT 652.380 1303.940 652.640 1304.200 ;
        RECT 652.840 1303.940 653.100 1304.200 ;
        RECT 652.840 1220.980 653.100 1221.240 ;
        RECT 654.220 1220.980 654.480 1221.240 ;
        RECT 652.840 1159.100 653.100 1159.360 ;
        RECT 654.220 1159.100 654.480 1159.360 ;
        RECT 652.840 1124.420 653.100 1124.680 ;
        RECT 654.220 1124.420 654.480 1124.680 ;
        RECT 652.840 1062.540 653.100 1062.800 ;
        RECT 654.220 1062.540 654.480 1062.800 ;
        RECT 652.380 1027.860 652.640 1028.120 ;
        RECT 654.220 1027.860 654.480 1028.120 ;
        RECT 652.380 965.980 652.640 966.240 ;
        RECT 654.220 965.980 654.480 966.240 ;
        RECT 651.920 930.960 652.180 931.220 ;
        RECT 654.220 931.300 654.480 931.560 ;
        RECT 651.920 869.420 652.180 869.680 ;
        RECT 654.220 869.420 654.480 869.680 ;
        RECT 652.380 834.740 652.640 835.000 ;
        RECT 654.220 834.740 654.480 835.000 ;
        RECT 652.380 737.500 652.640 737.760 ;
        RECT 654.220 737.500 654.480 737.760 ;
        RECT 653.300 641.280 653.560 641.540 ;
        RECT 654.220 641.280 654.480 641.540 ;
        RECT 651.920 627.680 652.180 627.940 ;
        RECT 653.300 627.680 653.560 627.940 ;
        RECT 651.920 587.900 652.180 588.160 ;
        RECT 678.140 587.900 678.400 588.160 ;
        RECT 679.520 587.900 679.780 588.160 ;
        RECT 794.980 587.900 795.240 588.160 ;
        RECT 246.660 22.140 246.920 22.400 ;
        RECT 651.920 22.140 652.180 22.400 ;
      LAYER met2 ;
        RECT 1554.900 2897.890 1555.160 2898.150 ;
        RECT 1556.210 2897.890 1556.490 2900.055 ;
        RECT 1554.900 2897.830 1556.490 2897.890 ;
        RECT 1554.960 2897.750 1556.490 2897.830 ;
        RECT 1556.210 2896.055 1556.490 2897.750 ;
        RECT 945.400 2895.450 945.660 2895.770 ;
        RECT 980.360 2895.450 980.620 2895.770 ;
        RECT 1495.560 2895.450 1495.820 2895.770 ;
        RECT 945.460 2895.090 945.600 2895.450 ;
        RECT 881.920 2894.770 882.180 2895.090 ;
        RECT 945.400 2894.770 945.660 2895.090 ;
        RECT 651.920 2894.090 652.180 2894.410 ;
        RECT 786.700 2894.090 786.960 2894.410 ;
        RECT 446.650 2600.660 446.930 2604.000 ;
        RECT 446.650 2600.000 446.960 2600.660 ;
        RECT 446.820 2594.530 446.960 2600.000 ;
        RECT 651.980 2594.530 652.120 2894.090 ;
        RECT 786.760 2893.390 786.900 2894.090 ;
        RECT 881.980 2893.730 882.120 2894.770 ;
        RECT 980.420 2894.070 980.560 2895.450 ;
        RECT 1186.900 2894.430 1187.160 2894.750 ;
        RECT 1234.740 2894.430 1235.000 2894.750 ;
        RECT 1186.960 2894.070 1187.100 2894.430 ;
        RECT 980.360 2893.750 980.620 2894.070 ;
        RECT 1000.600 2893.810 1000.860 2894.070 ;
        RECT 1000.200 2893.750 1000.860 2893.810 ;
        RECT 1076.960 2893.750 1077.220 2894.070 ;
        RECT 1097.200 2893.810 1097.460 2894.070 ;
        RECT 1096.800 2893.750 1097.460 2893.810 ;
        RECT 1173.560 2893.750 1173.820 2894.070 ;
        RECT 1186.900 2893.750 1187.160 2894.070 ;
        RECT 1000.200 2893.730 1000.800 2893.750 ;
        RECT 881.920 2893.410 882.180 2893.730 ;
        RECT 1000.140 2893.670 1000.800 2893.730 ;
        RECT 1000.140 2893.410 1000.400 2893.670 ;
        RECT 786.700 2893.070 786.960 2893.390 ;
        RECT 1076.040 2893.130 1076.300 2893.390 ;
        RECT 1077.020 2893.130 1077.160 2893.750 ;
        RECT 1096.800 2893.730 1097.400 2893.750 ;
        RECT 1096.740 2893.670 1097.400 2893.730 ;
        RECT 1096.740 2893.410 1097.000 2893.670 ;
        RECT 1076.040 2893.070 1077.160 2893.130 ;
        RECT 1172.640 2893.130 1172.900 2893.390 ;
        RECT 1173.620 2893.130 1173.760 2893.750 ;
        RECT 1234.800 2893.390 1234.940 2894.430 ;
        RECT 1249.460 2894.090 1249.720 2894.410 ;
        RECT 1249.520 2893.390 1249.660 2894.090 ;
        RECT 1495.620 2893.730 1495.760 2895.450 ;
        RECT 1439.900 2893.410 1440.160 2893.730 ;
        RECT 1495.560 2893.410 1495.820 2893.730 ;
        RECT 1172.640 2893.070 1173.760 2893.130 ;
        RECT 1234.740 2893.070 1235.000 2893.390 ;
        RECT 1249.460 2893.070 1249.720 2893.390 ;
        RECT 1400.800 2893.245 1401.060 2893.390 ;
        RECT 1439.960 2893.245 1440.100 2893.410 ;
        RECT 1076.100 2892.990 1077.160 2893.070 ;
        RECT 1172.700 2892.990 1173.760 2893.070 ;
        RECT 1400.790 2892.875 1401.070 2893.245 ;
        RECT 1439.890 2892.875 1440.170 2893.245 ;
        RECT 446.760 2594.210 447.020 2594.530 ;
        RECT 649.160 2594.210 649.420 2594.530 ;
        RECT 651.920 2594.210 652.180 2594.530 ;
        RECT 649.220 1756.090 649.360 2594.210 ;
        RECT 1908.170 1836.835 1908.450 1837.205 ;
        RECT 645.020 1755.770 645.280 1756.090 ;
        RECT 649.160 1755.770 649.420 1756.090 ;
        RECT 651.920 1755.770 652.180 1756.090 ;
        RECT 645.080 1754.925 645.220 1755.770 ;
        RECT 645.010 1754.555 645.290 1754.925 ;
        RECT 651.980 1703.390 652.120 1755.770 ;
        RECT 1908.240 1703.390 1908.380 1836.835 ;
        RECT 651.920 1703.070 652.180 1703.390 ;
        RECT 1908.180 1703.070 1908.440 1703.390 ;
        RECT 651.980 1642.530 652.120 1703.070 ;
        RECT 651.920 1642.210 652.180 1642.530 ;
        RECT 654.220 1642.210 654.480 1642.530 ;
        RECT 654.280 1607.850 654.420 1642.210 ;
        RECT 652.840 1607.530 653.100 1607.850 ;
        RECT 654.220 1607.530 654.480 1607.850 ;
        RECT 652.900 1559.570 653.040 1607.530 ;
        RECT 652.840 1559.250 653.100 1559.570 ;
        RECT 654.220 1559.250 654.480 1559.570 ;
        RECT 654.280 1510.950 654.420 1559.250 ;
        RECT 652.840 1510.630 653.100 1510.950 ;
        RECT 654.220 1510.630 654.480 1510.950 ;
        RECT 652.900 1497.350 653.040 1510.630 ;
        RECT 652.380 1497.030 652.640 1497.350 ;
        RECT 652.840 1497.030 653.100 1497.350 ;
        RECT 652.440 1449.410 652.580 1497.030 ;
        RECT 652.380 1449.090 652.640 1449.410 ;
        RECT 654.220 1449.090 654.480 1449.410 ;
        RECT 654.280 1414.390 654.420 1449.090 ;
        RECT 652.840 1414.070 653.100 1414.390 ;
        RECT 654.220 1414.070 654.480 1414.390 ;
        RECT 652.900 1400.790 653.040 1414.070 ;
        RECT 652.380 1400.470 652.640 1400.790 ;
        RECT 652.840 1400.470 653.100 1400.790 ;
        RECT 652.440 1352.850 652.580 1400.470 ;
        RECT 652.380 1352.530 652.640 1352.850 ;
        RECT 654.220 1352.530 654.480 1352.850 ;
        RECT 654.280 1317.830 654.420 1352.530 ;
        RECT 652.840 1317.510 653.100 1317.830 ;
        RECT 654.220 1317.510 654.480 1317.830 ;
        RECT 652.900 1304.230 653.040 1317.510 ;
        RECT 652.380 1303.910 652.640 1304.230 ;
        RECT 652.840 1303.910 653.100 1304.230 ;
        RECT 652.440 1256.485 652.580 1303.910 ;
        RECT 652.370 1256.115 652.650 1256.485 ;
        RECT 654.210 1256.115 654.490 1256.485 ;
        RECT 654.280 1221.270 654.420 1256.115 ;
        RECT 652.840 1220.950 653.100 1221.270 ;
        RECT 654.220 1220.950 654.480 1221.270 ;
        RECT 652.900 1159.390 653.040 1220.950 ;
        RECT 652.840 1159.070 653.100 1159.390 ;
        RECT 654.220 1159.070 654.480 1159.390 ;
        RECT 654.280 1124.710 654.420 1159.070 ;
        RECT 652.840 1124.390 653.100 1124.710 ;
        RECT 654.220 1124.390 654.480 1124.710 ;
        RECT 652.900 1062.830 653.040 1124.390 ;
        RECT 652.840 1062.510 653.100 1062.830 ;
        RECT 654.220 1062.510 654.480 1062.830 ;
        RECT 654.280 1028.150 654.420 1062.510 ;
        RECT 652.380 1027.830 652.640 1028.150 ;
        RECT 654.220 1027.830 654.480 1028.150 ;
        RECT 652.440 966.270 652.580 1027.830 ;
        RECT 652.380 965.950 652.640 966.270 ;
        RECT 654.220 965.950 654.480 966.270 ;
        RECT 654.280 931.590 654.420 965.950 ;
        RECT 654.220 931.270 654.480 931.590 ;
        RECT 651.920 930.930 652.180 931.250 ;
        RECT 651.980 869.710 652.120 930.930 ;
        RECT 651.920 869.390 652.180 869.710 ;
        RECT 654.220 869.390 654.480 869.710 ;
        RECT 654.280 835.030 654.420 869.390 ;
        RECT 652.380 834.710 652.640 835.030 ;
        RECT 654.220 834.710 654.480 835.030 ;
        RECT 652.440 773.005 652.580 834.710 ;
        RECT 652.370 772.635 652.650 773.005 ;
        RECT 654.210 772.635 654.490 773.005 ;
        RECT 654.280 737.790 654.420 772.635 ;
        RECT 652.380 737.470 652.640 737.790 ;
        RECT 654.220 737.470 654.480 737.790 ;
        RECT 652.440 676.445 652.580 737.470 ;
        RECT 652.370 676.075 652.650 676.445 ;
        RECT 654.210 676.075 654.490 676.445 ;
        RECT 654.280 641.570 654.420 676.075 ;
        RECT 653.300 641.250 653.560 641.570 ;
        RECT 654.220 641.250 654.480 641.570 ;
        RECT 653.360 627.970 653.500 641.250 ;
        RECT 651.920 627.650 652.180 627.970 ;
        RECT 653.300 627.650 653.560 627.970 ;
        RECT 651.980 588.190 652.120 627.650 ;
        RECT 796.590 600.170 796.870 604.000 ;
        RECT 795.040 600.030 796.870 600.170 ;
        RECT 795.040 588.190 795.180 600.030 ;
        RECT 796.590 600.000 796.870 600.030 ;
        RECT 651.920 587.870 652.180 588.190 ;
        RECT 678.140 587.870 678.400 588.190 ;
        RECT 679.520 587.870 679.780 588.190 ;
        RECT 794.980 587.870 795.240 588.190 ;
        RECT 651.980 22.430 652.120 587.870 ;
        RECT 678.200 587.365 678.340 587.870 ;
        RECT 679.580 587.365 679.720 587.870 ;
        RECT 678.130 586.995 678.410 587.365 ;
        RECT 679.510 586.995 679.790 587.365 ;
        RECT 246.660 22.110 246.920 22.430 ;
        RECT 651.920 22.110 652.180 22.430 ;
        RECT 246.720 2.400 246.860 22.110 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 1400.790 2892.920 1401.070 2893.200 ;
        RECT 1439.890 2892.920 1440.170 2893.200 ;
        RECT 1908.170 1836.880 1908.450 1837.160 ;
        RECT 645.010 1754.600 645.290 1754.880 ;
        RECT 652.370 1256.160 652.650 1256.440 ;
        RECT 654.210 1256.160 654.490 1256.440 ;
        RECT 652.370 772.680 652.650 772.960 ;
        RECT 654.210 772.680 654.490 772.960 ;
        RECT 652.370 676.120 652.650 676.400 ;
        RECT 654.210 676.120 654.490 676.400 ;
        RECT 678.130 587.040 678.410 587.320 ;
        RECT 679.510 587.040 679.790 587.320 ;
      LAYER met3 ;
        RECT 1400.765 2893.210 1401.095 2893.225 ;
        RECT 1439.865 2893.210 1440.195 2893.225 ;
        RECT 1400.765 2892.910 1440.195 2893.210 ;
        RECT 1400.765 2892.895 1401.095 2892.910 ;
        RECT 1439.865 2892.895 1440.195 2892.910 ;
        RECT 1920.000 1838.440 1924.000 1839.040 ;
        RECT 1908.145 1837.170 1908.475 1837.185 ;
        RECT 1920.350 1837.170 1920.650 1838.440 ;
        RECT 1908.145 1836.870 1920.650 1837.170 ;
        RECT 1908.145 1836.855 1908.475 1836.870 ;
        RECT 627.030 1754.890 631.030 1755.040 ;
        RECT 644.985 1754.890 645.315 1754.905 ;
        RECT 627.030 1754.590 645.315 1754.890 ;
        RECT 627.030 1754.440 631.030 1754.590 ;
        RECT 644.985 1754.575 645.315 1754.590 ;
        RECT 652.345 1256.450 652.675 1256.465 ;
        RECT 654.185 1256.450 654.515 1256.465 ;
        RECT 652.345 1256.150 654.515 1256.450 ;
        RECT 652.345 1256.135 652.675 1256.150 ;
        RECT 654.185 1256.135 654.515 1256.150 ;
        RECT 652.345 772.970 652.675 772.985 ;
        RECT 654.185 772.970 654.515 772.985 ;
        RECT 652.345 772.670 654.515 772.970 ;
        RECT 652.345 772.655 652.675 772.670 ;
        RECT 654.185 772.655 654.515 772.670 ;
        RECT 652.345 676.410 652.675 676.425 ;
        RECT 654.185 676.410 654.515 676.425 ;
        RECT 652.345 676.110 654.515 676.410 ;
        RECT 652.345 676.095 652.675 676.110 ;
        RECT 654.185 676.095 654.515 676.110 ;
        RECT 678.105 587.330 678.435 587.345 ;
        RECT 679.485 587.330 679.815 587.345 ;
        RECT 678.105 587.030 679.815 587.330 ;
        RECT 678.105 587.015 678.435 587.030 ;
        RECT 679.485 587.015 679.815 587.030 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1576.030 2897.720 1576.350 2897.780 ;
        RECT 1529.200 2897.580 1576.350 2897.720 ;
        RECT 1472.530 2895.000 1472.850 2895.060 ;
        RECT 1529.200 2895.000 1529.340 2897.580 ;
        RECT 1576.030 2897.520 1576.350 2897.580 ;
        RECT 1472.530 2894.860 1529.340 2895.000 ;
        RECT 1472.530 2894.800 1472.850 2894.860 ;
        RECT 676.270 2892.960 676.590 2893.020 ;
        RECT 627.600 2892.820 676.590 2892.960 ;
        RECT 613.710 2892.620 614.030 2892.680 ;
        RECT 627.600 2892.620 627.740 2892.820 ;
        RECT 676.270 2892.760 676.590 2892.820 ;
        RECT 724.110 2892.960 724.430 2893.020 ;
        RECT 772.870 2892.960 773.190 2893.020 ;
        RECT 724.110 2892.820 773.190 2892.960 ;
        RECT 724.110 2892.760 724.430 2892.820 ;
        RECT 772.870 2892.760 773.190 2892.820 ;
        RECT 820.710 2892.960 821.030 2893.020 ;
        RECT 950.890 2892.960 951.210 2893.020 ;
        RECT 820.710 2892.820 951.210 2892.960 ;
        RECT 820.710 2892.760 821.030 2892.820 ;
        RECT 950.890 2892.760 951.210 2892.820 ;
        RECT 951.350 2892.960 951.670 2893.020 ;
        RECT 1047.490 2892.960 1047.810 2893.020 ;
        RECT 951.350 2892.820 1047.810 2892.960 ;
        RECT 951.350 2892.760 951.670 2892.820 ;
        RECT 1047.490 2892.760 1047.810 2892.820 ;
        RECT 1047.950 2892.960 1048.270 2893.020 ;
        RECT 1144.090 2892.960 1144.410 2893.020 ;
        RECT 1047.950 2892.820 1144.410 2892.960 ;
        RECT 1047.950 2892.760 1048.270 2892.820 ;
        RECT 1144.090 2892.760 1144.410 2892.820 ;
        RECT 1144.550 2892.960 1144.870 2893.020 ;
        RECT 1248.970 2892.960 1249.290 2893.020 ;
        RECT 1144.550 2892.820 1249.290 2892.960 ;
        RECT 1144.550 2892.760 1144.870 2892.820 ;
        RECT 1248.970 2892.760 1249.290 2892.820 ;
        RECT 1249.890 2892.960 1250.210 2893.020 ;
        RECT 1449.070 2892.960 1449.390 2893.020 ;
        RECT 1249.890 2892.820 1449.390 2892.960 ;
        RECT 1249.890 2892.760 1250.210 2892.820 ;
        RECT 1449.070 2892.760 1449.390 2892.820 ;
        RECT 613.710 2892.480 627.740 2892.620 ;
        RECT 613.710 2892.420 614.030 2892.480 ;
        RECT 1449.070 2891.600 1449.390 2891.660 ;
        RECT 1472.530 2891.600 1472.850 2891.660 ;
        RECT 1449.070 2891.460 1472.850 2891.600 ;
        RECT 1449.070 2891.400 1449.390 2891.460 ;
        RECT 1472.530 2891.400 1472.850 2891.460 ;
        RECT 638.550 2594.100 638.870 2594.160 ;
        RECT 627.600 2593.960 638.870 2594.100 ;
        RECT 496.410 2593.760 496.730 2593.820 ;
        RECT 458.780 2593.620 496.730 2593.760 ;
        RECT 432.930 2593.420 433.250 2593.480 ;
        RECT 432.930 2593.280 447.880 2593.420 ;
        RECT 432.930 2593.220 433.250 2593.280 ;
        RECT 447.740 2593.080 447.880 2593.280 ;
        RECT 458.780 2593.080 458.920 2593.620 ;
        RECT 496.410 2593.560 496.730 2593.620 ;
        RECT 496.870 2593.760 497.190 2593.820 ;
        RECT 627.600 2593.760 627.740 2593.960 ;
        RECT 638.550 2593.900 638.870 2593.960 ;
        RECT 496.870 2593.620 531.140 2593.760 ;
        RECT 496.870 2593.560 497.190 2593.620 ;
        RECT 531.000 2593.420 531.140 2593.620 ;
        RECT 531.460 2593.620 573.000 2593.760 ;
        RECT 531.460 2593.420 531.600 2593.620 ;
        RECT 531.000 2593.280 531.600 2593.420 ;
        RECT 572.860 2593.420 573.000 2593.620 ;
        RECT 614.260 2593.620 627.740 2593.760 ;
        RECT 614.260 2593.480 614.400 2593.620 ;
        RECT 612.790 2593.420 613.110 2593.480 ;
        RECT 572.860 2593.280 613.110 2593.420 ;
        RECT 612.790 2593.220 613.110 2593.280 ;
        RECT 614.170 2593.220 614.490 2593.480 ;
        RECT 447.740 2592.940 458.920 2593.080 ;
        RECT 638.550 1703.640 638.870 1703.700 ;
        RECT 1908.610 1703.640 1908.930 1703.700 ;
        RECT 638.550 1703.500 1908.930 1703.640 ;
        RECT 638.550 1703.440 638.870 1703.500 ;
        RECT 1908.610 1703.440 1908.930 1703.500 ;
        RECT 613.250 1689.360 613.570 1689.420 ;
        RECT 638.550 1689.360 638.870 1689.420 ;
        RECT 613.250 1689.220 638.870 1689.360 ;
        RECT 613.250 1689.160 613.570 1689.220 ;
        RECT 638.550 1689.160 638.870 1689.220 ;
        RECT 612.790 1607.760 613.110 1607.820 ;
        RECT 613.710 1607.760 614.030 1607.820 ;
        RECT 612.790 1607.620 614.030 1607.760 ;
        RECT 612.790 1607.560 613.110 1607.620 ;
        RECT 613.710 1607.560 614.030 1607.620 ;
        RECT 612.330 1593.820 612.650 1593.880 ;
        RECT 613.710 1593.820 614.030 1593.880 ;
        RECT 612.330 1593.680 614.030 1593.820 ;
        RECT 612.330 1593.620 612.650 1593.680 ;
        RECT 613.710 1593.620 614.030 1593.680 ;
        RECT 612.330 1545.880 612.650 1545.940 ;
        RECT 613.250 1545.880 613.570 1545.940 ;
        RECT 612.330 1545.740 613.570 1545.880 ;
        RECT 612.330 1545.680 612.650 1545.740 ;
        RECT 613.250 1545.680 613.570 1545.740 ;
        RECT 613.710 883.560 614.030 883.620 ;
        RECT 613.340 883.420 614.030 883.560 ;
        RECT 613.340 882.940 613.480 883.420 ;
        RECT 613.710 883.360 614.030 883.420 ;
        RECT 613.250 882.680 613.570 882.940 ;
        RECT 613.250 821.000 613.570 821.060 ;
        RECT 613.710 821.000 614.030 821.060 ;
        RECT 613.250 820.860 614.030 821.000 ;
        RECT 613.250 820.800 613.570 820.860 ;
        RECT 613.710 820.800 614.030 820.860 ;
        RECT 613.250 786.660 613.570 786.720 ;
        RECT 613.710 786.660 614.030 786.720 ;
        RECT 613.250 786.520 614.030 786.660 ;
        RECT 613.250 786.460 613.570 786.520 ;
        RECT 613.710 786.460 614.030 786.520 ;
        RECT 613.710 739.060 614.030 739.120 ;
        RECT 613.340 738.920 614.030 739.060 ;
        RECT 613.340 738.440 613.480 738.920 ;
        RECT 613.710 738.860 614.030 738.920 ;
        RECT 613.250 738.180 613.570 738.440 ;
        RECT 613.250 689.900 613.570 690.160 ;
        RECT 613.340 689.480 613.480 689.900 ;
        RECT 613.250 689.220 613.570 689.480 ;
        RECT 610.490 590.480 610.810 590.540 ;
        RECT 613.250 590.480 613.570 590.540 ;
        RECT 610.490 590.340 613.570 590.480 ;
        RECT 610.490 590.280 610.810 590.340 ;
        RECT 613.250 590.280 613.570 590.340 ;
        RECT 614.170 589.120 614.490 589.180 ;
        RECT 804.150 589.120 804.470 589.180 ;
        RECT 614.170 588.980 804.470 589.120 ;
        RECT 614.170 588.920 614.490 588.980 ;
        RECT 804.150 588.920 804.470 588.980 ;
        RECT 264.110 22.000 264.430 22.060 ;
        RECT 610.490 22.000 610.810 22.060 ;
        RECT 264.110 21.860 610.810 22.000 ;
        RECT 264.110 21.800 264.430 21.860 ;
        RECT 610.490 21.800 610.810 21.860 ;
      LAYER via ;
        RECT 1472.560 2894.800 1472.820 2895.060 ;
        RECT 1576.060 2897.520 1576.320 2897.780 ;
        RECT 613.740 2892.420 614.000 2892.680 ;
        RECT 676.300 2892.760 676.560 2893.020 ;
        RECT 724.140 2892.760 724.400 2893.020 ;
        RECT 772.900 2892.760 773.160 2893.020 ;
        RECT 820.740 2892.760 821.000 2893.020 ;
        RECT 950.920 2892.760 951.180 2893.020 ;
        RECT 951.380 2892.760 951.640 2893.020 ;
        RECT 1047.520 2892.760 1047.780 2893.020 ;
        RECT 1047.980 2892.760 1048.240 2893.020 ;
        RECT 1144.120 2892.760 1144.380 2893.020 ;
        RECT 1144.580 2892.760 1144.840 2893.020 ;
        RECT 1249.000 2892.760 1249.260 2893.020 ;
        RECT 1249.920 2892.760 1250.180 2893.020 ;
        RECT 1449.100 2892.760 1449.360 2893.020 ;
        RECT 1449.100 2891.400 1449.360 2891.660 ;
        RECT 1472.560 2891.400 1472.820 2891.660 ;
        RECT 432.960 2593.220 433.220 2593.480 ;
        RECT 496.440 2593.560 496.700 2593.820 ;
        RECT 496.900 2593.560 497.160 2593.820 ;
        RECT 638.580 2593.900 638.840 2594.160 ;
        RECT 612.820 2593.220 613.080 2593.480 ;
        RECT 614.200 2593.220 614.460 2593.480 ;
        RECT 638.580 1703.440 638.840 1703.700 ;
        RECT 1908.640 1703.440 1908.900 1703.700 ;
        RECT 613.280 1689.160 613.540 1689.420 ;
        RECT 638.580 1689.160 638.840 1689.420 ;
        RECT 612.820 1607.560 613.080 1607.820 ;
        RECT 613.740 1607.560 614.000 1607.820 ;
        RECT 612.360 1593.620 612.620 1593.880 ;
        RECT 613.740 1593.620 614.000 1593.880 ;
        RECT 612.360 1545.680 612.620 1545.940 ;
        RECT 613.280 1545.680 613.540 1545.940 ;
        RECT 613.740 883.360 614.000 883.620 ;
        RECT 613.280 882.680 613.540 882.940 ;
        RECT 613.280 820.800 613.540 821.060 ;
        RECT 613.740 820.800 614.000 821.060 ;
        RECT 613.280 786.460 613.540 786.720 ;
        RECT 613.740 786.460 614.000 786.720 ;
        RECT 613.740 738.860 614.000 739.120 ;
        RECT 613.280 738.180 613.540 738.440 ;
        RECT 613.280 689.900 613.540 690.160 ;
        RECT 613.280 689.220 613.540 689.480 ;
        RECT 610.520 590.280 610.780 590.540 ;
        RECT 613.280 590.280 613.540 590.540 ;
        RECT 614.200 588.920 614.460 589.180 ;
        RECT 804.180 588.920 804.440 589.180 ;
        RECT 264.140 21.800 264.400 22.060 ;
        RECT 610.520 21.800 610.780 22.060 ;
      LAYER met2 ;
        RECT 1577.370 2897.890 1577.650 2900.055 ;
        RECT 1576.120 2897.810 1577.650 2897.890 ;
        RECT 1576.060 2897.750 1577.650 2897.810 ;
        RECT 1576.060 2897.490 1576.320 2897.750 ;
        RECT 1577.370 2896.055 1577.650 2897.750 ;
        RECT 1472.560 2894.770 1472.820 2895.090 ;
        RECT 676.290 2892.875 676.570 2893.245 ;
        RECT 724.130 2892.875 724.410 2893.245 ;
        RECT 772.890 2892.875 773.170 2893.245 ;
        RECT 820.730 2892.875 821.010 2893.245 ;
        RECT 950.980 2893.050 951.580 2893.130 ;
        RECT 1047.580 2893.050 1048.180 2893.130 ;
        RECT 1144.180 2893.050 1144.780 2893.130 ;
        RECT 950.920 2892.990 951.640 2893.050 ;
        RECT 676.300 2892.730 676.560 2892.875 ;
        RECT 724.140 2892.730 724.400 2892.875 ;
        RECT 772.900 2892.730 773.160 2892.875 ;
        RECT 820.740 2892.730 821.000 2892.875 ;
        RECT 950.920 2892.730 951.180 2892.990 ;
        RECT 951.380 2892.730 951.640 2892.990 ;
        RECT 1047.520 2892.990 1048.240 2893.050 ;
        RECT 1047.520 2892.730 1047.780 2892.990 ;
        RECT 1047.980 2892.730 1048.240 2892.990 ;
        RECT 1144.120 2892.990 1144.840 2893.050 ;
        RECT 1144.120 2892.730 1144.380 2892.990 ;
        RECT 1144.580 2892.730 1144.840 2892.990 ;
        RECT 1248.990 2892.875 1249.270 2893.245 ;
        RECT 1249.910 2892.875 1250.190 2893.245 ;
        RECT 1249.000 2892.730 1249.260 2892.875 ;
        RECT 1249.920 2892.730 1250.180 2892.875 ;
        RECT 1449.100 2892.730 1449.360 2893.050 ;
        RECT 613.740 2892.390 614.000 2892.710 ;
        RECT 432.850 2600.660 433.130 2604.000 ;
        RECT 432.850 2600.000 433.160 2600.660 ;
        RECT 433.020 2593.510 433.160 2600.000 ;
        RECT 496.500 2593.850 497.100 2593.930 ;
        RECT 496.440 2593.790 497.160 2593.850 ;
        RECT 496.440 2593.530 496.700 2593.790 ;
        RECT 496.900 2593.530 497.160 2593.790 ;
        RECT 432.960 2593.190 433.220 2593.510 ;
        RECT 612.820 2593.250 613.080 2593.510 ;
        RECT 613.800 2593.250 613.940 2892.390 ;
        RECT 1449.160 2891.690 1449.300 2892.730 ;
        RECT 1472.620 2891.690 1472.760 2894.770 ;
        RECT 1449.100 2891.370 1449.360 2891.690 ;
        RECT 1472.560 2891.370 1472.820 2891.690 ;
        RECT 638.580 2593.870 638.840 2594.190 ;
        RECT 614.200 2593.250 614.460 2593.510 ;
        RECT 612.820 2593.190 614.460 2593.250 ;
        RECT 612.880 2593.110 614.400 2593.190 ;
        RECT 613.090 1700.410 613.370 1704.000 ;
        RECT 638.640 1703.730 638.780 2593.870 ;
        RECT 1908.630 1801.475 1908.910 1801.845 ;
        RECT 1908.700 1703.730 1908.840 1801.475 ;
        RECT 638.580 1703.410 638.840 1703.730 ;
        RECT 1908.640 1703.410 1908.900 1703.730 ;
        RECT 613.090 1700.000 613.480 1700.410 ;
        RECT 613.340 1689.450 613.480 1700.000 ;
        RECT 638.640 1689.450 638.780 1703.410 ;
        RECT 613.280 1689.130 613.540 1689.450 ;
        RECT 638.580 1689.130 638.840 1689.450 ;
        RECT 613.340 1607.930 613.480 1689.130 ;
        RECT 612.880 1607.850 613.480 1607.930 ;
        RECT 612.820 1607.790 613.480 1607.850 ;
        RECT 612.820 1607.530 613.080 1607.790 ;
        RECT 613.740 1607.530 614.000 1607.850 ;
        RECT 612.880 1607.375 613.020 1607.530 ;
        RECT 613.800 1593.910 613.940 1607.530 ;
        RECT 612.360 1593.590 612.620 1593.910 ;
        RECT 613.740 1593.590 614.000 1593.910 ;
        RECT 612.420 1545.970 612.560 1593.590 ;
        RECT 612.360 1545.650 612.620 1545.970 ;
        RECT 613.280 1545.650 613.540 1545.970 ;
        RECT 613.340 1511.370 613.480 1545.650 ;
        RECT 612.880 1511.230 613.480 1511.370 ;
        RECT 612.880 1510.690 613.020 1511.230 ;
        RECT 612.880 1510.550 613.480 1510.690 ;
        RECT 613.340 1463.090 613.480 1510.550 ;
        RECT 613.340 1462.950 613.940 1463.090 ;
        RECT 613.800 1462.410 613.940 1462.950 ;
        RECT 613.340 1462.270 613.940 1462.410 ;
        RECT 613.340 1414.810 613.480 1462.270 ;
        RECT 612.880 1414.670 613.480 1414.810 ;
        RECT 612.880 1414.130 613.020 1414.670 ;
        RECT 612.880 1413.990 613.480 1414.130 ;
        RECT 613.340 1366.530 613.480 1413.990 ;
        RECT 613.340 1366.390 613.940 1366.530 ;
        RECT 613.800 1365.850 613.940 1366.390 ;
        RECT 613.340 1365.710 613.940 1365.850 ;
        RECT 613.340 1318.250 613.480 1365.710 ;
        RECT 612.880 1318.110 613.480 1318.250 ;
        RECT 612.880 1317.570 613.020 1318.110 ;
        RECT 612.880 1317.430 613.480 1317.570 ;
        RECT 613.340 1269.970 613.480 1317.430 ;
        RECT 613.340 1269.830 613.940 1269.970 ;
        RECT 613.800 1269.290 613.940 1269.830 ;
        RECT 613.340 1269.150 613.940 1269.290 ;
        RECT 613.340 1221.690 613.480 1269.150 ;
        RECT 612.880 1221.550 613.480 1221.690 ;
        RECT 612.880 1221.010 613.020 1221.550 ;
        RECT 612.880 1220.870 613.480 1221.010 ;
        RECT 613.340 1173.410 613.480 1220.870 ;
        RECT 613.340 1173.270 613.940 1173.410 ;
        RECT 613.800 1172.730 613.940 1173.270 ;
        RECT 613.340 1172.590 613.940 1172.730 ;
        RECT 613.340 1125.130 613.480 1172.590 ;
        RECT 612.880 1124.990 613.480 1125.130 ;
        RECT 612.880 1124.450 613.020 1124.990 ;
        RECT 612.880 1124.310 613.480 1124.450 ;
        RECT 613.340 1076.850 613.480 1124.310 ;
        RECT 613.340 1076.710 613.940 1076.850 ;
        RECT 613.800 1076.170 613.940 1076.710 ;
        RECT 613.340 1076.030 613.940 1076.170 ;
        RECT 613.340 1028.570 613.480 1076.030 ;
        RECT 612.880 1028.430 613.480 1028.570 ;
        RECT 612.880 1027.890 613.020 1028.430 ;
        RECT 612.880 1027.750 613.480 1027.890 ;
        RECT 613.340 980.290 613.480 1027.750 ;
        RECT 613.340 980.150 613.940 980.290 ;
        RECT 613.800 979.610 613.940 980.150 ;
        RECT 613.340 979.470 613.940 979.610 ;
        RECT 613.340 932.010 613.480 979.470 ;
        RECT 612.880 931.870 613.480 932.010 ;
        RECT 612.880 931.330 613.020 931.870 ;
        RECT 612.880 931.190 613.480 931.330 ;
        RECT 613.340 917.730 613.480 931.190 ;
        RECT 613.340 917.590 613.940 917.730 ;
        RECT 613.800 883.650 613.940 917.590 ;
        RECT 613.740 883.330 614.000 883.650 ;
        RECT 613.280 882.650 613.540 882.970 ;
        RECT 613.340 835.450 613.480 882.650 ;
        RECT 612.880 835.310 613.480 835.450 ;
        RECT 612.880 834.770 613.020 835.310 ;
        RECT 612.880 834.630 613.480 834.770 ;
        RECT 613.340 821.090 613.480 834.630 ;
        RECT 613.280 820.770 613.540 821.090 ;
        RECT 613.740 820.770 614.000 821.090 ;
        RECT 613.800 786.750 613.940 820.770 ;
        RECT 613.280 786.430 613.540 786.750 ;
        RECT 613.740 786.430 614.000 786.750 ;
        RECT 613.340 772.890 613.480 786.430 ;
        RECT 613.340 772.750 613.940 772.890 ;
        RECT 613.800 739.150 613.940 772.750 ;
        RECT 613.740 738.830 614.000 739.150 ;
        RECT 613.280 738.150 613.540 738.470 ;
        RECT 613.340 690.190 613.480 738.150 ;
        RECT 613.280 689.870 613.540 690.190 ;
        RECT 613.280 689.190 613.540 689.510 ;
        RECT 613.340 590.570 613.480 689.190 ;
        RECT 805.790 600.170 806.070 604.000 ;
        RECT 804.240 600.030 806.070 600.170 ;
        RECT 610.520 590.250 610.780 590.570 ;
        RECT 613.280 590.250 613.540 590.570 ;
        RECT 610.580 22.090 610.720 590.250 ;
        RECT 613.340 589.290 613.480 590.250 ;
        RECT 613.340 589.210 614.400 589.290 ;
        RECT 804.240 589.210 804.380 600.030 ;
        RECT 805.790 600.000 806.070 600.030 ;
        RECT 613.340 589.150 614.460 589.210 ;
        RECT 614.200 588.890 614.460 589.150 ;
        RECT 804.180 588.890 804.440 589.210 ;
        RECT 264.140 21.770 264.400 22.090 ;
        RECT 610.520 21.770 610.780 22.090 ;
        RECT 264.200 2.400 264.340 21.770 ;
        RECT 263.990 -4.800 264.550 2.400 ;
      LAYER via2 ;
        RECT 676.290 2892.920 676.570 2893.200 ;
        RECT 724.130 2892.920 724.410 2893.200 ;
        RECT 772.890 2892.920 773.170 2893.200 ;
        RECT 820.730 2892.920 821.010 2893.200 ;
        RECT 1248.990 2892.920 1249.270 2893.200 ;
        RECT 1249.910 2892.920 1250.190 2893.200 ;
        RECT 1908.630 1801.520 1908.910 1801.800 ;
      LAYER met3 ;
        RECT 676.265 2893.210 676.595 2893.225 ;
        RECT 724.105 2893.210 724.435 2893.225 ;
        RECT 676.265 2892.910 724.435 2893.210 ;
        RECT 676.265 2892.895 676.595 2892.910 ;
        RECT 724.105 2892.895 724.435 2892.910 ;
        RECT 772.865 2893.210 773.195 2893.225 ;
        RECT 820.705 2893.210 821.035 2893.225 ;
        RECT 772.865 2892.910 821.035 2893.210 ;
        RECT 772.865 2892.895 773.195 2892.910 ;
        RECT 820.705 2892.895 821.035 2892.910 ;
        RECT 1248.965 2893.210 1249.295 2893.225 ;
        RECT 1249.885 2893.210 1250.215 2893.225 ;
        RECT 1248.965 2892.910 1250.215 2893.210 ;
        RECT 1248.965 2892.895 1249.295 2892.910 ;
        RECT 1249.885 2892.895 1250.215 2892.910 ;
        RECT 1920.000 1804.440 1924.000 1805.040 ;
        RECT 1908.605 1801.810 1908.935 1801.825 ;
        RECT 1920.350 1801.810 1920.650 1804.440 ;
        RECT 1908.605 1801.510 1920.650 1801.810 ;
        RECT 1908.605 1801.495 1908.935 1801.510 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 2767.160 562.050 2767.220 ;
        RECT 580.130 2767.160 580.450 2767.220 ;
        RECT 561.730 2767.020 580.450 2767.160 ;
        RECT 561.730 2766.960 562.050 2767.020 ;
        RECT 580.130 2766.960 580.450 2767.020 ;
        RECT 580.130 2490.400 580.450 2490.460 ;
        RECT 1736.570 2490.400 1736.890 2490.460 ;
        RECT 580.130 2490.260 1736.890 2490.400 ;
        RECT 580.130 2490.200 580.450 2490.260 ;
        RECT 1736.570 2490.200 1736.890 2490.260 ;
        RECT 544.710 2488.020 545.030 2488.080 ;
        RECT 580.130 2488.020 580.450 2488.080 ;
        RECT 544.710 2487.880 580.450 2488.020 ;
        RECT 544.710 2487.820 545.030 2487.880 ;
        RECT 580.130 2487.820 580.450 2487.880 ;
        RECT 419.680 1978.900 421.200 1979.040 ;
        RECT 419.680 1978.700 419.820 1978.900 ;
        RECT 396.680 1978.560 419.820 1978.700 ;
        RECT 350.130 1978.360 350.450 1978.420 ;
        RECT 396.680 1978.360 396.820 1978.560 ;
        RECT 350.130 1978.220 396.820 1978.360 ;
        RECT 421.060 1978.360 421.200 1978.900 ;
        RECT 544.710 1978.360 545.030 1978.420 ;
        RECT 628.890 1978.360 629.210 1978.420 ;
        RECT 421.060 1978.220 629.210 1978.360 ;
        RECT 350.130 1978.160 350.450 1978.220 ;
        RECT 544.710 1978.160 545.030 1978.220 ;
        RECT 628.890 1978.160 629.210 1978.220 ;
        RECT 282.510 591.840 282.830 591.900 ;
        RECT 628.890 591.840 629.210 591.900 ;
        RECT 282.510 591.700 629.210 591.840 ;
        RECT 282.510 591.640 282.830 591.700 ;
        RECT 628.890 591.640 629.210 591.700 ;
        RECT 628.890 588.780 629.210 588.840 ;
        RECT 814.270 588.780 814.590 588.840 ;
        RECT 628.890 588.640 814.590 588.780 ;
        RECT 628.890 588.580 629.210 588.640 ;
        RECT 814.270 588.580 814.590 588.640 ;
      LAYER via ;
        RECT 561.760 2766.960 562.020 2767.220 ;
        RECT 580.160 2766.960 580.420 2767.220 ;
        RECT 580.160 2490.200 580.420 2490.460 ;
        RECT 1736.600 2490.200 1736.860 2490.460 ;
        RECT 544.740 2487.820 545.000 2488.080 ;
        RECT 580.160 2487.820 580.420 2488.080 ;
        RECT 350.160 1978.160 350.420 1978.420 ;
        RECT 544.740 1978.160 545.000 1978.420 ;
        RECT 628.920 1978.160 629.180 1978.420 ;
        RECT 282.540 591.640 282.800 591.900 ;
        RECT 628.920 591.640 629.180 591.900 ;
        RECT 628.920 588.580 629.180 588.840 ;
        RECT 814.300 588.580 814.560 588.840 ;
      LAYER met2 ;
        RECT 561.760 2766.930 562.020 2767.250 ;
        RECT 580.160 2766.930 580.420 2767.250 ;
        RECT 561.820 2759.520 561.960 2766.930 ;
        RECT 561.650 2759.100 561.960 2759.520 ;
        RECT 561.650 2755.520 561.930 2759.100 ;
        RECT 580.220 2490.490 580.360 2766.930 ;
        RECT 1736.530 2500.000 1736.810 2504.000 ;
        RECT 1736.660 2490.490 1736.800 2500.000 ;
        RECT 580.160 2490.170 580.420 2490.490 ;
        RECT 1736.600 2490.170 1736.860 2490.490 ;
        RECT 580.220 2488.110 580.360 2490.170 ;
        RECT 544.740 2487.790 545.000 2488.110 ;
        RECT 580.160 2487.790 580.420 2488.110 ;
        RECT 544.800 1978.450 544.940 2487.790 ;
        RECT 350.160 1978.130 350.420 1978.450 ;
        RECT 544.740 1978.130 545.000 1978.450 ;
        RECT 628.920 1978.130 629.180 1978.450 ;
        RECT 350.220 1814.765 350.360 1978.130 ;
        RECT 350.150 1814.395 350.430 1814.765 ;
        RECT 628.980 591.930 629.120 1978.130 ;
        RECT 814.990 600.170 815.270 604.000 ;
        RECT 814.360 600.030 815.270 600.170 ;
        RECT 282.540 591.610 282.800 591.930 ;
        RECT 628.920 591.610 629.180 591.930 ;
        RECT 282.600 24.210 282.740 591.610 ;
        RECT 628.980 588.870 629.120 591.610 ;
        RECT 814.360 588.870 814.500 600.030 ;
        RECT 814.990 600.000 815.270 600.030 ;
        RECT 628.920 588.550 629.180 588.870 ;
        RECT 814.300 588.550 814.560 588.870 ;
        RECT 282.140 24.070 282.740 24.210 ;
        RECT 282.140 2.400 282.280 24.070 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 350.150 1814.440 350.430 1814.720 ;
      LAYER met3 ;
        RECT 350.125 1814.730 350.455 1814.745 ;
        RECT 360.000 1814.730 364.000 1814.880 ;
        RECT 350.125 1814.430 364.000 1814.730 ;
        RECT 350.125 1814.415 350.455 1814.430 ;
        RECT 360.000 1814.280 364.000 1814.430 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.970 2487.340 559.290 2487.400 ;
        RECT 629.350 2487.340 629.670 2487.400 ;
        RECT 1863.530 2487.340 1863.850 2487.400 ;
        RECT 558.970 2487.200 1863.850 2487.340 ;
        RECT 558.970 2487.140 559.290 2487.200 ;
        RECT 629.350 2487.140 629.670 2487.200 ;
        RECT 1863.530 2487.140 1863.850 2487.200 ;
        RECT 413.610 1683.580 413.930 1683.640 ;
        RECT 629.350 1683.580 629.670 1683.640 ;
        RECT 413.610 1683.440 629.670 1683.580 ;
        RECT 413.610 1683.380 413.930 1683.440 ;
        RECT 629.350 1683.380 629.670 1683.440 ;
        RECT 413.610 592.520 413.930 592.580 ;
        RECT 822.550 592.520 822.870 592.580 ;
        RECT 413.610 592.380 822.870 592.520 ;
        RECT 413.610 592.320 413.930 592.380 ;
        RECT 822.550 592.320 822.870 592.380 ;
        RECT 303.210 590.140 303.530 590.200 ;
        RECT 413.610 590.140 413.930 590.200 ;
        RECT 303.210 590.000 413.930 590.140 ;
        RECT 303.210 589.940 303.530 590.000 ;
        RECT 413.610 589.940 413.930 590.000 ;
        RECT 299.990 16.220 300.310 16.280 ;
        RECT 303.210 16.220 303.530 16.280 ;
        RECT 299.990 16.080 303.530 16.220 ;
        RECT 299.990 16.020 300.310 16.080 ;
        RECT 303.210 16.020 303.530 16.080 ;
      LAYER via ;
        RECT 559.000 2487.140 559.260 2487.400 ;
        RECT 629.380 2487.140 629.640 2487.400 ;
        RECT 1863.560 2487.140 1863.820 2487.400 ;
        RECT 413.640 1683.380 413.900 1683.640 ;
        RECT 629.380 1683.380 629.640 1683.640 ;
        RECT 413.640 592.320 413.900 592.580 ;
        RECT 822.580 592.320 822.840 592.580 ;
        RECT 303.240 589.940 303.500 590.200 ;
        RECT 413.640 589.940 413.900 590.200 ;
        RECT 300.020 16.020 300.280 16.280 ;
        RECT 303.240 16.020 303.500 16.280 ;
      LAYER met2 ;
        RECT 562.570 2600.730 562.850 2604.000 ;
        RECT 559.060 2600.590 562.850 2600.730 ;
        RECT 559.060 2487.430 559.200 2600.590 ;
        RECT 562.570 2600.000 562.850 2600.590 ;
        RECT 1863.490 2500.000 1863.770 2504.000 ;
        RECT 1863.620 2487.430 1863.760 2500.000 ;
        RECT 559.000 2487.110 559.260 2487.430 ;
        RECT 629.380 2487.110 629.640 2487.430 ;
        RECT 1863.560 2487.110 1863.820 2487.430 ;
        RECT 412.530 1700.410 412.810 1704.000 ;
        RECT 412.530 1700.270 413.840 1700.410 ;
        RECT 412.530 1700.000 412.810 1700.270 ;
        RECT 413.700 1683.670 413.840 1700.270 ;
        RECT 629.440 1683.670 629.580 2487.110 ;
        RECT 413.640 1683.350 413.900 1683.670 ;
        RECT 629.380 1683.350 629.640 1683.670 ;
        RECT 413.700 592.610 413.840 1683.350 ;
        RECT 824.190 600.170 824.470 604.000 ;
        RECT 822.640 600.030 824.470 600.170 ;
        RECT 822.640 592.610 822.780 600.030 ;
        RECT 824.190 600.000 824.470 600.030 ;
        RECT 413.640 592.290 413.900 592.610 ;
        RECT 822.580 592.290 822.840 592.610 ;
        RECT 413.700 590.230 413.840 592.290 ;
        RECT 303.240 589.910 303.500 590.230 ;
        RECT 413.640 589.910 413.900 590.230 ;
        RECT 303.300 16.310 303.440 589.910 ;
        RECT 300.020 15.990 300.280 16.310 ;
        RECT 303.240 15.990 303.500 16.310 ;
        RECT 300.080 2.400 300.220 15.990 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1574.650 2898.060 1574.970 2898.120 ;
        RECT 1578.330 2898.060 1578.650 2898.120 ;
        RECT 1574.650 2897.920 1578.650 2898.060 ;
        RECT 1574.650 2897.860 1574.970 2897.920 ;
        RECT 1578.330 2897.860 1578.650 2897.920 ;
        RECT 1666.190 2897.720 1666.510 2897.780 ;
        RECT 1690.110 2897.720 1690.430 2897.780 ;
        RECT 1666.190 2897.580 1690.430 2897.720 ;
        RECT 1666.190 2897.520 1666.510 2897.580 ;
        RECT 1690.110 2897.520 1690.430 2897.580 ;
        RECT 1574.650 2896.500 1574.970 2896.760 ;
        RECT 1578.330 2896.500 1578.650 2896.760 ;
        RECT 1666.190 2896.500 1666.510 2896.760 ;
        RECT 1690.110 2896.500 1690.430 2896.760 ;
        RECT 1821.210 2896.500 1821.530 2896.760 ;
        RECT 1440.330 2893.980 1440.650 2894.040 ;
        RECT 1488.630 2893.980 1488.950 2894.040 ;
        RECT 1440.330 2893.840 1488.950 2893.980 ;
        RECT 1440.330 2893.780 1440.650 2893.840 ;
        RECT 1488.630 2893.780 1488.950 2893.840 ;
        RECT 1574.740 2893.640 1574.880 2896.500 ;
        RECT 1539.320 2893.500 1574.880 2893.640 ;
        RECT 1539.320 2892.620 1539.460 2893.500 ;
        RECT 1538.860 2892.480 1539.460 2892.620 ;
        RECT 1578.420 2892.620 1578.560 2896.500 ;
        RECT 1666.280 2892.620 1666.420 2896.500 ;
        RECT 1578.420 2892.480 1666.420 2892.620 ;
        RECT 1538.860 2892.280 1539.000 2892.480 ;
        RECT 1508.040 2892.140 1539.000 2892.280 ;
        RECT 1488.630 2891.940 1488.950 2892.000 ;
        RECT 1508.040 2891.940 1508.180 2892.140 ;
        RECT 1488.630 2891.800 1508.180 2891.940 ;
        RECT 1690.200 2891.940 1690.340 2896.500 ;
        RECT 1821.300 2892.620 1821.440 2896.500 ;
        RECT 1787.720 2892.480 1821.440 2892.620 ;
        RECT 1690.200 2891.800 1751.980 2891.940 ;
        RECT 1488.630 2891.740 1488.950 2891.800 ;
        RECT 1751.840 2891.600 1751.980 2891.800 ;
        RECT 1787.720 2891.600 1787.860 2892.480 ;
        RECT 1751.840 2891.460 1787.860 2891.600 ;
        RECT 645.910 2891.260 646.230 2891.320 ;
        RECT 1440.330 2891.260 1440.650 2891.320 ;
        RECT 645.910 2891.120 1440.650 2891.260 ;
        RECT 645.910 2891.060 646.230 2891.120 ;
        RECT 1440.330 2891.060 1440.650 2891.120 ;
        RECT 586.570 2625.380 586.890 2625.440 ;
        RECT 645.910 2625.380 646.230 2625.440 ;
        RECT 586.570 2625.240 646.230 2625.380 ;
        RECT 586.570 2625.180 586.890 2625.240 ;
        RECT 645.910 2625.180 646.230 2625.240 ;
        RECT 644.530 2608.380 644.850 2608.440 ;
        RECT 645.910 2608.380 646.230 2608.440 ;
        RECT 644.530 2608.240 646.230 2608.380 ;
        RECT 644.530 2608.180 644.850 2608.240 ;
        RECT 645.910 2608.180 646.230 2608.240 ;
        RECT 642.690 2511.820 643.010 2511.880 ;
        RECT 644.070 2511.820 644.390 2511.880 ;
        RECT 642.690 2511.680 644.390 2511.820 ;
        RECT 642.690 2511.620 643.010 2511.680 ;
        RECT 644.070 2511.620 644.390 2511.680 ;
        RECT 642.690 2463.200 643.010 2463.260 ;
        RECT 643.610 2463.200 643.930 2463.260 ;
        RECT 642.690 2463.060 643.930 2463.200 ;
        RECT 642.690 2463.000 643.010 2463.060 ;
        RECT 643.610 2463.000 643.930 2463.060 ;
        RECT 643.150 2076.960 643.470 2077.020 ;
        RECT 644.070 2076.960 644.390 2077.020 ;
        RECT 643.150 2076.820 644.390 2076.960 ;
        RECT 643.150 2076.760 643.470 2076.820 ;
        RECT 644.070 2076.760 644.390 2076.820 ;
        RECT 642.690 2028.680 643.010 2028.740 ;
        RECT 644.070 2028.680 644.390 2028.740 ;
        RECT 642.690 2028.540 644.390 2028.680 ;
        RECT 642.690 2028.480 643.010 2028.540 ;
        RECT 644.070 2028.480 644.390 2028.540 ;
        RECT 642.690 1980.740 643.010 1980.800 ;
        RECT 643.150 1980.740 643.470 1980.800 ;
        RECT 642.690 1980.600 643.470 1980.740 ;
        RECT 642.690 1980.540 643.010 1980.600 ;
        RECT 643.150 1980.540 643.470 1980.600 ;
        RECT 643.150 1973.260 643.470 1973.320 ;
        RECT 644.070 1973.260 644.390 1973.320 ;
        RECT 643.150 1973.120 644.390 1973.260 ;
        RECT 643.150 1973.060 643.470 1973.120 ;
        RECT 644.070 1973.060 644.390 1973.120 ;
        RECT 643.150 1945.720 643.470 1945.780 ;
        RECT 644.070 1945.720 644.390 1945.780 ;
        RECT 643.150 1945.580 644.390 1945.720 ;
        RECT 643.150 1945.520 643.470 1945.580 ;
        RECT 644.070 1945.520 644.390 1945.580 ;
        RECT 644.070 1859.360 644.390 1859.420 ;
        RECT 644.990 1859.360 645.310 1859.420 ;
        RECT 644.070 1859.220 645.310 1859.360 ;
        RECT 644.070 1859.160 644.390 1859.220 ;
        RECT 644.990 1859.160 645.310 1859.220 ;
        RECT 644.530 1594.160 644.850 1594.220 ;
        RECT 644.990 1594.160 645.310 1594.220 ;
        RECT 644.530 1594.020 645.310 1594.160 ;
        RECT 644.530 1593.960 644.850 1594.020 ;
        RECT 644.990 1593.960 645.310 1594.020 ;
        RECT 644.070 1511.200 644.390 1511.260 ;
        RECT 644.990 1511.200 645.310 1511.260 ;
        RECT 644.070 1511.060 645.310 1511.200 ;
        RECT 644.070 1511.000 644.390 1511.060 ;
        RECT 644.990 1511.000 645.310 1511.060 ;
        RECT 644.070 1414.640 644.390 1414.700 ;
        RECT 644.990 1414.640 645.310 1414.700 ;
        RECT 644.070 1414.500 645.310 1414.640 ;
        RECT 644.070 1414.440 644.390 1414.500 ;
        RECT 644.990 1414.440 645.310 1414.500 ;
        RECT 644.070 1318.080 644.390 1318.140 ;
        RECT 644.990 1318.080 645.310 1318.140 ;
        RECT 644.070 1317.940 645.310 1318.080 ;
        RECT 644.070 1317.880 644.390 1317.940 ;
        RECT 644.990 1317.880 645.310 1317.940 ;
        RECT 644.070 1221.520 644.390 1221.580 ;
        RECT 644.990 1221.520 645.310 1221.580 ;
        RECT 644.070 1221.380 645.310 1221.520 ;
        RECT 644.070 1221.320 644.390 1221.380 ;
        RECT 644.990 1221.320 645.310 1221.380 ;
        RECT 644.070 1124.960 644.390 1125.020 ;
        RECT 644.990 1124.960 645.310 1125.020 ;
        RECT 644.070 1124.820 645.310 1124.960 ;
        RECT 644.070 1124.760 644.390 1124.820 ;
        RECT 644.990 1124.760 645.310 1124.820 ;
        RECT 643.150 1007.320 643.470 1007.380 ;
        RECT 643.610 1007.320 643.930 1007.380 ;
        RECT 643.150 1007.180 643.930 1007.320 ;
        RECT 643.150 1007.120 643.470 1007.180 ;
        RECT 643.610 1007.120 643.930 1007.180 ;
        RECT 642.690 959.380 643.010 959.440 ;
        RECT 643.150 959.380 643.470 959.440 ;
        RECT 642.690 959.240 643.470 959.380 ;
        RECT 642.690 959.180 643.010 959.240 ;
        RECT 643.150 959.180 643.470 959.240 ;
        RECT 642.690 917.900 643.010 917.960 ;
        RECT 644.530 917.900 644.850 917.960 ;
        RECT 642.690 917.760 644.850 917.900 ;
        RECT 642.690 917.700 643.010 917.760 ;
        RECT 644.530 917.700 644.850 917.760 ;
        RECT 644.070 893.760 644.390 893.820 ;
        RECT 644.990 893.760 645.310 893.820 ;
        RECT 644.070 893.620 645.310 893.760 ;
        RECT 644.070 893.560 644.390 893.620 ;
        RECT 644.990 893.560 645.310 893.620 ;
        RECT 643.150 821.000 643.470 821.060 ;
        RECT 644.070 821.000 644.390 821.060 ;
        RECT 643.150 820.860 644.390 821.000 ;
        RECT 643.150 820.800 643.470 820.860 ;
        RECT 644.070 820.800 644.390 820.860 ;
        RECT 644.070 724.440 644.390 724.500 ;
        RECT 644.530 724.440 644.850 724.500 ;
        RECT 644.070 724.300 644.850 724.440 ;
        RECT 644.070 724.240 644.390 724.300 ;
        RECT 644.530 724.240 644.850 724.300 ;
        RECT 644.070 717.640 644.390 717.700 ;
        RECT 644.990 717.640 645.310 717.700 ;
        RECT 644.070 717.500 645.310 717.640 ;
        RECT 644.070 717.440 644.390 717.500 ;
        RECT 644.990 717.440 645.310 717.500 ;
        RECT 644.070 669.700 644.390 669.760 ;
        RECT 644.990 669.700 645.310 669.760 ;
        RECT 644.070 669.560 645.310 669.700 ;
        RECT 644.070 669.500 644.390 669.560 ;
        RECT 644.990 669.500 645.310 669.560 ;
        RECT 644.070 641.960 644.390 642.220 ;
        RECT 644.160 641.540 644.300 641.960 ;
        RECT 644.070 641.280 644.390 641.540 ;
        RECT 644.070 613.940 644.390 614.000 ;
        RECT 649.590 613.940 649.910 614.000 ;
        RECT 644.070 613.800 649.910 613.940 ;
        RECT 644.070 613.740 644.390 613.800 ;
        RECT 649.590 613.740 649.910 613.800 ;
        RECT 686.390 588.440 686.710 588.500 ;
        RECT 831.750 588.440 832.070 588.500 ;
        RECT 686.390 588.300 832.070 588.440 ;
        RECT 686.390 588.240 686.710 588.300 ;
        RECT 831.750 588.240 832.070 588.300 ;
        RECT 643.150 587.760 643.470 587.820 ;
        RECT 649.590 587.760 649.910 587.820 ;
        RECT 677.190 587.760 677.510 587.820 ;
        RECT 643.150 587.620 677.510 587.760 ;
        RECT 643.150 587.560 643.470 587.620 ;
        RECT 649.590 587.560 649.910 587.620 ;
        RECT 677.190 587.560 677.510 587.620 ;
        RECT 677.190 586.060 677.510 586.120 ;
        RECT 686.390 586.060 686.710 586.120 ;
        RECT 677.190 585.920 686.710 586.060 ;
        RECT 677.190 585.860 677.510 585.920 ;
        RECT 686.390 585.860 686.710 585.920 ;
        RECT 643.150 524.520 643.470 524.580 ;
        RECT 644.990 524.520 645.310 524.580 ;
        RECT 643.150 524.380 645.310 524.520 ;
        RECT 643.150 524.320 643.470 524.380 ;
        RECT 644.990 524.320 645.310 524.380 ;
        RECT 644.990 496.780 645.310 497.040 ;
        RECT 644.530 496.640 644.850 496.700 ;
        RECT 645.080 496.640 645.220 496.780 ;
        RECT 644.530 496.500 645.220 496.640 ;
        RECT 644.530 496.440 644.850 496.500 ;
        RECT 644.530 483.040 644.850 483.100 ;
        RECT 644.990 483.040 645.310 483.100 ;
        RECT 644.530 482.900 645.310 483.040 ;
        RECT 644.530 482.840 644.850 482.900 ;
        RECT 644.990 482.840 645.310 482.900 ;
        RECT 643.610 434.760 643.930 434.820 ;
        RECT 644.530 434.760 644.850 434.820 ;
        RECT 643.610 434.620 644.850 434.760 ;
        RECT 643.610 434.560 643.930 434.620 ;
        RECT 644.530 434.560 644.850 434.620 ;
        RECT 642.690 427.620 643.010 427.680 ;
        RECT 643.610 427.620 643.930 427.680 ;
        RECT 642.690 427.480 643.930 427.620 ;
        RECT 642.690 427.420 643.010 427.480 ;
        RECT 643.610 427.420 643.930 427.480 ;
        RECT 643.150 331.060 643.470 331.120 ;
        RECT 644.070 331.060 644.390 331.120 ;
        RECT 643.150 330.920 644.390 331.060 ;
        RECT 643.150 330.860 643.470 330.920 ;
        RECT 644.070 330.860 644.390 330.920 ;
        RECT 643.150 283.120 643.470 283.180 ;
        RECT 644.530 283.120 644.850 283.180 ;
        RECT 643.150 282.980 644.850 283.120 ;
        RECT 643.150 282.920 643.470 282.980 ;
        RECT 644.530 282.920 644.850 282.980 ;
        RECT 644.530 255.040 644.850 255.300 ;
        RECT 644.620 254.900 644.760 255.040 ;
        RECT 644.990 254.900 645.310 254.960 ;
        RECT 644.620 254.760 645.310 254.900 ;
        RECT 644.990 254.700 645.310 254.760 ;
        RECT 644.990 159.020 645.310 159.080 ;
        RECT 644.620 158.880 645.310 159.020 ;
        RECT 644.620 158.740 644.760 158.880 ;
        RECT 644.990 158.820 645.310 158.880 ;
        RECT 644.530 158.480 644.850 158.740 ;
        RECT 644.530 144.540 644.850 144.800 ;
        RECT 644.620 144.400 644.760 144.540 ;
        RECT 644.990 144.400 645.310 144.460 ;
        RECT 644.620 144.260 645.310 144.400 ;
        RECT 644.990 144.200 645.310 144.260 ;
        RECT 317.930 21.660 318.250 21.720 ;
        RECT 644.070 21.660 644.390 21.720 ;
        RECT 317.930 21.520 644.390 21.660 ;
        RECT 317.930 21.460 318.250 21.520 ;
        RECT 644.070 21.460 644.390 21.520 ;
      LAYER via ;
        RECT 1574.680 2897.860 1574.940 2898.120 ;
        RECT 1578.360 2897.860 1578.620 2898.120 ;
        RECT 1666.220 2897.520 1666.480 2897.780 ;
        RECT 1690.140 2897.520 1690.400 2897.780 ;
        RECT 1574.680 2896.500 1574.940 2896.760 ;
        RECT 1578.360 2896.500 1578.620 2896.760 ;
        RECT 1666.220 2896.500 1666.480 2896.760 ;
        RECT 1690.140 2896.500 1690.400 2896.760 ;
        RECT 1821.240 2896.500 1821.500 2896.760 ;
        RECT 1440.360 2893.780 1440.620 2894.040 ;
        RECT 1488.660 2893.780 1488.920 2894.040 ;
        RECT 1488.660 2891.740 1488.920 2892.000 ;
        RECT 645.940 2891.060 646.200 2891.320 ;
        RECT 1440.360 2891.060 1440.620 2891.320 ;
        RECT 586.600 2625.180 586.860 2625.440 ;
        RECT 645.940 2625.180 646.200 2625.440 ;
        RECT 644.560 2608.180 644.820 2608.440 ;
        RECT 645.940 2608.180 646.200 2608.440 ;
        RECT 642.720 2511.620 642.980 2511.880 ;
        RECT 644.100 2511.620 644.360 2511.880 ;
        RECT 642.720 2463.000 642.980 2463.260 ;
        RECT 643.640 2463.000 643.900 2463.260 ;
        RECT 643.180 2076.760 643.440 2077.020 ;
        RECT 644.100 2076.760 644.360 2077.020 ;
        RECT 642.720 2028.480 642.980 2028.740 ;
        RECT 644.100 2028.480 644.360 2028.740 ;
        RECT 642.720 1980.540 642.980 1980.800 ;
        RECT 643.180 1980.540 643.440 1980.800 ;
        RECT 643.180 1973.060 643.440 1973.320 ;
        RECT 644.100 1973.060 644.360 1973.320 ;
        RECT 643.180 1945.520 643.440 1945.780 ;
        RECT 644.100 1945.520 644.360 1945.780 ;
        RECT 644.100 1859.160 644.360 1859.420 ;
        RECT 645.020 1859.160 645.280 1859.420 ;
        RECT 644.560 1593.960 644.820 1594.220 ;
        RECT 645.020 1593.960 645.280 1594.220 ;
        RECT 644.100 1511.000 644.360 1511.260 ;
        RECT 645.020 1511.000 645.280 1511.260 ;
        RECT 644.100 1414.440 644.360 1414.700 ;
        RECT 645.020 1414.440 645.280 1414.700 ;
        RECT 644.100 1317.880 644.360 1318.140 ;
        RECT 645.020 1317.880 645.280 1318.140 ;
        RECT 644.100 1221.320 644.360 1221.580 ;
        RECT 645.020 1221.320 645.280 1221.580 ;
        RECT 644.100 1124.760 644.360 1125.020 ;
        RECT 645.020 1124.760 645.280 1125.020 ;
        RECT 643.180 1007.120 643.440 1007.380 ;
        RECT 643.640 1007.120 643.900 1007.380 ;
        RECT 642.720 959.180 642.980 959.440 ;
        RECT 643.180 959.180 643.440 959.440 ;
        RECT 642.720 917.700 642.980 917.960 ;
        RECT 644.560 917.700 644.820 917.960 ;
        RECT 644.100 893.560 644.360 893.820 ;
        RECT 645.020 893.560 645.280 893.820 ;
        RECT 643.180 820.800 643.440 821.060 ;
        RECT 644.100 820.800 644.360 821.060 ;
        RECT 644.100 724.240 644.360 724.500 ;
        RECT 644.560 724.240 644.820 724.500 ;
        RECT 644.100 717.440 644.360 717.700 ;
        RECT 645.020 717.440 645.280 717.700 ;
        RECT 644.100 669.500 644.360 669.760 ;
        RECT 645.020 669.500 645.280 669.760 ;
        RECT 644.100 641.960 644.360 642.220 ;
        RECT 644.100 641.280 644.360 641.540 ;
        RECT 644.100 613.740 644.360 614.000 ;
        RECT 649.620 613.740 649.880 614.000 ;
        RECT 686.420 588.240 686.680 588.500 ;
        RECT 831.780 588.240 832.040 588.500 ;
        RECT 643.180 587.560 643.440 587.820 ;
        RECT 649.620 587.560 649.880 587.820 ;
        RECT 677.220 587.560 677.480 587.820 ;
        RECT 677.220 585.860 677.480 586.120 ;
        RECT 686.420 585.860 686.680 586.120 ;
        RECT 643.180 524.320 643.440 524.580 ;
        RECT 645.020 524.320 645.280 524.580 ;
        RECT 645.020 496.780 645.280 497.040 ;
        RECT 644.560 496.440 644.820 496.700 ;
        RECT 644.560 482.840 644.820 483.100 ;
        RECT 645.020 482.840 645.280 483.100 ;
        RECT 643.640 434.560 643.900 434.820 ;
        RECT 644.560 434.560 644.820 434.820 ;
        RECT 642.720 427.420 642.980 427.680 ;
        RECT 643.640 427.420 643.900 427.680 ;
        RECT 643.180 330.860 643.440 331.120 ;
        RECT 644.100 330.860 644.360 331.120 ;
        RECT 643.180 282.920 643.440 283.180 ;
        RECT 644.560 282.920 644.820 283.180 ;
        RECT 644.560 255.040 644.820 255.300 ;
        RECT 645.020 254.700 645.280 254.960 ;
        RECT 645.020 158.820 645.280 159.080 ;
        RECT 644.560 158.480 644.820 158.740 ;
        RECT 644.560 144.540 644.820 144.800 ;
        RECT 645.020 144.200 645.280 144.460 ;
        RECT 317.960 21.460 318.220 21.720 ;
        RECT 644.100 21.460 644.360 21.720 ;
      LAYER met2 ;
        RECT 1574.680 2897.830 1574.940 2898.150 ;
        RECT 1578.360 2897.830 1578.620 2898.150 ;
        RECT 1574.740 2896.790 1574.880 2897.830 ;
        RECT 1578.420 2896.790 1578.560 2897.830 ;
        RECT 1666.220 2897.490 1666.480 2897.810 ;
        RECT 1690.140 2897.490 1690.400 2897.810 ;
        RECT 1666.280 2896.790 1666.420 2897.490 ;
        RECT 1690.200 2896.790 1690.340 2897.490 ;
        RECT 1574.680 2896.470 1574.940 2896.790 ;
        RECT 1578.360 2896.470 1578.620 2896.790 ;
        RECT 1666.220 2896.470 1666.480 2896.790 ;
        RECT 1690.140 2896.470 1690.400 2896.790 ;
        RECT 1821.240 2896.530 1821.500 2896.790 ;
        RECT 1822.090 2896.530 1822.370 2900.055 ;
        RECT 1821.240 2896.470 1822.370 2896.530 ;
        RECT 1821.300 2896.390 1822.370 2896.470 ;
        RECT 1822.090 2896.055 1822.370 2896.390 ;
        RECT 1440.360 2893.750 1440.620 2894.070 ;
        RECT 1488.660 2893.750 1488.920 2894.070 ;
        RECT 1440.420 2891.350 1440.560 2893.750 ;
        RECT 1488.720 2892.030 1488.860 2893.750 ;
        RECT 1488.660 2891.710 1488.920 2892.030 ;
        RECT 645.940 2891.030 646.200 2891.350 ;
        RECT 1440.360 2891.030 1440.620 2891.350 ;
        RECT 586.590 2625.635 586.870 2626.005 ;
        RECT 586.660 2625.470 586.800 2625.635 ;
        RECT 646.000 2625.470 646.140 2891.030 ;
        RECT 586.600 2625.150 586.860 2625.470 ;
        RECT 645.940 2625.150 646.200 2625.470 ;
        RECT 646.000 2608.470 646.140 2625.150 ;
        RECT 644.560 2608.150 644.820 2608.470 ;
        RECT 645.940 2608.150 646.200 2608.470 ;
        RECT 644.620 2573.530 644.760 2608.150 ;
        RECT 643.700 2573.390 644.760 2573.530 ;
        RECT 643.700 2560.045 643.840 2573.390 ;
        RECT 642.710 2559.675 642.990 2560.045 ;
        RECT 643.630 2559.675 643.910 2560.045 ;
        RECT 642.780 2511.910 642.920 2559.675 ;
        RECT 642.720 2511.590 642.980 2511.910 ;
        RECT 644.100 2511.590 644.360 2511.910 ;
        RECT 644.160 2476.970 644.300 2511.590 ;
        RECT 643.700 2476.830 644.300 2476.970 ;
        RECT 643.700 2463.290 643.840 2476.830 ;
        RECT 642.720 2462.970 642.980 2463.290 ;
        RECT 643.640 2462.970 643.900 2463.290 ;
        RECT 642.780 2415.205 642.920 2462.970 ;
        RECT 642.710 2414.835 642.990 2415.205 ;
        RECT 644.090 2414.835 644.370 2415.205 ;
        RECT 644.160 2380.410 644.300 2414.835 ;
        RECT 643.700 2380.270 644.300 2380.410 ;
        RECT 643.700 2342.330 643.840 2380.270 ;
        RECT 642.780 2342.190 643.840 2342.330 ;
        RECT 642.780 2318.645 642.920 2342.190 ;
        RECT 642.710 2318.275 642.990 2318.645 ;
        RECT 644.090 2318.275 644.370 2318.645 ;
        RECT 644.160 2283.850 644.300 2318.275 ;
        RECT 643.700 2283.710 644.300 2283.850 ;
        RECT 643.700 2245.770 643.840 2283.710 ;
        RECT 642.780 2245.630 643.840 2245.770 ;
        RECT 642.780 2222.085 642.920 2245.630 ;
        RECT 642.710 2221.715 642.990 2222.085 ;
        RECT 644.090 2221.715 644.370 2222.085 ;
        RECT 644.160 2187.290 644.300 2221.715 ;
        RECT 643.700 2187.150 644.300 2187.290 ;
        RECT 643.700 2149.210 643.840 2187.150 ;
        RECT 642.780 2149.070 643.840 2149.210 ;
        RECT 642.780 2125.525 642.920 2149.070 ;
        RECT 642.710 2125.155 642.990 2125.525 ;
        RECT 644.090 2125.155 644.370 2125.525 ;
        RECT 644.160 2090.730 644.300 2125.155 ;
        RECT 643.240 2090.590 644.300 2090.730 ;
        RECT 643.240 2077.050 643.380 2090.590 ;
        RECT 643.180 2076.730 643.440 2077.050 ;
        RECT 644.100 2076.730 644.360 2077.050 ;
        RECT 644.160 2028.770 644.300 2076.730 ;
        RECT 642.720 2028.450 642.980 2028.770 ;
        RECT 644.100 2028.450 644.360 2028.770 ;
        RECT 642.780 1980.830 642.920 2028.450 ;
        RECT 642.720 1980.510 642.980 1980.830 ;
        RECT 643.180 1980.510 643.440 1980.830 ;
        RECT 643.240 1973.350 643.380 1980.510 ;
        RECT 643.180 1973.030 643.440 1973.350 ;
        RECT 644.100 1973.030 644.360 1973.350 ;
        RECT 644.160 1945.810 644.300 1973.030 ;
        RECT 643.180 1945.490 643.440 1945.810 ;
        RECT 644.100 1945.490 644.360 1945.810 ;
        RECT 643.240 1939.885 643.380 1945.490 ;
        RECT 643.170 1939.515 643.450 1939.885 ;
        RECT 643.240 1895.570 643.380 1939.515 ;
        RECT 643.240 1895.430 644.300 1895.570 ;
        RECT 644.160 1859.450 644.300 1895.430 ;
        RECT 644.100 1859.130 644.360 1859.450 ;
        RECT 645.020 1859.130 645.280 1859.450 ;
        RECT 645.080 1801.050 645.220 1859.130 ;
        RECT 644.160 1800.910 645.220 1801.050 ;
        RECT 644.160 1800.370 644.300 1800.910 ;
        RECT 644.160 1800.230 644.760 1800.370 ;
        RECT 644.620 1707.890 644.760 1800.230 ;
        RECT 644.620 1707.750 645.220 1707.890 ;
        RECT 645.080 1594.250 645.220 1707.750 ;
        RECT 644.560 1593.930 644.820 1594.250 ;
        RECT 645.020 1593.930 645.280 1594.250 ;
        RECT 644.620 1559.650 644.760 1593.930 ;
        RECT 644.620 1559.510 645.220 1559.650 ;
        RECT 645.080 1511.290 645.220 1559.510 ;
        RECT 644.100 1510.970 644.360 1511.290 ;
        RECT 645.020 1510.970 645.280 1511.290 ;
        RECT 644.160 1510.690 644.300 1510.970 ;
        RECT 644.160 1510.550 644.760 1510.690 ;
        RECT 644.620 1463.090 644.760 1510.550 ;
        RECT 644.620 1462.950 645.220 1463.090 ;
        RECT 645.080 1414.730 645.220 1462.950 ;
        RECT 644.100 1414.410 644.360 1414.730 ;
        RECT 645.020 1414.410 645.280 1414.730 ;
        RECT 644.160 1414.130 644.300 1414.410 ;
        RECT 644.160 1413.990 644.760 1414.130 ;
        RECT 644.620 1366.530 644.760 1413.990 ;
        RECT 644.620 1366.390 645.220 1366.530 ;
        RECT 645.080 1318.170 645.220 1366.390 ;
        RECT 644.100 1317.850 644.360 1318.170 ;
        RECT 645.020 1317.850 645.280 1318.170 ;
        RECT 644.160 1317.570 644.300 1317.850 ;
        RECT 644.160 1317.430 644.760 1317.570 ;
        RECT 644.620 1269.970 644.760 1317.430 ;
        RECT 644.620 1269.830 645.220 1269.970 ;
        RECT 645.080 1221.610 645.220 1269.830 ;
        RECT 644.100 1221.290 644.360 1221.610 ;
        RECT 645.020 1221.290 645.280 1221.610 ;
        RECT 644.160 1221.010 644.300 1221.290 ;
        RECT 644.160 1220.870 644.760 1221.010 ;
        RECT 644.620 1173.410 644.760 1220.870 ;
        RECT 644.620 1173.270 645.220 1173.410 ;
        RECT 645.080 1125.050 645.220 1173.270 ;
        RECT 644.100 1124.730 644.360 1125.050 ;
        RECT 645.020 1124.730 645.280 1125.050 ;
        RECT 644.160 1124.450 644.300 1124.730 ;
        RECT 644.160 1124.310 644.760 1124.450 ;
        RECT 644.620 1076.850 644.760 1124.310 ;
        RECT 644.620 1076.710 645.220 1076.850 ;
        RECT 645.080 1062.685 645.220 1076.710 ;
        RECT 643.630 1062.315 643.910 1062.685 ;
        RECT 645.010 1062.315 645.290 1062.685 ;
        RECT 643.700 1028.060 643.840 1062.315 ;
        RECT 643.700 1027.920 644.760 1028.060 ;
        RECT 644.620 1014.290 644.760 1027.920 ;
        RECT 643.700 1014.150 644.760 1014.290 ;
        RECT 643.700 1007.410 643.840 1014.150 ;
        RECT 643.180 1007.090 643.440 1007.410 ;
        RECT 643.640 1007.090 643.900 1007.410 ;
        RECT 643.240 959.470 643.380 1007.090 ;
        RECT 642.720 959.150 642.980 959.470 ;
        RECT 643.180 959.150 643.440 959.470 ;
        RECT 642.780 917.990 642.920 959.150 ;
        RECT 644.620 917.990 644.760 918.145 ;
        RECT 642.720 917.670 642.980 917.990 ;
        RECT 644.560 917.730 644.820 917.990 ;
        RECT 644.160 917.670 644.820 917.730 ;
        RECT 644.160 917.590 644.760 917.670 ;
        RECT 644.160 893.850 644.300 917.590 ;
        RECT 644.100 893.530 644.360 893.850 ;
        RECT 645.020 893.530 645.280 893.850 ;
        RECT 645.080 821.285 645.220 893.530 ;
        RECT 643.180 820.770 643.440 821.090 ;
        RECT 644.090 820.915 644.370 821.285 ;
        RECT 645.010 820.915 645.290 821.285 ;
        RECT 644.100 820.770 644.360 820.915 ;
        RECT 643.240 773.005 643.380 820.770 ;
        RECT 643.170 772.635 643.450 773.005 ;
        RECT 644.090 772.635 644.370 773.005 ;
        RECT 644.160 738.040 644.300 772.635 ;
        RECT 644.160 737.900 644.760 738.040 ;
        RECT 644.620 724.530 644.760 737.900 ;
        RECT 644.100 724.210 644.360 724.530 ;
        RECT 644.560 724.210 644.820 724.530 ;
        RECT 644.160 717.730 644.300 724.210 ;
        RECT 644.100 717.410 644.360 717.730 ;
        RECT 645.020 717.410 645.280 717.730 ;
        RECT 645.080 669.790 645.220 717.410 ;
        RECT 644.100 669.470 644.360 669.790 ;
        RECT 645.020 669.470 645.280 669.790 ;
        RECT 644.160 642.250 644.300 669.470 ;
        RECT 644.100 641.930 644.360 642.250 ;
        RECT 644.100 641.250 644.360 641.570 ;
        RECT 644.160 614.030 644.300 641.250 ;
        RECT 644.100 613.710 644.360 614.030 ;
        RECT 649.620 613.710 649.880 614.030 ;
        RECT 649.680 587.850 649.820 613.710 ;
        RECT 833.390 600.170 833.670 604.000 ;
        RECT 831.840 600.030 833.670 600.170 ;
        RECT 831.840 588.530 831.980 600.030 ;
        RECT 833.390 600.000 833.670 600.030 ;
        RECT 686.420 588.210 686.680 588.530 ;
        RECT 831.780 588.210 832.040 588.530 ;
        RECT 643.180 587.530 643.440 587.850 ;
        RECT 649.620 587.530 649.880 587.850 ;
        RECT 677.220 587.530 677.480 587.850 ;
        RECT 643.240 524.610 643.380 587.530 ;
        RECT 677.280 586.150 677.420 587.530 ;
        RECT 686.480 586.150 686.620 588.210 ;
        RECT 677.220 585.830 677.480 586.150 ;
        RECT 686.420 585.830 686.680 586.150 ;
        RECT 643.180 524.290 643.440 524.610 ;
        RECT 645.020 524.290 645.280 524.610 ;
        RECT 645.080 497.070 645.220 524.290 ;
        RECT 645.020 496.750 645.280 497.070 ;
        RECT 644.560 496.410 644.820 496.730 ;
        RECT 644.620 483.210 644.760 496.410 ;
        RECT 644.620 483.130 645.220 483.210 ;
        RECT 644.560 483.070 645.280 483.130 ;
        RECT 644.560 482.810 644.820 483.070 ;
        RECT 645.020 482.810 645.280 483.070 ;
        RECT 644.620 434.850 644.760 482.810 ;
        RECT 645.080 482.655 645.220 482.810 ;
        RECT 643.640 434.530 643.900 434.850 ;
        RECT 644.560 434.530 644.820 434.850 ;
        RECT 643.700 427.710 643.840 434.530 ;
        RECT 642.720 427.390 642.980 427.710 ;
        RECT 643.640 427.390 643.900 427.710 ;
        RECT 642.780 385.970 642.920 427.390 ;
        RECT 642.780 385.830 643.840 385.970 ;
        RECT 643.700 362.170 643.840 385.830 ;
        RECT 643.240 362.030 643.840 362.170 ;
        RECT 643.240 338.485 643.380 362.030 ;
        RECT 643.170 338.115 643.450 338.485 ;
        RECT 644.090 338.115 644.370 338.485 ;
        RECT 644.160 331.150 644.300 338.115 ;
        RECT 643.180 330.830 643.440 331.150 ;
        RECT 644.100 330.830 644.360 331.150 ;
        RECT 643.240 283.210 643.380 330.830 ;
        RECT 643.180 282.890 643.440 283.210 ;
        RECT 644.560 282.890 644.820 283.210 ;
        RECT 644.620 255.330 644.760 282.890 ;
        RECT 644.560 255.010 644.820 255.330 ;
        RECT 645.020 254.670 645.280 254.990 ;
        RECT 645.080 159.110 645.220 254.670 ;
        RECT 645.020 158.790 645.280 159.110 ;
        RECT 644.560 158.450 644.820 158.770 ;
        RECT 644.620 144.830 644.760 158.450 ;
        RECT 644.560 144.510 644.820 144.830 ;
        RECT 645.020 144.170 645.280 144.490 ;
        RECT 645.080 62.970 645.220 144.170 ;
        RECT 644.620 62.830 645.220 62.970 ;
        RECT 644.620 62.290 644.760 62.830 ;
        RECT 644.160 62.150 644.760 62.290 ;
        RECT 644.160 21.750 644.300 62.150 ;
        RECT 317.960 21.430 318.220 21.750 ;
        RECT 644.100 21.430 644.360 21.750 ;
        RECT 318.020 2.400 318.160 21.430 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 586.590 2625.680 586.870 2625.960 ;
        RECT 642.710 2559.720 642.990 2560.000 ;
        RECT 643.630 2559.720 643.910 2560.000 ;
        RECT 642.710 2414.880 642.990 2415.160 ;
        RECT 644.090 2414.880 644.370 2415.160 ;
        RECT 642.710 2318.320 642.990 2318.600 ;
        RECT 644.090 2318.320 644.370 2318.600 ;
        RECT 642.710 2221.760 642.990 2222.040 ;
        RECT 644.090 2221.760 644.370 2222.040 ;
        RECT 642.710 2125.200 642.990 2125.480 ;
        RECT 644.090 2125.200 644.370 2125.480 ;
        RECT 643.170 1939.560 643.450 1939.840 ;
        RECT 643.630 1062.360 643.910 1062.640 ;
        RECT 645.010 1062.360 645.290 1062.640 ;
        RECT 644.090 820.960 644.370 821.240 ;
        RECT 645.010 820.960 645.290 821.240 ;
        RECT 643.170 772.680 643.450 772.960 ;
        RECT 644.090 772.680 644.370 772.960 ;
        RECT 643.170 338.160 643.450 338.440 ;
        RECT 644.090 338.160 644.370 338.440 ;
      LAYER met3 ;
        RECT 574.800 2625.970 578.800 2626.480 ;
        RECT 586.565 2625.970 586.895 2625.985 ;
        RECT 574.800 2625.880 586.895 2625.970 ;
        RECT 578.070 2625.670 586.895 2625.880 ;
        RECT 586.565 2625.655 586.895 2625.670 ;
        RECT 642.685 2560.010 643.015 2560.025 ;
        RECT 643.605 2560.010 643.935 2560.025 ;
        RECT 642.685 2559.710 643.935 2560.010 ;
        RECT 642.685 2559.695 643.015 2559.710 ;
        RECT 643.605 2559.695 643.935 2559.710 ;
        RECT 642.685 2415.170 643.015 2415.185 ;
        RECT 644.065 2415.170 644.395 2415.185 ;
        RECT 642.685 2414.870 644.395 2415.170 ;
        RECT 642.685 2414.855 643.015 2414.870 ;
        RECT 644.065 2414.855 644.395 2414.870 ;
        RECT 642.685 2318.610 643.015 2318.625 ;
        RECT 644.065 2318.610 644.395 2318.625 ;
        RECT 642.685 2318.310 644.395 2318.610 ;
        RECT 642.685 2318.295 643.015 2318.310 ;
        RECT 644.065 2318.295 644.395 2318.310 ;
        RECT 642.685 2222.050 643.015 2222.065 ;
        RECT 644.065 2222.050 644.395 2222.065 ;
        RECT 642.685 2221.750 644.395 2222.050 ;
        RECT 642.685 2221.735 643.015 2221.750 ;
        RECT 644.065 2221.735 644.395 2221.750 ;
        RECT 642.685 2125.490 643.015 2125.505 ;
        RECT 644.065 2125.490 644.395 2125.505 ;
        RECT 642.685 2125.190 644.395 2125.490 ;
        RECT 642.685 2125.175 643.015 2125.190 ;
        RECT 644.065 2125.175 644.395 2125.190 ;
        RECT 627.030 1939.850 631.030 1940.000 ;
        RECT 643.145 1939.850 643.475 1939.865 ;
        RECT 627.030 1939.550 643.475 1939.850 ;
        RECT 627.030 1939.400 631.030 1939.550 ;
        RECT 643.145 1939.535 643.475 1939.550 ;
        RECT 643.605 1062.650 643.935 1062.665 ;
        RECT 644.985 1062.650 645.315 1062.665 ;
        RECT 643.605 1062.350 645.315 1062.650 ;
        RECT 643.605 1062.335 643.935 1062.350 ;
        RECT 644.985 1062.335 645.315 1062.350 ;
        RECT 644.065 821.250 644.395 821.265 ;
        RECT 644.985 821.250 645.315 821.265 ;
        RECT 644.065 820.950 645.315 821.250 ;
        RECT 644.065 820.935 644.395 820.950 ;
        RECT 644.985 820.935 645.315 820.950 ;
        RECT 643.145 772.970 643.475 772.985 ;
        RECT 644.065 772.970 644.395 772.985 ;
        RECT 643.145 772.670 644.395 772.970 ;
        RECT 643.145 772.655 643.475 772.670 ;
        RECT 644.065 772.655 644.395 772.670 ;
        RECT 643.145 338.450 643.475 338.465 ;
        RECT 644.065 338.450 644.395 338.465 ;
        RECT 643.145 338.150 644.395 338.450 ;
        RECT 643.145 338.135 643.475 338.150 ;
        RECT 644.065 338.135 644.395 338.150 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 2504.680 482.930 2504.740 ;
        RECT 1902.170 2504.680 1902.490 2504.740 ;
        RECT 482.610 2504.540 1902.490 2504.680 ;
        RECT 482.610 2504.480 482.930 2504.540 ;
        RECT 1902.170 2504.480 1902.490 2504.540 ;
        RECT 351.050 2501.280 351.370 2501.340 ;
        RECT 476.170 2501.280 476.490 2501.340 ;
        RECT 482.610 2501.280 482.930 2501.340 ;
        RECT 351.050 2501.140 482.930 2501.280 ;
        RECT 351.050 2501.080 351.370 2501.140 ;
        RECT 476.170 2501.080 476.490 2501.140 ;
        RECT 482.610 2501.080 482.930 2501.140 ;
        RECT 337.710 587.080 338.030 587.140 ;
        RECT 355.190 587.080 355.510 587.140 ;
        RECT 841.870 587.080 842.190 587.140 ;
        RECT 337.710 586.940 842.190 587.080 ;
        RECT 337.710 586.880 338.030 586.940 ;
        RECT 355.190 586.880 355.510 586.940 ;
        RECT 841.870 586.880 842.190 586.940 ;
      LAYER via ;
        RECT 482.640 2504.480 482.900 2504.740 ;
        RECT 1902.200 2504.480 1902.460 2504.740 ;
        RECT 351.080 2501.080 351.340 2501.340 ;
        RECT 476.200 2501.080 476.460 2501.340 ;
        RECT 482.640 2501.080 482.900 2501.340 ;
        RECT 337.740 586.880 338.000 587.140 ;
        RECT 355.220 586.880 355.480 587.140 ;
        RECT 841.900 586.880 842.160 587.140 ;
      LAYER met2 ;
        RECT 476.090 2600.660 476.370 2604.000 ;
        RECT 476.090 2600.000 476.400 2600.660 ;
        RECT 476.260 2501.370 476.400 2600.000 ;
        RECT 1902.190 2532.475 1902.470 2532.845 ;
        RECT 1902.260 2504.770 1902.400 2532.475 ;
        RECT 482.640 2504.450 482.900 2504.770 ;
        RECT 1902.200 2504.450 1902.460 2504.770 ;
        RECT 482.700 2501.370 482.840 2504.450 ;
        RECT 351.080 2501.050 351.340 2501.370 ;
        RECT 476.200 2501.050 476.460 2501.370 ;
        RECT 482.640 2501.050 482.900 2501.370 ;
        RECT 351.140 1889.565 351.280 2501.050 ;
        RECT 351.070 1889.195 351.350 1889.565 ;
        RECT 355.210 1889.195 355.490 1889.565 ;
        RECT 355.280 587.170 355.420 1889.195 ;
        RECT 842.590 600.170 842.870 604.000 ;
        RECT 841.960 600.030 842.870 600.170 ;
        RECT 841.960 587.170 842.100 600.030 ;
        RECT 842.590 600.000 842.870 600.030 ;
        RECT 337.740 586.850 338.000 587.170 ;
        RECT 355.220 586.850 355.480 587.170 ;
        RECT 841.900 586.850 842.160 587.170 ;
        RECT 337.800 17.410 337.940 586.850 ;
        RECT 335.960 17.270 337.940 17.410 ;
        RECT 335.960 2.400 336.100 17.270 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 1902.190 2532.520 1902.470 2532.800 ;
        RECT 351.070 1889.240 351.350 1889.520 ;
        RECT 355.210 1889.240 355.490 1889.520 ;
      LAYER met3 ;
        RECT 1885.335 2534.360 1889.335 2534.640 ;
        RECT 1885.335 2534.040 1889.370 2534.360 ;
        RECT 1889.070 2532.810 1889.370 2534.040 ;
        RECT 1902.165 2532.810 1902.495 2532.825 ;
        RECT 1889.070 2532.510 1902.495 2532.810 ;
        RECT 1902.165 2532.495 1902.495 2532.510 ;
        RECT 351.045 1889.530 351.375 1889.545 ;
        RECT 355.185 1889.530 355.515 1889.545 ;
        RECT 360.000 1889.530 364.000 1889.680 ;
        RECT 351.045 1889.230 364.000 1889.530 ;
        RECT 351.045 1889.215 351.375 1889.230 ;
        RECT 355.185 1889.215 355.515 1889.230 ;
        RECT 360.000 1889.080 364.000 1889.230 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 475.250 2768.860 475.570 2768.920 ;
        RECT 603.590 2768.860 603.910 2768.920 ;
        RECT 475.250 2768.720 603.910 2768.860 ;
        RECT 475.250 2768.660 475.570 2768.720 ;
        RECT 603.590 2768.660 603.910 2768.720 ;
        RECT 603.590 2490.060 603.910 2490.120 ;
        RECT 606.810 2490.060 607.130 2490.120 ;
        RECT 1694.250 2490.060 1694.570 2490.120 ;
        RECT 603.590 2489.920 1694.570 2490.060 ;
        RECT 603.590 2489.860 603.910 2489.920 ;
        RECT 606.810 2489.860 607.130 2489.920 ;
        RECT 1694.250 2489.860 1694.570 2489.920 ;
        RECT 604.510 1994.340 604.830 1994.400 ;
        RECT 606.810 1994.340 607.130 1994.400 ;
        RECT 628.430 1994.340 628.750 1994.400 ;
        RECT 604.510 1994.200 628.750 1994.340 ;
        RECT 604.510 1994.140 604.830 1994.200 ;
        RECT 606.810 1994.140 607.130 1994.200 ;
        RECT 628.430 1994.140 628.750 1994.200 ;
        RECT 628.430 590.480 628.750 590.540 ;
        RECT 850.150 590.480 850.470 590.540 ;
        RECT 628.430 590.340 850.470 590.480 ;
        RECT 628.430 590.280 628.750 590.340 ;
        RECT 850.150 590.280 850.470 590.340 ;
        RECT 603.590 587.760 603.910 587.820 ;
        RECT 628.430 587.760 628.750 587.820 ;
        RECT 603.590 587.620 628.750 587.760 ;
        RECT 603.590 587.560 603.910 587.620 ;
        RECT 628.430 587.560 628.750 587.620 ;
        RECT 353.350 21.320 353.670 21.380 ;
        RECT 603.590 21.320 603.910 21.380 ;
        RECT 353.350 21.180 603.910 21.320 ;
        RECT 353.350 21.120 353.670 21.180 ;
        RECT 603.590 21.120 603.910 21.180 ;
      LAYER via ;
        RECT 475.280 2768.660 475.540 2768.920 ;
        RECT 603.620 2768.660 603.880 2768.920 ;
        RECT 603.620 2489.860 603.880 2490.120 ;
        RECT 606.840 2489.860 607.100 2490.120 ;
        RECT 1694.280 2489.860 1694.540 2490.120 ;
        RECT 604.540 1994.140 604.800 1994.400 ;
        RECT 606.840 1994.140 607.100 1994.400 ;
        RECT 628.460 1994.140 628.720 1994.400 ;
        RECT 628.460 590.280 628.720 590.540 ;
        RECT 850.180 590.280 850.440 590.540 ;
        RECT 603.620 587.560 603.880 587.820 ;
        RECT 628.460 587.560 628.720 587.820 ;
        RECT 353.380 21.120 353.640 21.380 ;
        RECT 603.620 21.120 603.880 21.380 ;
      LAYER met2 ;
        RECT 475.280 2768.630 475.540 2768.950 ;
        RECT 603.620 2768.630 603.880 2768.950 ;
        RECT 475.340 2759.520 475.480 2768.630 ;
        RECT 475.170 2759.100 475.480 2759.520 ;
        RECT 475.170 2755.520 475.450 2759.100 ;
        RECT 603.680 2490.150 603.820 2768.630 ;
        RECT 1694.210 2500.000 1694.490 2504.000 ;
        RECT 1694.340 2490.150 1694.480 2500.000 ;
        RECT 603.620 2489.830 603.880 2490.150 ;
        RECT 606.840 2489.830 607.100 2490.150 ;
        RECT 1694.280 2489.830 1694.540 2490.150 ;
        RECT 606.900 1994.430 607.040 2489.830 ;
        RECT 604.540 1994.110 604.800 1994.430 ;
        RECT 606.840 1994.110 607.100 1994.430 ;
        RECT 628.460 1994.110 628.720 1994.430 ;
        RECT 602.970 1981.250 603.250 1981.750 ;
        RECT 604.600 1981.250 604.740 1994.110 ;
        RECT 602.970 1981.110 604.740 1981.250 ;
        RECT 602.970 1977.750 603.250 1981.110 ;
        RECT 628.520 590.570 628.660 1994.110 ;
        RECT 851.790 600.170 852.070 604.000 ;
        RECT 850.240 600.030 852.070 600.170 ;
        RECT 850.240 590.570 850.380 600.030 ;
        RECT 851.790 600.000 852.070 600.030 ;
        RECT 628.460 590.250 628.720 590.570 ;
        RECT 850.180 590.250 850.440 590.570 ;
        RECT 628.520 587.850 628.660 590.250 ;
        RECT 603.620 587.530 603.880 587.850 ;
        RECT 628.460 587.530 628.720 587.850 ;
        RECT 603.680 21.410 603.820 587.530 ;
        RECT 353.380 21.090 353.640 21.410 ;
        RECT 603.620 21.090 603.880 21.410 ;
        RECT 353.440 2.400 353.580 21.090 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1529.570 2897.380 1529.890 2897.440 ;
        RECT 1587.070 2897.380 1587.390 2897.440 ;
        RECT 1529.570 2897.240 1587.390 2897.380 ;
        RECT 1529.570 2897.180 1529.890 2897.240 ;
        RECT 1587.070 2897.180 1587.390 2897.240 ;
        RECT 738.370 2894.320 738.690 2894.380 ;
        RECT 786.210 2894.320 786.530 2894.380 ;
        RECT 738.370 2894.180 786.530 2894.320 ;
        RECT 738.370 2894.120 738.690 2894.180 ;
        RECT 786.210 2894.120 786.530 2894.180 ;
        RECT 834.970 2894.320 835.290 2894.380 ;
        RECT 882.350 2894.320 882.670 2894.380 ;
        RECT 834.970 2894.180 882.670 2894.320 ;
        RECT 834.970 2894.120 835.290 2894.180 ;
        RECT 882.350 2894.120 882.670 2894.180 ;
        RECT 1317.970 2894.320 1318.290 2894.380 ;
        RECT 1365.810 2894.320 1366.130 2894.380 ;
        RECT 1317.970 2894.180 1366.130 2894.320 ;
        RECT 1317.970 2894.120 1318.290 2894.180 ;
        RECT 1365.810 2894.120 1366.130 2894.180 ;
        RECT 616.930 2893.980 617.250 2894.040 ;
        RECT 616.930 2893.840 676.500 2893.980 ;
        RECT 616.930 2893.780 617.250 2893.840 ;
        RECT 676.360 2893.700 676.500 2893.840 ;
        RECT 676.270 2893.440 676.590 2893.700 ;
        RECT 1464.250 2892.960 1464.570 2893.020 ;
        RECT 1501.050 2892.960 1501.370 2893.020 ;
        RECT 1464.250 2892.820 1501.370 2892.960 ;
        RECT 1464.250 2892.760 1464.570 2892.820 ;
        RECT 1501.050 2892.760 1501.370 2892.820 ;
        RECT 1438.950 2892.620 1439.270 2892.680 ;
        RECT 1449.530 2892.620 1449.850 2892.680 ;
        RECT 1438.950 2892.480 1449.850 2892.620 ;
        RECT 1438.950 2892.420 1439.270 2892.480 ;
        RECT 1449.530 2892.420 1449.850 2892.480 ;
        RECT 677.650 2892.280 677.970 2892.340 ;
        RECT 738.370 2892.280 738.690 2892.340 ;
        RECT 677.650 2892.140 738.690 2892.280 ;
        RECT 677.650 2892.080 677.970 2892.140 ;
        RECT 738.370 2892.080 738.690 2892.140 ;
        RECT 786.210 2892.280 786.530 2892.340 ;
        RECT 834.970 2892.280 835.290 2892.340 ;
        RECT 786.210 2892.140 835.290 2892.280 ;
        RECT 786.210 2892.080 786.530 2892.140 ;
        RECT 834.970 2892.080 835.290 2892.140 ;
        RECT 882.350 2892.280 882.670 2892.340 ;
        RECT 927.430 2892.280 927.750 2892.340 ;
        RECT 882.350 2892.140 927.750 2892.280 ;
        RECT 882.350 2892.080 882.670 2892.140 ;
        RECT 927.430 2892.080 927.750 2892.140 ;
        RECT 951.350 2892.280 951.670 2892.340 ;
        RECT 1015.750 2892.280 1016.070 2892.340 ;
        RECT 951.350 2892.140 1016.070 2892.280 ;
        RECT 951.350 2892.080 951.670 2892.140 ;
        RECT 1015.750 2892.080 1016.070 2892.140 ;
        RECT 1047.950 2892.280 1048.270 2892.340 ;
        RECT 1112.350 2892.280 1112.670 2892.340 ;
        RECT 1047.950 2892.140 1112.670 2892.280 ;
        RECT 1047.950 2892.080 1048.270 2892.140 ;
        RECT 1112.350 2892.080 1112.670 2892.140 ;
        RECT 1144.550 2892.280 1144.870 2892.340 ;
        RECT 1317.970 2892.280 1318.290 2892.340 ;
        RECT 1144.550 2892.140 1318.290 2892.280 ;
        RECT 1144.550 2892.080 1144.870 2892.140 ;
        RECT 1317.970 2892.080 1318.290 2892.140 ;
        RECT 1365.810 2892.280 1366.130 2892.340 ;
        RECT 1400.770 2892.280 1401.090 2892.340 ;
        RECT 1365.810 2892.140 1401.090 2892.280 ;
        RECT 1365.810 2892.080 1366.130 2892.140 ;
        RECT 1400.770 2892.080 1401.090 2892.140 ;
        RECT 576.910 2891.600 577.230 2891.660 ;
        RECT 616.930 2891.600 617.250 2891.660 ;
        RECT 576.910 2891.460 617.250 2891.600 ;
        RECT 576.910 2891.400 577.230 2891.460 ;
        RECT 616.930 2891.400 617.250 2891.460 ;
        RECT 427.410 2749.480 427.730 2749.540 ;
        RECT 432.010 2749.480 432.330 2749.540 ;
        RECT 576.910 2749.480 577.230 2749.540 ;
        RECT 427.410 2749.340 577.230 2749.480 ;
        RECT 427.410 2749.280 427.730 2749.340 ;
        RECT 432.010 2749.280 432.330 2749.340 ;
        RECT 576.910 2749.280 577.230 2749.340 ;
        RECT 358.410 1994.340 358.730 1994.400 ;
        RECT 427.410 1994.340 427.730 1994.400 ;
        RECT 358.410 1994.200 427.730 1994.340 ;
        RECT 358.410 1994.140 358.730 1994.200 ;
        RECT 427.410 1994.140 427.730 1994.200 ;
        RECT 427.410 1993.660 427.730 1993.720 ;
        RECT 451.330 1993.660 451.650 1993.720 ;
        RECT 427.410 1993.520 451.650 1993.660 ;
        RECT 427.410 1993.460 427.730 1993.520 ;
        RECT 451.330 1993.460 451.650 1993.520 ;
        RECT 358.410 590.480 358.730 590.540 ;
        RECT 368.990 590.480 369.310 590.540 ;
        RECT 369.910 590.480 370.230 590.540 ;
        RECT 358.410 590.340 370.230 590.480 ;
        RECT 358.410 590.280 358.730 590.340 ;
        RECT 368.990 590.280 369.310 590.340 ;
        RECT 369.910 590.280 370.230 590.340 ;
        RECT 369.910 589.800 370.230 589.860 ;
        RECT 448.570 589.800 448.890 589.860 ;
        RECT 369.910 589.660 448.890 589.800 ;
        RECT 369.910 589.600 370.230 589.660 ;
        RECT 448.570 589.600 448.890 589.660 ;
        RECT 587.950 589.800 588.270 589.860 ;
        RECT 689.610 589.800 689.930 589.860 ;
        RECT 587.950 589.660 689.930 589.800 ;
        RECT 587.950 589.600 588.270 589.660 ;
        RECT 689.610 589.600 689.930 589.660 ;
        RECT 690.070 589.800 690.390 589.860 ;
        RECT 738.370 589.800 738.690 589.860 ;
        RECT 690.070 589.660 738.690 589.800 ;
        RECT 690.070 589.600 690.390 589.660 ;
        RECT 738.370 589.600 738.690 589.660 ;
        RECT 820.710 589.800 821.030 589.860 ;
        RECT 859.350 589.800 859.670 589.860 ;
        RECT 820.710 589.660 859.670 589.800 ;
        RECT 820.710 589.600 821.030 589.660 ;
        RECT 859.350 589.600 859.670 589.660 ;
        RECT 762.290 589.460 762.610 589.520 ;
        RECT 772.870 589.460 773.190 589.520 ;
        RECT 762.290 589.320 773.190 589.460 ;
        RECT 762.290 589.260 762.610 589.320 ;
        RECT 772.870 589.260 773.190 589.320 ;
        RECT 448.570 588.780 448.890 588.840 ;
        RECT 587.950 588.780 588.270 588.840 ;
        RECT 448.570 588.640 496.180 588.780 ;
        RECT 448.570 588.580 448.890 588.640 ;
        RECT 496.040 587.760 496.180 588.640 ;
        RECT 569.180 588.640 588.270 588.780 ;
        RECT 497.420 587.960 544.940 588.100 ;
        RECT 497.420 587.760 497.560 587.960 ;
        RECT 496.040 587.620 497.560 587.760 ;
        RECT 544.800 587.760 544.940 587.960 ;
        RECT 569.180 587.760 569.320 588.640 ;
        RECT 587.950 588.580 588.270 588.640 ;
        RECT 544.800 587.620 569.320 587.760 ;
        RECT 738.370 587.420 738.690 587.480 ;
        RECT 762.290 587.420 762.610 587.480 ;
        RECT 738.370 587.280 762.610 587.420 ;
        RECT 738.370 587.220 738.690 587.280 ;
        RECT 762.290 587.220 762.610 587.280 ;
        RECT 689.610 586.400 689.930 586.460 ;
        RECT 690.070 586.400 690.390 586.460 ;
        RECT 689.610 586.260 690.390 586.400 ;
        RECT 689.610 586.200 689.930 586.260 ;
        RECT 690.070 586.200 690.390 586.260 ;
        RECT 368.990 16.220 369.310 16.280 ;
        RECT 371.290 16.220 371.610 16.280 ;
        RECT 368.990 16.080 371.610 16.220 ;
        RECT 368.990 16.020 369.310 16.080 ;
        RECT 371.290 16.020 371.610 16.080 ;
      LAYER via ;
        RECT 1529.600 2897.180 1529.860 2897.440 ;
        RECT 1587.100 2897.180 1587.360 2897.440 ;
        RECT 738.400 2894.120 738.660 2894.380 ;
        RECT 786.240 2894.120 786.500 2894.380 ;
        RECT 835.000 2894.120 835.260 2894.380 ;
        RECT 882.380 2894.120 882.640 2894.380 ;
        RECT 1318.000 2894.120 1318.260 2894.380 ;
        RECT 1365.840 2894.120 1366.100 2894.380 ;
        RECT 616.960 2893.780 617.220 2894.040 ;
        RECT 676.300 2893.440 676.560 2893.700 ;
        RECT 1464.280 2892.760 1464.540 2893.020 ;
        RECT 1501.080 2892.760 1501.340 2893.020 ;
        RECT 1438.980 2892.420 1439.240 2892.680 ;
        RECT 1449.560 2892.420 1449.820 2892.680 ;
        RECT 677.680 2892.080 677.940 2892.340 ;
        RECT 738.400 2892.080 738.660 2892.340 ;
        RECT 786.240 2892.080 786.500 2892.340 ;
        RECT 835.000 2892.080 835.260 2892.340 ;
        RECT 882.380 2892.080 882.640 2892.340 ;
        RECT 927.460 2892.080 927.720 2892.340 ;
        RECT 951.380 2892.080 951.640 2892.340 ;
        RECT 1015.780 2892.080 1016.040 2892.340 ;
        RECT 1047.980 2892.080 1048.240 2892.340 ;
        RECT 1112.380 2892.080 1112.640 2892.340 ;
        RECT 1144.580 2892.080 1144.840 2892.340 ;
        RECT 1318.000 2892.080 1318.260 2892.340 ;
        RECT 1365.840 2892.080 1366.100 2892.340 ;
        RECT 1400.800 2892.080 1401.060 2892.340 ;
        RECT 576.940 2891.400 577.200 2891.660 ;
        RECT 616.960 2891.400 617.220 2891.660 ;
        RECT 427.440 2749.280 427.700 2749.540 ;
        RECT 432.040 2749.280 432.300 2749.540 ;
        RECT 576.940 2749.280 577.200 2749.540 ;
        RECT 358.440 1994.140 358.700 1994.400 ;
        RECT 427.440 1994.140 427.700 1994.400 ;
        RECT 427.440 1993.460 427.700 1993.720 ;
        RECT 451.360 1993.460 451.620 1993.720 ;
        RECT 358.440 590.280 358.700 590.540 ;
        RECT 369.020 590.280 369.280 590.540 ;
        RECT 369.940 590.280 370.200 590.540 ;
        RECT 369.940 589.600 370.200 589.860 ;
        RECT 448.600 589.600 448.860 589.860 ;
        RECT 587.980 589.600 588.240 589.860 ;
        RECT 689.640 589.600 689.900 589.860 ;
        RECT 690.100 589.600 690.360 589.860 ;
        RECT 738.400 589.600 738.660 589.860 ;
        RECT 820.740 589.600 821.000 589.860 ;
        RECT 859.380 589.600 859.640 589.860 ;
        RECT 762.320 589.260 762.580 589.520 ;
        RECT 772.900 589.260 773.160 589.520 ;
        RECT 448.600 588.580 448.860 588.840 ;
        RECT 587.980 588.580 588.240 588.840 ;
        RECT 738.400 587.220 738.660 587.480 ;
        RECT 762.320 587.220 762.580 587.480 ;
        RECT 689.640 586.200 689.900 586.460 ;
        RECT 690.100 586.200 690.360 586.460 ;
        RECT 369.020 16.020 369.280 16.280 ;
        RECT 371.320 16.020 371.580 16.280 ;
      LAYER met2 ;
        RECT 1529.600 2897.150 1529.860 2897.470 ;
        RECT 1587.100 2897.210 1587.360 2897.470 ;
        RECT 1588.410 2897.210 1588.690 2900.055 ;
        RECT 1587.100 2897.150 1588.690 2897.210 ;
        RECT 1529.660 2896.645 1529.800 2897.150 ;
        RECT 1587.160 2897.070 1588.690 2897.150 ;
        RECT 1501.070 2896.275 1501.350 2896.645 ;
        RECT 1529.590 2896.275 1529.870 2896.645 ;
        RECT 738.400 2894.090 738.660 2894.410 ;
        RECT 786.240 2894.090 786.500 2894.410 ;
        RECT 835.000 2894.090 835.260 2894.410 ;
        RECT 882.380 2894.090 882.640 2894.410 ;
        RECT 1318.000 2894.090 1318.260 2894.410 ;
        RECT 1365.840 2894.090 1366.100 2894.410 ;
        RECT 616.960 2893.750 617.220 2894.070 ;
        RECT 617.020 2891.690 617.160 2893.750 ;
        RECT 676.300 2893.640 676.560 2893.730 ;
        RECT 676.300 2893.500 676.960 2893.640 ;
        RECT 676.300 2893.410 676.560 2893.500 ;
        RECT 676.820 2892.280 676.960 2893.500 ;
        RECT 738.460 2892.370 738.600 2894.090 ;
        RECT 786.300 2892.370 786.440 2894.090 ;
        RECT 835.060 2892.370 835.200 2894.090 ;
        RECT 882.440 2892.370 882.580 2894.090 ;
        RECT 677.680 2892.280 677.940 2892.370 ;
        RECT 676.820 2892.140 677.940 2892.280 ;
        RECT 677.680 2892.050 677.940 2892.140 ;
        RECT 738.400 2892.050 738.660 2892.370 ;
        RECT 786.240 2892.050 786.500 2892.370 ;
        RECT 835.000 2892.050 835.260 2892.370 ;
        RECT 882.380 2892.050 882.640 2892.370 ;
        RECT 927.450 2892.195 927.730 2892.565 ;
        RECT 951.370 2892.195 951.650 2892.565 ;
        RECT 1015.770 2892.195 1016.050 2892.565 ;
        RECT 1047.970 2892.195 1048.250 2892.565 ;
        RECT 1112.370 2892.195 1112.650 2892.565 ;
        RECT 1144.570 2892.195 1144.850 2892.565 ;
        RECT 1318.060 2892.370 1318.200 2894.090 ;
        RECT 1365.900 2892.370 1366.040 2894.090 ;
        RECT 1449.550 2892.875 1449.830 2893.245 ;
        RECT 1464.270 2892.875 1464.550 2893.245 ;
        RECT 1501.140 2893.050 1501.280 2896.275 ;
        RECT 1588.410 2896.055 1588.690 2897.070 ;
        RECT 1449.620 2892.710 1449.760 2892.875 ;
        RECT 1464.280 2892.730 1464.540 2892.875 ;
        RECT 1501.080 2892.730 1501.340 2893.050 ;
        RECT 1438.980 2892.565 1439.240 2892.710 ;
        RECT 927.460 2892.050 927.720 2892.195 ;
        RECT 951.380 2892.050 951.640 2892.195 ;
        RECT 1015.780 2892.050 1016.040 2892.195 ;
        RECT 1047.980 2892.050 1048.240 2892.195 ;
        RECT 1112.380 2892.050 1112.640 2892.195 ;
        RECT 1144.580 2892.050 1144.840 2892.195 ;
        RECT 1318.000 2892.050 1318.260 2892.370 ;
        RECT 1365.840 2892.050 1366.100 2892.370 ;
        RECT 1400.790 2892.025 1401.070 2892.395 ;
        RECT 1438.970 2892.195 1439.250 2892.565 ;
        RECT 1449.560 2892.390 1449.820 2892.710 ;
        RECT 576.940 2891.370 577.200 2891.690 ;
        RECT 616.960 2891.370 617.220 2891.690 ;
        RECT 427.440 2749.250 427.700 2749.570 ;
        RECT 432.030 2749.395 432.310 2749.765 ;
        RECT 577.000 2749.570 577.140 2891.370 ;
        RECT 432.040 2749.250 432.300 2749.395 ;
        RECT 576.940 2749.250 577.200 2749.570 ;
        RECT 427.500 1994.430 427.640 2749.250 ;
        RECT 358.440 1994.110 358.700 1994.430 ;
        RECT 427.440 1994.110 427.700 1994.430 ;
        RECT 358.500 590.570 358.640 1994.110 ;
        RECT 427.500 1993.750 427.640 1994.110 ;
        RECT 427.440 1993.430 427.700 1993.750 ;
        RECT 451.360 1993.430 451.620 1993.750 ;
        RECT 451.420 1981.250 451.560 1993.430 ;
        RECT 453.010 1981.250 453.290 1981.750 ;
        RECT 451.420 1981.110 453.290 1981.250 ;
        RECT 453.010 1977.750 453.290 1981.110 ;
        RECT 860.990 600.170 861.270 604.000 ;
        RECT 859.440 600.030 861.270 600.170 ;
        RECT 358.440 590.250 358.700 590.570 ;
        RECT 369.020 590.250 369.280 590.570 ;
        RECT 369.940 590.250 370.200 590.570 ;
        RECT 369.080 16.310 369.220 590.250 ;
        RECT 370.000 589.890 370.140 590.250 ;
        RECT 859.440 589.890 859.580 600.030 ;
        RECT 860.990 600.000 861.270 600.030 ;
        RECT 369.940 589.570 370.200 589.890 ;
        RECT 448.600 589.570 448.860 589.890 ;
        RECT 587.980 589.570 588.240 589.890 ;
        RECT 689.640 589.570 689.900 589.890 ;
        RECT 690.100 589.570 690.360 589.890 ;
        RECT 738.400 589.570 738.660 589.890 ;
        RECT 820.740 589.570 821.000 589.890 ;
        RECT 859.380 589.570 859.640 589.890 ;
        RECT 448.660 588.870 448.800 589.570 ;
        RECT 588.040 588.870 588.180 589.570 ;
        RECT 448.600 588.550 448.860 588.870 ;
        RECT 587.980 588.550 588.240 588.870 ;
        RECT 689.700 586.490 689.840 589.570 ;
        RECT 690.160 586.490 690.300 589.570 ;
        RECT 738.460 587.510 738.600 589.570 ;
        RECT 762.320 589.230 762.580 589.550 ;
        RECT 772.900 589.230 773.160 589.550 ;
        RECT 762.380 587.510 762.520 589.230 ;
        RECT 772.960 588.725 773.100 589.230 ;
        RECT 820.800 588.725 820.940 589.570 ;
        RECT 772.890 588.355 773.170 588.725 ;
        RECT 820.730 588.355 821.010 588.725 ;
        RECT 738.400 587.190 738.660 587.510 ;
        RECT 762.320 587.190 762.580 587.510 ;
        RECT 689.640 586.170 689.900 586.490 ;
        RECT 690.100 586.170 690.360 586.490 ;
        RECT 369.020 15.990 369.280 16.310 ;
        RECT 371.320 15.990 371.580 16.310 ;
        RECT 371.380 2.400 371.520 15.990 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 1501.070 2896.320 1501.350 2896.600 ;
        RECT 1529.590 2896.320 1529.870 2896.600 ;
        RECT 927.450 2892.240 927.730 2892.520 ;
        RECT 951.370 2892.240 951.650 2892.520 ;
        RECT 1015.770 2892.240 1016.050 2892.520 ;
        RECT 1047.970 2892.240 1048.250 2892.520 ;
        RECT 1112.370 2892.240 1112.650 2892.520 ;
        RECT 1144.570 2892.240 1144.850 2892.520 ;
        RECT 1449.550 2892.920 1449.830 2893.200 ;
        RECT 1464.270 2892.920 1464.550 2893.200 ;
        RECT 1400.790 2892.070 1401.070 2892.350 ;
        RECT 1438.970 2892.240 1439.250 2892.520 ;
        RECT 432.030 2749.440 432.310 2749.720 ;
        RECT 772.890 588.400 773.170 588.680 ;
        RECT 820.730 588.400 821.010 588.680 ;
      LAYER met3 ;
        RECT 1501.045 2896.610 1501.375 2896.625 ;
        RECT 1529.565 2896.610 1529.895 2896.625 ;
        RECT 1501.045 2896.310 1529.895 2896.610 ;
        RECT 1501.045 2896.295 1501.375 2896.310 ;
        RECT 1529.565 2896.295 1529.895 2896.310 ;
        RECT 1449.525 2893.210 1449.855 2893.225 ;
        RECT 1464.245 2893.210 1464.575 2893.225 ;
        RECT 1449.525 2892.910 1464.575 2893.210 ;
        RECT 1449.525 2892.895 1449.855 2892.910 ;
        RECT 1464.245 2892.895 1464.575 2892.910 ;
        RECT 927.425 2892.530 927.755 2892.545 ;
        RECT 951.345 2892.530 951.675 2892.545 ;
        RECT 927.425 2892.230 951.675 2892.530 ;
        RECT 927.425 2892.215 927.755 2892.230 ;
        RECT 951.345 2892.215 951.675 2892.230 ;
        RECT 1015.745 2892.530 1016.075 2892.545 ;
        RECT 1047.945 2892.530 1048.275 2892.545 ;
        RECT 1015.745 2892.230 1048.275 2892.530 ;
        RECT 1015.745 2892.215 1016.075 2892.230 ;
        RECT 1047.945 2892.215 1048.275 2892.230 ;
        RECT 1112.345 2892.530 1112.675 2892.545 ;
        RECT 1144.545 2892.530 1144.875 2892.545 ;
        RECT 1438.945 2892.530 1439.275 2892.545 ;
        RECT 1112.345 2892.230 1144.875 2892.530 ;
        RECT 1112.345 2892.215 1112.675 2892.230 ;
        RECT 1144.545 2892.215 1144.875 2892.230 ;
        RECT 1400.550 2892.230 1439.275 2892.530 ;
        RECT 1400.550 2892.060 1401.095 2892.230 ;
        RECT 1438.945 2892.215 1439.275 2892.230 ;
        RECT 1400.765 2892.045 1401.095 2892.060 ;
        RECT 430.000 2752.360 434.000 2752.960 ;
        RECT 431.790 2749.745 432.090 2752.360 ;
        RECT 431.790 2749.430 432.335 2749.745 ;
        RECT 432.005 2749.415 432.335 2749.430 ;
        RECT 772.865 588.690 773.195 588.705 ;
        RECT 820.705 588.690 821.035 588.705 ;
        RECT 772.865 588.390 821.035 588.690 ;
        RECT 772.865 588.375 773.195 588.390 ;
        RECT 820.705 588.375 821.035 588.390 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 503.770 2768.520 504.090 2768.580 ;
        RECT 645.450 2768.520 645.770 2768.580 ;
        RECT 503.770 2768.380 645.770 2768.520 ;
        RECT 503.770 2768.320 504.090 2768.380 ;
        RECT 645.450 2768.320 645.770 2768.380 ;
        RECT 645.450 2490.740 645.770 2490.800 ;
        RECT 1821.210 2490.740 1821.530 2490.800 ;
        RECT 645.450 2490.600 1821.530 2490.740 ;
        RECT 645.450 2490.540 645.770 2490.600 ;
        RECT 1821.210 2490.540 1821.530 2490.600 ;
        RECT 645.450 590.820 645.770 590.880 ;
        RECT 869.470 590.820 869.790 590.880 ;
        RECT 645.450 590.680 869.790 590.820 ;
        RECT 645.450 590.620 645.770 590.680 ;
        RECT 869.470 590.620 869.790 590.680 ;
        RECT 593.010 36.620 593.330 36.680 ;
        RECT 434.400 36.480 593.330 36.620 ;
        RECT 389.230 36.280 389.550 36.340 ;
        RECT 434.400 36.280 434.540 36.480 ;
        RECT 593.010 36.420 593.330 36.480 ;
        RECT 389.230 36.140 434.540 36.280 ;
        RECT 389.230 36.080 389.550 36.140 ;
        RECT 617.850 35.940 618.170 36.000 ;
        RECT 645.450 35.940 645.770 36.000 ;
        RECT 617.850 35.800 645.770 35.940 ;
        RECT 617.850 35.740 618.170 35.800 ;
        RECT 645.450 35.740 645.770 35.800 ;
      LAYER via ;
        RECT 503.800 2768.320 504.060 2768.580 ;
        RECT 645.480 2768.320 645.740 2768.580 ;
        RECT 645.480 2490.540 645.740 2490.800 ;
        RECT 1821.240 2490.540 1821.500 2490.800 ;
        RECT 645.480 590.620 645.740 590.880 ;
        RECT 869.500 590.620 869.760 590.880 ;
        RECT 389.260 36.080 389.520 36.340 ;
        RECT 593.040 36.420 593.300 36.680 ;
        RECT 617.880 35.740 618.140 36.000 ;
        RECT 645.480 35.740 645.740 36.000 ;
      LAYER met2 ;
        RECT 503.800 2768.290 504.060 2768.610 ;
        RECT 645.480 2768.290 645.740 2768.610 ;
        RECT 503.860 2759.520 504.000 2768.290 ;
        RECT 503.690 2759.100 504.000 2759.520 ;
        RECT 503.690 2755.520 503.970 2759.100 ;
        RECT 645.540 2490.830 645.680 2768.290 ;
        RECT 1821.170 2500.000 1821.450 2504.000 ;
        RECT 1821.300 2490.830 1821.440 2500.000 ;
        RECT 645.480 2490.510 645.740 2490.830 ;
        RECT 1821.240 2490.510 1821.500 2490.830 ;
        RECT 645.540 1903.165 645.680 2490.510 ;
        RECT 645.470 1902.795 645.750 1903.165 ;
        RECT 645.540 590.910 645.680 1902.795 ;
        RECT 870.190 600.170 870.470 604.000 ;
        RECT 869.560 600.030 870.470 600.170 ;
        RECT 869.560 590.910 869.700 600.030 ;
        RECT 870.190 600.000 870.470 600.030 ;
        RECT 645.480 590.590 645.740 590.910 ;
        RECT 869.500 590.590 869.760 590.910 ;
        RECT 593.040 36.565 593.300 36.710 ;
        RECT 389.260 36.050 389.520 36.370 ;
        RECT 593.030 36.195 593.310 36.565 ;
        RECT 617.870 36.195 618.150 36.565 ;
        RECT 389.320 2.400 389.460 36.050 ;
        RECT 617.940 36.030 618.080 36.195 ;
        RECT 645.540 36.030 645.680 590.590 ;
        RECT 617.880 35.710 618.140 36.030 ;
        RECT 645.480 35.710 645.740 36.030 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 645.470 1902.840 645.750 1903.120 ;
        RECT 593.030 36.240 593.310 36.520 ;
        RECT 617.870 36.240 618.150 36.520 ;
      LAYER met3 ;
        RECT 627.030 1903.130 631.030 1903.280 ;
        RECT 645.445 1903.130 645.775 1903.145 ;
        RECT 627.030 1902.830 645.775 1903.130 ;
        RECT 627.030 1902.680 631.030 1902.830 ;
        RECT 645.445 1902.815 645.775 1902.830 ;
        RECT 593.005 36.530 593.335 36.545 ;
        RECT 617.845 36.530 618.175 36.545 ;
        RECT 593.005 36.230 618.175 36.530 ;
        RECT 593.005 36.215 593.335 36.230 ;
        RECT 617.845 36.215 618.175 36.230 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.590 2487.680 419.910 2487.740 ;
        RECT 635.330 2487.680 635.650 2487.740 ;
        RECT 1800.050 2487.680 1800.370 2487.740 ;
        RECT 419.590 2487.540 1800.370 2487.680 ;
        RECT 419.590 2487.480 419.910 2487.540 ;
        RECT 635.330 2487.480 635.650 2487.540 ;
        RECT 1800.050 2487.480 1800.370 2487.540 ;
        RECT 564.030 1689.700 564.350 1689.760 ;
        RECT 565.410 1689.700 565.730 1689.760 ;
        RECT 635.330 1689.700 635.650 1689.760 ;
        RECT 564.030 1689.560 635.650 1689.700 ;
        RECT 564.030 1689.500 564.350 1689.560 ;
        RECT 565.410 1689.500 565.730 1689.560 ;
        RECT 635.330 1689.500 635.650 1689.560 ;
        RECT 565.410 591.500 565.730 591.560 ;
        RECT 878.210 591.500 878.530 591.560 ;
        RECT 565.410 591.360 878.530 591.500 ;
        RECT 565.410 591.300 565.730 591.360 ;
        RECT 878.210 591.300 878.530 591.360 ;
        RECT 506.990 589.800 507.310 589.860 ;
        RECT 483.160 589.660 507.310 589.800 ;
        RECT 413.610 589.120 413.930 589.180 ;
        RECT 483.160 589.120 483.300 589.660 ;
        RECT 506.990 589.600 507.310 589.660 ;
        RECT 413.610 588.980 483.300 589.120 ;
        RECT 413.610 588.920 413.930 588.980 ;
        RECT 506.990 588.780 507.310 588.840 ;
        RECT 565.410 588.780 565.730 588.840 ;
        RECT 506.990 588.640 565.730 588.780 ;
        RECT 506.990 588.580 507.310 588.640 ;
        RECT 565.410 588.580 565.730 588.640 ;
        RECT 407.170 16.220 407.490 16.280 ;
        RECT 413.610 16.220 413.930 16.280 ;
        RECT 407.170 16.080 413.930 16.220 ;
        RECT 407.170 16.020 407.490 16.080 ;
        RECT 413.610 16.020 413.930 16.080 ;
      LAYER via ;
        RECT 419.620 2487.480 419.880 2487.740 ;
        RECT 635.360 2487.480 635.620 2487.740 ;
        RECT 1800.080 2487.480 1800.340 2487.740 ;
        RECT 564.060 1689.500 564.320 1689.760 ;
        RECT 565.440 1689.500 565.700 1689.760 ;
        RECT 635.360 1689.500 635.620 1689.760 ;
        RECT 565.440 591.300 565.700 591.560 ;
        RECT 878.240 591.300 878.500 591.560 ;
        RECT 413.640 588.920 413.900 589.180 ;
        RECT 507.020 589.600 507.280 589.860 ;
        RECT 507.020 588.580 507.280 588.840 ;
        RECT 565.440 588.580 565.700 588.840 ;
        RECT 407.200 16.020 407.460 16.280 ;
        RECT 413.640 16.020 413.900 16.280 ;
      LAYER met2 ;
        RECT 419.610 2643.315 419.890 2643.685 ;
        RECT 419.680 2487.770 419.820 2643.315 ;
        RECT 1800.010 2500.000 1800.290 2504.000 ;
        RECT 1800.140 2487.770 1800.280 2500.000 ;
        RECT 419.620 2487.450 419.880 2487.770 ;
        RECT 635.360 2487.450 635.620 2487.770 ;
        RECT 1800.080 2487.450 1800.340 2487.770 ;
        RECT 562.490 1700.410 562.770 1704.000 ;
        RECT 562.490 1700.270 564.260 1700.410 ;
        RECT 562.490 1700.000 562.770 1700.270 ;
        RECT 564.120 1689.790 564.260 1700.270 ;
        RECT 635.420 1689.790 635.560 2487.450 ;
        RECT 564.060 1689.470 564.320 1689.790 ;
        RECT 565.440 1689.470 565.700 1689.790 ;
        RECT 635.360 1689.470 635.620 1689.790 ;
        RECT 565.500 591.590 565.640 1689.470 ;
        RECT 879.390 600.170 879.670 604.000 ;
        RECT 878.300 600.030 879.670 600.170 ;
        RECT 878.300 591.590 878.440 600.030 ;
        RECT 879.390 600.000 879.670 600.030 ;
        RECT 565.440 591.270 565.700 591.590 ;
        RECT 878.240 591.270 878.500 591.590 ;
        RECT 507.020 589.570 507.280 589.890 ;
        RECT 413.640 588.890 413.900 589.210 ;
        RECT 413.700 16.310 413.840 588.890 ;
        RECT 507.080 588.870 507.220 589.570 ;
        RECT 565.500 588.870 565.640 591.270 ;
        RECT 507.020 588.550 507.280 588.870 ;
        RECT 565.440 588.550 565.700 588.870 ;
        RECT 407.200 15.990 407.460 16.310 ;
        RECT 413.640 15.990 413.900 16.310 ;
        RECT 407.260 2.400 407.400 15.990 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 419.610 2643.360 419.890 2643.640 ;
      LAYER met3 ;
        RECT 430.000 2646.560 434.000 2646.880 ;
        RECT 429.950 2646.280 434.000 2646.560 ;
        RECT 419.585 2643.650 419.915 2643.665 ;
        RECT 429.950 2643.650 430.250 2646.280 ;
        RECT 419.585 2643.350 430.250 2643.650 ;
        RECT 419.585 2643.335 419.915 2643.350 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1575.110 2898.400 1575.430 2898.460 ;
        RECT 1577.870 2898.400 1578.190 2898.460 ;
        RECT 1575.110 2898.260 1578.190 2898.400 ;
        RECT 1575.110 2898.200 1575.430 2898.260 ;
        RECT 1577.870 2898.200 1578.190 2898.260 ;
        RECT 1575.110 2896.500 1575.430 2896.760 ;
        RECT 1577.870 2896.500 1578.190 2896.760 ;
        RECT 1683.210 2896.500 1683.530 2896.760 ;
        RECT 1575.200 2895.000 1575.340 2896.500 ;
        RECT 1575.200 2894.860 1576.260 2895.000 ;
        RECT 1576.120 2894.320 1576.260 2894.860 ;
        RECT 1575.200 2894.180 1576.260 2894.320 ;
        RECT 618.860 2891.800 1476.900 2891.940 ;
        RECT 596.690 2891.260 597.010 2891.320 ;
        RECT 618.860 2891.260 619.000 2891.800 ;
        RECT 596.690 2891.120 619.000 2891.260 ;
        RECT 596.690 2891.060 597.010 2891.120 ;
        RECT 1476.760 2890.240 1476.900 2891.800 ;
        RECT 1529.660 2891.800 1545.900 2891.940 ;
        RECT 1501.970 2891.260 1502.290 2891.320 ;
        RECT 1529.660 2891.260 1529.800 2891.800 ;
        RECT 1501.970 2891.120 1529.800 2891.260 ;
        RECT 1545.760 2891.260 1545.900 2891.800 ;
        RECT 1575.200 2891.260 1575.340 2894.180 ;
        RECT 1545.760 2891.120 1546.820 2891.260 ;
        RECT 1501.970 2891.060 1502.290 2891.120 ;
        RECT 1546.680 2890.920 1546.820 2891.120 ;
        RECT 1547.140 2891.120 1575.340 2891.260 ;
        RECT 1547.140 2890.920 1547.280 2891.120 ;
        RECT 1546.680 2890.780 1547.280 2890.920 ;
        RECT 1501.970 2890.240 1502.290 2890.300 ;
        RECT 1476.760 2890.100 1502.290 2890.240 ;
        RECT 1577.960 2890.240 1578.100 2896.500 ;
        RECT 1683.300 2890.240 1683.440 2896.500 ;
        RECT 1577.960 2890.100 1683.440 2890.240 ;
        RECT 1501.970 2890.040 1502.290 2890.100 ;
        RECT 589.790 2649.520 590.110 2649.580 ;
        RECT 596.690 2649.520 597.010 2649.580 ;
        RECT 589.790 2649.380 597.010 2649.520 ;
        RECT 589.790 2649.320 590.110 2649.380 ;
        RECT 596.690 2649.320 597.010 2649.380 ;
        RECT 349.670 1983.800 349.990 1983.860 ;
        RECT 589.790 1983.800 590.110 1983.860 ;
        RECT 632.570 1983.800 632.890 1983.860 ;
        RECT 349.670 1983.660 632.890 1983.800 ;
        RECT 349.670 1983.600 349.990 1983.660 ;
        RECT 589.790 1983.600 590.110 1983.660 ;
        RECT 632.570 1983.600 632.890 1983.660 ;
        RECT 632.570 1921.580 632.890 1921.640 ;
        RECT 703.870 1921.580 704.190 1921.640 ;
        RECT 632.570 1921.440 704.190 1921.580 ;
        RECT 632.570 1921.380 632.890 1921.440 ;
        RECT 703.870 1921.380 704.190 1921.440 ;
        RECT 703.870 1702.960 704.190 1703.020 ;
        RECT 1918.270 1702.960 1918.590 1703.020 ;
        RECT 703.870 1702.820 1918.590 1702.960 ;
        RECT 703.870 1702.760 704.190 1702.820 ;
        RECT 1918.270 1702.760 1918.590 1702.820 ;
        RECT 653.730 1700.920 654.050 1700.980 ;
        RECT 703.870 1700.920 704.190 1700.980 ;
        RECT 653.730 1700.780 704.190 1700.920 ;
        RECT 653.730 1700.720 654.050 1700.780 ;
        RECT 703.870 1700.720 704.190 1700.780 ;
        RECT 653.730 594.900 654.050 594.960 ;
        RECT 703.870 594.900 704.190 594.960 ;
        RECT 653.730 594.760 704.190 594.900 ;
        RECT 653.730 594.700 654.050 594.760 ;
        RECT 703.870 594.700 704.190 594.760 ;
        RECT 704.790 497.320 705.110 497.380 ;
        RECT 704.420 497.180 705.110 497.320 ;
        RECT 704.420 497.040 704.560 497.180 ;
        RECT 704.790 497.120 705.110 497.180 ;
        RECT 704.330 496.780 704.650 497.040 ;
        RECT 703.410 475.900 703.730 475.960 ;
        RECT 704.330 475.900 704.650 475.960 ;
        RECT 703.410 475.760 704.650 475.900 ;
        RECT 703.410 475.700 703.730 475.760 ;
        RECT 704.330 475.700 704.650 475.760 ;
        RECT 703.410 428.300 703.730 428.360 ;
        RECT 704.790 428.300 705.110 428.360 ;
        RECT 703.410 428.160 705.110 428.300 ;
        RECT 703.410 428.100 703.730 428.160 ;
        RECT 704.790 428.100 705.110 428.160 ;
        RECT 704.790 427.620 705.110 427.680 ;
        RECT 705.250 427.620 705.570 427.680 ;
        RECT 704.790 427.480 705.570 427.620 ;
        RECT 704.790 427.420 705.110 427.480 ;
        RECT 705.250 427.420 705.570 427.480 ;
        RECT 704.330 379.680 704.650 379.740 ;
        RECT 705.250 379.680 705.570 379.740 ;
        RECT 704.330 379.540 705.570 379.680 ;
        RECT 704.330 379.480 704.650 379.540 ;
        RECT 705.250 379.480 705.570 379.540 ;
        RECT 704.330 379.000 704.650 379.060 ;
        RECT 705.250 379.000 705.570 379.060 ;
        RECT 704.330 378.860 705.570 379.000 ;
        RECT 704.330 378.800 704.650 378.860 ;
        RECT 705.250 378.800 705.570 378.860 ;
        RECT 704.330 289.920 704.650 289.980 ;
        RECT 705.250 289.920 705.570 289.980 ;
        RECT 704.330 289.780 705.570 289.920 ;
        RECT 704.330 289.720 704.650 289.780 ;
        RECT 705.250 289.720 705.570 289.780 ;
        RECT 704.790 241.640 705.110 241.700 ;
        RECT 706.170 241.640 706.490 241.700 ;
        RECT 704.790 241.500 706.490 241.640 ;
        RECT 704.790 241.440 705.110 241.500 ;
        RECT 706.170 241.440 706.490 241.500 ;
        RECT 704.330 193.360 704.650 193.420 ;
        RECT 705.250 193.360 705.570 193.420 ;
        RECT 704.330 193.220 705.570 193.360 ;
        RECT 704.330 193.160 704.650 193.220 ;
        RECT 705.250 193.160 705.570 193.220 ;
        RECT 703.410 144.740 703.730 144.800 ;
        RECT 704.790 144.740 705.110 144.800 ;
        RECT 703.410 144.600 705.110 144.740 ;
        RECT 703.410 144.540 703.730 144.600 ;
        RECT 704.790 144.540 705.110 144.600 ;
        RECT 703.410 97.140 703.730 97.200 ;
        RECT 704.330 97.140 704.650 97.200 ;
        RECT 703.410 97.000 704.650 97.140 ;
        RECT 703.410 96.940 703.730 97.000 ;
        RECT 704.330 96.940 704.650 97.000 ;
        RECT 703.410 96.460 703.730 96.520 ;
        RECT 704.330 96.460 704.650 96.520 ;
        RECT 703.410 96.320 704.650 96.460 ;
        RECT 703.410 96.260 703.730 96.320 ;
        RECT 704.330 96.260 704.650 96.320 ;
        RECT 703.410 48.520 703.730 48.580 ;
        RECT 705.250 48.520 705.570 48.580 ;
        RECT 703.410 48.380 705.570 48.520 ;
        RECT 703.410 48.320 703.730 48.380 ;
        RECT 705.250 48.320 705.570 48.380 ;
        RECT 68.150 39.680 68.470 39.740 ;
        RECT 705.250 39.680 705.570 39.740 ;
        RECT 68.150 39.540 705.570 39.680 ;
        RECT 68.150 39.480 68.470 39.540 ;
        RECT 705.250 39.480 705.570 39.540 ;
      LAYER via ;
        RECT 1575.140 2898.200 1575.400 2898.460 ;
        RECT 1577.900 2898.200 1578.160 2898.460 ;
        RECT 1575.140 2896.500 1575.400 2896.760 ;
        RECT 1577.900 2896.500 1578.160 2896.760 ;
        RECT 1683.240 2896.500 1683.500 2896.760 ;
        RECT 596.720 2891.060 596.980 2891.320 ;
        RECT 1502.000 2891.060 1502.260 2891.320 ;
        RECT 1502.000 2890.040 1502.260 2890.300 ;
        RECT 589.820 2649.320 590.080 2649.580 ;
        RECT 596.720 2649.320 596.980 2649.580 ;
        RECT 349.700 1983.600 349.960 1983.860 ;
        RECT 589.820 1983.600 590.080 1983.860 ;
        RECT 632.600 1983.600 632.860 1983.860 ;
        RECT 632.600 1921.380 632.860 1921.640 ;
        RECT 703.900 1921.380 704.160 1921.640 ;
        RECT 703.900 1702.760 704.160 1703.020 ;
        RECT 1918.300 1702.760 1918.560 1703.020 ;
        RECT 653.760 1700.720 654.020 1700.980 ;
        RECT 703.900 1700.720 704.160 1700.980 ;
        RECT 653.760 594.700 654.020 594.960 ;
        RECT 703.900 594.700 704.160 594.960 ;
        RECT 704.820 497.120 705.080 497.380 ;
        RECT 704.360 496.780 704.620 497.040 ;
        RECT 703.440 475.700 703.700 475.960 ;
        RECT 704.360 475.700 704.620 475.960 ;
        RECT 703.440 428.100 703.700 428.360 ;
        RECT 704.820 428.100 705.080 428.360 ;
        RECT 704.820 427.420 705.080 427.680 ;
        RECT 705.280 427.420 705.540 427.680 ;
        RECT 704.360 379.480 704.620 379.740 ;
        RECT 705.280 379.480 705.540 379.740 ;
        RECT 704.360 378.800 704.620 379.060 ;
        RECT 705.280 378.800 705.540 379.060 ;
        RECT 704.360 289.720 704.620 289.980 ;
        RECT 705.280 289.720 705.540 289.980 ;
        RECT 704.820 241.440 705.080 241.700 ;
        RECT 706.200 241.440 706.460 241.700 ;
        RECT 704.360 193.160 704.620 193.420 ;
        RECT 705.280 193.160 705.540 193.420 ;
        RECT 703.440 144.540 703.700 144.800 ;
        RECT 704.820 144.540 705.080 144.800 ;
        RECT 703.440 96.940 703.700 97.200 ;
        RECT 704.360 96.940 704.620 97.200 ;
        RECT 703.440 96.260 703.700 96.520 ;
        RECT 704.360 96.260 704.620 96.520 ;
        RECT 703.440 48.320 703.700 48.580 ;
        RECT 705.280 48.320 705.540 48.580 ;
        RECT 68.180 39.480 68.440 39.740 ;
        RECT 705.280 39.480 705.540 39.740 ;
      LAYER met2 ;
        RECT 1575.140 2898.170 1575.400 2898.490 ;
        RECT 1577.900 2898.170 1578.160 2898.490 ;
        RECT 1575.200 2896.790 1575.340 2898.170 ;
        RECT 1577.960 2896.790 1578.100 2898.170 ;
        RECT 1575.140 2896.470 1575.400 2896.790 ;
        RECT 1577.900 2896.470 1578.160 2896.790 ;
        RECT 1683.240 2896.530 1683.500 2896.790 ;
        RECT 1684.090 2896.530 1684.370 2900.055 ;
        RECT 1683.240 2896.470 1684.370 2896.530 ;
        RECT 1683.300 2896.390 1684.370 2896.470 ;
        RECT 1684.090 2896.055 1684.370 2896.390 ;
        RECT 596.720 2891.030 596.980 2891.350 ;
        RECT 1502.000 2891.030 1502.260 2891.350 ;
        RECT 596.780 2649.610 596.920 2891.030 ;
        RECT 1502.060 2890.330 1502.200 2891.030 ;
        RECT 1502.000 2890.010 1502.260 2890.330 ;
        RECT 589.820 2649.290 590.080 2649.610 ;
        RECT 596.720 2649.290 596.980 2649.610 ;
        RECT 589.880 2647.765 590.020 2649.290 ;
        RECT 589.810 2647.395 590.090 2647.765 ;
        RECT 589.880 1983.890 590.020 2647.395 ;
        RECT 349.700 1983.570 349.960 1983.890 ;
        RECT 589.820 1983.570 590.080 1983.890 ;
        RECT 632.600 1983.570 632.860 1983.890 ;
        RECT 349.760 1926.285 349.900 1983.570 ;
        RECT 349.690 1925.915 349.970 1926.285 ;
        RECT 632.660 1921.670 632.800 1983.570 ;
        RECT 632.600 1921.350 632.860 1921.670 ;
        RECT 703.900 1921.350 704.160 1921.670 ;
        RECT 703.960 1703.050 704.100 1921.350 ;
        RECT 1922.850 1750.730 1923.130 1754.000 ;
        RECT 1918.360 1750.590 1923.130 1750.730 ;
        RECT 1918.360 1703.050 1918.500 1750.590 ;
        RECT 1922.850 1750.000 1923.130 1750.590 ;
        RECT 703.900 1702.730 704.160 1703.050 ;
        RECT 1918.300 1702.730 1918.560 1703.050 ;
        RECT 703.960 1701.010 704.100 1702.730 ;
        RECT 653.760 1700.690 654.020 1701.010 ;
        RECT 703.900 1700.690 704.160 1701.010 ;
        RECT 653.820 594.990 653.960 1700.690 ;
        RECT 705.050 600.170 705.330 604.000 ;
        RECT 703.960 600.030 705.330 600.170 ;
        RECT 703.960 594.990 704.100 600.030 ;
        RECT 705.050 600.000 705.330 600.030 ;
        RECT 653.760 594.670 654.020 594.990 ;
        RECT 703.900 594.670 704.160 594.990 ;
        RECT 703.960 569.570 704.100 594.670 ;
        RECT 703.960 569.430 705.020 569.570 ;
        RECT 704.880 497.410 705.020 569.430 ;
        RECT 704.820 497.090 705.080 497.410 ;
        RECT 704.360 496.750 704.620 497.070 ;
        RECT 704.420 475.990 704.560 496.750 ;
        RECT 703.440 475.670 703.700 475.990 ;
        RECT 704.360 475.670 704.620 475.990 ;
        RECT 703.500 428.390 703.640 475.670 ;
        RECT 703.440 428.070 703.700 428.390 ;
        RECT 704.820 428.070 705.080 428.390 ;
        RECT 704.880 427.710 705.020 428.070 ;
        RECT 704.820 427.390 705.080 427.710 ;
        RECT 705.280 427.390 705.540 427.710 ;
        RECT 705.340 379.770 705.480 427.390 ;
        RECT 704.360 379.450 704.620 379.770 ;
        RECT 705.280 379.450 705.540 379.770 ;
        RECT 704.420 379.090 704.560 379.450 ;
        RECT 704.360 378.770 704.620 379.090 ;
        RECT 705.280 378.770 705.540 379.090 ;
        RECT 705.340 290.010 705.480 378.770 ;
        RECT 704.360 289.690 704.620 290.010 ;
        RECT 705.280 289.690 705.540 290.010 ;
        RECT 704.420 289.525 704.560 289.690 ;
        RECT 704.350 289.155 704.630 289.525 ;
        RECT 706.190 289.155 706.470 289.525 ;
        RECT 706.260 241.730 706.400 289.155 ;
        RECT 704.820 241.410 705.080 241.730 ;
        RECT 706.200 241.410 706.460 241.730 ;
        RECT 704.880 241.130 705.020 241.410 ;
        RECT 704.880 240.990 705.480 241.130 ;
        RECT 705.340 193.450 705.480 240.990 ;
        RECT 704.360 193.130 704.620 193.450 ;
        RECT 705.280 193.130 705.540 193.450 ;
        RECT 704.420 192.965 704.560 193.130 ;
        RECT 704.350 192.595 704.630 192.965 ;
        RECT 704.810 144.995 705.090 145.365 ;
        RECT 704.880 144.830 705.020 144.995 ;
        RECT 703.440 144.510 703.700 144.830 ;
        RECT 704.820 144.510 705.080 144.830 ;
        RECT 703.500 97.230 703.640 144.510 ;
        RECT 703.440 96.910 703.700 97.230 ;
        RECT 704.360 96.910 704.620 97.230 ;
        RECT 704.420 96.550 704.560 96.910 ;
        RECT 703.440 96.230 703.700 96.550 ;
        RECT 704.360 96.230 704.620 96.550 ;
        RECT 703.500 48.610 703.640 96.230 ;
        RECT 703.440 48.290 703.700 48.610 ;
        RECT 705.280 48.290 705.540 48.610 ;
        RECT 705.340 39.770 705.480 48.290 ;
        RECT 68.180 39.450 68.440 39.770 ;
        RECT 705.280 39.450 705.540 39.770 ;
        RECT 68.240 2.400 68.380 39.450 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 589.810 2647.440 590.090 2647.720 ;
        RECT 349.690 1925.960 349.970 1926.240 ;
        RECT 704.350 289.200 704.630 289.480 ;
        RECT 706.190 289.200 706.470 289.480 ;
        RECT 704.350 192.640 704.630 192.920 ;
        RECT 704.810 145.040 705.090 145.320 ;
      LAYER met3 ;
        RECT 574.800 2647.730 578.800 2648.240 ;
        RECT 589.785 2647.730 590.115 2647.745 ;
        RECT 574.800 2647.640 590.115 2647.730 ;
        RECT 578.070 2647.430 590.115 2647.640 ;
        RECT 589.785 2647.415 590.115 2647.430 ;
        RECT 349.665 1926.250 349.995 1926.265 ;
        RECT 360.000 1926.250 364.000 1926.400 ;
        RECT 349.665 1925.950 364.000 1926.250 ;
        RECT 349.665 1925.935 349.995 1925.950 ;
        RECT 360.000 1925.800 364.000 1925.950 ;
        RECT 704.325 289.490 704.655 289.505 ;
        RECT 706.165 289.490 706.495 289.505 ;
        RECT 704.325 289.190 706.495 289.490 ;
        RECT 704.325 289.175 704.655 289.190 ;
        RECT 706.165 289.175 706.495 289.190 ;
        RECT 704.325 192.940 704.655 192.945 ;
        RECT 704.070 192.930 704.655 192.940 ;
        RECT 704.070 192.630 704.880 192.930 ;
        RECT 704.070 192.620 704.655 192.630 ;
        RECT 704.325 192.615 704.655 192.620 ;
        RECT 704.070 145.330 704.450 145.340 ;
        RECT 704.785 145.330 705.115 145.345 ;
        RECT 704.070 145.030 705.115 145.330 ;
        RECT 704.070 145.020 704.450 145.030 ;
        RECT 704.785 145.015 705.115 145.030 ;
      LAYER via3 ;
        RECT 704.100 192.620 704.420 192.940 ;
        RECT 704.100 145.020 704.420 145.340 ;
      LAYER met4 ;
        RECT 704.095 192.615 704.425 192.945 ;
        RECT 704.110 145.345 704.410 192.615 ;
        RECT 704.095 145.015 704.425 145.345 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1650.550 2897.040 1650.870 2897.100 ;
        RECT 1565.080 2896.900 1650.870 2897.040 ;
        RECT 1565.080 2895.000 1565.220 2896.900 ;
        RECT 1650.550 2896.840 1650.870 2896.900 ;
        RECT 1561.860 2894.860 1565.220 2895.000 ;
        RECT 1501.970 2894.660 1502.290 2894.720 ;
        RECT 1501.970 2894.520 1539.000 2894.660 ;
        RECT 1501.970 2894.460 1502.290 2894.520 ;
        RECT 1438.030 2894.320 1438.350 2894.380 ;
        RECT 1491.850 2894.320 1492.170 2894.380 ;
        RECT 1438.030 2894.180 1492.170 2894.320 ;
        RECT 1438.030 2894.120 1438.350 2894.180 ;
        RECT 1491.850 2894.120 1492.170 2894.180 ;
        RECT 1538.860 2893.980 1539.000 2894.520 ;
        RECT 1561.860 2894.320 1562.000 2894.860 ;
        RECT 1545.760 2894.180 1562.000 2894.320 ;
        RECT 1545.760 2893.980 1545.900 2894.180 ;
        RECT 1538.860 2893.840 1545.900 2893.980 ;
        RECT 644.990 2892.620 645.310 2892.680 ;
        RECT 678.570 2892.620 678.890 2892.680 ;
        RECT 928.350 2892.620 928.670 2892.680 ;
        RECT 644.990 2892.480 676.500 2892.620 ;
        RECT 644.990 2892.420 645.310 2892.480 ;
        RECT 676.360 2892.340 676.500 2892.480 ;
        RECT 678.570 2892.480 928.670 2892.620 ;
        RECT 678.570 2892.420 678.890 2892.480 ;
        RECT 928.350 2892.420 928.670 2892.480 ;
        RECT 951.810 2892.620 952.130 2892.680 ;
        RECT 1047.030 2892.620 1047.350 2892.680 ;
        RECT 951.810 2892.480 1047.350 2892.620 ;
        RECT 951.810 2892.420 952.130 2892.480 ;
        RECT 1047.030 2892.420 1047.350 2892.480 ;
        RECT 1048.410 2892.620 1048.730 2892.680 ;
        RECT 1143.630 2892.620 1143.950 2892.680 ;
        RECT 1048.410 2892.480 1143.950 2892.620 ;
        RECT 1048.410 2892.420 1048.730 2892.480 ;
        RECT 1143.630 2892.420 1143.950 2892.480 ;
        RECT 1145.010 2892.620 1145.330 2892.680 ;
        RECT 1438.030 2892.620 1438.350 2892.680 ;
        RECT 1145.010 2892.480 1438.350 2892.620 ;
        RECT 1145.010 2892.420 1145.330 2892.480 ;
        RECT 1438.030 2892.420 1438.350 2892.480 ;
        RECT 676.270 2892.080 676.590 2892.340 ;
        RECT 1491.850 2892.280 1492.170 2892.340 ;
        RECT 1501.970 2892.280 1502.290 2892.340 ;
        RECT 1491.850 2892.140 1502.290 2892.280 ;
        RECT 1491.850 2892.080 1492.170 2892.140 ;
        RECT 1501.970 2892.080 1502.290 2892.140 ;
        RECT 586.570 2604.640 586.890 2604.700 ;
        RECT 642.230 2604.640 642.550 2604.700 ;
        RECT 644.990 2604.640 645.310 2604.700 ;
        RECT 586.570 2604.500 645.310 2604.640 ;
        RECT 586.570 2604.440 586.890 2604.500 ;
        RECT 642.230 2604.440 642.550 2604.500 ;
        RECT 644.990 2604.440 645.310 2604.500 ;
        RECT 645.910 591.160 646.230 591.220 ;
        RECT 886.950 591.160 887.270 591.220 ;
        RECT 645.910 591.020 887.270 591.160 ;
        RECT 645.910 590.960 646.230 591.020 ;
        RECT 886.950 590.960 887.270 591.020 ;
        RECT 424.650 35.940 424.970 36.000 ;
        RECT 424.650 35.800 617.620 35.940 ;
        RECT 424.650 35.740 424.970 35.800 ;
        RECT 617.480 35.600 617.620 35.800 ;
        RECT 645.910 35.600 646.230 35.660 ;
        RECT 617.480 35.460 646.230 35.600 ;
        RECT 645.910 35.400 646.230 35.460 ;
      LAYER via ;
        RECT 1650.580 2896.840 1650.840 2897.100 ;
        RECT 1502.000 2894.460 1502.260 2894.720 ;
        RECT 1438.060 2894.120 1438.320 2894.380 ;
        RECT 1491.880 2894.120 1492.140 2894.380 ;
        RECT 645.020 2892.420 645.280 2892.680 ;
        RECT 678.600 2892.420 678.860 2892.680 ;
        RECT 928.380 2892.420 928.640 2892.680 ;
        RECT 951.840 2892.420 952.100 2892.680 ;
        RECT 1047.060 2892.420 1047.320 2892.680 ;
        RECT 1048.440 2892.420 1048.700 2892.680 ;
        RECT 1143.660 2892.420 1143.920 2892.680 ;
        RECT 1145.040 2892.420 1145.300 2892.680 ;
        RECT 1438.060 2892.420 1438.320 2892.680 ;
        RECT 676.300 2892.080 676.560 2892.340 ;
        RECT 1491.880 2892.080 1492.140 2892.340 ;
        RECT 1502.000 2892.080 1502.260 2892.340 ;
        RECT 586.600 2604.440 586.860 2604.700 ;
        RECT 642.260 2604.440 642.520 2604.700 ;
        RECT 645.020 2604.440 645.280 2604.700 ;
        RECT 645.940 590.960 646.200 591.220 ;
        RECT 886.980 590.960 887.240 591.220 ;
        RECT 424.680 35.740 424.940 36.000 ;
        RECT 645.940 35.400 646.200 35.660 ;
      LAYER met2 ;
        RECT 1651.890 2897.210 1652.170 2900.055 ;
        RECT 1650.640 2897.130 1652.170 2897.210 ;
        RECT 1650.580 2897.070 1652.170 2897.130 ;
        RECT 1650.580 2896.810 1650.840 2897.070 ;
        RECT 1651.890 2896.055 1652.170 2897.070 ;
        RECT 1502.000 2894.430 1502.260 2894.750 ;
        RECT 1438.060 2894.090 1438.320 2894.410 ;
        RECT 1491.880 2894.090 1492.140 2894.410 ;
        RECT 1047.120 2893.500 1048.640 2893.640 ;
        RECT 928.370 2892.875 928.650 2893.245 ;
        RECT 951.830 2892.875 952.110 2893.245 ;
        RECT 928.440 2892.710 928.580 2892.875 ;
        RECT 951.900 2892.710 952.040 2892.875 ;
        RECT 1047.120 2892.710 1047.260 2893.500 ;
        RECT 1048.500 2892.710 1048.640 2893.500 ;
        RECT 1143.720 2893.500 1145.240 2893.640 ;
        RECT 1143.720 2892.710 1143.860 2893.500 ;
        RECT 1145.100 2892.710 1145.240 2893.500 ;
        RECT 1438.120 2892.710 1438.260 2894.090 ;
        RECT 645.020 2892.390 645.280 2892.710 ;
        RECT 678.600 2892.390 678.860 2892.710 ;
        RECT 928.380 2892.390 928.640 2892.710 ;
        RECT 951.840 2892.390 952.100 2892.710 ;
        RECT 1047.060 2892.390 1047.320 2892.710 ;
        RECT 1048.440 2892.390 1048.700 2892.710 ;
        RECT 1143.660 2892.390 1143.920 2892.710 ;
        RECT 1145.040 2892.390 1145.300 2892.710 ;
        RECT 1438.060 2892.390 1438.320 2892.710 ;
        RECT 586.590 2605.235 586.870 2605.605 ;
        RECT 586.660 2604.730 586.800 2605.235 ;
        RECT 645.080 2604.730 645.220 2892.390 ;
        RECT 676.300 2892.050 676.560 2892.370 ;
        RECT 676.360 2891.885 676.500 2892.050 ;
        RECT 678.660 2891.885 678.800 2892.390 ;
        RECT 1491.940 2892.370 1492.080 2894.090 ;
        RECT 1502.060 2892.370 1502.200 2894.430 ;
        RECT 1491.880 2892.050 1492.140 2892.370 ;
        RECT 1502.000 2892.050 1502.260 2892.370 ;
        RECT 676.290 2891.515 676.570 2891.885 ;
        RECT 678.590 2891.515 678.870 2891.885 ;
        RECT 586.600 2604.410 586.860 2604.730 ;
        RECT 642.260 2604.410 642.520 2604.730 ;
        RECT 645.020 2604.410 645.280 2604.730 ;
        RECT 642.320 1866.445 642.460 2604.410 ;
        RECT 642.250 1866.075 642.530 1866.445 ;
        RECT 645.930 1866.075 646.210 1866.445 ;
        RECT 646.000 591.250 646.140 1866.075 ;
        RECT 888.590 600.170 888.870 604.000 ;
        RECT 887.040 600.030 888.870 600.170 ;
        RECT 887.040 591.250 887.180 600.030 ;
        RECT 888.590 600.000 888.870 600.030 ;
        RECT 645.940 590.930 646.200 591.250 ;
        RECT 886.980 590.930 887.240 591.250 ;
        RECT 424.680 35.710 424.940 36.030 ;
        RECT 424.740 2.400 424.880 35.710 ;
        RECT 646.000 35.690 646.140 590.930 ;
        RECT 645.940 35.370 646.200 35.690 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 928.370 2892.920 928.650 2893.200 ;
        RECT 951.830 2892.920 952.110 2893.200 ;
        RECT 586.590 2605.280 586.870 2605.560 ;
        RECT 676.290 2891.560 676.570 2891.840 ;
        RECT 678.590 2891.560 678.870 2891.840 ;
        RECT 642.250 1866.120 642.530 1866.400 ;
        RECT 645.930 1866.120 646.210 1866.400 ;
      LAYER met3 ;
        RECT 928.345 2893.210 928.675 2893.225 ;
        RECT 951.805 2893.210 952.135 2893.225 ;
        RECT 928.345 2892.910 952.135 2893.210 ;
        RECT 928.345 2892.895 928.675 2892.910 ;
        RECT 951.805 2892.895 952.135 2892.910 ;
        RECT 676.265 2891.850 676.595 2891.865 ;
        RECT 678.565 2891.850 678.895 2891.865 ;
        RECT 676.265 2891.550 678.895 2891.850 ;
        RECT 676.265 2891.535 676.595 2891.550 ;
        RECT 678.565 2891.535 678.895 2891.550 ;
        RECT 574.800 2605.570 578.800 2606.080 ;
        RECT 586.565 2605.570 586.895 2605.585 ;
        RECT 574.800 2605.480 586.895 2605.570 ;
        RECT 578.070 2605.270 586.895 2605.480 ;
        RECT 586.565 2605.255 586.895 2605.270 ;
        RECT 627.030 1866.410 631.030 1866.560 ;
        RECT 642.225 1866.410 642.555 1866.425 ;
        RECT 645.905 1866.410 646.235 1866.425 ;
        RECT 627.030 1866.110 646.235 1866.410 ;
        RECT 627.030 1865.960 631.030 1866.110 ;
        RECT 642.225 1866.095 642.555 1866.110 ;
        RECT 645.905 1866.095 646.235 1866.110 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 426.950 2916.760 427.270 2916.820 ;
        RECT 1673.090 2916.760 1673.410 2916.820 ;
        RECT 426.950 2916.620 1673.410 2916.760 ;
        RECT 426.950 2916.560 427.270 2916.620 ;
        RECT 1673.090 2916.560 1673.410 2916.620 ;
        RECT 351.510 2622.320 351.830 2622.380 ;
        RECT 414.070 2622.320 414.390 2622.380 ;
        RECT 351.510 2622.180 414.390 2622.320 ;
        RECT 351.510 2622.120 351.830 2622.180 ;
        RECT 414.070 2622.120 414.390 2622.180 ;
        RECT 357.490 592.180 357.810 592.240 ;
        RECT 441.670 592.180 441.990 592.240 ;
        RECT 357.490 592.040 441.990 592.180 ;
        RECT 357.490 591.980 357.810 592.040 ;
        RECT 441.670 591.980 441.990 592.040 ;
        RECT 441.670 590.140 441.990 590.200 ;
        RECT 897.070 590.140 897.390 590.200 ;
        RECT 441.670 590.000 897.390 590.140 ;
        RECT 441.670 589.940 441.990 590.000 ;
        RECT 897.070 589.940 897.390 590.000 ;
      LAYER via ;
        RECT 426.980 2916.560 427.240 2916.820 ;
        RECT 1673.120 2916.560 1673.380 2916.820 ;
        RECT 351.540 2622.120 351.800 2622.380 ;
        RECT 414.100 2622.120 414.360 2622.380 ;
        RECT 357.520 591.980 357.780 592.240 ;
        RECT 441.700 591.980 441.960 592.240 ;
        RECT 441.700 589.940 441.960 590.200 ;
        RECT 897.100 589.940 897.360 590.200 ;
      LAYER met2 ;
        RECT 426.980 2916.530 427.240 2916.850 ;
        RECT 1673.120 2916.530 1673.380 2916.850 ;
        RECT 427.040 2628.045 427.180 2916.530 ;
        RECT 1673.180 2900.055 1673.320 2916.530 ;
        RECT 1673.050 2896.055 1673.330 2900.055 ;
        RECT 426.970 2627.675 427.250 2628.045 ;
        RECT 414.090 2624.275 414.370 2624.645 ;
        RECT 414.160 2622.410 414.300 2624.275 ;
        RECT 351.540 2622.090 351.800 2622.410 ;
        RECT 414.100 2622.090 414.360 2622.410 ;
        RECT 351.600 1741.325 351.740 2622.090 ;
        RECT 351.530 1740.955 351.810 1741.325 ;
        RECT 357.510 1740.955 357.790 1741.325 ;
        RECT 357.580 592.270 357.720 1740.955 ;
        RECT 897.790 600.170 898.070 604.000 ;
        RECT 897.160 600.030 898.070 600.170 ;
        RECT 357.520 591.950 357.780 592.270 ;
        RECT 441.700 591.950 441.960 592.270 ;
        RECT 441.760 590.230 441.900 591.950 ;
        RECT 897.160 590.230 897.300 600.030 ;
        RECT 897.790 600.000 898.070 600.030 ;
        RECT 441.700 589.910 441.960 590.230 ;
        RECT 897.100 589.910 897.360 590.230 ;
        RECT 441.760 17.410 441.900 589.910 ;
        RECT 441.760 17.270 442.820 17.410 ;
        RECT 442.680 2.400 442.820 17.270 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 426.970 2627.720 427.250 2628.000 ;
        RECT 414.090 2624.320 414.370 2624.600 ;
        RECT 351.530 1741.000 351.810 1741.280 ;
        RECT 357.510 1741.000 357.790 1741.280 ;
      LAYER met3 ;
        RECT 426.945 2628.010 427.275 2628.025 ;
        RECT 426.945 2627.710 430.250 2628.010 ;
        RECT 426.945 2627.695 427.275 2627.710 ;
        RECT 429.950 2625.120 430.250 2627.710 ;
        RECT 414.065 2624.610 414.395 2624.625 ;
        RECT 429.950 2624.610 434.000 2625.120 ;
        RECT 414.065 2624.520 434.000 2624.610 ;
        RECT 414.065 2624.310 430.250 2624.520 ;
        RECT 414.065 2624.295 414.395 2624.310 ;
        RECT 351.505 1741.290 351.835 1741.305 ;
        RECT 357.485 1741.290 357.815 1741.305 ;
        RECT 360.000 1741.290 364.000 1741.440 ;
        RECT 351.505 1740.990 364.000 1741.290 ;
        RECT 351.505 1740.975 351.835 1740.990 ;
        RECT 357.485 1740.975 357.815 1740.990 ;
        RECT 360.000 1740.840 364.000 1740.990 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.450 2591.040 461.770 2591.100 ;
        RECT 634.870 2591.040 635.190 2591.100 ;
        RECT 1487.250 2591.040 1487.570 2591.100 ;
        RECT 461.450 2590.900 1487.570 2591.040 ;
        RECT 461.450 2590.840 461.770 2590.900 ;
        RECT 634.870 2590.840 635.190 2590.900 ;
        RECT 1487.250 2590.840 1487.570 2590.900 ;
        RECT 489.510 1690.040 489.830 1690.100 ;
        RECT 634.870 1690.040 635.190 1690.100 ;
        RECT 489.510 1689.900 635.190 1690.040 ;
        RECT 489.510 1689.840 489.830 1689.900 ;
        RECT 634.870 1689.840 635.190 1689.900 ;
        RECT 489.510 592.860 489.830 592.920 ;
        RECT 905.350 592.860 905.670 592.920 ;
        RECT 489.510 592.720 905.670 592.860 ;
        RECT 489.510 592.660 489.830 592.720 ;
        RECT 905.350 592.660 905.670 592.720 ;
        RECT 486.290 586.740 486.610 586.800 ;
        RECT 489.510 586.740 489.830 586.800 ;
        RECT 486.290 586.600 489.830 586.740 ;
        RECT 486.290 586.540 486.610 586.600 ;
        RECT 489.510 586.540 489.830 586.600 ;
        RECT 486.290 15.880 486.610 15.940 ;
        RECT 477.640 15.740 486.610 15.880 ;
        RECT 460.530 15.540 460.850 15.600 ;
        RECT 477.640 15.540 477.780 15.740 ;
        RECT 486.290 15.680 486.610 15.740 ;
        RECT 460.530 15.400 477.780 15.540 ;
        RECT 460.530 15.340 460.850 15.400 ;
      LAYER via ;
        RECT 461.480 2590.840 461.740 2591.100 ;
        RECT 634.900 2590.840 635.160 2591.100 ;
        RECT 1487.280 2590.840 1487.540 2591.100 ;
        RECT 489.540 1689.840 489.800 1690.100 ;
        RECT 634.900 1689.840 635.160 1690.100 ;
        RECT 489.540 592.660 489.800 592.920 ;
        RECT 905.380 592.660 905.640 592.920 ;
        RECT 486.320 586.540 486.580 586.800 ;
        RECT 489.540 586.540 489.800 586.800 ;
        RECT 460.560 15.340 460.820 15.600 ;
        RECT 486.320 15.680 486.580 15.940 ;
      LAYER met2 ;
        RECT 1487.270 2642.635 1487.550 2643.005 ;
        RECT 461.370 2600.660 461.650 2604.000 ;
        RECT 461.370 2600.000 461.680 2600.660 ;
        RECT 461.540 2591.130 461.680 2600.000 ;
        RECT 1487.340 2591.130 1487.480 2642.635 ;
        RECT 461.480 2590.810 461.740 2591.130 ;
        RECT 634.900 2590.810 635.160 2591.130 ;
        RECT 1487.280 2590.810 1487.540 2591.130 ;
        RECT 487.970 1700.410 488.250 1704.000 ;
        RECT 487.970 1700.270 489.740 1700.410 ;
        RECT 487.970 1700.000 488.250 1700.270 ;
        RECT 489.600 1690.130 489.740 1700.270 ;
        RECT 634.960 1690.130 635.100 2590.810 ;
        RECT 489.540 1689.810 489.800 1690.130 ;
        RECT 634.900 1689.810 635.160 1690.130 ;
        RECT 489.600 592.950 489.740 1689.810 ;
        RECT 906.990 600.170 907.270 604.000 ;
        RECT 905.440 600.030 907.270 600.170 ;
        RECT 905.440 592.950 905.580 600.030 ;
        RECT 906.990 600.000 907.270 600.030 ;
        RECT 489.540 592.630 489.800 592.950 ;
        RECT 905.380 592.630 905.640 592.950 ;
        RECT 489.600 586.830 489.740 592.630 ;
        RECT 486.320 586.510 486.580 586.830 ;
        RECT 489.540 586.510 489.800 586.830 ;
        RECT 486.380 15.970 486.520 586.510 ;
        RECT 486.320 15.650 486.580 15.970 ;
        RECT 460.560 15.310 460.820 15.630 ;
        RECT 460.620 2.400 460.760 15.310 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 1487.270 2642.680 1487.550 2642.960 ;
      LAYER met3 ;
        RECT 1500.000 2645.880 1504.000 2646.160 ;
        RECT 1499.910 2645.560 1504.000 2645.880 ;
        RECT 1487.245 2642.970 1487.575 2642.985 ;
        RECT 1499.910 2642.970 1500.210 2645.560 ;
        RECT 1487.245 2642.670 1500.210 2642.970 ;
        RECT 1487.245 2642.655 1487.575 2642.670 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 646.370 2917.440 646.690 2917.500 ;
        RECT 1737.490 2917.440 1737.810 2917.500 ;
        RECT 646.370 2917.300 1737.810 2917.440 ;
        RECT 646.370 2917.240 646.690 2917.300 ;
        RECT 1737.490 2917.240 1737.810 2917.300 ;
        RECT 575.530 2769.200 575.850 2769.260 ;
        RECT 641.770 2769.200 642.090 2769.260 ;
        RECT 646.370 2769.200 646.690 2769.260 ;
        RECT 575.530 2769.060 646.690 2769.200 ;
        RECT 575.530 2769.000 575.850 2769.060 ;
        RECT 641.770 2769.000 642.090 2769.060 ;
        RECT 646.370 2769.000 646.690 2769.060 ;
        RECT 646.370 591.840 646.690 591.900 ;
        RECT 914.550 591.840 914.870 591.900 ;
        RECT 646.370 591.700 914.870 591.840 ;
        RECT 646.370 591.640 646.690 591.700 ;
        RECT 914.550 591.640 914.870 591.700 ;
        RECT 478.470 35.600 478.790 35.660 ;
        RECT 478.470 35.460 603.360 35.600 ;
        RECT 478.470 35.400 478.790 35.460 ;
        RECT 603.220 34.580 603.360 35.460 ;
        RECT 646.370 34.580 646.690 34.640 ;
        RECT 603.220 34.440 646.690 34.580 ;
        RECT 646.370 34.380 646.690 34.440 ;
      LAYER via ;
        RECT 646.400 2917.240 646.660 2917.500 ;
        RECT 1737.520 2917.240 1737.780 2917.500 ;
        RECT 575.560 2769.000 575.820 2769.260 ;
        RECT 641.800 2769.000 642.060 2769.260 ;
        RECT 646.400 2769.000 646.660 2769.260 ;
        RECT 646.400 591.640 646.660 591.900 ;
        RECT 914.580 591.640 914.840 591.900 ;
        RECT 478.500 35.400 478.760 35.660 ;
        RECT 646.400 34.380 646.660 34.640 ;
      LAYER met2 ;
        RECT 646.400 2917.210 646.660 2917.530 ;
        RECT 1737.520 2917.210 1737.780 2917.530 ;
        RECT 646.460 2769.290 646.600 2917.210 ;
        RECT 1737.580 2900.055 1737.720 2917.210 ;
        RECT 1737.450 2896.055 1737.730 2900.055 ;
        RECT 575.560 2768.970 575.820 2769.290 ;
        RECT 641.800 2768.970 642.060 2769.290 ;
        RECT 646.400 2768.970 646.660 2769.290 ;
        RECT 575.620 2759.520 575.760 2768.970 ;
        RECT 575.450 2759.100 575.760 2759.520 ;
        RECT 575.450 2755.520 575.730 2759.100 ;
        RECT 641.860 1791.645 642.000 2768.970 ;
        RECT 641.790 1791.275 642.070 1791.645 ;
        RECT 646.390 1791.275 646.670 1791.645 ;
        RECT 646.460 591.930 646.600 1791.275 ;
        RECT 916.190 600.170 916.470 604.000 ;
        RECT 914.640 600.030 916.470 600.170 ;
        RECT 914.640 591.930 914.780 600.030 ;
        RECT 916.190 600.000 916.470 600.030 ;
        RECT 646.400 591.610 646.660 591.930 ;
        RECT 914.580 591.610 914.840 591.930 ;
        RECT 478.500 35.370 478.760 35.690 ;
        RECT 478.560 2.400 478.700 35.370 ;
        RECT 646.460 34.670 646.600 591.610 ;
        RECT 646.400 34.350 646.660 34.670 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 641.790 1791.320 642.070 1791.600 ;
        RECT 646.390 1791.320 646.670 1791.600 ;
      LAYER met3 ;
        RECT 627.030 1791.610 631.030 1791.760 ;
        RECT 641.765 1791.610 642.095 1791.625 ;
        RECT 646.365 1791.610 646.695 1791.625 ;
        RECT 627.030 1791.310 646.695 1791.610 ;
        RECT 627.030 1791.160 631.030 1791.310 ;
        RECT 641.765 1791.295 642.095 1791.310 ;
        RECT 646.365 1791.295 646.695 1791.310 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 1687.320 389.550 1687.380 ;
        RECT 496.410 1687.320 496.730 1687.380 ;
        RECT 1649.170 1687.320 1649.490 1687.380 ;
        RECT 389.230 1687.180 1649.490 1687.320 ;
        RECT 389.230 1687.120 389.550 1687.180 ;
        RECT 496.410 1687.120 496.730 1687.180 ;
        RECT 1649.170 1687.120 1649.490 1687.180 ;
        RECT 489.970 15.880 490.290 15.940 ;
        RECT 496.410 15.880 496.730 15.940 ;
        RECT 489.970 15.740 496.730 15.880 ;
        RECT 489.970 15.680 490.290 15.740 ;
        RECT 496.410 15.680 496.730 15.740 ;
      LAYER via ;
        RECT 389.260 1687.120 389.520 1687.380 ;
        RECT 496.440 1687.120 496.700 1687.380 ;
        RECT 1649.200 1687.120 1649.460 1687.380 ;
        RECT 490.000 15.680 490.260 15.940 ;
        RECT 496.440 15.680 496.700 15.940 ;
      LAYER met2 ;
        RECT 1650.970 2500.090 1651.250 2504.000 ;
        RECT 1649.260 2500.000 1651.250 2500.090 ;
        RECT 1649.260 2499.950 1651.170 2500.000 ;
        RECT 387.690 1700.410 387.970 1704.000 ;
        RECT 387.690 1700.270 389.460 1700.410 ;
        RECT 387.690 1700.000 387.970 1700.270 ;
        RECT 389.320 1687.410 389.460 1700.270 ;
        RECT 1649.260 1687.410 1649.400 2499.950 ;
        RECT 389.260 1687.090 389.520 1687.410 ;
        RECT 496.440 1687.090 496.700 1687.410 ;
        RECT 1649.200 1687.090 1649.460 1687.410 ;
        RECT 496.500 593.485 496.640 1687.090 ;
        RECT 925.390 600.170 925.670 604.000 ;
        RECT 924.760 600.030 925.670 600.170 ;
        RECT 924.760 593.485 924.900 600.030 ;
        RECT 925.390 600.000 925.670 600.030 ;
        RECT 496.430 593.115 496.710 593.485 ;
        RECT 924.690 593.115 924.970 593.485 ;
        RECT 496.500 586.685 496.640 593.115 ;
        RECT 489.990 586.315 490.270 586.685 ;
        RECT 496.430 586.315 496.710 586.685 ;
        RECT 490.060 15.970 490.200 586.315 ;
        RECT 490.000 15.650 490.260 15.970 ;
        RECT 496.440 15.650 496.700 15.970 ;
        RECT 496.500 2.400 496.640 15.650 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 496.430 593.160 496.710 593.440 ;
        RECT 924.690 593.160 924.970 593.440 ;
        RECT 489.990 586.360 490.270 586.640 ;
        RECT 496.430 586.360 496.710 586.640 ;
      LAYER met3 ;
        RECT 496.405 593.450 496.735 593.465 ;
        RECT 924.665 593.450 924.995 593.465 ;
        RECT 496.405 593.150 924.995 593.450 ;
        RECT 496.405 593.135 496.735 593.150 ;
        RECT 924.665 593.135 924.995 593.150 ;
        RECT 489.965 586.650 490.295 586.665 ;
        RECT 496.405 586.650 496.735 586.665 ;
        RECT 489.965 586.350 496.735 586.650 ;
        RECT 489.965 586.335 490.295 586.350 ;
        RECT 496.405 586.335 496.735 586.350 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1499.670 2429.200 1499.990 2429.260 ;
        RECT 1502.890 2429.200 1503.210 2429.260 ;
        RECT 1499.670 2429.060 1503.210 2429.200 ;
        RECT 1499.670 2429.000 1499.990 2429.060 ;
        RECT 1502.890 2429.000 1503.210 2429.060 ;
        RECT 1498.750 2380.580 1499.070 2380.640 ;
        RECT 1499.670 2380.580 1499.990 2380.640 ;
        RECT 1498.750 2380.440 1499.990 2380.580 ;
        RECT 1498.750 2380.380 1499.070 2380.440 ;
        RECT 1499.670 2380.380 1499.990 2380.440 ;
        RECT 1499.210 2366.640 1499.530 2366.700 ;
        RECT 1499.670 2366.640 1499.990 2366.700 ;
        RECT 1499.210 2366.500 1499.990 2366.640 ;
        RECT 1499.210 2366.440 1499.530 2366.500 ;
        RECT 1499.670 2366.440 1499.990 2366.500 ;
        RECT 1499.670 2332.300 1499.990 2332.360 ;
        RECT 1499.300 2332.160 1499.990 2332.300 ;
        RECT 1499.300 2332.020 1499.440 2332.160 ;
        RECT 1499.670 2332.100 1499.990 2332.160 ;
        RECT 1499.210 2331.760 1499.530 2332.020 ;
        RECT 1498.750 2284.020 1499.070 2284.080 ;
        RECT 1499.670 2284.020 1499.990 2284.080 ;
        RECT 1498.750 2283.880 1499.990 2284.020 ;
        RECT 1498.750 2283.820 1499.070 2283.880 ;
        RECT 1499.670 2283.820 1499.990 2283.880 ;
        RECT 1499.210 2270.080 1499.530 2270.140 ;
        RECT 1499.670 2270.080 1499.990 2270.140 ;
        RECT 1499.210 2269.940 1499.990 2270.080 ;
        RECT 1499.210 2269.880 1499.530 2269.940 ;
        RECT 1499.670 2269.880 1499.990 2269.940 ;
        RECT 1499.670 2235.740 1499.990 2235.800 ;
        RECT 1499.300 2235.600 1499.990 2235.740 ;
        RECT 1499.300 2235.460 1499.440 2235.600 ;
        RECT 1499.670 2235.540 1499.990 2235.600 ;
        RECT 1499.210 2235.200 1499.530 2235.460 ;
        RECT 1498.750 2187.460 1499.070 2187.520 ;
        RECT 1499.670 2187.460 1499.990 2187.520 ;
        RECT 1498.750 2187.320 1499.990 2187.460 ;
        RECT 1498.750 2187.260 1499.070 2187.320 ;
        RECT 1499.670 2187.260 1499.990 2187.320 ;
        RECT 1499.210 2173.520 1499.530 2173.580 ;
        RECT 1499.670 2173.520 1499.990 2173.580 ;
        RECT 1499.210 2173.380 1499.990 2173.520 ;
        RECT 1499.210 2173.320 1499.530 2173.380 ;
        RECT 1499.670 2173.320 1499.990 2173.380 ;
        RECT 1499.670 2139.180 1499.990 2139.240 ;
        RECT 1499.300 2139.040 1499.990 2139.180 ;
        RECT 1499.300 2138.900 1499.440 2139.040 ;
        RECT 1499.670 2138.980 1499.990 2139.040 ;
        RECT 1499.210 2138.640 1499.530 2138.900 ;
        RECT 1498.750 2090.900 1499.070 2090.960 ;
        RECT 1499.670 2090.900 1499.990 2090.960 ;
        RECT 1498.750 2090.760 1499.990 2090.900 ;
        RECT 1498.750 2090.700 1499.070 2090.760 ;
        RECT 1499.670 2090.700 1499.990 2090.760 ;
        RECT 1499.210 2076.960 1499.530 2077.020 ;
        RECT 1500.590 2076.960 1500.910 2077.020 ;
        RECT 1499.210 2076.820 1500.910 2076.960 ;
        RECT 1499.210 2076.760 1499.530 2076.820 ;
        RECT 1500.590 2076.760 1500.910 2076.820 ;
        RECT 1499.670 2028.680 1499.990 2028.740 ;
        RECT 1500.590 2028.680 1500.910 2028.740 ;
        RECT 1499.670 2028.540 1500.910 2028.680 ;
        RECT 1499.670 2028.480 1499.990 2028.540 ;
        RECT 1500.590 2028.480 1500.910 2028.540 ;
        RECT 1499.210 1980.400 1499.530 1980.460 ;
        RECT 1499.670 1980.400 1499.990 1980.460 ;
        RECT 1499.210 1980.260 1499.990 1980.400 ;
        RECT 1499.210 1980.200 1499.530 1980.260 ;
        RECT 1499.670 1980.200 1499.990 1980.260 ;
        RECT 1499.210 1883.840 1499.530 1883.900 ;
        RECT 1499.670 1883.840 1499.990 1883.900 ;
        RECT 1499.210 1883.700 1499.990 1883.840 ;
        RECT 1499.210 1883.640 1499.530 1883.700 ;
        RECT 1499.670 1883.640 1499.990 1883.700 ;
        RECT 1499.210 1752.400 1499.530 1752.660 ;
        RECT 1499.300 1752.260 1499.440 1752.400 ;
        RECT 1499.670 1752.260 1499.990 1752.320 ;
        RECT 1499.300 1752.120 1499.990 1752.260 ;
        RECT 1499.670 1752.060 1499.990 1752.120 ;
        RECT 364.390 1688.000 364.710 1688.060 ;
        RECT 670.290 1688.000 670.610 1688.060 ;
        RECT 1499.670 1688.000 1499.990 1688.060 ;
        RECT 364.390 1687.860 1499.990 1688.000 ;
        RECT 364.390 1687.800 364.710 1687.860 ;
        RECT 670.290 1687.800 670.610 1687.860 ;
        RECT 1499.670 1687.800 1499.990 1687.860 ;
        RECT 668.910 615.300 669.230 615.360 ;
        RECT 670.290 615.300 670.610 615.360 ;
        RECT 668.910 615.160 670.610 615.300 ;
        RECT 668.910 615.100 669.230 615.160 ;
        RECT 670.290 615.100 670.610 615.160 ;
        RECT 710.400 602.580 737.220 602.720 ;
        RECT 668.910 602.380 669.230 602.440 ;
        RECT 710.400 602.380 710.540 602.580 ;
        RECT 668.910 602.240 710.540 602.380 ;
        RECT 737.080 602.380 737.220 602.580 ;
        RECT 737.080 602.240 759.300 602.380 ;
        RECT 668.910 602.180 669.230 602.240 ;
        RECT 759.160 601.760 759.300 602.240 ;
        RECT 807.000 602.240 855.900 602.380 ;
        RECT 807.000 601.760 807.140 602.240 ;
        RECT 855.760 601.760 855.900 602.240 ;
        RECT 903.600 602.240 911.560 602.380 ;
        RECT 759.070 601.500 759.390 601.760 ;
        RECT 806.910 601.500 807.230 601.760 ;
        RECT 855.670 601.500 855.990 601.760 ;
        RECT 759.070 601.020 759.390 601.080 ;
        RECT 806.910 601.020 807.230 601.080 ;
        RECT 759.070 600.880 807.230 601.020 ;
        RECT 759.070 600.820 759.390 600.880 ;
        RECT 806.910 600.820 807.230 600.880 ;
        RECT 855.670 601.020 855.990 601.080 ;
        RECT 903.600 601.020 903.740 602.240 ;
        RECT 911.420 601.700 911.560 602.240 ;
        RECT 932.950 601.700 933.270 601.760 ;
        RECT 911.420 601.560 933.270 601.700 ;
        RECT 932.950 601.500 933.270 601.560 ;
        RECT 855.670 600.880 903.740 601.020 ;
        RECT 855.670 600.820 855.990 600.880 ;
        RECT 932.030 569.400 932.350 569.460 ;
        RECT 932.950 569.400 933.270 569.460 ;
        RECT 932.030 569.260 933.270 569.400 ;
        RECT 932.030 569.200 932.350 569.260 ;
        RECT 932.950 569.200 933.270 569.260 ;
      LAYER via ;
        RECT 1499.700 2429.000 1499.960 2429.260 ;
        RECT 1502.920 2429.000 1503.180 2429.260 ;
        RECT 1498.780 2380.380 1499.040 2380.640 ;
        RECT 1499.700 2380.380 1499.960 2380.640 ;
        RECT 1499.240 2366.440 1499.500 2366.700 ;
        RECT 1499.700 2366.440 1499.960 2366.700 ;
        RECT 1499.700 2332.100 1499.960 2332.360 ;
        RECT 1499.240 2331.760 1499.500 2332.020 ;
        RECT 1498.780 2283.820 1499.040 2284.080 ;
        RECT 1499.700 2283.820 1499.960 2284.080 ;
        RECT 1499.240 2269.880 1499.500 2270.140 ;
        RECT 1499.700 2269.880 1499.960 2270.140 ;
        RECT 1499.700 2235.540 1499.960 2235.800 ;
        RECT 1499.240 2235.200 1499.500 2235.460 ;
        RECT 1498.780 2187.260 1499.040 2187.520 ;
        RECT 1499.700 2187.260 1499.960 2187.520 ;
        RECT 1499.240 2173.320 1499.500 2173.580 ;
        RECT 1499.700 2173.320 1499.960 2173.580 ;
        RECT 1499.700 2138.980 1499.960 2139.240 ;
        RECT 1499.240 2138.640 1499.500 2138.900 ;
        RECT 1498.780 2090.700 1499.040 2090.960 ;
        RECT 1499.700 2090.700 1499.960 2090.960 ;
        RECT 1499.240 2076.760 1499.500 2077.020 ;
        RECT 1500.620 2076.760 1500.880 2077.020 ;
        RECT 1499.700 2028.480 1499.960 2028.740 ;
        RECT 1500.620 2028.480 1500.880 2028.740 ;
        RECT 1499.240 1980.200 1499.500 1980.460 ;
        RECT 1499.700 1980.200 1499.960 1980.460 ;
        RECT 1499.240 1883.640 1499.500 1883.900 ;
        RECT 1499.700 1883.640 1499.960 1883.900 ;
        RECT 1499.240 1752.400 1499.500 1752.660 ;
        RECT 1499.700 1752.060 1499.960 1752.320 ;
        RECT 364.420 1687.800 364.680 1688.060 ;
        RECT 670.320 1687.800 670.580 1688.060 ;
        RECT 1499.700 1687.800 1499.960 1688.060 ;
        RECT 668.940 615.100 669.200 615.360 ;
        RECT 670.320 615.100 670.580 615.360 ;
        RECT 668.940 602.180 669.200 602.440 ;
        RECT 759.100 601.500 759.360 601.760 ;
        RECT 806.940 601.500 807.200 601.760 ;
        RECT 855.700 601.500 855.960 601.760 ;
        RECT 759.100 600.820 759.360 601.080 ;
        RECT 806.940 600.820 807.200 601.080 ;
        RECT 855.700 600.820 855.960 601.080 ;
        RECT 932.980 601.500 933.240 601.760 ;
        RECT 932.060 569.200 932.320 569.460 ;
        RECT 932.980 569.200 933.240 569.460 ;
      LAYER met2 ;
        RECT 1502.850 2500.770 1503.130 2504.000 ;
        RECT 1502.850 2500.630 1503.580 2500.770 ;
        RECT 1502.850 2500.000 1503.130 2500.630 ;
        RECT 1503.440 2476.970 1503.580 2500.630 ;
        RECT 1502.980 2476.830 1503.580 2476.970 ;
        RECT 1502.980 2429.290 1503.120 2476.830 ;
        RECT 1499.700 2428.970 1499.960 2429.290 ;
        RECT 1502.920 2428.970 1503.180 2429.290 ;
        RECT 1499.760 2380.670 1499.900 2428.970 ;
        RECT 1498.780 2380.410 1499.040 2380.670 ;
        RECT 1498.780 2380.350 1499.440 2380.410 ;
        RECT 1499.700 2380.350 1499.960 2380.670 ;
        RECT 1498.840 2380.270 1499.440 2380.350 ;
        RECT 1499.300 2366.730 1499.440 2380.270 ;
        RECT 1499.240 2366.410 1499.500 2366.730 ;
        RECT 1499.700 2366.410 1499.960 2366.730 ;
        RECT 1499.760 2332.390 1499.900 2366.410 ;
        RECT 1499.700 2332.070 1499.960 2332.390 ;
        RECT 1499.240 2331.730 1499.500 2332.050 ;
        RECT 1499.300 2318.530 1499.440 2331.730 ;
        RECT 1499.300 2318.390 1499.900 2318.530 ;
        RECT 1499.760 2284.110 1499.900 2318.390 ;
        RECT 1498.780 2283.850 1499.040 2284.110 ;
        RECT 1498.780 2283.790 1499.440 2283.850 ;
        RECT 1499.700 2283.790 1499.960 2284.110 ;
        RECT 1498.840 2283.710 1499.440 2283.790 ;
        RECT 1499.300 2270.170 1499.440 2283.710 ;
        RECT 1499.240 2269.850 1499.500 2270.170 ;
        RECT 1499.700 2269.850 1499.960 2270.170 ;
        RECT 1499.760 2235.830 1499.900 2269.850 ;
        RECT 1499.700 2235.510 1499.960 2235.830 ;
        RECT 1499.240 2235.170 1499.500 2235.490 ;
        RECT 1499.300 2221.970 1499.440 2235.170 ;
        RECT 1499.300 2221.830 1499.900 2221.970 ;
        RECT 1499.760 2187.550 1499.900 2221.830 ;
        RECT 1498.780 2187.290 1499.040 2187.550 ;
        RECT 1498.780 2187.230 1499.440 2187.290 ;
        RECT 1499.700 2187.230 1499.960 2187.550 ;
        RECT 1498.840 2187.150 1499.440 2187.230 ;
        RECT 1499.300 2173.610 1499.440 2187.150 ;
        RECT 1499.240 2173.290 1499.500 2173.610 ;
        RECT 1499.700 2173.290 1499.960 2173.610 ;
        RECT 1499.760 2139.270 1499.900 2173.290 ;
        RECT 1499.700 2138.950 1499.960 2139.270 ;
        RECT 1499.240 2138.610 1499.500 2138.930 ;
        RECT 1499.300 2125.410 1499.440 2138.610 ;
        RECT 1499.300 2125.270 1499.900 2125.410 ;
        RECT 1499.760 2090.990 1499.900 2125.270 ;
        RECT 1498.780 2090.730 1499.040 2090.990 ;
        RECT 1498.780 2090.670 1499.440 2090.730 ;
        RECT 1499.700 2090.670 1499.960 2090.990 ;
        RECT 1498.840 2090.590 1499.440 2090.670 ;
        RECT 1499.300 2077.050 1499.440 2090.590 ;
        RECT 1499.240 2076.730 1499.500 2077.050 ;
        RECT 1500.620 2076.730 1500.880 2077.050 ;
        RECT 1500.680 2028.770 1500.820 2076.730 ;
        RECT 1499.700 2028.450 1499.960 2028.770 ;
        RECT 1500.620 2028.450 1500.880 2028.770 ;
        RECT 1499.760 1980.490 1499.900 2028.450 ;
        RECT 1499.240 1980.170 1499.500 1980.490 ;
        RECT 1499.700 1980.170 1499.960 1980.490 ;
        RECT 1499.300 1945.890 1499.440 1980.170 ;
        RECT 1499.300 1945.750 1499.900 1945.890 ;
        RECT 1499.760 1883.930 1499.900 1945.750 ;
        RECT 1499.240 1883.610 1499.500 1883.930 ;
        RECT 1499.700 1883.610 1499.960 1883.930 ;
        RECT 1499.300 1849.330 1499.440 1883.610 ;
        RECT 1499.300 1849.190 1499.900 1849.330 ;
        RECT 1499.760 1801.050 1499.900 1849.190 ;
        RECT 1498.840 1800.910 1499.900 1801.050 ;
        RECT 1498.840 1800.370 1498.980 1800.910 ;
        RECT 1498.840 1800.230 1499.440 1800.370 ;
        RECT 1499.300 1752.690 1499.440 1800.230 ;
        RECT 1499.240 1752.370 1499.500 1752.690 ;
        RECT 1499.700 1752.030 1499.960 1752.350 ;
        RECT 362.850 1700.410 363.130 1704.000 ;
        RECT 362.850 1700.270 364.620 1700.410 ;
        RECT 362.850 1700.000 363.130 1700.270 ;
        RECT 364.480 1688.090 364.620 1700.270 ;
        RECT 1499.760 1688.090 1499.900 1752.030 ;
        RECT 364.420 1687.770 364.680 1688.090 ;
        RECT 670.320 1687.770 670.580 1688.090 ;
        RECT 1499.700 1687.770 1499.960 1688.090 ;
        RECT 670.380 615.390 670.520 1687.770 ;
        RECT 668.940 615.070 669.200 615.390 ;
        RECT 670.320 615.070 670.580 615.390 ;
        RECT 669.000 602.470 669.140 615.070 ;
        RECT 668.940 602.150 669.200 602.470 ;
        RECT 759.100 601.470 759.360 601.790 ;
        RECT 806.940 601.470 807.200 601.790 ;
        RECT 855.700 601.470 855.960 601.790 ;
        RECT 932.980 601.530 933.240 601.790 ;
        RECT 934.590 601.530 934.870 604.000 ;
        RECT 932.980 601.470 934.870 601.530 ;
        RECT 759.160 601.110 759.300 601.470 ;
        RECT 807.000 601.110 807.140 601.470 ;
        RECT 855.760 601.110 855.900 601.470 ;
        RECT 933.040 601.390 934.870 601.470 ;
        RECT 759.100 600.790 759.360 601.110 ;
        RECT 806.940 600.790 807.200 601.110 ;
        RECT 855.700 600.790 855.960 601.110 ;
        RECT 933.040 569.490 933.180 601.390 ;
        RECT 934.590 600.000 934.870 601.390 ;
        RECT 932.060 569.170 932.320 569.490 ;
        RECT 932.980 569.170 933.240 569.490 ;
        RECT 932.120 31.125 932.260 569.170 ;
        RECT 513.910 30.755 514.190 31.125 ;
        RECT 932.050 30.755 932.330 31.125 ;
        RECT 513.980 2.400 514.120 30.755 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 513.910 30.800 514.190 31.080 ;
        RECT 932.050 30.800 932.330 31.080 ;
      LAYER met3 ;
        RECT 513.885 31.090 514.215 31.105 ;
        RECT 932.025 31.090 932.355 31.105 ;
        RECT 513.885 30.790 932.355 31.090 ;
        RECT 513.885 30.775 514.215 30.790 ;
        RECT 932.025 30.775 932.355 30.790 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 665.230 2039.560 665.550 2039.620 ;
        RECT 1903.090 2039.560 1903.410 2039.620 ;
        RECT 665.230 2039.420 1903.410 2039.560 ;
        RECT 665.230 2039.360 665.550 2039.420 ;
        RECT 1903.090 2039.360 1903.410 2039.420 ;
        RECT 664.310 2021.880 664.630 2021.940 ;
        RECT 665.230 2021.880 665.550 2021.940 ;
        RECT 664.310 2021.740 665.550 2021.880 ;
        RECT 664.310 2021.680 664.630 2021.740 ;
        RECT 665.230 2021.680 665.550 2021.740 ;
        RECT 663.390 1994.000 663.710 1994.060 ;
        RECT 664.310 1994.000 664.630 1994.060 ;
        RECT 663.390 1993.860 664.630 1994.000 ;
        RECT 663.390 1993.800 663.710 1993.860 ;
        RECT 664.310 1993.800 664.630 1993.860 ;
        RECT 662.010 1973.260 662.330 1973.320 ;
        RECT 664.310 1973.260 664.630 1973.320 ;
        RECT 662.010 1973.120 664.630 1973.260 ;
        RECT 662.010 1973.060 662.330 1973.120 ;
        RECT 664.310 1973.060 664.630 1973.120 ;
        RECT 662.010 1897.440 662.330 1897.500 ;
        RECT 663.390 1897.440 663.710 1897.500 ;
        RECT 662.010 1897.300 663.710 1897.440 ;
        RECT 662.010 1897.240 662.330 1897.300 ;
        RECT 663.390 1897.240 663.710 1897.300 ;
        RECT 663.850 1780.480 664.170 1780.540 ;
        RECT 664.310 1780.480 664.630 1780.540 ;
        RECT 663.850 1780.340 664.630 1780.480 ;
        RECT 663.850 1780.280 664.170 1780.340 ;
        RECT 664.310 1780.280 664.630 1780.340 ;
        RECT 663.850 1752.940 664.170 1753.000 ;
        RECT 663.480 1752.800 664.170 1752.940 ;
        RECT 663.480 1752.660 663.620 1752.800 ;
        RECT 663.850 1752.740 664.170 1752.800 ;
        RECT 663.390 1752.400 663.710 1752.660 ;
        RECT 663.390 1541.460 663.710 1541.520 ;
        RECT 664.310 1541.460 664.630 1541.520 ;
        RECT 663.390 1541.320 664.630 1541.460 ;
        RECT 663.390 1541.260 663.710 1541.320 ;
        RECT 664.310 1541.260 664.630 1541.320 ;
        RECT 663.390 1480.600 663.710 1480.660 ;
        RECT 664.310 1480.600 664.630 1480.660 ;
        RECT 663.390 1480.460 664.630 1480.600 ;
        RECT 663.390 1480.400 663.710 1480.460 ;
        RECT 664.310 1480.400 664.630 1480.460 ;
        RECT 663.390 1444.900 663.710 1444.960 ;
        RECT 664.310 1444.900 664.630 1444.960 ;
        RECT 663.390 1444.760 664.630 1444.900 ;
        RECT 663.390 1444.700 663.710 1444.760 ;
        RECT 664.310 1444.700 664.630 1444.760 ;
        RECT 664.310 1390.500 664.630 1390.560 ;
        RECT 667.530 1390.500 667.850 1390.560 ;
        RECT 664.310 1390.360 667.850 1390.500 ;
        RECT 664.310 1390.300 664.630 1390.360 ;
        RECT 667.530 1390.300 667.850 1390.360 ;
        RECT 664.310 1342.220 664.630 1342.280 ;
        RECT 667.530 1342.220 667.850 1342.280 ;
        RECT 664.310 1342.080 667.850 1342.220 ;
        RECT 664.310 1342.020 664.630 1342.080 ;
        RECT 667.530 1342.020 667.850 1342.080 ;
        RECT 664.310 1293.940 664.630 1294.000 ;
        RECT 667.530 1293.940 667.850 1294.000 ;
        RECT 664.310 1293.800 667.850 1293.940 ;
        RECT 664.310 1293.740 664.630 1293.800 ;
        RECT 667.530 1293.740 667.850 1293.800 ;
        RECT 664.310 1245.660 664.630 1245.720 ;
        RECT 667.530 1245.660 667.850 1245.720 ;
        RECT 664.310 1245.520 667.850 1245.660 ;
        RECT 664.310 1245.460 664.630 1245.520 ;
        RECT 667.530 1245.460 667.850 1245.520 ;
        RECT 664.310 1197.380 664.630 1197.440 ;
        RECT 667.530 1197.380 667.850 1197.440 ;
        RECT 664.310 1197.240 667.850 1197.380 ;
        RECT 664.310 1197.180 664.630 1197.240 ;
        RECT 667.530 1197.180 667.850 1197.240 ;
        RECT 664.310 1148.760 664.630 1148.820 ;
        RECT 667.530 1148.760 667.850 1148.820 ;
        RECT 664.310 1148.620 667.850 1148.760 ;
        RECT 664.310 1148.560 664.630 1148.620 ;
        RECT 667.530 1148.560 667.850 1148.620 ;
        RECT 664.310 1100.480 664.630 1100.540 ;
        RECT 667.530 1100.480 667.850 1100.540 ;
        RECT 664.310 1100.340 667.850 1100.480 ;
        RECT 664.310 1100.280 664.630 1100.340 ;
        RECT 667.530 1100.280 667.850 1100.340 ;
        RECT 664.310 1052.200 664.630 1052.260 ;
        RECT 667.530 1052.200 667.850 1052.260 ;
        RECT 664.310 1052.060 667.850 1052.200 ;
        RECT 664.310 1052.000 664.630 1052.060 ;
        RECT 667.530 1052.000 667.850 1052.060 ;
        RECT 664.310 907.360 664.630 907.420 ;
        RECT 666.610 907.360 666.930 907.420 ;
        RECT 664.310 907.220 666.930 907.360 ;
        RECT 664.310 907.160 664.630 907.220 ;
        RECT 666.610 907.160 666.930 907.220 ;
        RECT 664.770 834.600 665.090 834.660 ;
        RECT 666.610 834.600 666.930 834.660 ;
        RECT 664.770 834.460 666.930 834.600 ;
        RECT 664.770 834.400 665.090 834.460 ;
        RECT 666.610 834.400 666.930 834.460 ;
        RECT 664.310 821.000 664.630 821.060 ;
        RECT 664.770 821.000 665.090 821.060 ;
        RECT 664.310 820.860 665.090 821.000 ;
        RECT 664.310 820.800 664.630 820.860 ;
        RECT 664.770 820.800 665.090 820.860 ;
        RECT 663.390 814.200 663.710 814.260 ;
        RECT 664.310 814.200 664.630 814.260 ;
        RECT 663.390 814.060 664.630 814.200 ;
        RECT 663.390 814.000 663.710 814.060 ;
        RECT 664.310 814.000 664.630 814.060 ;
        RECT 663.390 766.260 663.710 766.320 ;
        RECT 664.310 766.260 664.630 766.320 ;
        RECT 663.390 766.120 664.630 766.260 ;
        RECT 663.390 766.060 663.710 766.120 ;
        RECT 664.310 766.060 664.630 766.120 ;
        RECT 664.310 738.520 664.630 738.780 ;
        RECT 664.400 738.100 664.540 738.520 ;
        RECT 664.310 737.840 664.630 738.100 ;
        RECT 663.850 628.220 664.170 628.280 ;
        RECT 664.310 628.220 664.630 628.280 ;
        RECT 663.850 628.080 664.630 628.220 ;
        RECT 663.850 628.020 664.170 628.080 ;
        RECT 664.310 628.020 664.630 628.080 ;
        RECT 663.850 595.240 664.170 595.300 ;
        RECT 670.750 595.240 671.070 595.300 ;
        RECT 663.850 595.100 671.070 595.240 ;
        RECT 663.850 595.040 664.170 595.100 ;
        RECT 670.750 595.040 671.070 595.100 ;
        RECT 665.690 234.500 666.010 234.560 ;
        RECT 666.610 234.500 666.930 234.560 ;
        RECT 665.690 234.360 666.930 234.500 ;
        RECT 665.690 234.300 666.010 234.360 ;
        RECT 666.610 234.300 666.930 234.360 ;
        RECT 665.690 186.560 666.010 186.620 ;
        RECT 667.530 186.560 667.850 186.620 ;
        RECT 665.690 186.420 667.850 186.560 ;
        RECT 665.690 186.360 666.010 186.420 ;
        RECT 667.530 186.360 667.850 186.420 ;
        RECT 666.610 145.080 666.930 145.140 ;
        RECT 667.530 145.080 667.850 145.140 ;
        RECT 666.610 144.940 667.850 145.080 ;
        RECT 666.610 144.880 666.930 144.940 ;
        RECT 667.530 144.880 667.850 144.940 ;
        RECT 665.690 137.940 666.010 138.000 ;
        RECT 666.610 137.940 666.930 138.000 ;
        RECT 665.690 137.800 666.930 137.940 ;
        RECT 665.690 137.740 666.010 137.800 ;
        RECT 666.610 137.740 666.930 137.800 ;
        RECT 665.690 90.000 666.010 90.060 ;
        RECT 666.610 90.000 666.930 90.060 ;
        RECT 665.690 89.860 666.930 90.000 ;
        RECT 665.690 89.800 666.010 89.860 ;
        RECT 666.610 89.800 666.930 89.860 ;
        RECT 665.690 48.520 666.010 48.580 ;
        RECT 666.610 48.520 666.930 48.580 ;
        RECT 665.690 48.380 666.930 48.520 ;
        RECT 665.690 48.320 666.010 48.380 ;
        RECT 666.610 48.320 666.930 48.380 ;
        RECT 531.830 43.080 532.150 43.140 ;
        RECT 665.690 43.080 666.010 43.140 ;
        RECT 531.830 42.940 666.010 43.080 ;
        RECT 531.830 42.880 532.150 42.940 ;
        RECT 665.690 42.880 666.010 42.940 ;
      LAYER via ;
        RECT 665.260 2039.360 665.520 2039.620 ;
        RECT 1903.120 2039.360 1903.380 2039.620 ;
        RECT 664.340 2021.680 664.600 2021.940 ;
        RECT 665.260 2021.680 665.520 2021.940 ;
        RECT 663.420 1993.800 663.680 1994.060 ;
        RECT 664.340 1993.800 664.600 1994.060 ;
        RECT 662.040 1973.060 662.300 1973.320 ;
        RECT 664.340 1973.060 664.600 1973.320 ;
        RECT 662.040 1897.240 662.300 1897.500 ;
        RECT 663.420 1897.240 663.680 1897.500 ;
        RECT 663.880 1780.280 664.140 1780.540 ;
        RECT 664.340 1780.280 664.600 1780.540 ;
        RECT 663.880 1752.740 664.140 1753.000 ;
        RECT 663.420 1752.400 663.680 1752.660 ;
        RECT 663.420 1541.260 663.680 1541.520 ;
        RECT 664.340 1541.260 664.600 1541.520 ;
        RECT 663.420 1480.400 663.680 1480.660 ;
        RECT 664.340 1480.400 664.600 1480.660 ;
        RECT 663.420 1444.700 663.680 1444.960 ;
        RECT 664.340 1444.700 664.600 1444.960 ;
        RECT 664.340 1390.300 664.600 1390.560 ;
        RECT 667.560 1390.300 667.820 1390.560 ;
        RECT 664.340 1342.020 664.600 1342.280 ;
        RECT 667.560 1342.020 667.820 1342.280 ;
        RECT 664.340 1293.740 664.600 1294.000 ;
        RECT 667.560 1293.740 667.820 1294.000 ;
        RECT 664.340 1245.460 664.600 1245.720 ;
        RECT 667.560 1245.460 667.820 1245.720 ;
        RECT 664.340 1197.180 664.600 1197.440 ;
        RECT 667.560 1197.180 667.820 1197.440 ;
        RECT 664.340 1148.560 664.600 1148.820 ;
        RECT 667.560 1148.560 667.820 1148.820 ;
        RECT 664.340 1100.280 664.600 1100.540 ;
        RECT 667.560 1100.280 667.820 1100.540 ;
        RECT 664.340 1052.000 664.600 1052.260 ;
        RECT 667.560 1052.000 667.820 1052.260 ;
        RECT 664.340 907.160 664.600 907.420 ;
        RECT 666.640 907.160 666.900 907.420 ;
        RECT 664.800 834.400 665.060 834.660 ;
        RECT 666.640 834.400 666.900 834.660 ;
        RECT 664.340 820.800 664.600 821.060 ;
        RECT 664.800 820.800 665.060 821.060 ;
        RECT 663.420 814.000 663.680 814.260 ;
        RECT 664.340 814.000 664.600 814.260 ;
        RECT 663.420 766.060 663.680 766.320 ;
        RECT 664.340 766.060 664.600 766.320 ;
        RECT 664.340 738.520 664.600 738.780 ;
        RECT 664.340 737.840 664.600 738.100 ;
        RECT 663.880 628.020 664.140 628.280 ;
        RECT 664.340 628.020 664.600 628.280 ;
        RECT 663.880 595.040 664.140 595.300 ;
        RECT 670.780 595.040 671.040 595.300 ;
        RECT 665.720 234.300 665.980 234.560 ;
        RECT 666.640 234.300 666.900 234.560 ;
        RECT 665.720 186.360 665.980 186.620 ;
        RECT 667.560 186.360 667.820 186.620 ;
        RECT 666.640 144.880 666.900 145.140 ;
        RECT 667.560 144.880 667.820 145.140 ;
        RECT 665.720 137.740 665.980 138.000 ;
        RECT 666.640 137.740 666.900 138.000 ;
        RECT 665.720 89.800 665.980 90.060 ;
        RECT 666.640 89.800 666.900 90.060 ;
        RECT 665.720 48.320 665.980 48.580 ;
        RECT 666.640 48.320 666.900 48.580 ;
        RECT 531.860 42.880 532.120 43.140 ;
        RECT 665.720 42.880 665.980 43.140 ;
      LAYER met2 ;
        RECT 1903.110 2877.235 1903.390 2877.605 ;
        RECT 1903.180 2039.650 1903.320 2877.235 ;
        RECT 665.260 2039.330 665.520 2039.650 ;
        RECT 1903.120 2039.330 1903.380 2039.650 ;
        RECT 665.320 2021.970 665.460 2039.330 ;
        RECT 664.340 2021.650 664.600 2021.970 ;
        RECT 665.260 2021.650 665.520 2021.970 ;
        RECT 664.400 1994.170 664.540 2021.650 ;
        RECT 663.480 1994.090 664.540 1994.170 ;
        RECT 663.420 1994.030 664.600 1994.090 ;
        RECT 663.420 1993.770 663.680 1994.030 ;
        RECT 664.340 1993.770 664.600 1994.030 ;
        RECT 663.480 1993.615 663.620 1993.770 ;
        RECT 664.400 1973.350 664.540 1993.770 ;
        RECT 662.040 1973.030 662.300 1973.350 ;
        RECT 664.340 1973.030 664.600 1973.350 ;
        RECT 662.100 1897.530 662.240 1973.030 ;
        RECT 662.040 1897.210 662.300 1897.530 ;
        RECT 663.420 1897.210 663.680 1897.530 ;
        RECT 663.480 1849.330 663.620 1897.210 ;
        RECT 663.480 1849.190 664.540 1849.330 ;
        RECT 664.400 1780.570 664.540 1849.190 ;
        RECT 663.880 1780.250 664.140 1780.570 ;
        RECT 664.340 1780.250 664.600 1780.570 ;
        RECT 351.070 1777.675 351.350 1778.045 ;
        RECT 351.140 1710.045 351.280 1777.675 ;
        RECT 663.940 1753.030 664.080 1780.250 ;
        RECT 663.880 1752.710 664.140 1753.030 ;
        RECT 663.420 1752.370 663.680 1752.690 ;
        RECT 663.480 1710.045 663.620 1752.370 ;
        RECT 351.070 1709.675 351.350 1710.045 ;
        RECT 663.410 1709.675 663.690 1710.045 ;
        RECT 663.480 1703.810 663.620 1709.675 ;
        RECT 663.480 1703.670 664.080 1703.810 ;
        RECT 663.940 1608.610 664.080 1703.670 ;
        RECT 663.480 1608.470 664.080 1608.610 ;
        RECT 663.480 1541.550 663.620 1608.470 ;
        RECT 663.420 1541.230 663.680 1541.550 ;
        RECT 664.340 1541.230 664.600 1541.550 ;
        RECT 664.400 1480.690 664.540 1541.230 ;
        RECT 663.420 1480.370 663.680 1480.690 ;
        RECT 664.340 1480.370 664.600 1480.690 ;
        RECT 663.480 1444.990 663.620 1480.370 ;
        RECT 663.420 1444.670 663.680 1444.990 ;
        RECT 664.340 1444.670 664.600 1444.990 ;
        RECT 664.400 1390.590 664.540 1444.670 ;
        RECT 664.340 1390.270 664.600 1390.590 ;
        RECT 667.560 1390.270 667.820 1390.590 ;
        RECT 667.620 1342.310 667.760 1390.270 ;
        RECT 664.340 1341.990 664.600 1342.310 ;
        RECT 667.560 1341.990 667.820 1342.310 ;
        RECT 664.400 1294.030 664.540 1341.990 ;
        RECT 664.340 1293.710 664.600 1294.030 ;
        RECT 667.560 1293.710 667.820 1294.030 ;
        RECT 667.620 1245.750 667.760 1293.710 ;
        RECT 664.340 1245.430 664.600 1245.750 ;
        RECT 667.560 1245.430 667.820 1245.750 ;
        RECT 664.400 1197.470 664.540 1245.430 ;
        RECT 664.340 1197.150 664.600 1197.470 ;
        RECT 667.560 1197.150 667.820 1197.470 ;
        RECT 667.620 1148.850 667.760 1197.150 ;
        RECT 664.340 1148.530 664.600 1148.850 ;
        RECT 667.560 1148.530 667.820 1148.850 ;
        RECT 664.400 1100.570 664.540 1148.530 ;
        RECT 664.340 1100.250 664.600 1100.570 ;
        RECT 667.560 1100.250 667.820 1100.570 ;
        RECT 667.620 1052.290 667.760 1100.250 ;
        RECT 664.340 1051.970 664.600 1052.290 ;
        RECT 667.560 1051.970 667.820 1052.290 ;
        RECT 664.400 980.405 664.540 1051.970 ;
        RECT 664.330 980.035 664.610 980.405 ;
        RECT 664.330 979.355 664.610 979.725 ;
        RECT 664.400 907.450 664.540 979.355 ;
        RECT 664.340 907.130 664.600 907.450 ;
        RECT 666.640 907.130 666.900 907.450 ;
        RECT 666.700 834.690 666.840 907.130 ;
        RECT 664.800 834.370 665.060 834.690 ;
        RECT 666.640 834.370 666.900 834.690 ;
        RECT 664.860 821.090 665.000 834.370 ;
        RECT 664.340 820.770 664.600 821.090 ;
        RECT 664.800 820.770 665.060 821.090 ;
        RECT 664.400 814.290 664.540 820.770 ;
        RECT 663.420 813.970 663.680 814.290 ;
        RECT 664.340 813.970 664.600 814.290 ;
        RECT 663.480 766.350 663.620 813.970 ;
        RECT 663.420 766.030 663.680 766.350 ;
        RECT 664.340 766.030 664.600 766.350 ;
        RECT 664.400 738.810 664.540 766.030 ;
        RECT 664.340 738.490 664.600 738.810 ;
        RECT 664.340 737.810 664.600 738.130 ;
        RECT 664.400 677.125 664.540 737.810 ;
        RECT 664.330 676.755 664.610 677.125 ;
        RECT 664.330 676.075 664.610 676.445 ;
        RECT 664.400 628.310 664.540 676.075 ;
        RECT 663.880 627.990 664.140 628.310 ;
        RECT 664.340 627.990 664.600 628.310 ;
        RECT 663.940 595.330 664.080 627.990 ;
        RECT 943.790 600.170 944.070 604.000 ;
        RECT 942.240 600.030 944.070 600.170 ;
        RECT 663.880 595.010 664.140 595.330 ;
        RECT 670.780 595.010 671.040 595.330 ;
        RECT 663.940 579.885 664.080 595.010 ;
        RECT 670.840 590.765 670.980 595.010 ;
        RECT 942.240 590.765 942.380 600.030 ;
        RECT 943.790 600.000 944.070 600.030 ;
        RECT 670.770 590.395 671.050 590.765 ;
        RECT 942.170 590.395 942.450 590.765 ;
        RECT 663.870 579.515 664.150 579.885 ;
        RECT 666.630 579.515 666.910 579.885 ;
        RECT 666.700 303.690 666.840 579.515 ;
        RECT 666.240 303.550 666.840 303.690 ;
        RECT 666.240 303.010 666.380 303.550 ;
        RECT 666.240 302.870 666.840 303.010 ;
        RECT 666.700 234.590 666.840 302.870 ;
        RECT 665.720 234.270 665.980 234.590 ;
        RECT 666.640 234.270 666.900 234.590 ;
        RECT 665.780 186.650 665.920 234.270 ;
        RECT 665.720 186.330 665.980 186.650 ;
        RECT 667.560 186.330 667.820 186.650 ;
        RECT 667.620 145.170 667.760 186.330 ;
        RECT 666.640 144.850 666.900 145.170 ;
        RECT 667.560 144.850 667.820 145.170 ;
        RECT 666.700 138.030 666.840 144.850 ;
        RECT 665.720 137.710 665.980 138.030 ;
        RECT 666.640 137.710 666.900 138.030 ;
        RECT 665.780 90.090 665.920 137.710 ;
        RECT 665.720 89.770 665.980 90.090 ;
        RECT 666.640 89.770 666.900 90.090 ;
        RECT 666.700 48.610 666.840 89.770 ;
        RECT 665.720 48.290 665.980 48.610 ;
        RECT 666.640 48.290 666.900 48.610 ;
        RECT 665.780 43.170 665.920 48.290 ;
        RECT 531.860 42.850 532.120 43.170 ;
        RECT 665.720 42.850 665.980 43.170 ;
        RECT 531.920 2.400 532.060 42.850 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 1903.110 2877.280 1903.390 2877.560 ;
        RECT 351.070 1777.720 351.350 1778.000 ;
        RECT 351.070 1709.720 351.350 1710.000 ;
        RECT 663.410 1709.720 663.690 1710.000 ;
        RECT 664.330 980.080 664.610 980.360 ;
        RECT 664.330 979.400 664.610 979.680 ;
        RECT 664.330 676.800 664.610 677.080 ;
        RECT 664.330 676.120 664.610 676.400 ;
        RECT 670.770 590.440 671.050 590.720 ;
        RECT 942.170 590.440 942.450 590.720 ;
        RECT 663.870 579.560 664.150 579.840 ;
        RECT 666.630 579.560 666.910 579.840 ;
      LAYER met3 ;
        RECT 1885.335 2879.800 1889.335 2880.080 ;
        RECT 1885.335 2879.480 1889.370 2879.800 ;
        RECT 1889.070 2877.570 1889.370 2879.480 ;
        RECT 1903.085 2877.570 1903.415 2877.585 ;
        RECT 1889.070 2877.270 1903.415 2877.570 ;
        RECT 1903.085 2877.255 1903.415 2877.270 ;
        RECT 351.045 1778.010 351.375 1778.025 ;
        RECT 360.000 1778.010 364.000 1778.160 ;
        RECT 351.045 1777.710 364.000 1778.010 ;
        RECT 351.045 1777.695 351.375 1777.710 ;
        RECT 360.000 1777.560 364.000 1777.710 ;
        RECT 351.045 1710.010 351.375 1710.025 ;
        RECT 663.385 1710.010 663.715 1710.025 ;
        RECT 351.045 1709.710 663.715 1710.010 ;
        RECT 351.045 1709.695 351.375 1709.710 ;
        RECT 663.385 1709.695 663.715 1709.710 ;
        RECT 663.590 980.370 663.970 980.380 ;
        RECT 664.305 980.370 664.635 980.385 ;
        RECT 663.590 980.070 664.635 980.370 ;
        RECT 663.590 980.060 663.970 980.070 ;
        RECT 664.305 980.055 664.635 980.070 ;
        RECT 663.590 979.690 663.970 979.700 ;
        RECT 664.305 979.690 664.635 979.705 ;
        RECT 663.590 979.390 664.635 979.690 ;
        RECT 663.590 979.380 663.970 979.390 ;
        RECT 664.305 979.375 664.635 979.390 ;
        RECT 664.305 677.090 664.635 677.105 ;
        RECT 664.305 676.775 664.850 677.090 ;
        RECT 664.550 676.425 664.850 676.775 ;
        RECT 664.305 676.110 664.850 676.425 ;
        RECT 664.305 676.095 664.635 676.110 ;
        RECT 670.745 590.730 671.075 590.745 ;
        RECT 942.145 590.730 942.475 590.745 ;
        RECT 670.745 590.430 942.475 590.730 ;
        RECT 670.745 590.415 671.075 590.430 ;
        RECT 942.145 590.415 942.475 590.430 ;
        RECT 663.845 579.850 664.175 579.865 ;
        RECT 666.605 579.850 666.935 579.865 ;
        RECT 663.845 579.550 666.935 579.850 ;
        RECT 663.845 579.535 664.175 579.550 ;
        RECT 666.605 579.535 666.935 579.550 ;
      LAYER via3 ;
        RECT 663.620 980.060 663.940 980.380 ;
        RECT 663.620 979.380 663.940 979.700 ;
      LAYER met4 ;
        RECT 663.615 980.055 663.945 980.385 ;
        RECT 663.630 979.705 663.930 980.055 ;
        RECT 663.615 979.375 663.945 979.705 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 589.790 1687.660 590.110 1687.720 ;
        RECT 620.610 1687.660 620.930 1687.720 ;
        RECT 1486.790 1687.660 1487.110 1687.720 ;
        RECT 589.790 1687.520 1487.110 1687.660 ;
        RECT 589.790 1687.460 590.110 1687.520 ;
        RECT 620.610 1687.460 620.930 1687.520 ;
        RECT 1486.790 1687.460 1487.110 1687.520 ;
        RECT 620.610 592.180 620.930 592.240 ;
        RECT 952.270 592.180 952.590 592.240 ;
        RECT 620.610 592.040 952.590 592.180 ;
        RECT 620.610 591.980 620.930 592.040 ;
        RECT 952.270 591.980 952.590 592.040 ;
        RECT 617.390 587.420 617.710 587.480 ;
        RECT 620.610 587.420 620.930 587.480 ;
        RECT 617.390 587.280 620.930 587.420 ;
        RECT 617.390 587.220 617.710 587.280 ;
        RECT 620.610 587.220 620.930 587.280 ;
        RECT 617.390 21.120 617.710 21.380 ;
        RECT 549.770 20.980 550.090 21.040 ;
        RECT 617.480 20.980 617.620 21.120 ;
        RECT 549.770 20.840 617.620 20.980 ;
        RECT 549.770 20.780 550.090 20.840 ;
      LAYER via ;
        RECT 589.820 1687.460 590.080 1687.720 ;
        RECT 620.640 1687.460 620.900 1687.720 ;
        RECT 1486.820 1687.460 1487.080 1687.720 ;
        RECT 620.640 591.980 620.900 592.240 ;
        RECT 952.300 591.980 952.560 592.240 ;
        RECT 617.420 587.220 617.680 587.480 ;
        RECT 620.640 587.220 620.900 587.480 ;
        RECT 617.420 21.120 617.680 21.380 ;
        RECT 549.800 20.780 550.060 21.040 ;
      LAYER met2 ;
        RECT 1486.810 2705.195 1487.090 2705.565 ;
        RECT 588.250 1700.410 588.530 1704.000 ;
        RECT 588.250 1700.270 590.020 1700.410 ;
        RECT 588.250 1700.000 588.530 1700.270 ;
        RECT 589.880 1687.750 590.020 1700.270 ;
        RECT 1486.880 1687.750 1487.020 2705.195 ;
        RECT 589.820 1687.430 590.080 1687.750 ;
        RECT 620.640 1687.430 620.900 1687.750 ;
        RECT 1486.820 1687.430 1487.080 1687.750 ;
        RECT 620.700 592.270 620.840 1687.430 ;
        RECT 952.990 600.170 953.270 604.000 ;
        RECT 952.360 600.030 953.270 600.170 ;
        RECT 952.360 592.270 952.500 600.030 ;
        RECT 952.990 600.000 953.270 600.030 ;
        RECT 620.640 591.950 620.900 592.270 ;
        RECT 952.300 591.950 952.560 592.270 ;
        RECT 620.700 587.510 620.840 591.950 ;
        RECT 617.420 587.190 617.680 587.510 ;
        RECT 620.640 587.190 620.900 587.510 ;
        RECT 617.480 21.410 617.620 587.190 ;
        RECT 617.420 21.090 617.680 21.410 ;
        RECT 549.800 20.750 550.060 21.070 ;
        RECT 549.860 2.400 550.000 20.750 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 1486.810 2705.240 1487.090 2705.520 ;
      LAYER met3 ;
        RECT 1500.000 2708.440 1504.000 2708.720 ;
        RECT 1499.910 2708.120 1504.000 2708.440 ;
        RECT 1486.785 2705.530 1487.115 2705.545 ;
        RECT 1499.910 2705.530 1500.210 2708.120 ;
        RECT 1486.785 2705.230 1500.210 2705.530 ;
        RECT 1486.785 2705.215 1487.115 2705.230 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 962.390 2532.560 962.710 2532.620 ;
        RECT 1483.570 2532.560 1483.890 2532.620 ;
        RECT 962.390 2532.420 1483.890 2532.560 ;
        RECT 962.390 2532.360 962.710 2532.420 ;
        RECT 1483.570 2532.360 1483.890 2532.420 ;
        RECT 644.990 1714.520 645.310 1714.580 ;
        RECT 653.270 1714.520 653.590 1714.580 ;
        RECT 962.390 1714.520 962.710 1714.580 ;
        RECT 644.990 1714.380 962.710 1714.520 ;
        RECT 644.990 1714.320 645.310 1714.380 ;
        RECT 653.270 1714.320 653.590 1714.380 ;
        RECT 962.390 1714.320 962.710 1714.380 ;
        RECT 653.270 677.860 653.590 677.920 ;
        RECT 661.550 677.860 661.870 677.920 ;
        RECT 653.270 677.720 661.870 677.860 ;
        RECT 653.270 677.660 653.590 677.720 ;
        RECT 661.550 677.660 661.870 677.720 ;
        RECT 661.550 662.220 661.870 662.280 ;
        RECT 665.690 662.220 666.010 662.280 ;
        RECT 661.550 662.080 666.010 662.220 ;
        RECT 661.550 662.020 661.870 662.080 ;
        RECT 665.690 662.020 666.010 662.080 ;
        RECT 665.690 601.700 666.010 601.760 ;
        RECT 675.810 601.700 676.130 601.760 ;
        RECT 665.690 601.560 676.130 601.700 ;
        RECT 665.690 601.500 666.010 601.560 ;
        RECT 675.810 601.500 676.130 601.560 ;
        RECT 675.810 596.940 676.130 597.000 ;
        RECT 960.090 596.940 960.410 597.000 ;
        RECT 675.810 596.800 960.410 596.940 ;
        RECT 675.810 596.740 676.130 596.800 ;
        RECT 960.090 596.740 960.410 596.800 ;
        RECT 960.090 531.460 960.410 531.720 ;
        RECT 960.180 530.980 960.320 531.460 ;
        RECT 961.010 530.980 961.330 531.040 ;
        RECT 960.180 530.840 961.330 530.980 ;
        RECT 961.010 530.780 961.330 530.840 ;
        RECT 961.010 517.380 961.330 517.440 ;
        RECT 961.930 517.380 962.250 517.440 ;
        RECT 961.010 517.240 962.250 517.380 ;
        RECT 961.010 517.180 961.330 517.240 ;
        RECT 961.930 517.180 962.250 517.240 ;
        RECT 961.930 435.240 962.250 435.500 ;
        RECT 962.020 434.820 962.160 435.240 ;
        RECT 961.930 434.560 962.250 434.820 ;
        RECT 960.090 420.820 960.410 420.880 ;
        RECT 961.930 420.820 962.250 420.880 ;
        RECT 960.090 420.680 962.250 420.820 ;
        RECT 960.090 420.620 960.410 420.680 ;
        RECT 961.930 420.620 962.250 420.680 ;
        RECT 960.090 372.880 960.410 372.940 ;
        RECT 961.010 372.880 961.330 372.940 ;
        RECT 960.090 372.740 961.330 372.880 ;
        RECT 960.090 372.680 960.410 372.740 ;
        RECT 961.010 372.680 961.330 372.740 ;
        RECT 961.010 352.480 961.330 352.540 ;
        RECT 960.640 352.340 961.330 352.480 ;
        RECT 960.640 351.860 960.780 352.340 ;
        RECT 961.010 352.280 961.330 352.340 ;
        RECT 960.550 351.600 960.870 351.860 ;
        RECT 960.550 304.000 960.870 304.260 ;
        RECT 960.640 303.580 960.780 304.000 ;
        RECT 960.550 303.320 960.870 303.580 ;
        RECT 960.550 282.780 960.870 282.840 ;
        RECT 961.470 282.780 961.790 282.840 ;
        RECT 960.550 282.640 961.790 282.780 ;
        RECT 960.550 282.580 960.870 282.640 ;
        RECT 961.470 282.580 961.790 282.640 ;
        RECT 961.010 275.980 961.330 276.040 ;
        RECT 961.470 275.980 961.790 276.040 ;
        RECT 961.010 275.840 961.790 275.980 ;
        RECT 961.010 275.780 961.330 275.840 ;
        RECT 961.470 275.780 961.790 275.840 ;
        RECT 960.550 227.700 960.870 227.760 ;
        RECT 961.010 227.700 961.330 227.760 ;
        RECT 960.550 227.560 961.330 227.700 ;
        RECT 960.550 227.500 960.870 227.560 ;
        RECT 961.010 227.500 961.330 227.560 ;
        RECT 960.090 172.620 960.410 172.680 ;
        RECT 961.010 172.620 961.330 172.680 ;
        RECT 960.090 172.480 961.330 172.620 ;
        RECT 960.090 172.420 960.410 172.480 ;
        RECT 961.010 172.420 961.330 172.480 ;
        RECT 961.010 158.820 961.330 159.080 ;
        RECT 960.550 158.680 960.870 158.740 ;
        RECT 961.100 158.680 961.240 158.820 ;
        RECT 960.550 158.540 961.240 158.680 ;
        RECT 960.550 158.480 960.870 158.540 ;
        RECT 960.090 131.820 960.410 131.880 ;
        RECT 960.550 131.820 960.870 131.880 ;
        RECT 960.090 131.680 960.870 131.820 ;
        RECT 960.090 131.620 960.410 131.680 ;
        RECT 960.550 131.620 960.870 131.680 ;
        RECT 960.090 131.140 960.410 131.200 ;
        RECT 961.930 131.140 962.250 131.200 ;
        RECT 960.090 131.000 962.250 131.140 ;
        RECT 960.090 130.940 960.410 131.000 ;
        RECT 961.930 130.940 962.250 131.000 ;
        RECT 961.010 83.200 961.330 83.260 ;
        RECT 961.930 83.200 962.250 83.260 ;
        RECT 961.010 83.060 962.250 83.200 ;
        RECT 961.010 83.000 961.330 83.060 ;
        RECT 961.930 83.000 962.250 83.060 ;
        RECT 567.710 29.140 568.030 29.200 ;
        RECT 961.010 29.140 961.330 29.200 ;
        RECT 567.710 29.000 961.330 29.140 ;
        RECT 567.710 28.940 568.030 29.000 ;
        RECT 961.010 28.940 961.330 29.000 ;
      LAYER via ;
        RECT 962.420 2532.360 962.680 2532.620 ;
        RECT 1483.600 2532.360 1483.860 2532.620 ;
        RECT 645.020 1714.320 645.280 1714.580 ;
        RECT 653.300 1714.320 653.560 1714.580 ;
        RECT 962.420 1714.320 962.680 1714.580 ;
        RECT 653.300 677.660 653.560 677.920 ;
        RECT 661.580 677.660 661.840 677.920 ;
        RECT 661.580 662.020 661.840 662.280 ;
        RECT 665.720 662.020 665.980 662.280 ;
        RECT 665.720 601.500 665.980 601.760 ;
        RECT 675.840 601.500 676.100 601.760 ;
        RECT 675.840 596.740 676.100 597.000 ;
        RECT 960.120 596.740 960.380 597.000 ;
        RECT 960.120 531.460 960.380 531.720 ;
        RECT 961.040 530.780 961.300 531.040 ;
        RECT 961.040 517.180 961.300 517.440 ;
        RECT 961.960 517.180 962.220 517.440 ;
        RECT 961.960 435.240 962.220 435.500 ;
        RECT 961.960 434.560 962.220 434.820 ;
        RECT 960.120 420.620 960.380 420.880 ;
        RECT 961.960 420.620 962.220 420.880 ;
        RECT 960.120 372.680 960.380 372.940 ;
        RECT 961.040 372.680 961.300 372.940 ;
        RECT 961.040 352.280 961.300 352.540 ;
        RECT 960.580 351.600 960.840 351.860 ;
        RECT 960.580 304.000 960.840 304.260 ;
        RECT 960.580 303.320 960.840 303.580 ;
        RECT 960.580 282.580 960.840 282.840 ;
        RECT 961.500 282.580 961.760 282.840 ;
        RECT 961.040 275.780 961.300 276.040 ;
        RECT 961.500 275.780 961.760 276.040 ;
        RECT 960.580 227.500 960.840 227.760 ;
        RECT 961.040 227.500 961.300 227.760 ;
        RECT 960.120 172.420 960.380 172.680 ;
        RECT 961.040 172.420 961.300 172.680 ;
        RECT 961.040 158.820 961.300 159.080 ;
        RECT 960.580 158.480 960.840 158.740 ;
        RECT 960.120 131.620 960.380 131.880 ;
        RECT 960.580 131.620 960.840 131.880 ;
        RECT 960.120 130.940 960.380 131.200 ;
        RECT 961.960 130.940 962.220 131.200 ;
        RECT 961.040 83.000 961.300 83.260 ;
        RECT 961.960 83.000 962.220 83.260 ;
        RECT 567.740 28.940 568.000 29.200 ;
        RECT 961.040 28.940 961.300 29.200 ;
      LAYER met2 ;
        RECT 1483.590 2533.155 1483.870 2533.525 ;
        RECT 1483.660 2532.650 1483.800 2533.155 ;
        RECT 962.420 2532.330 962.680 2532.650 ;
        RECT 1483.600 2532.330 1483.860 2532.650 ;
        RECT 645.010 1717.835 645.290 1718.205 ;
        RECT 645.080 1714.610 645.220 1717.835 ;
        RECT 962.480 1714.610 962.620 2532.330 ;
        RECT 645.020 1714.290 645.280 1714.610 ;
        RECT 653.300 1714.290 653.560 1714.610 ;
        RECT 962.420 1714.290 962.680 1714.610 ;
        RECT 653.360 677.950 653.500 1714.290 ;
        RECT 653.300 677.630 653.560 677.950 ;
        RECT 661.580 677.630 661.840 677.950 ;
        RECT 661.640 662.310 661.780 677.630 ;
        RECT 661.580 661.990 661.840 662.310 ;
        RECT 665.720 661.990 665.980 662.310 ;
        RECT 665.780 601.790 665.920 661.990 ;
        RECT 665.720 601.470 665.980 601.790 ;
        RECT 675.840 601.470 676.100 601.790 ;
        RECT 962.190 601.530 962.470 604.000 ;
        RECT 675.900 597.030 676.040 601.470 ;
        RECT 960.180 601.390 962.470 601.530 ;
        RECT 960.180 597.030 960.320 601.390 ;
        RECT 962.190 600.000 962.470 601.390 ;
        RECT 675.840 596.710 676.100 597.030 ;
        RECT 960.120 596.710 960.380 597.030 ;
        RECT 960.180 531.750 960.320 596.710 ;
        RECT 960.120 531.430 960.380 531.750 ;
        RECT 961.040 530.750 961.300 531.070 ;
        RECT 961.100 517.470 961.240 530.750 ;
        RECT 961.040 517.150 961.300 517.470 ;
        RECT 961.960 517.150 962.220 517.470 ;
        RECT 962.020 435.530 962.160 517.150 ;
        RECT 961.960 435.210 962.220 435.530 ;
        RECT 961.960 434.530 962.220 434.850 ;
        RECT 962.020 420.910 962.160 434.530 ;
        RECT 960.120 420.590 960.380 420.910 ;
        RECT 961.960 420.590 962.220 420.910 ;
        RECT 960.180 372.970 960.320 420.590 ;
        RECT 960.120 372.650 960.380 372.970 ;
        RECT 961.040 372.650 961.300 372.970 ;
        RECT 961.100 352.570 961.240 372.650 ;
        RECT 961.040 352.250 961.300 352.570 ;
        RECT 960.580 351.570 960.840 351.890 ;
        RECT 960.640 304.290 960.780 351.570 ;
        RECT 960.580 303.970 960.840 304.290 ;
        RECT 960.580 303.290 960.840 303.610 ;
        RECT 960.640 282.870 960.780 303.290 ;
        RECT 960.580 282.550 960.840 282.870 ;
        RECT 961.500 282.550 961.760 282.870 ;
        RECT 961.560 276.070 961.700 282.550 ;
        RECT 961.040 275.750 961.300 276.070 ;
        RECT 961.500 275.750 961.760 276.070 ;
        RECT 961.100 228.210 961.240 275.750 ;
        RECT 960.640 228.070 961.240 228.210 ;
        RECT 960.640 227.790 960.780 228.070 ;
        RECT 960.580 227.470 960.840 227.790 ;
        RECT 961.040 227.470 961.300 227.790 ;
        RECT 961.100 220.845 961.240 227.470 ;
        RECT 960.110 220.475 960.390 220.845 ;
        RECT 961.030 220.475 961.310 220.845 ;
        RECT 960.180 172.710 960.320 220.475 ;
        RECT 960.120 172.390 960.380 172.710 ;
        RECT 961.040 172.390 961.300 172.710 ;
        RECT 961.100 159.110 961.240 172.390 ;
        RECT 961.040 158.790 961.300 159.110 ;
        RECT 960.580 158.450 960.840 158.770 ;
        RECT 960.640 131.910 960.780 158.450 ;
        RECT 960.120 131.590 960.380 131.910 ;
        RECT 960.580 131.590 960.840 131.910 ;
        RECT 960.180 131.230 960.320 131.590 ;
        RECT 960.120 130.910 960.380 131.230 ;
        RECT 961.960 130.910 962.220 131.230 ;
        RECT 962.020 83.290 962.160 130.910 ;
        RECT 961.040 82.970 961.300 83.290 ;
        RECT 961.960 82.970 962.220 83.290 ;
        RECT 961.100 29.230 961.240 82.970 ;
        RECT 567.740 28.910 568.000 29.230 ;
        RECT 961.040 28.910 961.300 29.230 ;
        RECT 567.800 2.400 567.940 28.910 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1483.590 2533.200 1483.870 2533.480 ;
        RECT 645.010 1717.880 645.290 1718.160 ;
        RECT 960.110 220.520 960.390 220.800 ;
        RECT 961.030 220.520 961.310 220.800 ;
      LAYER met3 ;
        RECT 1500.000 2535.720 1504.000 2536.000 ;
        RECT 1499.910 2535.400 1504.000 2535.720 ;
        RECT 1483.565 2533.490 1483.895 2533.505 ;
        RECT 1499.910 2533.490 1500.210 2535.400 ;
        RECT 1483.565 2533.190 1500.210 2533.490 ;
        RECT 1483.565 2533.175 1483.895 2533.190 ;
        RECT 627.030 1718.170 631.030 1718.320 ;
        RECT 644.985 1718.170 645.315 1718.185 ;
        RECT 627.030 1717.870 645.315 1718.170 ;
        RECT 627.030 1717.720 631.030 1717.870 ;
        RECT 644.985 1717.855 645.315 1717.870 ;
        RECT 960.085 220.810 960.415 220.825 ;
        RECT 961.005 220.810 961.335 220.825 ;
        RECT 960.085 220.510 961.335 220.810 ;
        RECT 960.085 220.495 960.415 220.510 ;
        RECT 961.005 220.495 961.335 220.510 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 438.910 1686.980 439.230 1687.040 ;
        RECT 641.310 1686.980 641.630 1687.040 ;
        RECT 1902.630 1686.980 1902.950 1687.040 ;
        RECT 438.910 1686.840 1902.950 1686.980 ;
        RECT 438.910 1686.780 439.230 1686.840 ;
        RECT 641.310 1686.780 641.630 1686.840 ;
        RECT 1902.630 1686.780 1902.950 1686.840 ;
        RECT 593.560 36.480 618.540 36.620 ;
        RECT 585.650 36.280 585.970 36.340 ;
        RECT 593.560 36.280 593.700 36.480 ;
        RECT 585.650 36.140 593.700 36.280 ;
        RECT 618.400 36.280 618.540 36.480 ;
        RECT 638.090 36.280 638.410 36.340 ;
        RECT 618.400 36.140 638.410 36.280 ;
        RECT 585.650 36.080 585.970 36.140 ;
        RECT 638.090 36.080 638.410 36.140 ;
      LAYER via ;
        RECT 438.940 1686.780 439.200 1687.040 ;
        RECT 641.340 1686.780 641.600 1687.040 ;
        RECT 1902.660 1686.780 1902.920 1687.040 ;
        RECT 585.680 36.080 585.940 36.340 ;
        RECT 638.120 36.080 638.380 36.340 ;
      LAYER met2 ;
        RECT 1902.650 2643.315 1902.930 2643.685 ;
        RECT 437.370 1700.410 437.650 1704.000 ;
        RECT 437.370 1700.270 439.140 1700.410 ;
        RECT 437.370 1700.000 437.650 1700.270 ;
        RECT 439.000 1687.070 439.140 1700.270 ;
        RECT 1902.720 1687.070 1902.860 2643.315 ;
        RECT 438.940 1686.750 439.200 1687.070 ;
        RECT 641.340 1686.750 641.600 1687.070 ;
        RECT 1902.660 1686.750 1902.920 1687.070 ;
        RECT 641.400 591.445 641.540 1686.750 ;
        RECT 971.390 600.170 971.670 604.000 ;
        RECT 969.840 600.030 971.670 600.170 ;
        RECT 969.840 591.445 969.980 600.030 ;
        RECT 971.390 600.000 971.670 600.030 ;
        RECT 641.330 591.075 641.610 591.445 ;
        RECT 969.770 591.075 970.050 591.445 ;
        RECT 641.400 586.685 641.540 591.075 ;
        RECT 638.110 586.315 638.390 586.685 ;
        RECT 641.330 586.315 641.610 586.685 ;
        RECT 638.180 36.370 638.320 586.315 ;
        RECT 585.680 36.050 585.940 36.370 ;
        RECT 638.120 36.050 638.380 36.370 ;
        RECT 585.740 2.400 585.880 36.050 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 1902.650 2643.360 1902.930 2643.640 ;
        RECT 641.330 591.120 641.610 591.400 ;
        RECT 969.770 591.120 970.050 591.400 ;
        RECT 638.110 586.360 638.390 586.640 ;
        RECT 641.330 586.360 641.610 586.640 ;
      LAYER met3 ;
        RECT 1885.335 2644.520 1889.335 2644.800 ;
        RECT 1885.335 2644.200 1889.370 2644.520 ;
        RECT 1889.070 2643.650 1889.370 2644.200 ;
        RECT 1902.625 2643.650 1902.955 2643.665 ;
        RECT 1889.070 2643.350 1902.955 2643.650 ;
        RECT 1902.625 2643.335 1902.955 2643.350 ;
        RECT 641.305 591.410 641.635 591.425 ;
        RECT 969.745 591.410 970.075 591.425 ;
        RECT 641.305 591.110 970.075 591.410 ;
        RECT 641.305 591.095 641.635 591.110 ;
        RECT 969.745 591.095 970.075 591.110 ;
        RECT 638.085 586.650 638.415 586.665 ;
        RECT 641.305 586.650 641.635 586.665 ;
        RECT 638.085 586.350 641.635 586.650 ;
        RECT 638.085 586.335 638.415 586.350 ;
        RECT 641.305 586.335 641.635 586.350 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1479.890 2663.800 1480.210 2663.860 ;
        RECT 1487.250 2663.800 1487.570 2663.860 ;
        RECT 1479.890 2663.660 1487.570 2663.800 ;
        RECT 1479.890 2663.600 1480.210 2663.660 ;
        RECT 1487.250 2663.600 1487.570 2663.660 ;
        RECT 1476.670 2608.040 1476.990 2608.100 ;
        RECT 1479.890 2608.040 1480.210 2608.100 ;
        RECT 1476.670 2607.900 1480.210 2608.040 ;
        RECT 1476.670 2607.840 1476.990 2607.900 ;
        RECT 1479.890 2607.840 1480.210 2607.900 ;
        RECT 426.490 2606.340 426.810 2606.400 ;
        RECT 1476.670 2606.340 1476.990 2606.400 ;
        RECT 426.490 2606.200 1476.990 2606.340 ;
        RECT 426.490 2606.140 426.810 2606.200 ;
        RECT 1476.670 2606.140 1476.990 2606.200 ;
        RECT 1014.460 2034.660 1062.440 2034.800 ;
        RECT 988.610 2032.760 988.930 2032.820 ;
        RECT 1014.460 2032.760 1014.600 2034.660 ;
        RECT 1062.300 2033.100 1062.440 2034.660 ;
        RECT 1330.390 2033.780 1330.710 2033.840 ;
        RECT 1172.700 2033.640 1222.520 2033.780 ;
        RECT 1172.700 2033.440 1172.840 2033.640 ;
        RECT 1111.060 2033.300 1124.540 2033.440 ;
        RECT 1062.300 2032.960 1076.240 2033.100 ;
        RECT 988.610 2032.620 1014.600 2032.760 ;
        RECT 1076.100 2032.760 1076.240 2032.960 ;
        RECT 1111.060 2032.760 1111.200 2033.300 ;
        RECT 1076.100 2032.620 1111.200 2032.760 ;
        RECT 1124.400 2032.760 1124.540 2033.300 ;
        RECT 1158.900 2033.300 1172.840 2033.440 ;
        RECT 1222.380 2033.440 1222.520 2033.640 ;
        RECT 1269.300 2033.640 1330.710 2033.780 ;
        RECT 1269.300 2033.440 1269.440 2033.640 ;
        RECT 1330.390 2033.580 1330.710 2033.640 ;
        RECT 1222.380 2033.300 1269.440 2033.440 ;
        RECT 1158.900 2032.760 1159.040 2033.300 ;
        RECT 1330.390 2033.100 1330.710 2033.160 ;
        RECT 1366.270 2033.100 1366.590 2033.160 ;
        RECT 1330.390 2032.960 1366.590 2033.100 ;
        RECT 1330.390 2032.900 1330.710 2032.960 ;
        RECT 1366.270 2032.900 1366.590 2032.960 ;
        RECT 1366.730 2033.100 1367.050 2033.160 ;
        RECT 1366.730 2032.960 1400.540 2033.100 ;
        RECT 1366.730 2032.900 1367.050 2032.960 ;
        RECT 1124.400 2032.620 1159.040 2032.760 ;
        RECT 1400.400 2032.760 1400.540 2032.960 ;
        RECT 1400.400 2032.620 1414.340 2032.760 ;
        RECT 988.610 2032.560 988.930 2032.620 ;
        RECT 1414.200 2032.080 1414.340 2032.620 ;
        RECT 1449.070 2032.080 1449.390 2032.140 ;
        RECT 1414.200 2031.940 1449.390 2032.080 ;
        RECT 1449.070 2031.880 1449.390 2031.940 ;
        RECT 1476.670 2030.040 1476.990 2030.100 ;
        RECT 1479.890 2030.040 1480.210 2030.100 ;
        RECT 1476.670 2029.900 1480.210 2030.040 ;
        RECT 1476.670 2029.840 1476.990 2029.900 ;
        RECT 1479.890 2029.840 1480.210 2029.900 ;
        RECT 1479.890 1928.720 1480.210 1928.780 ;
        RECT 1941.270 1928.720 1941.590 1928.780 ;
        RECT 1479.890 1928.580 1941.590 1928.720 ;
        RECT 1479.890 1928.520 1480.210 1928.580 ;
        RECT 1941.270 1928.520 1941.590 1928.580 ;
        RECT 646.830 1828.420 647.150 1828.480 ;
        RECT 988.610 1828.420 988.930 1828.480 ;
        RECT 646.830 1828.280 988.930 1828.420 ;
        RECT 646.830 1828.220 647.150 1828.280 ;
        RECT 988.610 1828.220 988.930 1828.280 ;
        RECT 646.830 588.440 647.150 588.500 ;
        RECT 676.270 588.440 676.590 588.500 ;
        RECT 646.830 588.300 676.590 588.440 ;
        RECT 646.830 588.240 647.150 588.300 ;
        RECT 676.270 588.240 676.590 588.300 ;
        RECT 683.170 587.760 683.490 587.820 ;
        RECT 714.910 587.760 715.230 587.820 ;
        RECT 683.170 587.620 715.230 587.760 ;
        RECT 683.170 587.560 683.490 587.620 ;
        RECT 714.910 587.560 715.230 587.620 ;
        RECT 676.270 586.400 676.590 586.460 ;
        RECT 683.170 586.400 683.490 586.460 ;
        RECT 676.270 586.260 683.490 586.400 ;
        RECT 676.270 586.200 676.590 586.260 ;
        RECT 676.820 585.380 676.960 586.260 ;
        RECT 683.170 586.200 683.490 586.260 ;
        RECT 677.190 585.380 677.510 585.440 ;
        RECT 676.820 585.240 677.510 585.380 ;
        RECT 677.190 585.180 677.510 585.240 ;
        RECT 91.610 45.800 91.930 45.860 ;
        RECT 677.190 45.800 677.510 45.860 ;
        RECT 91.610 45.660 677.510 45.800 ;
        RECT 91.610 45.600 91.930 45.660 ;
        RECT 677.190 45.600 677.510 45.660 ;
      LAYER via ;
        RECT 1479.920 2663.600 1480.180 2663.860 ;
        RECT 1487.280 2663.600 1487.540 2663.860 ;
        RECT 1476.700 2607.840 1476.960 2608.100 ;
        RECT 1479.920 2607.840 1480.180 2608.100 ;
        RECT 426.520 2606.140 426.780 2606.400 ;
        RECT 1476.700 2606.140 1476.960 2606.400 ;
        RECT 988.640 2032.560 988.900 2032.820 ;
        RECT 1330.420 2033.580 1330.680 2033.840 ;
        RECT 1330.420 2032.900 1330.680 2033.160 ;
        RECT 1366.300 2032.900 1366.560 2033.160 ;
        RECT 1366.760 2032.900 1367.020 2033.160 ;
        RECT 1449.100 2031.880 1449.360 2032.140 ;
        RECT 1476.700 2029.840 1476.960 2030.100 ;
        RECT 1479.920 2029.840 1480.180 2030.100 ;
        RECT 1479.920 1928.520 1480.180 1928.780 ;
        RECT 1941.300 1928.520 1941.560 1928.780 ;
        RECT 646.860 1828.220 647.120 1828.480 ;
        RECT 988.640 1828.220 988.900 1828.480 ;
        RECT 646.860 588.240 647.120 588.500 ;
        RECT 676.300 588.240 676.560 588.500 ;
        RECT 683.200 587.560 683.460 587.820 ;
        RECT 714.940 587.560 715.200 587.820 ;
        RECT 676.300 586.200 676.560 586.460 ;
        RECT 683.200 586.200 683.460 586.460 ;
        RECT 677.220 585.180 677.480 585.440 ;
        RECT 91.640 45.600 91.900 45.860 ;
        RECT 677.220 45.600 677.480 45.860 ;
      LAYER met2 ;
        RECT 1487.270 2864.315 1487.550 2864.685 ;
        RECT 426.510 2665.075 426.790 2665.445 ;
        RECT 426.580 2606.430 426.720 2665.075 ;
        RECT 1487.340 2663.890 1487.480 2864.315 ;
        RECT 1479.920 2663.570 1480.180 2663.890 ;
        RECT 1487.280 2663.570 1487.540 2663.890 ;
        RECT 1479.980 2608.130 1480.120 2663.570 ;
        RECT 1476.700 2607.810 1476.960 2608.130 ;
        RECT 1479.920 2607.810 1480.180 2608.130 ;
        RECT 1476.760 2606.430 1476.900 2607.810 ;
        RECT 426.520 2606.110 426.780 2606.430 ;
        RECT 1476.700 2606.110 1476.960 2606.430 ;
        RECT 1330.420 2033.550 1330.680 2033.870 ;
        RECT 1330.480 2033.190 1330.620 2033.550 ;
        RECT 1330.420 2032.870 1330.680 2033.190 ;
        RECT 1366.300 2032.930 1366.560 2033.190 ;
        RECT 1366.760 2032.930 1367.020 2033.190 ;
        RECT 1366.300 2032.870 1367.020 2032.930 ;
        RECT 988.640 2032.530 988.900 2032.850 ;
        RECT 1366.360 2032.790 1366.960 2032.870 ;
        RECT 646.850 1829.355 647.130 1829.725 ;
        RECT 646.920 1828.510 647.060 1829.355 ;
        RECT 988.700 1828.510 988.840 2032.530 ;
        RECT 1476.760 2032.365 1476.900 2606.110 ;
        RECT 1449.090 2031.995 1449.370 2032.365 ;
        RECT 1476.690 2031.995 1476.970 2032.365 ;
        RECT 1449.100 2031.850 1449.360 2031.995 ;
        RECT 1476.760 2030.130 1476.900 2031.995 ;
        RECT 1476.700 2029.810 1476.960 2030.130 ;
        RECT 1479.920 2029.810 1480.180 2030.130 ;
        RECT 1479.980 1928.810 1480.120 2029.810 ;
        RECT 1479.920 1928.490 1480.180 1928.810 ;
        RECT 1941.300 1928.490 1941.560 1928.810 ;
        RECT 1941.360 1917.095 1941.500 1928.490 ;
        RECT 1941.250 1913.095 1941.530 1917.095 ;
        RECT 646.860 1828.190 647.120 1828.510 ;
        RECT 988.640 1828.190 988.900 1828.510 ;
        RECT 646.920 588.530 647.060 1828.190 ;
        RECT 717.010 600.170 717.290 604.000 ;
        RECT 715.460 600.030 717.290 600.170 ;
        RECT 646.860 588.210 647.120 588.530 ;
        RECT 676.300 588.210 676.560 588.530 ;
        RECT 676.360 586.490 676.500 588.210 ;
        RECT 715.460 587.930 715.600 600.030 ;
        RECT 717.010 600.000 717.290 600.030 ;
        RECT 715.000 587.850 715.600 587.930 ;
        RECT 683.200 587.530 683.460 587.850 ;
        RECT 714.940 587.790 715.600 587.850 ;
        RECT 714.940 587.530 715.200 587.790 ;
        RECT 683.260 586.490 683.400 587.530 ;
        RECT 676.300 586.170 676.560 586.490 ;
        RECT 683.200 586.170 683.460 586.490 ;
        RECT 677.220 585.150 677.480 585.470 ;
        RECT 677.280 45.890 677.420 585.150 ;
        RECT 91.640 45.570 91.900 45.890 ;
        RECT 677.220 45.570 677.480 45.890 ;
        RECT 91.700 2.400 91.840 45.570 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 1487.270 2864.360 1487.550 2864.640 ;
        RECT 426.510 2665.120 426.790 2665.400 ;
        RECT 646.850 1829.400 647.130 1829.680 ;
        RECT 1449.090 2032.040 1449.370 2032.320 ;
        RECT 1476.690 2032.040 1476.970 2032.320 ;
      LAYER met3 ;
        RECT 1500.000 2864.840 1504.000 2865.120 ;
        RECT 1487.245 2864.650 1487.575 2864.665 ;
        RECT 1499.910 2864.650 1504.000 2864.840 ;
        RECT 1487.245 2864.520 1504.000 2864.650 ;
        RECT 1487.245 2864.350 1500.210 2864.520 ;
        RECT 1487.245 2864.335 1487.575 2864.350 ;
        RECT 430.000 2668.320 434.000 2668.640 ;
        RECT 429.950 2668.040 434.000 2668.320 ;
        RECT 426.485 2665.410 426.815 2665.425 ;
        RECT 429.950 2665.410 430.250 2668.040 ;
        RECT 426.485 2665.110 430.250 2665.410 ;
        RECT 426.485 2665.095 426.815 2665.110 ;
        RECT 1449.065 2032.330 1449.395 2032.345 ;
        RECT 1476.665 2032.330 1476.995 2032.345 ;
        RECT 1449.065 2032.030 1476.995 2032.330 ;
        RECT 1449.065 2032.015 1449.395 2032.030 ;
        RECT 1476.665 2032.015 1476.995 2032.030 ;
        RECT 627.030 1829.690 631.030 1829.840 ;
        RECT 646.825 1829.690 647.155 1829.705 ;
        RECT 627.030 1829.390 647.155 1829.690 ;
        RECT 627.030 1829.240 631.030 1829.390 ;
        RECT 646.825 1829.375 647.155 1829.390 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 879.590 2918.460 879.910 2918.520 ;
        RECT 1513.930 2918.460 1514.250 2918.520 ;
        RECT 879.590 2918.320 1514.250 2918.460 ;
        RECT 879.590 2918.260 879.910 2918.320 ;
        RECT 1513.930 2918.260 1514.250 2918.320 ;
        RECT 665.230 1990.600 665.550 1990.660 ;
        RECT 879.590 1990.600 879.910 1990.660 ;
        RECT 665.230 1990.460 879.910 1990.600 ;
        RECT 665.230 1990.400 665.550 1990.460 ;
        RECT 879.590 1990.400 879.910 1990.460 ;
        RECT 479.390 1987.880 479.710 1987.940 ;
        RECT 665.230 1987.880 665.550 1987.940 ;
        RECT 479.390 1987.740 665.550 1987.880 ;
        RECT 479.390 1987.680 479.710 1987.740 ;
        RECT 665.230 1987.680 665.550 1987.740 ;
        RECT 876.370 588.440 876.690 588.500 ;
        RECT 877.290 588.440 877.610 588.500 ;
        RECT 979.870 588.440 980.190 588.500 ;
        RECT 876.370 588.300 980.190 588.440 ;
        RECT 876.370 588.240 876.690 588.300 ;
        RECT 877.290 588.240 877.610 588.300 ;
        RECT 979.870 588.240 980.190 588.300 ;
        RECT 603.130 43.420 603.450 43.480 ;
        RECT 877.290 43.420 877.610 43.480 ;
        RECT 603.130 43.280 877.610 43.420 ;
        RECT 603.130 43.220 603.450 43.280 ;
        RECT 877.290 43.220 877.610 43.280 ;
      LAYER via ;
        RECT 879.620 2918.260 879.880 2918.520 ;
        RECT 1513.960 2918.260 1514.220 2918.520 ;
        RECT 665.260 1990.400 665.520 1990.660 ;
        RECT 879.620 1990.400 879.880 1990.660 ;
        RECT 479.420 1987.680 479.680 1987.940 ;
        RECT 665.260 1987.680 665.520 1987.940 ;
        RECT 876.400 588.240 876.660 588.500 ;
        RECT 877.320 588.240 877.580 588.500 ;
        RECT 979.900 588.240 980.160 588.500 ;
        RECT 603.160 43.220 603.420 43.480 ;
        RECT 877.320 43.220 877.580 43.480 ;
      LAYER met2 ;
        RECT 879.620 2918.230 879.880 2918.550 ;
        RECT 1513.960 2918.230 1514.220 2918.550 ;
        RECT 879.680 1990.690 879.820 2918.230 ;
        RECT 1514.020 2900.055 1514.160 2918.230 ;
        RECT 1513.890 2896.055 1514.170 2900.055 ;
        RECT 665.260 1990.370 665.520 1990.690 ;
        RECT 879.620 1990.370 879.880 1990.690 ;
        RECT 665.320 1987.970 665.460 1990.370 ;
        RECT 479.420 1987.650 479.680 1987.970 ;
        RECT 665.260 1987.650 665.520 1987.970 ;
        RECT 477.850 1981.250 478.130 1981.750 ;
        RECT 479.480 1981.250 479.620 1987.650 ;
        RECT 477.850 1981.110 479.620 1981.250 ;
        RECT 477.850 1977.750 478.130 1981.110 ;
        RECT 665.320 590.085 665.460 1987.650 ;
        RECT 980.590 600.170 980.870 604.000 ;
        RECT 979.960 600.030 980.870 600.170 ;
        RECT 665.250 589.715 665.530 590.085 ;
        RECT 876.390 589.715 876.670 590.085 ;
        RECT 876.460 588.530 876.600 589.715 ;
        RECT 979.960 588.530 980.100 600.030 ;
        RECT 980.590 600.000 980.870 600.030 ;
        RECT 876.400 588.210 876.660 588.530 ;
        RECT 877.320 588.210 877.580 588.530 ;
        RECT 979.900 588.210 980.160 588.530 ;
        RECT 877.380 43.510 877.520 588.210 ;
        RECT 603.160 43.190 603.420 43.510 ;
        RECT 877.320 43.190 877.580 43.510 ;
        RECT 603.220 2.400 603.360 43.190 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 665.250 589.760 665.530 590.040 ;
        RECT 876.390 589.760 876.670 590.040 ;
      LAYER met3 ;
        RECT 665.225 590.050 665.555 590.065 ;
        RECT 876.365 590.050 876.695 590.065 ;
        RECT 665.225 589.750 876.695 590.050 ;
        RECT 665.225 589.735 665.555 589.750 ;
        RECT 876.365 589.735 876.695 589.750 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 631.650 2917.100 631.970 2917.160 ;
        RECT 1620.650 2917.100 1620.970 2917.160 ;
        RECT 631.650 2916.960 1620.970 2917.100 ;
        RECT 631.650 2916.900 631.970 2916.960 ;
        RECT 1620.650 2916.900 1620.970 2916.960 ;
        RECT 403.950 1989.240 404.270 1989.300 ;
        RECT 630.730 1989.240 631.050 1989.300 ;
        RECT 631.650 1989.240 631.970 1989.300 ;
        RECT 403.950 1989.100 631.970 1989.240 ;
        RECT 403.950 1989.040 404.270 1989.100 ;
        RECT 630.730 1989.040 631.050 1989.100 ;
        RECT 631.650 1989.040 631.970 1989.100 ;
        RECT 630.730 1918.520 631.050 1918.580 ;
        RECT 631.650 1918.520 631.970 1918.580 ;
        RECT 630.730 1918.380 631.970 1918.520 ;
        RECT 630.730 1918.320 631.050 1918.380 ;
        RECT 631.650 1918.320 631.970 1918.380 ;
        RECT 631.650 1870.580 631.970 1870.640 ;
        RECT 630.820 1870.440 631.970 1870.580 ;
        RECT 630.820 1870.300 630.960 1870.440 ;
        RECT 631.650 1870.380 631.970 1870.440 ;
        RECT 630.730 1870.040 631.050 1870.300 ;
        RECT 630.730 1821.960 631.050 1822.020 ;
        RECT 631.650 1821.960 631.970 1822.020 ;
        RECT 630.730 1821.820 631.970 1821.960 ;
        RECT 630.730 1821.760 631.050 1821.820 ;
        RECT 631.650 1821.760 631.970 1821.820 ;
        RECT 631.650 1774.020 631.970 1774.080 ;
        RECT 630.820 1773.880 631.970 1774.020 ;
        RECT 630.820 1773.740 630.960 1773.880 ;
        RECT 631.650 1773.820 631.970 1773.880 ;
        RECT 630.730 1773.480 631.050 1773.740 ;
        RECT 630.730 1725.400 631.050 1725.460 ;
        RECT 631.650 1725.400 631.970 1725.460 ;
        RECT 630.730 1725.260 631.970 1725.400 ;
        RECT 630.730 1725.200 631.050 1725.260 ;
        RECT 631.650 1725.200 631.970 1725.260 ;
        RECT 630.270 1642.440 630.590 1642.500 ;
        RECT 631.650 1642.440 631.970 1642.500 ;
        RECT 630.270 1642.300 631.970 1642.440 ;
        RECT 630.270 1642.240 630.590 1642.300 ;
        RECT 631.650 1642.240 631.970 1642.300 ;
        RECT 629.350 1641.760 629.670 1641.820 ;
        RECT 630.270 1641.760 630.590 1641.820 ;
        RECT 629.350 1641.620 630.590 1641.760 ;
        RECT 629.350 1641.560 629.670 1641.620 ;
        RECT 630.270 1641.560 630.590 1641.620 ;
        RECT 629.350 1594.160 629.670 1594.220 ;
        RECT 630.730 1594.160 631.050 1594.220 ;
        RECT 629.350 1594.020 631.050 1594.160 ;
        RECT 629.350 1593.960 629.670 1594.020 ;
        RECT 630.730 1593.960 631.050 1594.020 ;
        RECT 629.810 1545.540 630.130 1545.600 ;
        RECT 630.270 1545.540 630.590 1545.600 ;
        RECT 629.810 1545.400 630.590 1545.540 ;
        RECT 629.810 1545.340 630.130 1545.400 ;
        RECT 630.270 1545.340 630.590 1545.400 ;
        RECT 629.810 1497.600 630.130 1497.660 ;
        RECT 630.730 1497.600 631.050 1497.660 ;
        RECT 629.810 1497.460 631.050 1497.600 ;
        RECT 629.810 1497.400 630.130 1497.460 ;
        RECT 630.730 1497.400 631.050 1497.460 ;
        RECT 629.810 1448.980 630.130 1449.040 ;
        RECT 630.270 1448.980 630.590 1449.040 ;
        RECT 629.810 1448.840 630.590 1448.980 ;
        RECT 629.810 1448.780 630.130 1448.840 ;
        RECT 630.270 1448.780 630.590 1448.840 ;
        RECT 629.810 1401.040 630.130 1401.100 ;
        RECT 630.730 1401.040 631.050 1401.100 ;
        RECT 629.810 1400.900 631.050 1401.040 ;
        RECT 629.810 1400.840 630.130 1400.900 ;
        RECT 630.730 1400.840 631.050 1400.900 ;
        RECT 629.810 1352.420 630.130 1352.480 ;
        RECT 630.270 1352.420 630.590 1352.480 ;
        RECT 629.810 1352.280 630.590 1352.420 ;
        RECT 629.810 1352.220 630.130 1352.280 ;
        RECT 630.270 1352.220 630.590 1352.280 ;
        RECT 629.810 1304.480 630.130 1304.540 ;
        RECT 630.730 1304.480 631.050 1304.540 ;
        RECT 629.810 1304.340 631.050 1304.480 ;
        RECT 629.810 1304.280 630.130 1304.340 ;
        RECT 630.730 1304.280 631.050 1304.340 ;
        RECT 629.810 1255.860 630.130 1255.920 ;
        RECT 630.270 1255.860 630.590 1255.920 ;
        RECT 629.810 1255.720 630.590 1255.860 ;
        RECT 629.810 1255.660 630.130 1255.720 ;
        RECT 630.270 1255.660 630.590 1255.720 ;
        RECT 629.810 1207.580 630.130 1207.640 ;
        RECT 630.730 1207.580 631.050 1207.640 ;
        RECT 629.810 1207.440 631.050 1207.580 ;
        RECT 629.810 1207.380 630.130 1207.440 ;
        RECT 630.730 1207.380 631.050 1207.440 ;
        RECT 629.810 1158.960 630.130 1159.020 ;
        RECT 630.270 1158.960 630.590 1159.020 ;
        RECT 629.810 1158.820 630.590 1158.960 ;
        RECT 629.810 1158.760 630.130 1158.820 ;
        RECT 630.270 1158.760 630.590 1158.820 ;
        RECT 629.810 1111.020 630.130 1111.080 ;
        RECT 630.730 1111.020 631.050 1111.080 ;
        RECT 629.810 1110.880 631.050 1111.020 ;
        RECT 629.810 1110.820 630.130 1110.880 ;
        RECT 630.730 1110.820 631.050 1110.880 ;
        RECT 630.270 1014.460 630.590 1014.520 ;
        RECT 633.030 1014.460 633.350 1014.520 ;
        RECT 630.270 1014.320 633.350 1014.460 ;
        RECT 630.270 1014.260 630.590 1014.320 ;
        RECT 633.030 1014.260 633.350 1014.320 ;
        RECT 632.570 773.400 632.890 773.460 ;
        RECT 632.200 773.260 632.890 773.400 ;
        RECT 632.200 773.120 632.340 773.260 ;
        RECT 632.570 773.200 632.890 773.260 ;
        RECT 632.110 772.860 632.430 773.120 ;
        RECT 632.110 724.440 632.430 724.500 ;
        RECT 632.570 724.440 632.890 724.500 ;
        RECT 632.110 724.300 632.890 724.440 ;
        RECT 632.110 724.240 632.430 724.300 ;
        RECT 632.570 724.240 632.890 724.300 ;
        RECT 632.110 593.880 632.430 593.940 ;
        RECT 631.740 593.740 632.430 593.880 ;
        RECT 631.740 593.600 631.880 593.740 ;
        RECT 632.110 593.680 632.430 593.740 ;
        RECT 631.650 593.340 631.970 593.600 ;
        RECT 630.270 448.700 630.590 448.760 ;
        RECT 631.190 448.700 631.510 448.760 ;
        RECT 630.270 448.560 631.510 448.700 ;
        RECT 630.270 448.500 630.590 448.560 ;
        RECT 631.190 448.500 631.510 448.560 ;
        RECT 631.190 386.480 631.510 386.540 ;
        RECT 631.650 386.480 631.970 386.540 ;
        RECT 631.190 386.340 631.970 386.480 ;
        RECT 631.190 386.280 631.510 386.340 ;
        RECT 631.650 386.280 631.970 386.340 ;
        RECT 631.190 283.260 631.510 283.520 ;
        RECT 630.730 283.120 631.050 283.180 ;
        RECT 631.280 283.120 631.420 283.260 ;
        RECT 630.730 282.980 631.420 283.120 ;
        RECT 630.730 282.920 631.050 282.980 ;
        RECT 629.810 234.840 630.130 234.900 ;
        RECT 630.730 234.840 631.050 234.900 ;
        RECT 629.810 234.700 631.050 234.840 ;
        RECT 629.810 234.640 630.130 234.700 ;
        RECT 630.730 234.640 631.050 234.700 ;
        RECT 629.810 234.160 630.130 234.220 ;
        RECT 630.730 234.160 631.050 234.220 ;
        RECT 629.810 234.020 631.050 234.160 ;
        RECT 629.810 233.960 630.130 234.020 ;
        RECT 630.730 233.960 631.050 234.020 ;
        RECT 629.350 137.940 629.670 138.000 ;
        RECT 630.270 137.940 630.590 138.000 ;
        RECT 629.350 137.800 630.590 137.940 ;
        RECT 629.350 137.740 629.670 137.800 ;
        RECT 630.270 137.740 630.590 137.800 ;
        RECT 628.890 90.000 629.210 90.060 ;
        RECT 629.350 90.000 629.670 90.060 ;
        RECT 628.890 89.860 629.670 90.000 ;
        RECT 628.890 89.800 629.210 89.860 ;
        RECT 629.350 89.800 629.670 89.860 ;
        RECT 628.890 48.520 629.210 48.580 ;
        RECT 629.810 48.520 630.130 48.580 ;
        RECT 628.890 48.380 630.130 48.520 ;
        RECT 628.890 48.320 629.210 48.380 ;
        RECT 629.810 48.320 630.130 48.380 ;
        RECT 621.070 22.000 621.390 22.060 ;
        RECT 629.810 22.000 630.130 22.060 ;
        RECT 621.070 21.860 630.130 22.000 ;
        RECT 621.070 21.800 621.390 21.860 ;
        RECT 629.810 21.800 630.130 21.860 ;
      LAYER via ;
        RECT 631.680 2916.900 631.940 2917.160 ;
        RECT 1620.680 2916.900 1620.940 2917.160 ;
        RECT 403.980 1989.040 404.240 1989.300 ;
        RECT 630.760 1989.040 631.020 1989.300 ;
        RECT 631.680 1989.040 631.940 1989.300 ;
        RECT 630.760 1918.320 631.020 1918.580 ;
        RECT 631.680 1918.320 631.940 1918.580 ;
        RECT 631.680 1870.380 631.940 1870.640 ;
        RECT 630.760 1870.040 631.020 1870.300 ;
        RECT 630.760 1821.760 631.020 1822.020 ;
        RECT 631.680 1821.760 631.940 1822.020 ;
        RECT 631.680 1773.820 631.940 1774.080 ;
        RECT 630.760 1773.480 631.020 1773.740 ;
        RECT 630.760 1725.200 631.020 1725.460 ;
        RECT 631.680 1725.200 631.940 1725.460 ;
        RECT 630.300 1642.240 630.560 1642.500 ;
        RECT 631.680 1642.240 631.940 1642.500 ;
        RECT 629.380 1641.560 629.640 1641.820 ;
        RECT 630.300 1641.560 630.560 1641.820 ;
        RECT 629.380 1593.960 629.640 1594.220 ;
        RECT 630.760 1593.960 631.020 1594.220 ;
        RECT 629.840 1545.340 630.100 1545.600 ;
        RECT 630.300 1545.340 630.560 1545.600 ;
        RECT 629.840 1497.400 630.100 1497.660 ;
        RECT 630.760 1497.400 631.020 1497.660 ;
        RECT 629.840 1448.780 630.100 1449.040 ;
        RECT 630.300 1448.780 630.560 1449.040 ;
        RECT 629.840 1400.840 630.100 1401.100 ;
        RECT 630.760 1400.840 631.020 1401.100 ;
        RECT 629.840 1352.220 630.100 1352.480 ;
        RECT 630.300 1352.220 630.560 1352.480 ;
        RECT 629.840 1304.280 630.100 1304.540 ;
        RECT 630.760 1304.280 631.020 1304.540 ;
        RECT 629.840 1255.660 630.100 1255.920 ;
        RECT 630.300 1255.660 630.560 1255.920 ;
        RECT 629.840 1207.380 630.100 1207.640 ;
        RECT 630.760 1207.380 631.020 1207.640 ;
        RECT 629.840 1158.760 630.100 1159.020 ;
        RECT 630.300 1158.760 630.560 1159.020 ;
        RECT 629.840 1110.820 630.100 1111.080 ;
        RECT 630.760 1110.820 631.020 1111.080 ;
        RECT 630.300 1014.260 630.560 1014.520 ;
        RECT 633.060 1014.260 633.320 1014.520 ;
        RECT 632.600 773.200 632.860 773.460 ;
        RECT 632.140 772.860 632.400 773.120 ;
        RECT 632.140 724.240 632.400 724.500 ;
        RECT 632.600 724.240 632.860 724.500 ;
        RECT 632.140 593.680 632.400 593.940 ;
        RECT 631.680 593.340 631.940 593.600 ;
        RECT 630.300 448.500 630.560 448.760 ;
        RECT 631.220 448.500 631.480 448.760 ;
        RECT 631.220 386.280 631.480 386.540 ;
        RECT 631.680 386.280 631.940 386.540 ;
        RECT 631.220 283.260 631.480 283.520 ;
        RECT 630.760 282.920 631.020 283.180 ;
        RECT 629.840 234.640 630.100 234.900 ;
        RECT 630.760 234.640 631.020 234.900 ;
        RECT 629.840 233.960 630.100 234.220 ;
        RECT 630.760 233.960 631.020 234.220 ;
        RECT 629.380 137.740 629.640 138.000 ;
        RECT 630.300 137.740 630.560 138.000 ;
        RECT 628.920 89.800 629.180 90.060 ;
        RECT 629.380 89.800 629.640 90.060 ;
        RECT 628.920 48.320 629.180 48.580 ;
        RECT 629.840 48.320 630.100 48.580 ;
        RECT 621.100 21.800 621.360 22.060 ;
        RECT 629.840 21.800 630.100 22.060 ;
      LAYER met2 ;
        RECT 631.680 2916.870 631.940 2917.190 ;
        RECT 1620.680 2916.870 1620.940 2917.190 ;
        RECT 631.740 1989.330 631.880 2916.870 ;
        RECT 1620.740 2900.055 1620.880 2916.870 ;
        RECT 1620.610 2896.055 1620.890 2900.055 ;
        RECT 403.980 1989.010 404.240 1989.330 ;
        RECT 630.760 1989.010 631.020 1989.330 ;
        RECT 631.680 1989.010 631.940 1989.330 ;
        RECT 402.410 1981.250 402.690 1981.750 ;
        RECT 404.040 1981.250 404.180 1989.010 ;
        RECT 402.410 1981.110 404.180 1981.250 ;
        RECT 402.410 1977.750 402.690 1981.110 ;
        RECT 630.820 1918.610 630.960 1989.010 ;
        RECT 630.760 1918.290 631.020 1918.610 ;
        RECT 631.680 1918.290 631.940 1918.610 ;
        RECT 631.740 1870.670 631.880 1918.290 ;
        RECT 631.680 1870.350 631.940 1870.670 ;
        RECT 630.760 1870.010 631.020 1870.330 ;
        RECT 630.820 1822.050 630.960 1870.010 ;
        RECT 630.760 1821.730 631.020 1822.050 ;
        RECT 631.680 1821.730 631.940 1822.050 ;
        RECT 631.740 1774.110 631.880 1821.730 ;
        RECT 631.680 1773.790 631.940 1774.110 ;
        RECT 630.760 1773.450 631.020 1773.770 ;
        RECT 630.820 1725.490 630.960 1773.450 ;
        RECT 630.760 1725.170 631.020 1725.490 ;
        RECT 631.680 1725.170 631.940 1725.490 ;
        RECT 631.740 1642.530 631.880 1725.170 ;
        RECT 630.300 1642.210 630.560 1642.530 ;
        RECT 631.680 1642.210 631.940 1642.530 ;
        RECT 630.360 1641.850 630.500 1642.210 ;
        RECT 629.380 1641.530 629.640 1641.850 ;
        RECT 630.300 1641.530 630.560 1641.850 ;
        RECT 629.440 1594.250 629.580 1641.530 ;
        RECT 629.380 1593.930 629.640 1594.250 ;
        RECT 630.760 1593.930 631.020 1594.250 ;
        RECT 630.820 1559.650 630.960 1593.930 ;
        RECT 630.360 1559.510 630.960 1559.650 ;
        RECT 630.360 1545.630 630.500 1559.510 ;
        RECT 629.840 1545.310 630.100 1545.630 ;
        RECT 630.300 1545.310 630.560 1545.630 ;
        RECT 629.900 1497.690 630.040 1545.310 ;
        RECT 629.840 1497.370 630.100 1497.690 ;
        RECT 630.760 1497.370 631.020 1497.690 ;
        RECT 630.820 1463.090 630.960 1497.370 ;
        RECT 630.360 1462.950 630.960 1463.090 ;
        RECT 630.360 1449.070 630.500 1462.950 ;
        RECT 629.840 1448.750 630.100 1449.070 ;
        RECT 630.300 1448.750 630.560 1449.070 ;
        RECT 629.900 1401.130 630.040 1448.750 ;
        RECT 629.840 1400.810 630.100 1401.130 ;
        RECT 630.760 1400.810 631.020 1401.130 ;
        RECT 630.820 1366.530 630.960 1400.810 ;
        RECT 630.360 1366.390 630.960 1366.530 ;
        RECT 630.360 1352.510 630.500 1366.390 ;
        RECT 629.840 1352.190 630.100 1352.510 ;
        RECT 630.300 1352.190 630.560 1352.510 ;
        RECT 629.900 1304.570 630.040 1352.190 ;
        RECT 629.840 1304.250 630.100 1304.570 ;
        RECT 630.760 1304.250 631.020 1304.570 ;
        RECT 630.820 1269.970 630.960 1304.250 ;
        RECT 630.360 1269.830 630.960 1269.970 ;
        RECT 630.360 1255.950 630.500 1269.830 ;
        RECT 629.840 1255.630 630.100 1255.950 ;
        RECT 630.300 1255.630 630.560 1255.950 ;
        RECT 629.900 1207.670 630.040 1255.630 ;
        RECT 629.840 1207.350 630.100 1207.670 ;
        RECT 630.760 1207.350 631.020 1207.670 ;
        RECT 630.820 1173.410 630.960 1207.350 ;
        RECT 630.360 1173.270 630.960 1173.410 ;
        RECT 630.360 1159.050 630.500 1173.270 ;
        RECT 629.840 1158.730 630.100 1159.050 ;
        RECT 630.300 1158.730 630.560 1159.050 ;
        RECT 629.900 1111.110 630.040 1158.730 ;
        RECT 629.840 1110.790 630.100 1111.110 ;
        RECT 630.760 1110.790 631.020 1111.110 ;
        RECT 630.820 1076.850 630.960 1110.790 ;
        RECT 630.360 1076.710 630.960 1076.850 ;
        RECT 630.360 1014.550 630.500 1076.710 ;
        RECT 633.120 1014.550 633.260 1014.705 ;
        RECT 630.300 1014.230 630.560 1014.550 ;
        RECT 633.060 1014.290 633.320 1014.550 ;
        RECT 632.660 1014.230 633.320 1014.290 ;
        RECT 632.660 1014.150 633.260 1014.230 ;
        RECT 632.660 990.490 632.800 1014.150 ;
        RECT 632.660 990.350 633.260 990.490 ;
        RECT 633.120 931.330 633.260 990.350 ;
        RECT 632.660 931.190 633.260 931.330 ;
        RECT 632.660 893.930 632.800 931.190 ;
        RECT 632.660 893.790 633.260 893.930 ;
        RECT 633.120 834.770 633.260 893.790 ;
        RECT 632.660 834.630 633.260 834.770 ;
        RECT 632.660 773.490 632.800 834.630 ;
        RECT 632.600 773.170 632.860 773.490 ;
        RECT 632.140 772.830 632.400 773.150 ;
        RECT 632.200 772.380 632.340 772.830 ;
        RECT 632.200 772.240 632.800 772.380 ;
        RECT 632.660 724.530 632.800 772.240 ;
        RECT 632.140 724.210 632.400 724.530 ;
        RECT 632.600 724.210 632.860 724.530 ;
        RECT 632.200 593.970 632.340 724.210 ;
        RECT 989.790 600.170 990.070 604.000 ;
        RECT 988.240 600.030 990.070 600.170 ;
        RECT 631.740 593.630 631.880 593.785 ;
        RECT 632.140 593.650 632.400 593.970 ;
        RECT 631.680 593.370 631.940 593.630 ;
        RECT 631.280 593.310 631.940 593.370 ;
        RECT 631.280 593.230 631.880 593.310 ;
        RECT 631.280 588.725 631.420 593.230 ;
        RECT 631.210 588.355 631.490 588.725 ;
        RECT 631.280 587.930 631.420 588.355 ;
        RECT 988.240 588.045 988.380 600.030 ;
        RECT 989.790 600.000 990.070 600.030 ;
        RECT 630.360 587.790 631.420 587.930 ;
        RECT 630.360 545.090 630.500 587.790 ;
        RECT 988.170 587.675 988.450 588.045 ;
        RECT 630.360 544.950 630.960 545.090 ;
        RECT 630.820 507.010 630.960 544.950 ;
        RECT 630.820 506.870 631.420 507.010 ;
        RECT 631.280 448.790 631.420 506.870 ;
        RECT 630.300 448.530 630.560 448.790 ;
        RECT 631.220 448.530 631.480 448.790 ;
        RECT 630.300 448.470 631.480 448.530 ;
        RECT 630.360 448.390 631.420 448.470 ;
        RECT 631.280 386.570 631.420 448.390 ;
        RECT 631.220 386.250 631.480 386.570 ;
        RECT 631.680 386.250 631.940 386.570 ;
        RECT 631.740 362.170 631.880 386.250 ;
        RECT 631.280 362.030 631.880 362.170 ;
        RECT 631.280 283.550 631.420 362.030 ;
        RECT 631.220 283.230 631.480 283.550 ;
        RECT 630.760 282.890 631.020 283.210 ;
        RECT 630.820 234.930 630.960 282.890 ;
        RECT 629.840 234.610 630.100 234.930 ;
        RECT 630.760 234.610 631.020 234.930 ;
        RECT 629.900 234.250 630.040 234.610 ;
        RECT 629.840 233.930 630.100 234.250 ;
        RECT 630.760 233.930 631.020 234.250 ;
        RECT 630.820 206.960 630.960 233.930 ;
        RECT 630.360 206.820 630.960 206.960 ;
        RECT 630.360 138.030 630.500 206.820 ;
        RECT 629.380 137.710 629.640 138.030 ;
        RECT 630.300 137.710 630.560 138.030 ;
        RECT 629.440 90.090 629.580 137.710 ;
        RECT 628.920 89.770 629.180 90.090 ;
        RECT 629.380 89.770 629.640 90.090 ;
        RECT 628.980 48.610 629.120 89.770 ;
        RECT 628.920 48.290 629.180 48.610 ;
        RECT 629.840 48.290 630.100 48.610 ;
        RECT 629.900 22.090 630.040 48.290 ;
        RECT 621.100 21.770 621.360 22.090 ;
        RECT 629.840 21.770 630.100 22.090 ;
        RECT 621.160 2.400 621.300 21.770 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 631.210 588.400 631.490 588.680 ;
        RECT 988.170 587.720 988.450 588.000 ;
      LAYER met3 ;
        RECT 631.185 588.690 631.515 588.705 ;
        RECT 631.185 588.390 665.770 588.690 ;
        RECT 631.185 588.375 631.515 588.390 ;
        RECT 665.470 588.010 665.770 588.390 ;
        RECT 988.145 588.010 988.475 588.025 ;
        RECT 665.470 587.710 988.475 588.010 ;
        RECT 988.145 587.695 988.475 587.710 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 2877.660 551.930 2877.720 ;
        RECT 1483.570 2877.660 1483.890 2877.720 ;
        RECT 551.610 2877.520 1483.890 2877.660 ;
        RECT 551.610 2877.460 551.930 2877.520 ;
        RECT 1483.570 2877.460 1483.890 2877.520 ;
        RECT 547.010 2773.960 547.330 2774.020 ;
        RECT 551.610 2773.960 551.930 2774.020 ;
        RECT 579.670 2773.960 579.990 2774.020 ;
        RECT 547.010 2773.820 579.990 2773.960 ;
        RECT 547.010 2773.760 547.330 2773.820 ;
        RECT 551.610 2773.760 551.930 2773.820 ;
        RECT 579.670 2773.760 579.990 2773.820 ;
        RECT 379.110 1990.600 379.430 1990.660 ;
        RECT 579.670 1990.600 579.990 1990.660 ;
        RECT 635.790 1990.600 636.110 1990.660 ;
        RECT 379.110 1990.460 636.110 1990.600 ;
        RECT 379.110 1990.400 379.430 1990.460 ;
        RECT 579.670 1990.400 579.990 1990.460 ;
        RECT 635.790 1990.400 636.110 1990.460 ;
        RECT 635.790 1703.980 636.110 1704.040 ;
        RECT 2021.770 1703.980 2022.090 1704.040 ;
        RECT 635.790 1703.840 2022.090 1703.980 ;
        RECT 635.790 1703.780 636.110 1703.840 ;
        RECT 2021.770 1703.780 2022.090 1703.840 ;
        RECT 551.610 1700.920 551.930 1700.980 ;
        RECT 635.790 1700.920 636.110 1700.980 ;
        RECT 551.610 1700.780 636.110 1700.920 ;
        RECT 551.610 1700.720 551.930 1700.780 ;
        RECT 635.790 1700.720 636.110 1700.780 ;
        RECT 116.910 590.820 117.230 590.880 ;
        RECT 551.610 590.820 551.930 590.880 ;
        RECT 116.910 590.680 551.930 590.820 ;
        RECT 116.910 590.620 117.230 590.680 ;
        RECT 551.610 590.620 551.930 590.680 ;
        RECT 115.530 2.960 115.850 3.020 ;
        RECT 116.910 2.960 117.230 3.020 ;
        RECT 115.530 2.820 117.230 2.960 ;
        RECT 115.530 2.760 115.850 2.820 ;
        RECT 116.910 2.760 117.230 2.820 ;
      LAYER via ;
        RECT 551.640 2877.460 551.900 2877.720 ;
        RECT 1483.600 2877.460 1483.860 2877.720 ;
        RECT 547.040 2773.760 547.300 2774.020 ;
        RECT 551.640 2773.760 551.900 2774.020 ;
        RECT 579.700 2773.760 579.960 2774.020 ;
        RECT 379.140 1990.400 379.400 1990.660 ;
        RECT 579.700 1990.400 579.960 1990.660 ;
        RECT 635.820 1990.400 636.080 1990.660 ;
        RECT 635.820 1703.780 636.080 1704.040 ;
        RECT 2021.800 1703.780 2022.060 1704.040 ;
        RECT 551.640 1700.720 551.900 1700.980 ;
        RECT 635.820 1700.720 636.080 1700.980 ;
        RECT 116.940 590.620 117.200 590.880 ;
        RECT 551.640 590.620 551.900 590.880 ;
        RECT 115.560 2.760 115.820 3.020 ;
        RECT 116.940 2.760 117.200 3.020 ;
      LAYER met2 ;
        RECT 1483.590 2878.595 1483.870 2878.965 ;
        RECT 1483.660 2877.750 1483.800 2878.595 ;
        RECT 551.640 2877.430 551.900 2877.750 ;
        RECT 1483.600 2877.430 1483.860 2877.750 ;
        RECT 551.700 2774.050 551.840 2877.430 ;
        RECT 547.040 2773.730 547.300 2774.050 ;
        RECT 551.640 2773.730 551.900 2774.050 ;
        RECT 579.700 2773.730 579.960 2774.050 ;
        RECT 547.100 2759.520 547.240 2773.730 ;
        RECT 546.930 2759.100 547.240 2759.520 ;
        RECT 546.930 2755.520 547.210 2759.100 ;
        RECT 579.760 1990.690 579.900 2773.730 ;
        RECT 379.140 1990.370 379.400 1990.690 ;
        RECT 579.700 1990.370 579.960 1990.690 ;
        RECT 635.820 1990.370 636.080 1990.690 ;
        RECT 377.570 1981.250 377.850 1981.750 ;
        RECT 379.200 1981.250 379.340 1990.370 ;
        RECT 377.570 1981.110 379.340 1981.250 ;
        RECT 377.570 1977.750 377.850 1981.110 ;
        RECT 635.880 1704.070 636.020 1990.370 ;
        RECT 2025.890 1750.730 2026.170 1754.000 ;
        RECT 2021.860 1750.590 2026.170 1750.730 ;
        RECT 2021.860 1704.070 2022.000 1750.590 ;
        RECT 2025.890 1750.000 2026.170 1750.590 ;
        RECT 635.820 1703.750 636.080 1704.070 ;
        RECT 2021.800 1703.750 2022.060 1704.070 ;
        RECT 635.880 1701.010 636.020 1703.750 ;
        RECT 551.640 1700.690 551.900 1701.010 ;
        RECT 635.820 1700.690 636.080 1701.010 ;
        RECT 551.700 592.125 551.840 1700.690 ;
        RECT 729.430 600.170 729.710 604.000 ;
        RECT 727.880 600.030 729.710 600.170 ;
        RECT 727.880 592.125 728.020 600.030 ;
        RECT 729.430 600.000 729.710 600.030 ;
        RECT 551.630 591.755 551.910 592.125 ;
        RECT 727.810 591.755 728.090 592.125 ;
        RECT 551.700 590.910 551.840 591.755 ;
        RECT 116.940 590.590 117.200 590.910 ;
        RECT 551.640 590.590 551.900 590.910 ;
        RECT 117.000 3.050 117.140 590.590 ;
        RECT 115.560 2.730 115.820 3.050 ;
        RECT 116.940 2.730 117.200 3.050 ;
        RECT 115.620 2.400 115.760 2.730 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 1483.590 2878.640 1483.870 2878.920 ;
        RECT 551.630 591.800 551.910 592.080 ;
        RECT 727.810 591.800 728.090 592.080 ;
      LAYER met3 ;
        RECT 1500.000 2881.160 1504.000 2881.440 ;
        RECT 1499.910 2880.840 1504.000 2881.160 ;
        RECT 1483.565 2878.930 1483.895 2878.945 ;
        RECT 1499.910 2878.930 1500.210 2880.840 ;
        RECT 1483.565 2878.630 1500.210 2878.930 ;
        RECT 1483.565 2878.615 1483.895 2878.630 ;
        RECT 551.605 592.090 551.935 592.105 ;
        RECT 727.785 592.090 728.115 592.105 ;
        RECT 551.605 591.790 728.115 592.090 ;
        RECT 551.605 591.775 551.935 591.790 ;
        RECT 727.785 591.775 728.115 591.790 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 460.530 2769.880 460.850 2769.940 ;
        RECT 576.450 2769.880 576.770 2769.940 ;
        RECT 460.530 2769.740 576.770 2769.880 ;
        RECT 460.530 2769.680 460.850 2769.740 ;
        RECT 576.450 2769.680 576.770 2769.740 ;
        RECT 558.510 2489.720 558.830 2489.780 ;
        RECT 576.450 2489.720 576.770 2489.780 ;
        RECT 1566.370 2489.720 1566.690 2489.780 ;
        RECT 558.510 2489.580 1566.690 2489.720 ;
        RECT 558.510 2489.520 558.830 2489.580 ;
        RECT 576.450 2489.520 576.770 2489.580 ;
        RECT 1566.370 2489.520 1566.690 2489.580 ;
        RECT 554.830 1988.560 555.150 1988.620 ;
        RECT 558.510 1988.560 558.830 1988.620 ;
        RECT 636.250 1988.560 636.570 1988.620 ;
        RECT 554.830 1988.420 636.570 1988.560 ;
        RECT 554.830 1988.360 555.150 1988.420 ;
        RECT 558.510 1988.360 558.830 1988.420 ;
        RECT 636.250 1988.360 636.570 1988.420 ;
        RECT 636.250 1704.320 636.570 1704.380 ;
        RECT 2042.470 1704.320 2042.790 1704.380 ;
        RECT 636.250 1704.180 2042.790 1704.320 ;
        RECT 636.250 1704.120 636.570 1704.180 ;
        RECT 2042.470 1704.120 2042.790 1704.180 ;
        RECT 558.510 1701.260 558.830 1701.320 ;
        RECT 636.250 1701.260 636.570 1701.320 ;
        RECT 558.510 1701.120 636.570 1701.260 ;
        RECT 558.510 1701.060 558.830 1701.120 ;
        RECT 636.250 1701.060 636.570 1701.120 ;
        RECT 144.510 591.160 144.830 591.220 ;
        RECT 558.510 591.160 558.830 591.220 ;
        RECT 144.510 591.020 558.830 591.160 ;
        RECT 144.510 590.960 144.830 591.020 ;
        RECT 558.510 590.960 558.830 591.020 ;
        RECT 558.510 586.740 558.830 586.800 ;
        RECT 740.210 586.740 740.530 586.800 ;
        RECT 558.510 586.600 740.530 586.740 ;
        RECT 558.510 586.540 558.830 586.600 ;
        RECT 740.210 586.540 740.530 586.600 ;
        RECT 139.450 16.900 139.770 16.960 ;
        RECT 144.510 16.900 144.830 16.960 ;
        RECT 139.450 16.760 144.830 16.900 ;
        RECT 139.450 16.700 139.770 16.760 ;
        RECT 144.510 16.700 144.830 16.760 ;
      LAYER via ;
        RECT 460.560 2769.680 460.820 2769.940 ;
        RECT 576.480 2769.680 576.740 2769.940 ;
        RECT 558.540 2489.520 558.800 2489.780 ;
        RECT 576.480 2489.520 576.740 2489.780 ;
        RECT 1566.400 2489.520 1566.660 2489.780 ;
        RECT 554.860 1988.360 555.120 1988.620 ;
        RECT 558.540 1988.360 558.800 1988.620 ;
        RECT 636.280 1988.360 636.540 1988.620 ;
        RECT 636.280 1704.120 636.540 1704.380 ;
        RECT 2042.500 1704.120 2042.760 1704.380 ;
        RECT 558.540 1701.060 558.800 1701.320 ;
        RECT 636.280 1701.060 636.540 1701.320 ;
        RECT 144.540 590.960 144.800 591.220 ;
        RECT 558.540 590.960 558.800 591.220 ;
        RECT 558.540 586.540 558.800 586.800 ;
        RECT 740.240 586.540 740.500 586.800 ;
        RECT 139.480 16.700 139.740 16.960 ;
        RECT 144.540 16.700 144.800 16.960 ;
      LAYER met2 ;
        RECT 460.560 2769.650 460.820 2769.970 ;
        RECT 576.480 2769.650 576.740 2769.970 ;
        RECT 460.620 2759.520 460.760 2769.650 ;
        RECT 460.450 2759.100 460.760 2759.520 ;
        RECT 460.450 2755.520 460.730 2759.100 ;
        RECT 576.540 2489.810 576.680 2769.650 ;
        RECT 1566.330 2500.000 1566.610 2504.000 ;
        RECT 1566.460 2489.810 1566.600 2500.000 ;
        RECT 558.540 2489.490 558.800 2489.810 ;
        RECT 576.480 2489.490 576.740 2489.810 ;
        RECT 1566.400 2489.490 1566.660 2489.810 ;
        RECT 558.600 1988.650 558.740 2489.490 ;
        RECT 554.860 1988.330 555.120 1988.650 ;
        RECT 558.540 1988.330 558.800 1988.650 ;
        RECT 636.280 1988.330 636.540 1988.650 ;
        RECT 553.290 1981.250 553.570 1981.750 ;
        RECT 554.920 1981.250 555.060 1988.330 ;
        RECT 553.290 1981.110 555.060 1981.250 ;
        RECT 553.290 1977.750 553.570 1981.110 ;
        RECT 636.340 1704.410 636.480 1988.330 ;
        RECT 2048.890 1750.730 2049.170 1754.000 ;
        RECT 2042.560 1750.590 2049.170 1750.730 ;
        RECT 2042.560 1704.410 2042.700 1750.590 ;
        RECT 2048.890 1750.000 2049.170 1750.590 ;
        RECT 636.280 1704.090 636.540 1704.410 ;
        RECT 2042.500 1704.090 2042.760 1704.410 ;
        RECT 636.340 1701.350 636.480 1704.090 ;
        RECT 558.540 1701.030 558.800 1701.350 ;
        RECT 636.280 1701.030 636.540 1701.350 ;
        RECT 558.600 591.250 558.740 1701.030 ;
        RECT 741.850 600.170 742.130 604.000 ;
        RECT 740.300 600.030 742.130 600.170 ;
        RECT 144.540 590.930 144.800 591.250 ;
        RECT 558.540 590.930 558.800 591.250 ;
        RECT 144.600 16.990 144.740 590.930 ;
        RECT 558.600 586.830 558.740 590.930 ;
        RECT 740.300 586.830 740.440 600.030 ;
        RECT 741.850 600.000 742.130 600.030 ;
        RECT 558.540 586.510 558.800 586.830 ;
        RECT 740.240 586.510 740.500 586.830 ;
        RECT 139.480 16.670 139.740 16.990 ;
        RECT 144.540 16.670 144.800 16.990 ;
        RECT 139.540 2.400 139.680 16.670 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 590.250 2488.020 590.570 2488.080 ;
        RECT 1513.010 2488.020 1513.330 2488.080 ;
        RECT 590.250 2487.880 1513.330 2488.020 ;
        RECT 590.250 2487.820 590.570 2487.880 ;
        RECT 1513.010 2487.820 1513.330 2487.880 ;
        RECT 1510.710 2484.280 1511.030 2484.340 ;
        RECT 1513.010 2484.280 1513.330 2484.340 ;
        RECT 1510.710 2484.140 1513.330 2484.280 ;
        RECT 1510.710 2484.080 1511.030 2484.140 ;
        RECT 1513.010 2484.080 1513.330 2484.140 ;
        RECT 1507.950 1907.640 1508.270 1907.700 ;
        RECT 1510.710 1907.640 1511.030 1907.700 ;
        RECT 1904.470 1907.640 1904.790 1907.700 ;
        RECT 1507.950 1907.500 1904.790 1907.640 ;
        RECT 1507.950 1907.440 1508.270 1907.500 ;
        RECT 1510.710 1907.440 1511.030 1907.500 ;
        RECT 1904.470 1907.440 1904.790 1907.500 ;
        RECT 537.810 1690.380 538.130 1690.440 ;
        RECT 1507.950 1690.380 1508.270 1690.440 ;
        RECT 537.810 1690.240 1508.270 1690.380 ;
        RECT 537.810 1690.180 538.130 1690.240 ;
        RECT 1507.950 1690.180 1508.270 1690.240 ;
        RECT 158.310 591.500 158.630 591.560 ;
        RECT 537.810 591.500 538.130 591.560 ;
        RECT 158.310 591.360 538.130 591.500 ;
        RECT 158.310 591.300 158.630 591.360 ;
        RECT 537.810 591.300 538.130 591.360 ;
        RECT 579.670 590.820 579.990 590.880 ;
        RECT 614.630 590.820 614.950 590.880 ;
        RECT 579.670 590.680 614.950 590.820 ;
        RECT 579.670 590.620 579.990 590.680 ;
        RECT 614.630 590.620 614.950 590.680 ;
        RECT 537.810 589.460 538.130 589.520 ;
        RECT 579.670 589.460 579.990 589.520 ;
        RECT 537.810 589.320 579.990 589.460 ;
        RECT 537.810 589.260 538.130 589.320 ;
        RECT 579.670 589.260 579.990 589.320 ;
        RECT 614.630 589.460 614.950 589.520 ;
        RECT 749.410 589.460 749.730 589.520 ;
        RECT 614.630 589.320 749.730 589.460 ;
        RECT 614.630 589.260 614.950 589.320 ;
        RECT 749.410 589.260 749.730 589.320 ;
      LAYER via ;
        RECT 590.280 2487.820 590.540 2488.080 ;
        RECT 1513.040 2487.820 1513.300 2488.080 ;
        RECT 1510.740 2484.080 1511.000 2484.340 ;
        RECT 1513.040 2484.080 1513.300 2484.340 ;
        RECT 1507.980 1907.440 1508.240 1907.700 ;
        RECT 1510.740 1907.440 1511.000 1907.700 ;
        RECT 1904.500 1907.440 1904.760 1907.700 ;
        RECT 537.840 1690.180 538.100 1690.440 ;
        RECT 1507.980 1690.180 1508.240 1690.440 ;
        RECT 158.340 591.300 158.600 591.560 ;
        RECT 537.840 591.300 538.100 591.560 ;
        RECT 579.700 590.620 579.960 590.880 ;
        RECT 614.660 590.620 614.920 590.880 ;
        RECT 537.840 589.260 538.100 589.520 ;
        RECT 579.700 589.260 579.960 589.520 ;
        RECT 614.660 589.260 614.920 589.520 ;
        RECT 749.440 589.260 749.700 589.520 ;
      LAYER met2 ;
        RECT 590.270 2732.395 590.550 2732.765 ;
        RECT 590.340 2488.110 590.480 2732.395 ;
        RECT 1512.970 2500.000 1513.250 2504.000 ;
        RECT 1513.100 2488.110 1513.240 2500.000 ;
        RECT 590.280 2487.790 590.540 2488.110 ;
        RECT 1513.040 2487.790 1513.300 2488.110 ;
        RECT 1513.100 2484.370 1513.240 2487.790 ;
        RECT 1510.740 2484.050 1511.000 2484.370 ;
        RECT 1513.040 2484.050 1513.300 2484.370 ;
        RECT 1510.800 1907.730 1510.940 2484.050 ;
        RECT 1507.980 1907.410 1508.240 1907.730 ;
        RECT 1510.740 1907.410 1511.000 1907.730 ;
        RECT 1904.500 1907.410 1904.760 1907.730 ;
        RECT 537.650 1700.410 537.930 1704.000 ;
        RECT 537.650 1700.000 538.040 1700.410 ;
        RECT 537.900 1690.470 538.040 1700.000 ;
        RECT 1508.040 1690.470 1508.180 1907.410 ;
        RECT 1904.560 1907.245 1904.700 1907.410 ;
        RECT 1904.490 1906.875 1904.770 1907.245 ;
        RECT 537.840 1690.150 538.100 1690.470 ;
        RECT 1507.980 1690.150 1508.240 1690.470 ;
        RECT 537.900 591.590 538.040 1690.150 ;
        RECT 751.050 600.170 751.330 604.000 ;
        RECT 749.500 600.030 751.330 600.170 ;
        RECT 158.340 591.270 158.600 591.590 ;
        RECT 537.840 591.270 538.100 591.590 ;
        RECT 158.400 17.410 158.540 591.270 ;
        RECT 537.900 589.550 538.040 591.270 ;
        RECT 579.700 590.590 579.960 590.910 ;
        RECT 614.660 590.590 614.920 590.910 ;
        RECT 579.760 589.550 579.900 590.590 ;
        RECT 614.720 589.550 614.860 590.590 ;
        RECT 749.500 589.550 749.640 600.030 ;
        RECT 751.050 600.000 751.330 600.030 ;
        RECT 537.840 589.230 538.100 589.550 ;
        RECT 579.700 589.230 579.960 589.550 ;
        RECT 614.660 589.230 614.920 589.550 ;
        RECT 749.440 589.230 749.700 589.550 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 590.270 2732.440 590.550 2732.720 ;
        RECT 1904.490 1906.920 1904.770 1907.200 ;
      LAYER met3 ;
        RECT 574.800 2733.320 578.800 2733.920 ;
        RECT 578.070 2732.730 578.370 2733.320 ;
        RECT 590.245 2732.730 590.575 2732.745 ;
        RECT 578.070 2732.430 590.575 2732.730 ;
        RECT 590.245 2732.415 590.575 2732.430 ;
        RECT 1904.465 1907.210 1904.795 1907.225 ;
        RECT 1904.465 1907.040 1920.650 1907.210 ;
        RECT 1904.465 1906.910 1924.000 1907.040 ;
        RECT 1904.465 1906.895 1904.795 1906.910 ;
        RECT 1920.000 1906.440 1924.000 1906.910 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1714.950 2897.380 1715.270 2897.440 ;
        RECT 1652.480 2897.240 1715.270 2897.380 ;
        RECT 1576.030 2896.700 1576.350 2896.760 ;
        RECT 1576.030 2896.560 1576.720 2896.700 ;
        RECT 1576.030 2896.500 1576.350 2896.560 ;
        RECT 1437.570 2894.660 1437.890 2894.720 ;
        RECT 1457.350 2894.660 1457.670 2894.720 ;
        RECT 1437.570 2894.520 1457.670 2894.660 ;
        RECT 1437.570 2894.460 1437.890 2894.520 ;
        RECT 1457.350 2894.460 1457.670 2894.520 ;
        RECT 713.990 2893.640 714.310 2893.700 ;
        RECT 738.830 2893.640 739.150 2893.700 ;
        RECT 713.990 2893.500 739.150 2893.640 ;
        RECT 713.990 2893.440 714.310 2893.500 ;
        RECT 738.830 2893.440 739.150 2893.500 ;
        RECT 810.590 2893.640 810.910 2893.700 ;
        RECT 835.430 2893.640 835.750 2893.700 ;
        RECT 810.590 2893.500 835.750 2893.640 ;
        RECT 810.590 2893.440 810.910 2893.500 ;
        RECT 835.430 2893.440 835.750 2893.500 ;
        RECT 886.490 2893.640 886.810 2893.700 ;
        RECT 927.890 2893.640 928.210 2893.700 ;
        RECT 886.490 2893.500 928.210 2893.640 ;
        RECT 886.490 2893.440 886.810 2893.500 ;
        RECT 927.890 2893.440 928.210 2893.500 ;
        RECT 1293.590 2893.640 1293.910 2893.700 ;
        RECT 1318.430 2893.640 1318.750 2893.700 ;
        RECT 1293.590 2893.500 1318.750 2893.640 ;
        RECT 1293.590 2893.440 1293.910 2893.500 ;
        RECT 1318.430 2893.440 1318.750 2893.500 ;
        RECT 575.990 2892.620 576.310 2892.680 ;
        RECT 579.670 2892.620 579.990 2892.680 ;
        RECT 575.990 2892.480 579.990 2892.620 ;
        RECT 575.990 2892.420 576.310 2892.480 ;
        RECT 579.670 2892.420 579.990 2892.480 ;
        RECT 1457.350 2892.620 1457.670 2892.680 ;
        RECT 1501.510 2892.620 1501.830 2892.680 ;
        RECT 1457.350 2892.480 1501.830 2892.620 ;
        RECT 1457.350 2892.420 1457.670 2892.480 ;
        RECT 1501.510 2892.420 1501.830 2892.480 ;
        RECT 619.690 2891.600 620.010 2891.660 ;
        RECT 713.990 2891.600 714.310 2891.660 ;
        RECT 619.690 2891.460 714.310 2891.600 ;
        RECT 619.690 2891.400 620.010 2891.460 ;
        RECT 713.990 2891.400 714.310 2891.460 ;
        RECT 738.830 2891.600 739.150 2891.660 ;
        RECT 810.590 2891.600 810.910 2891.660 ;
        RECT 738.830 2891.460 810.910 2891.600 ;
        RECT 738.830 2891.400 739.150 2891.460 ;
        RECT 810.590 2891.400 810.910 2891.460 ;
        RECT 835.430 2891.600 835.750 2891.660 ;
        RECT 886.490 2891.600 886.810 2891.660 ;
        RECT 835.430 2891.460 886.810 2891.600 ;
        RECT 835.430 2891.400 835.750 2891.460 ;
        RECT 886.490 2891.400 886.810 2891.460 ;
        RECT 927.890 2891.600 928.210 2891.660 ;
        RECT 1293.590 2891.600 1293.910 2891.660 ;
        RECT 927.890 2891.460 1293.910 2891.600 ;
        RECT 927.890 2891.400 928.210 2891.460 ;
        RECT 1293.590 2891.400 1293.910 2891.460 ;
        RECT 1318.430 2891.600 1318.750 2891.660 ;
        RECT 1437.570 2891.600 1437.890 2891.660 ;
        RECT 1318.430 2891.460 1437.890 2891.600 ;
        RECT 1318.430 2891.400 1318.750 2891.460 ;
        RECT 1437.570 2891.400 1437.890 2891.460 ;
        RECT 1576.580 2890.920 1576.720 2896.560 ;
        RECT 1601.790 2896.500 1602.110 2896.760 ;
        RECT 1601.880 2893.640 1602.020 2896.500 ;
        RECT 1652.480 2894.660 1652.620 2897.240 ;
        RECT 1714.950 2897.180 1715.270 2897.240 ;
        RECT 1628.560 2894.520 1652.620 2894.660 ;
        RECT 1628.560 2893.640 1628.700 2894.520 ;
        RECT 1601.880 2893.500 1628.700 2893.640 ;
        RECT 1575.660 2890.780 1576.720 2890.920 ;
        RECT 1575.660 2890.240 1575.800 2890.780 ;
        RECT 1574.740 2890.100 1575.800 2890.240 ;
        RECT 1501.510 2889.900 1501.830 2889.960 ;
        RECT 1574.740 2889.900 1574.880 2890.100 ;
        RECT 1501.510 2889.760 1574.880 2889.900 ;
        RECT 1501.510 2889.700 1501.830 2889.760 ;
        RECT 572.310 2594.100 572.630 2594.160 ;
        RECT 575.990 2594.100 576.310 2594.160 ;
        RECT 572.310 2593.960 576.310 2594.100 ;
        RECT 572.310 2593.900 572.630 2593.960 ;
        RECT 575.990 2593.900 576.310 2593.960 ;
        RECT 989.990 2036.160 990.310 2036.220 ;
        RECT 2056.270 2036.160 2056.590 2036.220 ;
        RECT 989.990 2036.020 2056.590 2036.160 ;
        RECT 989.990 2035.960 990.310 2036.020 ;
        RECT 2056.270 2035.960 2056.590 2036.020 ;
        RECT 503.310 1991.280 503.630 1991.340 ;
        RECT 569.090 1991.280 569.410 1991.340 ;
        RECT 647.290 1991.280 647.610 1991.340 ;
        RECT 503.310 1991.140 647.610 1991.280 ;
        RECT 503.310 1991.080 503.630 1991.140 ;
        RECT 569.090 1991.080 569.410 1991.140 ;
        RECT 647.290 1991.080 647.610 1991.140 ;
        RECT 647.290 1987.200 647.610 1987.260 ;
        RECT 989.990 1987.200 990.310 1987.260 ;
        RECT 647.290 1987.060 990.310 1987.200 ;
        RECT 647.290 1987.000 647.610 1987.060 ;
        RECT 989.990 1987.000 990.310 1987.060 ;
        RECT 174.870 19.960 175.190 20.020 ;
        RECT 759.530 19.960 759.850 20.020 ;
        RECT 174.870 19.820 759.850 19.960 ;
        RECT 174.870 19.760 175.190 19.820 ;
        RECT 759.530 19.760 759.850 19.820 ;
      LAYER via ;
        RECT 1576.060 2896.500 1576.320 2896.760 ;
        RECT 1437.600 2894.460 1437.860 2894.720 ;
        RECT 1457.380 2894.460 1457.640 2894.720 ;
        RECT 714.020 2893.440 714.280 2893.700 ;
        RECT 738.860 2893.440 739.120 2893.700 ;
        RECT 810.620 2893.440 810.880 2893.700 ;
        RECT 835.460 2893.440 835.720 2893.700 ;
        RECT 886.520 2893.440 886.780 2893.700 ;
        RECT 927.920 2893.440 928.180 2893.700 ;
        RECT 1293.620 2893.440 1293.880 2893.700 ;
        RECT 1318.460 2893.440 1318.720 2893.700 ;
        RECT 576.020 2892.420 576.280 2892.680 ;
        RECT 579.700 2892.420 579.960 2892.680 ;
        RECT 1457.380 2892.420 1457.640 2892.680 ;
        RECT 1501.540 2892.420 1501.800 2892.680 ;
        RECT 619.720 2891.400 619.980 2891.660 ;
        RECT 714.020 2891.400 714.280 2891.660 ;
        RECT 738.860 2891.400 739.120 2891.660 ;
        RECT 810.620 2891.400 810.880 2891.660 ;
        RECT 835.460 2891.400 835.720 2891.660 ;
        RECT 886.520 2891.400 886.780 2891.660 ;
        RECT 927.920 2891.400 928.180 2891.660 ;
        RECT 1293.620 2891.400 1293.880 2891.660 ;
        RECT 1318.460 2891.400 1318.720 2891.660 ;
        RECT 1437.600 2891.400 1437.860 2891.660 ;
        RECT 1601.820 2896.500 1602.080 2896.760 ;
        RECT 1714.980 2897.180 1715.240 2897.440 ;
        RECT 1501.540 2889.700 1501.800 2889.960 ;
        RECT 572.340 2593.900 572.600 2594.160 ;
        RECT 576.020 2593.900 576.280 2594.160 ;
        RECT 990.020 2035.960 990.280 2036.220 ;
        RECT 2056.300 2035.960 2056.560 2036.220 ;
        RECT 503.340 1991.080 503.600 1991.340 ;
        RECT 569.120 1991.080 569.380 1991.340 ;
        RECT 647.320 1991.080 647.580 1991.340 ;
        RECT 647.320 1987.000 647.580 1987.260 ;
        RECT 990.020 1987.000 990.280 1987.260 ;
        RECT 174.900 19.760 175.160 20.020 ;
        RECT 759.560 19.760 759.820 20.020 ;
      LAYER met2 ;
        RECT 1714.980 2897.210 1715.240 2897.470 ;
        RECT 1716.290 2897.210 1716.570 2900.055 ;
        RECT 1714.980 2897.150 1716.570 2897.210 ;
        RECT 1715.040 2897.070 1716.570 2897.150 ;
        RECT 1576.060 2896.645 1576.320 2896.790 ;
        RECT 1601.820 2896.645 1602.080 2896.790 ;
        RECT 1576.050 2896.275 1576.330 2896.645 ;
        RECT 1601.810 2896.275 1602.090 2896.645 ;
        RECT 1716.290 2896.055 1716.570 2897.070 ;
        RECT 1437.600 2894.430 1437.860 2894.750 ;
        RECT 1457.380 2894.430 1457.640 2894.750 ;
        RECT 714.020 2893.410 714.280 2893.730 ;
        RECT 738.860 2893.410 739.120 2893.730 ;
        RECT 810.620 2893.410 810.880 2893.730 ;
        RECT 835.460 2893.410 835.720 2893.730 ;
        RECT 886.520 2893.410 886.780 2893.730 ;
        RECT 927.920 2893.410 928.180 2893.730 ;
        RECT 1293.620 2893.410 1293.880 2893.730 ;
        RECT 1318.460 2893.410 1318.720 2893.730 ;
        RECT 576.020 2892.390 576.280 2892.710 ;
        RECT 579.700 2892.565 579.960 2892.710 ;
        RECT 547.850 2600.660 548.130 2604.000 ;
        RECT 547.850 2600.000 548.160 2600.660 ;
        RECT 548.020 2594.045 548.160 2600.000 ;
        RECT 547.950 2593.675 548.230 2594.045 ;
        RECT 569.110 2593.675 569.390 2594.045 ;
        RECT 572.330 2593.845 572.610 2594.215 ;
        RECT 576.080 2594.190 576.220 2892.390 ;
        RECT 579.690 2892.195 579.970 2892.565 ;
        RECT 619.710 2892.195 619.990 2892.565 ;
        RECT 619.780 2891.690 619.920 2892.195 ;
        RECT 714.080 2891.690 714.220 2893.410 ;
        RECT 738.920 2891.690 739.060 2893.410 ;
        RECT 810.680 2891.690 810.820 2893.410 ;
        RECT 835.520 2891.690 835.660 2893.410 ;
        RECT 886.580 2891.690 886.720 2893.410 ;
        RECT 927.980 2891.690 928.120 2893.410 ;
        RECT 1293.680 2891.690 1293.820 2893.410 ;
        RECT 1318.520 2891.690 1318.660 2893.410 ;
        RECT 1437.660 2891.690 1437.800 2894.430 ;
        RECT 1457.440 2892.710 1457.580 2894.430 ;
        RECT 1457.380 2892.390 1457.640 2892.710 ;
        RECT 1501.540 2892.390 1501.800 2892.710 ;
        RECT 619.720 2891.370 619.980 2891.690 ;
        RECT 714.020 2891.370 714.280 2891.690 ;
        RECT 738.860 2891.370 739.120 2891.690 ;
        RECT 810.620 2891.370 810.880 2891.690 ;
        RECT 835.460 2891.370 835.720 2891.690 ;
        RECT 886.520 2891.370 886.780 2891.690 ;
        RECT 927.920 2891.370 928.180 2891.690 ;
        RECT 1293.620 2891.370 1293.880 2891.690 ;
        RECT 1318.460 2891.370 1318.720 2891.690 ;
        RECT 1437.600 2891.370 1437.860 2891.690 ;
        RECT 1501.600 2889.990 1501.740 2892.390 ;
        RECT 1501.540 2889.670 1501.800 2889.990 ;
        RECT 576.020 2593.870 576.280 2594.190 ;
        RECT 569.180 1991.370 569.320 2593.675 ;
        RECT 990.020 2035.930 990.280 2036.250 ;
        RECT 2056.300 2035.930 2056.560 2036.250 ;
        RECT 503.340 1991.050 503.600 1991.370 ;
        RECT 569.120 1991.050 569.380 1991.370 ;
        RECT 647.320 1991.050 647.580 1991.370 ;
        RECT 502.690 1981.250 502.970 1981.750 ;
        RECT 503.400 1981.250 503.540 1991.050 ;
        RECT 647.380 1987.290 647.520 1991.050 ;
        RECT 990.080 1987.290 990.220 2035.930 ;
        RECT 647.320 1986.970 647.580 1987.290 ;
        RECT 990.020 1986.970 990.280 1987.290 ;
        RECT 502.690 1981.110 503.540 1981.250 ;
        RECT 502.690 1977.750 502.970 1981.110 ;
        RECT 647.380 590.765 647.520 1986.970 ;
        RECT 2056.360 1917.095 2056.500 2035.930 ;
        RECT 2056.250 1913.095 2056.530 1917.095 ;
        RECT 759.790 600.000 760.070 604.000 ;
        RECT 759.850 598.810 759.990 600.000 ;
        RECT 759.620 598.670 759.990 598.810 ;
        RECT 647.310 590.395 647.590 590.765 ;
        RECT 666.170 590.395 666.450 590.765 ;
        RECT 666.240 588.725 666.380 590.395 ;
        RECT 759.620 588.725 759.760 598.670 ;
        RECT 666.170 588.355 666.450 588.725 ;
        RECT 759.550 588.355 759.830 588.725 ;
        RECT 759.620 20.050 759.760 588.355 ;
        RECT 174.900 19.730 175.160 20.050 ;
        RECT 759.560 19.730 759.820 20.050 ;
        RECT 174.960 2.400 175.100 19.730 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 1576.050 2896.320 1576.330 2896.600 ;
        RECT 1601.810 2896.320 1602.090 2896.600 ;
        RECT 579.690 2892.240 579.970 2892.520 ;
        RECT 619.710 2892.240 619.990 2892.520 ;
        RECT 547.950 2593.720 548.230 2594.000 ;
        RECT 569.110 2593.720 569.390 2594.000 ;
        RECT 572.330 2593.890 572.610 2594.170 ;
        RECT 647.310 590.440 647.590 590.720 ;
        RECT 666.170 590.440 666.450 590.720 ;
        RECT 666.170 588.400 666.450 588.680 ;
        RECT 759.550 588.400 759.830 588.680 ;
      LAYER met3 ;
        RECT 1576.025 2896.610 1576.355 2896.625 ;
        RECT 1575.350 2896.310 1576.355 2896.610 ;
        RECT 579.665 2892.530 579.995 2892.545 ;
        RECT 619.685 2892.530 620.015 2892.545 ;
        RECT 579.665 2892.230 620.015 2892.530 ;
        RECT 579.665 2892.215 579.995 2892.230 ;
        RECT 619.685 2892.215 620.015 2892.230 ;
        RECT 1575.350 2890.490 1575.650 2896.310 ;
        RECT 1576.025 2896.295 1576.355 2896.310 ;
        RECT 1601.785 2896.295 1602.115 2896.625 ;
        RECT 1601.800 2890.490 1602.100 2896.295 ;
        RECT 1575.350 2890.190 1602.100 2890.490 ;
        RECT 572.305 2594.180 572.635 2594.195 ;
        RECT 547.925 2594.010 548.255 2594.025 ;
        RECT 569.085 2594.010 569.415 2594.025 ;
        RECT 571.630 2594.010 572.635 2594.180 ;
        RECT 547.925 2593.880 572.635 2594.010 ;
        RECT 547.925 2593.710 571.930 2593.880 ;
        RECT 572.305 2593.865 572.635 2593.880 ;
        RECT 547.925 2593.695 548.255 2593.710 ;
        RECT 569.085 2593.695 569.415 2593.710 ;
        RECT 647.285 590.730 647.615 590.745 ;
        RECT 666.145 590.730 666.475 590.745 ;
        RECT 647.285 590.430 666.475 590.730 ;
        RECT 647.285 590.415 647.615 590.430 ;
        RECT 666.145 590.415 666.475 590.430 ;
        RECT 666.145 588.690 666.475 588.705 ;
        RECT 759.525 588.690 759.855 588.705 ;
        RECT 666.145 588.390 759.855 588.690 ;
        RECT 666.145 588.375 666.475 588.390 ;
        RECT 759.525 588.375 759.855 588.390 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.870 2916.420 428.190 2916.480 ;
        RECT 1726.450 2916.420 1726.770 2916.480 ;
        RECT 427.870 2916.280 1726.770 2916.420 ;
        RECT 427.870 2916.220 428.190 2916.280 ;
        RECT 1726.450 2916.220 1726.770 2916.280 ;
        RECT 357.950 2038.880 358.270 2038.940 ;
        RECT 427.870 2038.880 428.190 2038.940 ;
        RECT 2014.870 2038.880 2015.190 2038.940 ;
        RECT 357.950 2038.740 2015.190 2038.880 ;
        RECT 357.950 2038.680 358.270 2038.740 ;
        RECT 427.870 2038.680 428.190 2038.740 ;
        RECT 2014.870 2038.680 2015.190 2038.740 ;
        RECT 2014.870 1966.460 2015.190 1966.520 ;
        RECT 2019.470 1966.460 2019.790 1966.520 ;
        RECT 2014.870 1966.320 2019.790 1966.460 ;
        RECT 2014.870 1966.260 2015.190 1966.320 ;
        RECT 2019.470 1966.260 2019.790 1966.320 ;
        RECT 348.290 1952.860 348.610 1952.920 ;
        RECT 357.950 1952.860 358.270 1952.920 ;
        RECT 348.290 1952.720 358.270 1952.860 ;
        RECT 348.290 1952.660 348.610 1952.720 ;
        RECT 357.950 1952.660 358.270 1952.720 ;
        RECT 192.350 589.800 192.670 589.860 ;
        RECT 348.290 589.800 348.610 589.860 ;
        RECT 192.350 589.660 348.610 589.800 ;
        RECT 192.350 589.600 192.670 589.660 ;
        RECT 348.290 589.600 348.610 589.660 ;
      LAYER via ;
        RECT 427.900 2916.220 428.160 2916.480 ;
        RECT 1726.480 2916.220 1726.740 2916.480 ;
        RECT 357.980 2038.680 358.240 2038.940 ;
        RECT 427.900 2038.680 428.160 2038.940 ;
        RECT 2014.900 2038.680 2015.160 2038.940 ;
        RECT 2014.900 1966.260 2015.160 1966.520 ;
        RECT 2019.500 1966.260 2019.760 1966.520 ;
        RECT 348.320 1952.660 348.580 1952.920 ;
        RECT 357.980 1952.660 358.240 1952.920 ;
        RECT 192.380 589.600 192.640 589.860 ;
        RECT 348.320 589.600 348.580 589.860 ;
      LAYER met2 ;
        RECT 427.900 2916.190 428.160 2916.510 ;
        RECT 1726.480 2916.190 1726.740 2916.510 ;
        RECT 427.960 2688.905 428.100 2916.190 ;
        RECT 1726.540 2900.055 1726.680 2916.190 ;
        RECT 1726.410 2896.055 1726.690 2900.055 ;
        RECT 427.890 2688.535 428.170 2688.905 ;
        RECT 427.960 2038.970 428.100 2688.535 ;
        RECT 357.980 2038.650 358.240 2038.970 ;
        RECT 427.900 2038.650 428.160 2038.970 ;
        RECT 2014.900 2038.650 2015.160 2038.970 ;
        RECT 358.040 1963.005 358.180 2038.650 ;
        RECT 2014.960 1966.550 2015.100 2038.650 ;
        RECT 2014.900 1966.230 2015.160 1966.550 ;
        RECT 2019.500 1966.230 2019.760 1966.550 ;
        RECT 357.970 1962.635 358.250 1963.005 ;
        RECT 358.040 1952.950 358.180 1962.635 ;
        RECT 348.320 1952.630 348.580 1952.950 ;
        RECT 357.980 1952.630 358.240 1952.950 ;
        RECT 348.380 592.805 348.520 1952.630 ;
        RECT 2019.560 1916.650 2019.700 1966.230 ;
        RECT 2021.290 1916.650 2021.570 1917.095 ;
        RECT 2019.560 1916.510 2021.570 1916.650 ;
        RECT 2021.290 1913.095 2021.570 1916.510 ;
        RECT 768.990 600.170 769.270 604.000 ;
        RECT 767.440 600.030 769.270 600.170 ;
        RECT 767.440 592.805 767.580 600.030 ;
        RECT 768.990 600.000 769.270 600.030 ;
        RECT 348.310 592.435 348.590 592.805 ;
        RECT 767.370 592.435 767.650 592.805 ;
        RECT 348.380 589.890 348.520 592.435 ;
        RECT 192.380 589.570 192.640 589.890 ;
        RECT 348.320 589.570 348.580 589.890 ;
        RECT 192.440 3.130 192.580 589.570 ;
        RECT 192.440 2.990 193.040 3.130 ;
        RECT 192.900 2.400 193.040 2.990 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 427.890 2688.580 428.170 2688.860 ;
        RECT 357.970 1962.680 358.250 1962.960 ;
        RECT 348.310 592.480 348.590 592.760 ;
        RECT 767.370 592.480 767.650 592.760 ;
      LAYER met3 ;
        RECT 427.865 2688.870 428.195 2688.885 ;
        RECT 430.000 2688.870 434.000 2689.040 ;
        RECT 427.865 2688.570 434.000 2688.870 ;
        RECT 427.865 2688.555 428.195 2688.570 ;
        RECT 430.000 2688.440 434.000 2688.570 ;
        RECT 357.945 1962.970 358.275 1962.985 ;
        RECT 360.000 1962.970 364.000 1963.120 ;
        RECT 357.945 1962.670 364.000 1962.970 ;
        RECT 357.945 1962.655 358.275 1962.670 ;
        RECT 360.000 1962.520 364.000 1962.670 ;
        RECT 348.285 592.770 348.615 592.785 ;
        RECT 767.345 592.770 767.675 592.785 ;
        RECT 348.285 592.470 767.675 592.770 ;
        RECT 348.285 592.455 348.615 592.470 ;
        RECT 767.345 592.455 767.675 592.470 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 591.170 2670.260 591.490 2670.320 ;
        RECT 592.550 2670.260 592.870 2670.320 ;
        RECT 591.170 2670.120 592.870 2670.260 ;
        RECT 591.170 2670.060 591.490 2670.120 ;
        RECT 592.550 2670.060 592.870 2670.120 ;
        RECT 592.550 2622.660 592.870 2622.720 ;
        RECT 592.180 2622.520 592.870 2622.660 ;
        RECT 592.180 2622.040 592.320 2622.520 ;
        RECT 592.550 2622.460 592.870 2622.520 ;
        RECT 592.090 2621.780 592.410 2622.040 ;
        RECT 591.170 2560.100 591.490 2560.160 ;
        RECT 592.550 2560.100 592.870 2560.160 ;
        RECT 591.170 2559.960 592.870 2560.100 ;
        RECT 591.170 2559.900 591.490 2559.960 ;
        RECT 592.550 2559.900 592.870 2559.960 ;
        RECT 591.630 2511.820 591.950 2511.880 ;
        RECT 592.550 2511.820 592.870 2511.880 ;
        RECT 591.630 2511.680 592.870 2511.820 ;
        RECT 591.630 2511.620 591.950 2511.680 ;
        RECT 592.550 2511.620 592.870 2511.680 ;
        RECT 592.090 2463.200 592.410 2463.260 ;
        RECT 592.550 2463.200 592.870 2463.260 ;
        RECT 592.090 2463.060 592.870 2463.200 ;
        RECT 592.090 2463.000 592.410 2463.060 ;
        RECT 592.550 2463.000 592.870 2463.060 ;
        RECT 592.090 2429.200 592.410 2429.260 ;
        RECT 592.090 2429.060 592.780 2429.200 ;
        RECT 592.090 2429.000 592.410 2429.060 ;
        RECT 592.640 2428.920 592.780 2429.060 ;
        RECT 592.550 2428.660 592.870 2428.920 ;
        RECT 592.090 2332.640 592.410 2332.700 ;
        RECT 591.720 2332.500 592.410 2332.640 ;
        RECT 591.720 2332.020 591.860 2332.500 ;
        RECT 592.090 2332.440 592.410 2332.500 ;
        RECT 591.630 2331.760 591.950 2332.020 ;
        RECT 590.250 2318.360 590.570 2318.420 ;
        RECT 591.630 2318.360 591.950 2318.420 ;
        RECT 590.250 2318.220 591.950 2318.360 ;
        RECT 590.250 2318.160 590.570 2318.220 ;
        RECT 591.630 2318.160 591.950 2318.220 ;
        RECT 591.170 2235.540 591.490 2235.800 ;
        RECT 591.260 2235.400 591.400 2235.540 ;
        RECT 591.630 2235.400 591.950 2235.460 ;
        RECT 591.260 2235.260 591.950 2235.400 ;
        RECT 591.630 2235.200 591.950 2235.260 ;
        RECT 590.250 2221.800 590.570 2221.860 ;
        RECT 591.630 2221.800 591.950 2221.860 ;
        RECT 590.250 2221.660 591.950 2221.800 ;
        RECT 590.250 2221.600 590.570 2221.660 ;
        RECT 591.630 2221.600 591.950 2221.660 ;
        RECT 591.170 2138.980 591.490 2139.240 ;
        RECT 591.260 2138.840 591.400 2138.980 ;
        RECT 591.630 2138.840 591.950 2138.900 ;
        RECT 591.260 2138.700 591.950 2138.840 ;
        RECT 591.630 2138.640 591.950 2138.700 ;
        RECT 591.170 2076.960 591.490 2077.020 ;
        RECT 592.090 2076.960 592.410 2077.020 ;
        RECT 591.170 2076.820 592.410 2076.960 ;
        RECT 591.170 2076.760 591.490 2076.820 ;
        RECT 592.090 2076.760 592.410 2076.820 ;
        RECT 651.890 2035.820 652.210 2035.880 ;
        RECT 2084.330 2035.820 2084.650 2035.880 ;
        RECT 651.890 2035.680 2084.650 2035.820 ;
        RECT 651.890 2035.620 652.210 2035.680 ;
        RECT 2084.330 2035.620 2084.650 2035.680 ;
        RECT 591.170 2028.680 591.490 2028.740 ;
        RECT 592.550 2028.680 592.870 2028.740 ;
        RECT 591.170 2028.540 592.870 2028.680 ;
        RECT 591.170 2028.480 591.490 2028.540 ;
        RECT 592.550 2028.480 592.870 2028.540 ;
        RECT 586.570 1994.000 586.890 1994.060 ;
        RECT 593.010 1994.000 593.330 1994.060 ;
        RECT 648.670 1994.000 648.990 1994.060 ;
        RECT 586.570 1993.860 648.990 1994.000 ;
        RECT 586.570 1993.800 586.890 1993.860 ;
        RECT 593.010 1993.800 593.330 1993.860 ;
        RECT 648.670 1993.800 648.990 1993.860 ;
        RECT 648.670 1991.620 648.990 1991.680 ;
        RECT 651.890 1991.620 652.210 1991.680 ;
        RECT 648.670 1991.480 652.210 1991.620 ;
        RECT 648.670 1991.420 648.990 1991.480 ;
        RECT 651.890 1991.420 652.210 1991.480 ;
        RECT 429.710 1990.940 430.030 1991.000 ;
        RECT 586.570 1990.940 586.890 1991.000 ;
        RECT 429.710 1990.800 586.890 1990.940 ;
        RECT 429.710 1990.740 430.030 1990.800 ;
        RECT 586.570 1990.740 586.890 1990.800 ;
        RECT 213.510 593.200 213.830 593.260 ;
        RECT 648.670 593.200 648.990 593.260 ;
        RECT 776.550 593.200 776.870 593.260 ;
        RECT 213.510 593.060 776.870 593.200 ;
        RECT 213.510 593.000 213.830 593.060 ;
        RECT 648.670 593.000 648.990 593.060 ;
        RECT 776.550 593.000 776.870 593.060 ;
        RECT 210.750 16.560 211.070 16.620 ;
        RECT 213.510 16.560 213.830 16.620 ;
        RECT 210.750 16.420 213.830 16.560 ;
        RECT 210.750 16.360 211.070 16.420 ;
        RECT 213.510 16.360 213.830 16.420 ;
      LAYER via ;
        RECT 591.200 2670.060 591.460 2670.320 ;
        RECT 592.580 2670.060 592.840 2670.320 ;
        RECT 592.580 2622.460 592.840 2622.720 ;
        RECT 592.120 2621.780 592.380 2622.040 ;
        RECT 591.200 2559.900 591.460 2560.160 ;
        RECT 592.580 2559.900 592.840 2560.160 ;
        RECT 591.660 2511.620 591.920 2511.880 ;
        RECT 592.580 2511.620 592.840 2511.880 ;
        RECT 592.120 2463.000 592.380 2463.260 ;
        RECT 592.580 2463.000 592.840 2463.260 ;
        RECT 592.120 2429.000 592.380 2429.260 ;
        RECT 592.580 2428.660 592.840 2428.920 ;
        RECT 592.120 2332.440 592.380 2332.700 ;
        RECT 591.660 2331.760 591.920 2332.020 ;
        RECT 590.280 2318.160 590.540 2318.420 ;
        RECT 591.660 2318.160 591.920 2318.420 ;
        RECT 591.200 2235.540 591.460 2235.800 ;
        RECT 591.660 2235.200 591.920 2235.460 ;
        RECT 590.280 2221.600 590.540 2221.860 ;
        RECT 591.660 2221.600 591.920 2221.860 ;
        RECT 591.200 2138.980 591.460 2139.240 ;
        RECT 591.660 2138.640 591.920 2138.900 ;
        RECT 591.200 2076.760 591.460 2077.020 ;
        RECT 592.120 2076.760 592.380 2077.020 ;
        RECT 651.920 2035.620 652.180 2035.880 ;
        RECT 2084.360 2035.620 2084.620 2035.880 ;
        RECT 591.200 2028.480 591.460 2028.740 ;
        RECT 592.580 2028.480 592.840 2028.740 ;
        RECT 586.600 1993.800 586.860 1994.060 ;
        RECT 593.040 1993.800 593.300 1994.060 ;
        RECT 648.700 1993.800 648.960 1994.060 ;
        RECT 648.700 1991.420 648.960 1991.680 ;
        RECT 651.920 1991.420 652.180 1991.680 ;
        RECT 429.740 1990.740 430.000 1991.000 ;
        RECT 586.600 1990.740 586.860 1991.000 ;
        RECT 213.540 593.000 213.800 593.260 ;
        RECT 648.700 593.000 648.960 593.260 ;
        RECT 776.580 593.000 776.840 593.260 ;
        RECT 210.780 16.360 211.040 16.620 ;
        RECT 213.540 16.360 213.800 16.620 ;
      LAYER met2 ;
        RECT 591.190 2711.995 591.470 2712.365 ;
        RECT 591.260 2670.350 591.400 2711.995 ;
        RECT 591.200 2670.030 591.460 2670.350 ;
        RECT 592.580 2670.030 592.840 2670.350 ;
        RECT 592.640 2622.750 592.780 2670.030 ;
        RECT 592.580 2622.430 592.840 2622.750 ;
        RECT 592.120 2621.750 592.380 2622.070 ;
        RECT 592.180 2608.325 592.320 2621.750 ;
        RECT 591.190 2607.955 591.470 2608.325 ;
        RECT 592.110 2607.955 592.390 2608.325 ;
        RECT 591.260 2560.190 591.400 2607.955 ;
        RECT 591.200 2559.870 591.460 2560.190 ;
        RECT 592.580 2559.870 592.840 2560.190 ;
        RECT 592.640 2511.910 592.780 2559.870 ;
        RECT 591.660 2511.650 591.920 2511.910 ;
        RECT 591.660 2511.590 592.320 2511.650 ;
        RECT 592.580 2511.590 592.840 2511.910 ;
        RECT 591.720 2511.510 592.320 2511.590 ;
        RECT 592.180 2490.685 592.320 2511.510 ;
        RECT 1598.530 2500.000 1598.810 2504.000 ;
        RECT 1598.660 2490.685 1598.800 2500.000 ;
        RECT 592.110 2490.315 592.390 2490.685 ;
        RECT 1598.590 2490.315 1598.870 2490.685 ;
        RECT 592.180 2463.370 592.320 2490.315 ;
        RECT 592.180 2463.290 592.780 2463.370 ;
        RECT 592.120 2463.230 592.840 2463.290 ;
        RECT 592.120 2462.970 592.380 2463.230 ;
        RECT 592.580 2462.970 592.840 2463.230 ;
        RECT 592.180 2429.290 592.320 2462.970 ;
        RECT 592.120 2428.970 592.380 2429.290 ;
        RECT 592.580 2428.630 592.840 2428.950 ;
        RECT 592.640 2415.090 592.780 2428.630 ;
        RECT 592.640 2414.950 593.240 2415.090 ;
        RECT 593.100 2380.410 593.240 2414.950 ;
        RECT 592.180 2380.270 593.240 2380.410 ;
        RECT 592.180 2332.730 592.320 2380.270 ;
        RECT 592.120 2332.410 592.380 2332.730 ;
        RECT 591.660 2331.730 591.920 2332.050 ;
        RECT 591.720 2318.450 591.860 2331.730 ;
        RECT 590.280 2318.130 590.540 2318.450 ;
        RECT 591.660 2318.130 591.920 2318.450 ;
        RECT 590.340 2270.365 590.480 2318.130 ;
        RECT 590.270 2269.995 590.550 2270.365 ;
        RECT 591.190 2269.995 591.470 2270.365 ;
        RECT 591.260 2235.830 591.400 2269.995 ;
        RECT 591.200 2235.510 591.460 2235.830 ;
        RECT 591.660 2235.170 591.920 2235.490 ;
        RECT 591.720 2221.890 591.860 2235.170 ;
        RECT 590.280 2221.570 590.540 2221.890 ;
        RECT 591.660 2221.570 591.920 2221.890 ;
        RECT 590.340 2173.805 590.480 2221.570 ;
        RECT 590.270 2173.435 590.550 2173.805 ;
        RECT 591.190 2173.435 591.470 2173.805 ;
        RECT 591.260 2139.270 591.400 2173.435 ;
        RECT 591.200 2138.950 591.460 2139.270 ;
        RECT 591.660 2138.610 591.920 2138.930 ;
        RECT 591.720 2090.730 591.860 2138.610 ;
        RECT 591.720 2090.590 592.320 2090.730 ;
        RECT 592.180 2077.050 592.320 2090.590 ;
        RECT 591.200 2076.730 591.460 2077.050 ;
        RECT 592.120 2076.730 592.380 2077.050 ;
        RECT 591.260 2028.770 591.400 2076.730 ;
        RECT 651.920 2035.590 652.180 2035.910 ;
        RECT 2084.360 2035.590 2084.620 2035.910 ;
        RECT 591.200 2028.450 591.460 2028.770 ;
        RECT 592.580 2028.450 592.840 2028.770 ;
        RECT 592.640 1994.170 592.780 2028.450 ;
        RECT 592.640 1994.090 593.240 1994.170 ;
        RECT 586.600 1993.770 586.860 1994.090 ;
        RECT 592.640 1994.030 593.300 1994.090 ;
        RECT 593.040 1993.770 593.300 1994.030 ;
        RECT 648.700 1993.770 648.960 1994.090 ;
        RECT 586.660 1991.030 586.800 1993.770 ;
        RECT 593.100 1993.615 593.240 1993.770 ;
        RECT 648.760 1991.710 648.900 1993.770 ;
        RECT 651.980 1991.710 652.120 2035.590 ;
        RECT 648.700 1991.390 648.960 1991.710 ;
        RECT 651.920 1991.390 652.180 1991.710 ;
        RECT 429.740 1990.710 430.000 1991.030 ;
        RECT 586.600 1990.710 586.860 1991.030 ;
        RECT 428.170 1981.250 428.450 1981.750 ;
        RECT 429.800 1981.250 429.940 1990.710 ;
        RECT 428.170 1981.110 429.940 1981.250 ;
        RECT 428.170 1977.750 428.450 1981.110 ;
        RECT 648.760 593.290 648.900 1991.390 ;
        RECT 2084.420 1904.525 2084.560 2035.590 ;
        RECT 2084.350 1904.155 2084.630 1904.525 ;
        RECT 778.190 600.170 778.470 604.000 ;
        RECT 776.640 600.030 778.470 600.170 ;
        RECT 776.640 593.290 776.780 600.030 ;
        RECT 778.190 600.000 778.470 600.030 ;
        RECT 213.540 592.970 213.800 593.290 ;
        RECT 648.700 592.970 648.960 593.290 ;
        RECT 776.580 592.970 776.840 593.290 ;
        RECT 213.600 16.650 213.740 592.970 ;
        RECT 210.780 16.330 211.040 16.650 ;
        RECT 213.540 16.330 213.800 16.650 ;
        RECT 210.840 2.400 210.980 16.330 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 591.190 2712.040 591.470 2712.320 ;
        RECT 591.190 2608.000 591.470 2608.280 ;
        RECT 592.110 2608.000 592.390 2608.280 ;
        RECT 592.110 2490.360 592.390 2490.640 ;
        RECT 1598.590 2490.360 1598.870 2490.640 ;
        RECT 590.270 2270.040 590.550 2270.320 ;
        RECT 591.190 2270.040 591.470 2270.320 ;
        RECT 590.270 2173.480 590.550 2173.760 ;
        RECT 591.190 2173.480 591.470 2173.760 ;
        RECT 2084.350 1904.200 2084.630 1904.480 ;
      LAYER met3 ;
        RECT 591.165 2712.330 591.495 2712.345 ;
        RECT 578.070 2712.160 591.495 2712.330 ;
        RECT 574.800 2712.030 591.495 2712.160 ;
        RECT 574.800 2711.560 578.800 2712.030 ;
        RECT 591.165 2712.015 591.495 2712.030 ;
        RECT 591.165 2608.290 591.495 2608.305 ;
        RECT 592.085 2608.290 592.415 2608.305 ;
        RECT 591.165 2607.990 592.415 2608.290 ;
        RECT 591.165 2607.975 591.495 2607.990 ;
        RECT 592.085 2607.975 592.415 2607.990 ;
        RECT 592.085 2490.650 592.415 2490.665 ;
        RECT 1598.565 2490.650 1598.895 2490.665 ;
        RECT 592.085 2490.350 1598.895 2490.650 ;
        RECT 592.085 2490.335 592.415 2490.350 ;
        RECT 1598.565 2490.335 1598.895 2490.350 ;
        RECT 590.245 2270.330 590.575 2270.345 ;
        RECT 591.165 2270.330 591.495 2270.345 ;
        RECT 590.245 2270.030 591.495 2270.330 ;
        RECT 590.245 2270.015 590.575 2270.030 ;
        RECT 591.165 2270.015 591.495 2270.030 ;
        RECT 590.245 2173.770 590.575 2173.785 ;
        RECT 591.165 2173.770 591.495 2173.785 ;
        RECT 590.245 2173.470 591.495 2173.770 ;
        RECT 590.245 2173.455 590.575 2173.470 ;
        RECT 591.165 2173.455 591.495 2173.470 ;
        RECT 2084.325 1904.490 2084.655 1904.505 ;
        RECT 2075.830 1904.320 2084.655 1904.490 ;
        RECT 2072.375 1904.190 2084.655 1904.320 ;
        RECT 2072.375 1903.720 2076.375 1904.190 ;
        RECT 2084.325 1904.175 2084.655 1904.190 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 489.970 2592.060 490.290 2592.120 ;
        RECT 720.890 2592.060 721.210 2592.120 ;
        RECT 489.970 2591.920 721.210 2592.060 ;
        RECT 489.970 2591.860 490.290 2591.920 ;
        RECT 720.890 2591.860 721.210 2591.920 ;
        RECT 720.890 2489.380 721.210 2489.440 ;
        RECT 1672.170 2489.380 1672.490 2489.440 ;
        RECT 720.890 2489.240 1672.490 2489.380 ;
        RECT 720.890 2489.180 721.210 2489.240 ;
        RECT 1672.170 2489.180 1672.490 2489.240 ;
        RECT 627.970 1987.540 628.290 1987.600 ;
        RECT 720.890 1987.540 721.210 1987.600 ;
        RECT 627.970 1987.400 721.210 1987.540 ;
        RECT 627.970 1987.340 628.290 1987.400 ;
        RECT 720.890 1987.340 721.210 1987.400 ;
        RECT 720.890 1786.940 721.210 1787.000 ;
        RECT 727.790 1786.940 728.110 1787.000 ;
        RECT 720.890 1786.800 728.110 1786.940 ;
        RECT 720.890 1786.740 721.210 1786.800 ;
        RECT 727.790 1786.740 728.110 1786.800 ;
        RECT 727.790 1702.620 728.110 1702.680 ;
        RECT 1909.070 1702.620 1909.390 1702.680 ;
        RECT 727.790 1702.480 1909.390 1702.620 ;
        RECT 727.790 1702.420 728.110 1702.480 ;
        RECT 1909.070 1702.420 1909.390 1702.480 ;
        RECT 652.810 1006.300 653.130 1006.360 ;
        RECT 727.790 1006.300 728.110 1006.360 ;
        RECT 652.810 1006.160 728.110 1006.300 ;
        RECT 652.810 1006.100 653.130 1006.160 ;
        RECT 727.790 1006.100 728.110 1006.160 ;
        RECT 718.590 587.760 718.910 587.820 ;
        RECT 786.670 587.760 786.990 587.820 ;
        RECT 715.460 587.620 786.990 587.760 ;
        RECT 652.810 587.420 653.130 587.480 ;
        RECT 715.460 587.420 715.600 587.620 ;
        RECT 718.590 587.560 718.910 587.620 ;
        RECT 786.670 587.560 786.990 587.620 ;
        RECT 652.810 587.280 715.600 587.420 ;
        RECT 652.810 587.220 653.130 587.280 ;
        RECT 228.690 16.560 229.010 16.620 ;
        RECT 718.590 16.560 718.910 16.620 ;
        RECT 228.690 16.420 718.910 16.560 ;
        RECT 228.690 16.360 229.010 16.420 ;
        RECT 718.590 16.360 718.910 16.420 ;
      LAYER via ;
        RECT 490.000 2591.860 490.260 2592.120 ;
        RECT 720.920 2591.860 721.180 2592.120 ;
        RECT 720.920 2489.180 721.180 2489.440 ;
        RECT 1672.200 2489.180 1672.460 2489.440 ;
        RECT 628.000 1987.340 628.260 1987.600 ;
        RECT 720.920 1987.340 721.180 1987.600 ;
        RECT 720.920 1786.740 721.180 1787.000 ;
        RECT 727.820 1786.740 728.080 1787.000 ;
        RECT 727.820 1702.420 728.080 1702.680 ;
        RECT 1909.100 1702.420 1909.360 1702.680 ;
        RECT 652.840 1006.100 653.100 1006.360 ;
        RECT 727.820 1006.100 728.080 1006.360 ;
        RECT 652.840 587.220 653.100 587.480 ;
        RECT 718.620 587.560 718.880 587.820 ;
        RECT 786.700 587.560 786.960 587.820 ;
        RECT 228.720 16.360 228.980 16.620 ;
        RECT 718.620 16.360 718.880 16.620 ;
      LAYER met2 ;
        RECT 489.890 2600.660 490.170 2604.000 ;
        RECT 489.890 2600.000 490.200 2600.660 ;
        RECT 490.060 2592.150 490.200 2600.000 ;
        RECT 490.000 2591.830 490.260 2592.150 ;
        RECT 720.920 2591.830 721.180 2592.150 ;
        RECT 720.980 2489.470 721.120 2591.830 ;
        RECT 1672.130 2500.000 1672.410 2504.000 ;
        RECT 1672.260 2489.470 1672.400 2500.000 ;
        RECT 720.920 2489.150 721.180 2489.470 ;
        RECT 1672.200 2489.150 1672.460 2489.470 ;
        RECT 720.980 1987.630 721.120 2489.150 ;
        RECT 628.000 1987.310 628.260 1987.630 ;
        RECT 720.920 1987.310 721.180 1987.630 ;
        RECT 628.060 1981.750 628.200 1987.310 ;
        RECT 627.810 1981.110 628.200 1981.750 ;
        RECT 627.810 1977.750 628.090 1981.110 ;
        RECT 720.980 1787.030 721.120 1987.310 ;
        RECT 720.920 1786.710 721.180 1787.030 ;
        RECT 727.820 1786.710 728.080 1787.030 ;
        RECT 727.880 1702.710 728.020 1786.710 ;
        RECT 1909.090 1783.795 1909.370 1784.165 ;
        RECT 1909.160 1702.710 1909.300 1783.795 ;
        RECT 727.820 1702.390 728.080 1702.710 ;
        RECT 1909.100 1702.390 1909.360 1702.710 ;
        RECT 727.880 1006.390 728.020 1702.390 ;
        RECT 652.840 1006.070 653.100 1006.390 ;
        RECT 727.820 1006.070 728.080 1006.390 ;
        RECT 652.900 587.510 653.040 1006.070 ;
        RECT 787.390 600.170 787.670 604.000 ;
        RECT 786.760 600.030 787.670 600.170 ;
        RECT 786.760 587.850 786.900 600.030 ;
        RECT 787.390 600.000 787.670 600.030 ;
        RECT 718.620 587.530 718.880 587.850 ;
        RECT 786.700 587.530 786.960 587.850 ;
        RECT 652.840 587.190 653.100 587.510 ;
        RECT 718.680 16.650 718.820 587.530 ;
        RECT 228.720 16.330 228.980 16.650 ;
        RECT 718.620 16.330 718.880 16.650 ;
        RECT 228.780 2.400 228.920 16.330 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 1909.090 1783.840 1909.370 1784.120 ;
      LAYER met3 ;
        RECT 1920.000 1786.760 1924.000 1787.360 ;
        RECT 1909.065 1784.130 1909.395 1784.145 ;
        RECT 1920.350 1784.130 1920.650 1786.760 ;
        RECT 1909.065 1783.830 1920.650 1784.130 ;
        RECT 1909.065 1783.815 1909.395 1783.830 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 691.450 596.600 691.770 596.660 ;
        RECT 694.210 596.600 694.530 596.660 ;
        RECT 691.450 596.460 694.530 596.600 ;
        RECT 691.450 596.400 691.770 596.460 ;
        RECT 694.210 596.400 694.530 596.460 ;
        RECT 689.610 483.040 689.930 483.100 ;
        RECT 690.070 483.040 690.390 483.100 ;
        RECT 689.610 482.900 690.390 483.040 ;
        RECT 689.610 482.840 689.930 482.900 ;
        RECT 690.070 482.840 690.390 482.900 ;
        RECT 689.610 448.360 689.930 448.420 ;
        RECT 690.530 448.360 690.850 448.420 ;
        RECT 689.610 448.220 690.850 448.360 ;
        RECT 689.610 448.160 689.930 448.220 ;
        RECT 690.530 448.160 690.850 448.220 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 690.070 17.580 690.390 17.640 ;
        RECT 50.210 17.440 690.390 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 690.070 17.380 690.390 17.440 ;
      LAYER via ;
        RECT 691.480 596.400 691.740 596.660 ;
        RECT 694.240 596.400 694.500 596.660 ;
        RECT 689.640 482.840 689.900 483.100 ;
        RECT 690.100 482.840 690.360 483.100 ;
        RECT 689.640 448.160 689.900 448.420 ;
        RECT 690.560 448.160 690.820 448.420 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 690.100 17.380 690.360 17.640 ;
      LAYER met2 ;
        RECT 695.850 600.170 696.130 604.000 ;
        RECT 694.300 600.030 696.130 600.170 ;
        RECT 694.300 596.690 694.440 600.030 ;
        RECT 695.850 600.000 696.130 600.030 ;
        RECT 691.480 596.370 691.740 596.690 ;
        RECT 694.240 596.370 694.500 596.690 ;
        RECT 691.540 569.570 691.680 596.370 ;
        RECT 690.620 569.430 691.680 569.570 ;
        RECT 690.620 497.490 690.760 569.430 ;
        RECT 690.160 497.350 690.760 497.490 ;
        RECT 690.160 483.130 690.300 497.350 ;
        RECT 689.640 482.810 689.900 483.130 ;
        RECT 690.100 482.810 690.360 483.130 ;
        RECT 689.700 448.450 689.840 482.810 ;
        RECT 689.640 448.130 689.900 448.450 ;
        RECT 690.560 448.130 690.820 448.450 ;
        RECT 690.620 434.930 690.760 448.130 ;
        RECT 690.620 434.790 691.220 434.930 ;
        RECT 691.080 62.290 691.220 434.790 ;
        RECT 690.160 62.150 691.220 62.290 ;
        RECT 690.160 17.670 690.300 62.150 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 690.100 17.350 690.360 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 252.610 16.900 252.930 16.960 ;
        RECT 794.490 16.900 794.810 16.960 ;
        RECT 252.610 16.760 794.810 16.900 ;
        RECT 252.610 16.700 252.930 16.760 ;
        RECT 794.490 16.700 794.810 16.760 ;
      LAYER via ;
        RECT 252.640 16.700 252.900 16.960 ;
        RECT 794.520 16.700 794.780 16.960 ;
      LAYER met2 ;
        RECT 799.810 600.850 800.090 604.000 ;
        RECT 797.340 600.710 800.090 600.850 ;
        RECT 797.340 596.770 797.480 600.710 ;
        RECT 799.810 600.000 800.090 600.710 ;
        RECT 795.500 596.630 797.480 596.770 ;
        RECT 795.500 569.400 795.640 596.630 ;
        RECT 794.580 569.260 795.640 569.400 ;
        RECT 794.580 16.990 794.720 569.260 ;
        RECT 252.640 16.670 252.900 16.990 ;
        RECT 794.520 16.670 794.780 16.990 ;
        RECT 252.700 2.400 252.840 16.670 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 807.370 483.180 807.690 483.440 ;
        RECT 807.460 482.760 807.600 483.180 ;
        RECT 807.370 482.500 807.690 482.760 ;
        RECT 270.090 31.180 270.410 31.240 ;
        RECT 807.370 31.180 807.690 31.240 ;
        RECT 270.090 31.040 807.690 31.180 ;
        RECT 270.090 30.980 270.410 31.040 ;
        RECT 807.370 30.980 807.690 31.040 ;
      LAYER via ;
        RECT 807.400 483.180 807.660 483.440 ;
        RECT 807.400 482.500 807.660 482.760 ;
        RECT 270.120 30.980 270.380 31.240 ;
        RECT 807.400 30.980 807.660 31.240 ;
      LAYER met2 ;
        RECT 809.010 600.170 809.290 604.000 ;
        RECT 807.460 600.030 809.290 600.170 ;
        RECT 807.460 483.470 807.600 600.030 ;
        RECT 809.010 600.000 809.290 600.030 ;
        RECT 807.400 483.150 807.660 483.470 ;
        RECT 807.400 482.470 807.660 482.790 ;
        RECT 807.460 31.270 807.600 482.470 ;
        RECT 270.120 30.950 270.380 31.270 ;
        RECT 807.400 30.950 807.660 31.270 ;
        RECT 270.180 2.400 270.320 30.950 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 814.730 524.180 815.050 524.240 ;
        RECT 815.650 524.180 815.970 524.240 ;
        RECT 814.730 524.040 815.970 524.180 ;
        RECT 814.730 523.980 815.050 524.040 ;
        RECT 815.650 523.980 815.970 524.040 ;
        RECT 814.730 476.240 815.050 476.300 ;
        RECT 815.650 476.240 815.970 476.300 ;
        RECT 814.730 476.100 815.970 476.240 ;
        RECT 814.730 476.040 815.050 476.100 ;
        RECT 815.650 476.040 815.970 476.100 ;
        RECT 814.730 427.620 815.050 427.680 ;
        RECT 815.650 427.620 815.970 427.680 ;
        RECT 814.730 427.480 815.970 427.620 ;
        RECT 814.730 427.420 815.050 427.480 ;
        RECT 815.650 427.420 815.970 427.480 ;
        RECT 814.730 379.680 815.050 379.740 ;
        RECT 815.650 379.680 815.970 379.740 ;
        RECT 814.730 379.540 815.970 379.680 ;
        RECT 814.730 379.480 815.050 379.540 ;
        RECT 815.650 379.480 815.970 379.540 ;
        RECT 814.730 331.060 815.050 331.120 ;
        RECT 815.650 331.060 815.970 331.120 ;
        RECT 814.730 330.920 815.970 331.060 ;
        RECT 814.730 330.860 815.050 330.920 ;
        RECT 815.650 330.860 815.970 330.920 ;
        RECT 814.730 283.120 815.050 283.180 ;
        RECT 815.650 283.120 815.970 283.180 ;
        RECT 814.730 282.980 815.970 283.120 ;
        RECT 814.730 282.920 815.050 282.980 ;
        RECT 815.650 282.920 815.970 282.980 ;
        RECT 814.730 234.500 815.050 234.560 ;
        RECT 815.650 234.500 815.970 234.560 ;
        RECT 814.730 234.360 815.970 234.500 ;
        RECT 814.730 234.300 815.050 234.360 ;
        RECT 815.650 234.300 815.970 234.360 ;
        RECT 814.730 137.940 815.050 138.000 ;
        RECT 815.650 137.940 815.970 138.000 ;
        RECT 814.730 137.800 815.970 137.940 ;
        RECT 814.730 137.740 815.050 137.800 ;
        RECT 815.650 137.740 815.970 137.800 ;
        RECT 814.730 90.000 815.050 90.060 ;
        RECT 815.650 90.000 815.970 90.060 ;
        RECT 814.730 89.860 815.970 90.000 ;
        RECT 814.730 89.800 815.050 89.860 ;
        RECT 815.650 89.800 815.970 89.860 ;
        RECT 814.730 62.460 815.050 62.520 ;
        RECT 814.360 62.320 815.050 62.460 ;
        RECT 814.360 62.180 814.500 62.320 ;
        RECT 814.730 62.260 815.050 62.320 ;
        RECT 814.270 61.920 814.590 62.180 ;
        RECT 288.030 48.180 288.350 48.240 ;
        RECT 814.270 48.180 814.590 48.240 ;
        RECT 288.030 48.040 814.590 48.180 ;
        RECT 288.030 47.980 288.350 48.040 ;
        RECT 814.270 47.980 814.590 48.040 ;
      LAYER via ;
        RECT 814.760 523.980 815.020 524.240 ;
        RECT 815.680 523.980 815.940 524.240 ;
        RECT 814.760 476.040 815.020 476.300 ;
        RECT 815.680 476.040 815.940 476.300 ;
        RECT 814.760 427.420 815.020 427.680 ;
        RECT 815.680 427.420 815.940 427.680 ;
        RECT 814.760 379.480 815.020 379.740 ;
        RECT 815.680 379.480 815.940 379.740 ;
        RECT 814.760 330.860 815.020 331.120 ;
        RECT 815.680 330.860 815.940 331.120 ;
        RECT 814.760 282.920 815.020 283.180 ;
        RECT 815.680 282.920 815.940 283.180 ;
        RECT 814.760 234.300 815.020 234.560 ;
        RECT 815.680 234.300 815.940 234.560 ;
        RECT 814.760 137.740 815.020 138.000 ;
        RECT 815.680 137.740 815.940 138.000 ;
        RECT 814.760 89.800 815.020 90.060 ;
        RECT 815.680 89.800 815.940 90.060 ;
        RECT 814.760 62.260 815.020 62.520 ;
        RECT 814.300 61.920 814.560 62.180 ;
        RECT 288.060 47.980 288.320 48.240 ;
        RECT 814.300 47.980 814.560 48.240 ;
      LAYER met2 ;
        RECT 818.210 600.170 818.490 604.000 ;
        RECT 816.660 600.030 818.490 600.170 ;
        RECT 816.660 596.770 816.800 600.030 ;
        RECT 818.210 600.000 818.490 600.030 ;
        RECT 814.820 596.630 816.800 596.770 ;
        RECT 814.820 524.270 814.960 596.630 ;
        RECT 814.760 523.950 815.020 524.270 ;
        RECT 815.680 523.950 815.940 524.270 ;
        RECT 815.740 476.330 815.880 523.950 ;
        RECT 814.760 476.010 815.020 476.330 ;
        RECT 815.680 476.010 815.940 476.330 ;
        RECT 814.820 427.710 814.960 476.010 ;
        RECT 814.760 427.390 815.020 427.710 ;
        RECT 815.680 427.390 815.940 427.710 ;
        RECT 815.740 379.770 815.880 427.390 ;
        RECT 814.760 379.450 815.020 379.770 ;
        RECT 815.680 379.450 815.940 379.770 ;
        RECT 814.820 331.150 814.960 379.450 ;
        RECT 814.760 330.830 815.020 331.150 ;
        RECT 815.680 330.830 815.940 331.150 ;
        RECT 815.740 283.210 815.880 330.830 ;
        RECT 814.760 282.890 815.020 283.210 ;
        RECT 815.680 282.890 815.940 283.210 ;
        RECT 814.820 234.590 814.960 282.890 ;
        RECT 814.760 234.270 815.020 234.590 ;
        RECT 815.680 234.270 815.940 234.590 ;
        RECT 815.740 145.365 815.880 234.270 ;
        RECT 814.750 144.995 815.030 145.365 ;
        RECT 815.670 144.995 815.950 145.365 ;
        RECT 814.820 138.030 814.960 144.995 ;
        RECT 814.760 137.710 815.020 138.030 ;
        RECT 815.680 137.710 815.940 138.030 ;
        RECT 815.740 90.090 815.880 137.710 ;
        RECT 814.760 89.770 815.020 90.090 ;
        RECT 815.680 89.770 815.940 90.090 ;
        RECT 814.820 62.550 814.960 89.770 ;
        RECT 814.760 62.230 815.020 62.550 ;
        RECT 814.300 61.890 814.560 62.210 ;
        RECT 814.360 48.270 814.500 61.890 ;
        RECT 288.060 47.950 288.320 48.270 ;
        RECT 814.300 47.950 814.560 48.270 ;
        RECT 288.120 2.400 288.260 47.950 ;
        RECT 287.910 -4.800 288.470 2.400 ;
      LAYER via2 ;
        RECT 814.750 145.040 815.030 145.320 ;
        RECT 815.670 145.040 815.950 145.320 ;
      LAYER met3 ;
        RECT 814.725 145.330 815.055 145.345 ;
        RECT 815.645 145.330 815.975 145.345 ;
        RECT 814.725 145.030 815.975 145.330 ;
        RECT 814.725 145.015 815.055 145.030 ;
        RECT 815.645 145.015 815.975 145.030 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 31.520 306.290 31.580 ;
        RECT 822.090 31.520 822.410 31.580 ;
        RECT 305.970 31.380 822.410 31.520 ;
        RECT 305.970 31.320 306.290 31.380 ;
        RECT 822.090 31.320 822.410 31.380 ;
      LAYER via ;
        RECT 306.000 31.320 306.260 31.580 ;
        RECT 822.120 31.320 822.380 31.580 ;
      LAYER met2 ;
        RECT 827.410 600.850 827.690 604.000 ;
        RECT 824.940 600.710 827.690 600.850 ;
        RECT 824.940 596.770 825.080 600.710 ;
        RECT 827.410 600.000 827.690 600.710 ;
        RECT 823.100 596.630 825.080 596.770 ;
        RECT 823.100 569.400 823.240 596.630 ;
        RECT 822.180 569.260 823.240 569.400 ;
        RECT 822.180 31.610 822.320 569.260 ;
        RECT 306.000 31.290 306.260 31.610 ;
        RECT 822.120 31.290 822.380 31.610 ;
        RECT 306.060 2.400 306.200 31.290 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 44.440 324.230 44.500 ;
        RECT 835.430 44.440 835.750 44.500 ;
        RECT 323.910 44.300 835.750 44.440 ;
        RECT 323.910 44.240 324.230 44.300 ;
        RECT 835.430 44.240 835.750 44.300 ;
      LAYER via ;
        RECT 323.940 44.240 324.200 44.500 ;
        RECT 835.460 44.240 835.720 44.500 ;
      LAYER met2 ;
        RECT 836.610 600.170 836.890 604.000 ;
        RECT 835.520 600.030 836.890 600.170 ;
        RECT 835.520 44.530 835.660 600.030 ;
        RECT 836.610 600.000 836.890 600.030 ;
        RECT 323.940 44.210 324.200 44.530 ;
        RECT 835.460 44.210 835.720 44.530 ;
        RECT 324.000 2.400 324.140 44.210 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 840.950 72.660 841.270 72.720 ;
        RECT 842.330 72.660 842.650 72.720 ;
        RECT 840.950 72.520 842.650 72.660 ;
        RECT 840.950 72.460 841.270 72.520 ;
        RECT 842.330 72.460 842.650 72.520 ;
        RECT 840.950 48.520 841.270 48.580 ;
        RECT 841.870 48.520 842.190 48.580 ;
        RECT 840.950 48.380 842.190 48.520 ;
        RECT 840.950 48.320 841.270 48.380 ;
        RECT 841.870 48.320 842.190 48.380 ;
        RECT 341.390 31.860 341.710 31.920 ;
        RECT 841.870 31.860 842.190 31.920 ;
        RECT 341.390 31.720 842.190 31.860 ;
        RECT 341.390 31.660 341.710 31.720 ;
        RECT 841.870 31.660 842.190 31.720 ;
      LAYER via ;
        RECT 840.980 72.460 841.240 72.720 ;
        RECT 842.360 72.460 842.620 72.720 ;
        RECT 840.980 48.320 841.240 48.580 ;
        RECT 841.900 48.320 842.160 48.580 ;
        RECT 341.420 31.660 341.680 31.920 ;
        RECT 841.900 31.660 842.160 31.920 ;
      LAYER met2 ;
        RECT 845.810 600.170 846.090 604.000 ;
        RECT 844.260 600.030 846.090 600.170 ;
        RECT 844.260 596.770 844.400 600.030 ;
        RECT 845.810 600.000 846.090 600.030 ;
        RECT 842.420 596.630 844.400 596.770 ;
        RECT 842.420 72.750 842.560 596.630 ;
        RECT 840.980 72.430 841.240 72.750 ;
        RECT 842.360 72.430 842.620 72.750 ;
        RECT 841.040 48.610 841.180 72.430 ;
        RECT 840.980 48.290 841.240 48.610 ;
        RECT 841.900 48.290 842.160 48.610 ;
        RECT 841.960 31.950 842.100 48.290 ;
        RECT 341.420 31.630 341.680 31.950 ;
        RECT 841.900 31.630 842.160 31.950 ;
        RECT 341.480 2.400 341.620 31.630 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 849.230 557.500 849.550 557.560 ;
        RECT 853.370 557.500 853.690 557.560 ;
        RECT 849.230 557.360 853.690 557.500 ;
        RECT 849.230 557.300 849.550 557.360 ;
        RECT 853.370 557.300 853.690 557.360 ;
        RECT 359.330 44.100 359.650 44.160 ;
        RECT 849.230 44.100 849.550 44.160 ;
        RECT 359.330 43.960 849.550 44.100 ;
        RECT 359.330 43.900 359.650 43.960 ;
        RECT 849.230 43.900 849.550 43.960 ;
      LAYER via ;
        RECT 849.260 557.300 849.520 557.560 ;
        RECT 853.400 557.300 853.660 557.560 ;
        RECT 359.360 43.900 359.620 44.160 ;
        RECT 849.260 43.900 849.520 44.160 ;
      LAYER met2 ;
        RECT 855.010 600.170 855.290 604.000 ;
        RECT 853.460 600.030 855.290 600.170 ;
        RECT 853.460 557.590 853.600 600.030 ;
        RECT 855.010 600.000 855.290 600.030 ;
        RECT 849.260 557.270 849.520 557.590 ;
        RECT 853.400 557.270 853.660 557.590 ;
        RECT 849.320 44.190 849.460 557.270 ;
        RECT 359.360 43.870 359.620 44.190 ;
        RECT 849.260 43.870 849.520 44.190 ;
        RECT 359.420 2.400 359.560 43.870 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 377.270 32.200 377.590 32.260 ;
        RECT 863.030 32.200 863.350 32.260 ;
        RECT 377.270 32.060 863.350 32.200 ;
        RECT 377.270 32.000 377.590 32.060 ;
        RECT 863.030 32.000 863.350 32.060 ;
      LAYER via ;
        RECT 377.300 32.000 377.560 32.260 ;
        RECT 863.060 32.000 863.320 32.260 ;
      LAYER met2 ;
        RECT 864.210 600.170 864.490 604.000 ;
        RECT 863.120 600.030 864.490 600.170 ;
        RECT 863.120 32.290 863.260 600.030 ;
        RECT 864.210 600.000 864.490 600.030 ;
        RECT 377.300 31.970 377.560 32.290 ;
        RECT 863.060 31.970 863.320 32.290 ;
        RECT 377.360 2.400 377.500 31.970 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 869.930 579.600 870.250 579.660 ;
        RECT 871.770 579.600 872.090 579.660 ;
        RECT 869.930 579.460 872.090 579.600 ;
        RECT 869.930 579.400 870.250 579.460 ;
        RECT 871.770 579.400 872.090 579.460 ;
        RECT 869.930 572.460 870.250 572.520 ;
        RECT 871.770 572.460 872.090 572.520 ;
        RECT 869.930 572.320 872.090 572.460 ;
        RECT 869.930 572.260 870.250 572.320 ;
        RECT 871.770 572.260 872.090 572.320 ;
        RECT 869.930 524.520 870.250 524.580 ;
        RECT 870.850 524.520 871.170 524.580 ;
        RECT 869.930 524.380 871.170 524.520 ;
        RECT 869.930 524.320 870.250 524.380 ;
        RECT 870.850 524.320 871.170 524.380 ;
        RECT 870.850 483.180 871.170 483.440 ;
        RECT 869.930 483.040 870.250 483.100 ;
        RECT 870.940 483.040 871.080 483.180 ;
        RECT 869.930 482.900 871.080 483.040 ;
        RECT 869.930 482.840 870.250 482.900 ;
        RECT 869.470 476.240 869.790 476.300 ;
        RECT 869.930 476.240 870.250 476.300 ;
        RECT 869.470 476.100 870.250 476.240 ;
        RECT 869.470 476.040 869.790 476.100 ;
        RECT 869.930 476.040 870.250 476.100 ;
        RECT 869.930 338.000 870.250 338.260 ;
        RECT 870.020 337.520 870.160 338.000 ;
        RECT 870.390 337.520 870.710 337.580 ;
        RECT 870.020 337.380 870.710 337.520 ;
        RECT 870.390 337.320 870.710 337.380 ;
        RECT 870.390 324.260 870.710 324.320 ;
        RECT 871.310 324.260 871.630 324.320 ;
        RECT 870.390 324.120 871.630 324.260 ;
        RECT 870.390 324.060 870.710 324.120 ;
        RECT 871.310 324.060 871.630 324.120 ;
        RECT 869.930 193.360 870.250 193.420 ;
        RECT 871.310 193.360 871.630 193.420 ;
        RECT 869.930 193.220 871.630 193.360 ;
        RECT 869.930 193.160 870.250 193.220 ;
        RECT 871.310 193.160 871.630 193.220 ;
        RECT 869.930 145.220 870.250 145.480 ;
        RECT 870.020 145.080 870.160 145.220 ;
        RECT 870.390 145.080 870.710 145.140 ;
        RECT 870.020 144.940 870.710 145.080 ;
        RECT 870.390 144.880 870.710 144.940 ;
        RECT 869.010 137.940 869.330 138.000 ;
        RECT 870.390 137.940 870.710 138.000 ;
        RECT 869.010 137.800 870.710 137.940 ;
        RECT 869.010 137.740 869.330 137.800 ;
        RECT 870.390 137.740 870.710 137.800 ;
        RECT 869.010 90.000 869.330 90.060 ;
        RECT 869.930 90.000 870.250 90.060 ;
        RECT 869.010 89.860 870.250 90.000 ;
        RECT 869.010 89.800 869.330 89.860 ;
        RECT 869.930 89.800 870.250 89.860 ;
        RECT 395.210 43.760 395.530 43.820 ;
        RECT 869.930 43.760 870.250 43.820 ;
        RECT 395.210 43.620 870.250 43.760 ;
        RECT 395.210 43.560 395.530 43.620 ;
        RECT 869.930 43.560 870.250 43.620 ;
      LAYER via ;
        RECT 869.960 579.400 870.220 579.660 ;
        RECT 871.800 579.400 872.060 579.660 ;
        RECT 869.960 572.260 870.220 572.520 ;
        RECT 871.800 572.260 872.060 572.520 ;
        RECT 869.960 524.320 870.220 524.580 ;
        RECT 870.880 524.320 871.140 524.580 ;
        RECT 870.880 483.180 871.140 483.440 ;
        RECT 869.960 482.840 870.220 483.100 ;
        RECT 869.500 476.040 869.760 476.300 ;
        RECT 869.960 476.040 870.220 476.300 ;
        RECT 869.960 338.000 870.220 338.260 ;
        RECT 870.420 337.320 870.680 337.580 ;
        RECT 870.420 324.060 870.680 324.320 ;
        RECT 871.340 324.060 871.600 324.320 ;
        RECT 869.960 193.160 870.220 193.420 ;
        RECT 871.340 193.160 871.600 193.420 ;
        RECT 869.960 145.220 870.220 145.480 ;
        RECT 870.420 144.880 870.680 145.140 ;
        RECT 869.040 137.740 869.300 138.000 ;
        RECT 870.420 137.740 870.680 138.000 ;
        RECT 869.040 89.800 869.300 90.060 ;
        RECT 869.960 89.800 870.220 90.060 ;
        RECT 395.240 43.560 395.500 43.820 ;
        RECT 869.960 43.560 870.220 43.820 ;
      LAYER met2 ;
        RECT 873.410 600.170 873.690 604.000 ;
        RECT 871.860 600.030 873.690 600.170 ;
        RECT 871.860 596.770 872.000 600.030 ;
        RECT 873.410 600.000 873.690 600.030 ;
        RECT 870.020 596.630 872.000 596.770 ;
        RECT 870.020 579.690 870.160 596.630 ;
        RECT 869.960 579.370 870.220 579.690 ;
        RECT 871.800 579.370 872.060 579.690 ;
        RECT 871.860 572.550 872.000 579.370 ;
        RECT 869.960 572.230 870.220 572.550 ;
        RECT 871.800 572.230 872.060 572.550 ;
        RECT 870.020 524.610 870.160 572.230 ;
        RECT 869.960 524.290 870.220 524.610 ;
        RECT 870.880 524.290 871.140 524.610 ;
        RECT 870.940 483.470 871.080 524.290 ;
        RECT 870.880 483.150 871.140 483.470 ;
        RECT 869.960 482.810 870.220 483.130 ;
        RECT 870.020 476.330 870.160 482.810 ;
        RECT 869.500 476.010 869.760 476.330 ;
        RECT 869.960 476.010 870.220 476.330 ;
        RECT 869.560 434.930 869.700 476.010 ;
        RECT 869.560 434.790 870.160 434.930 ;
        RECT 870.020 400.930 870.160 434.790 ;
        RECT 869.560 400.790 870.160 400.930 ;
        RECT 869.560 386.650 869.700 400.790 ;
        RECT 869.560 386.510 870.160 386.650 ;
        RECT 870.020 338.290 870.160 386.510 ;
        RECT 869.960 337.970 870.220 338.290 ;
        RECT 870.420 337.290 870.680 337.610 ;
        RECT 870.480 324.350 870.620 337.290 ;
        RECT 870.420 324.030 870.680 324.350 ;
        RECT 871.340 324.030 871.600 324.350 ;
        RECT 871.400 193.450 871.540 324.030 ;
        RECT 869.960 193.130 870.220 193.450 ;
        RECT 871.340 193.130 871.600 193.450 ;
        RECT 870.020 145.510 870.160 193.130 ;
        RECT 869.960 145.190 870.220 145.510 ;
        RECT 870.420 144.850 870.680 145.170 ;
        RECT 870.480 138.030 870.620 144.850 ;
        RECT 869.040 137.710 869.300 138.030 ;
        RECT 870.420 137.710 870.680 138.030 ;
        RECT 869.100 90.090 869.240 137.710 ;
        RECT 869.040 89.770 869.300 90.090 ;
        RECT 869.960 89.770 870.220 90.090 ;
        RECT 870.020 43.850 870.160 89.770 ;
        RECT 395.240 43.530 395.500 43.850 ;
        RECT 869.960 43.530 870.220 43.850 ;
        RECT 395.300 2.400 395.440 43.530 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 876.830 569.400 877.150 569.460 ;
        RECT 880.970 569.400 881.290 569.460 ;
        RECT 876.830 569.260 881.290 569.400 ;
        RECT 876.830 569.200 877.150 569.260 ;
        RECT 880.970 569.200 881.290 569.260 ;
        RECT 413.150 32.880 413.470 32.940 ;
        RECT 876.830 32.880 877.150 32.940 ;
        RECT 413.150 32.740 877.150 32.880 ;
        RECT 413.150 32.680 413.470 32.740 ;
        RECT 876.830 32.680 877.150 32.740 ;
      LAYER via ;
        RECT 876.860 569.200 877.120 569.460 ;
        RECT 881.000 569.200 881.260 569.460 ;
        RECT 413.180 32.680 413.440 32.940 ;
        RECT 876.860 32.680 877.120 32.940 ;
      LAYER met2 ;
        RECT 882.610 600.170 882.890 604.000 ;
        RECT 881.060 600.030 882.890 600.170 ;
        RECT 881.060 569.490 881.200 600.030 ;
        RECT 882.610 600.000 882.890 600.030 ;
        RECT 876.860 569.170 877.120 569.490 ;
        RECT 881.000 569.170 881.260 569.490 ;
        RECT 876.920 32.970 877.060 569.170 ;
        RECT 413.180 32.650 413.440 32.970 ;
        RECT 876.860 32.650 877.120 32.970 ;
        RECT 413.240 2.400 413.380 32.650 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 703.870 560.560 704.190 560.620 ;
        RECT 706.170 560.560 706.490 560.620 ;
        RECT 703.870 560.420 706.490 560.560 ;
        RECT 703.870 560.360 704.190 560.420 ;
        RECT 706.170 560.360 706.490 560.420 ;
        RECT 74.130 18.260 74.450 18.320 ;
        RECT 703.870 18.260 704.190 18.320 ;
        RECT 74.130 18.120 704.190 18.260 ;
        RECT 74.130 18.060 74.450 18.120 ;
        RECT 703.870 18.060 704.190 18.120 ;
      LAYER via ;
        RECT 703.900 560.360 704.160 560.620 ;
        RECT 706.200 560.360 706.460 560.620 ;
        RECT 74.160 18.060 74.420 18.320 ;
        RECT 703.900 18.060 704.160 18.320 ;
      LAYER met2 ;
        RECT 707.810 600.170 708.090 604.000 ;
        RECT 706.260 600.030 708.090 600.170 ;
        RECT 706.260 560.650 706.400 600.030 ;
        RECT 707.810 600.000 708.090 600.030 ;
        RECT 703.900 560.330 704.160 560.650 ;
        RECT 706.200 560.330 706.460 560.650 ;
        RECT 703.960 18.350 704.100 560.330 ;
        RECT 74.160 18.030 74.420 18.350 ;
        RECT 703.900 18.030 704.160 18.350 ;
        RECT 74.220 2.400 74.360 18.030 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 430.630 33.220 430.950 33.280 ;
        RECT 890.630 33.220 890.950 33.280 ;
        RECT 430.630 33.080 890.950 33.220 ;
        RECT 430.630 33.020 430.950 33.080 ;
        RECT 890.630 33.020 890.950 33.080 ;
      LAYER via ;
        RECT 430.660 33.020 430.920 33.280 ;
        RECT 890.660 33.020 890.920 33.280 ;
      LAYER met2 ;
        RECT 891.810 600.170 892.090 604.000 ;
        RECT 890.720 600.030 892.090 600.170 ;
        RECT 890.720 33.310 890.860 600.030 ;
        RECT 891.810 600.000 892.090 600.030 ;
        RECT 430.660 32.990 430.920 33.310 ;
        RECT 890.660 32.990 890.920 33.310 ;
        RECT 430.720 2.400 430.860 32.990 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 897.530 531.320 897.850 531.380 ;
        RECT 897.990 531.320 898.310 531.380 ;
        RECT 897.530 531.180 898.310 531.320 ;
        RECT 897.530 531.120 897.850 531.180 ;
        RECT 897.990 531.120 898.310 531.180 ;
        RECT 897.990 496.980 898.310 497.040 ;
        RECT 897.620 496.840 898.310 496.980 ;
        RECT 897.620 496.700 897.760 496.840 ;
        RECT 897.990 496.780 898.310 496.840 ;
        RECT 897.530 496.440 897.850 496.700 ;
        RECT 897.070 448.700 897.390 448.760 ;
        RECT 897.990 448.700 898.310 448.760 ;
        RECT 897.070 448.560 898.310 448.700 ;
        RECT 897.070 448.500 897.390 448.560 ;
        RECT 897.990 448.500 898.310 448.560 ;
        RECT 898.450 352.480 898.770 352.540 ;
        RECT 898.080 352.340 898.770 352.480 ;
        RECT 898.080 351.860 898.220 352.340 ;
        RECT 898.450 352.280 898.770 352.340 ;
        RECT 897.990 351.600 898.310 351.860 ;
        RECT 896.150 265.780 896.470 265.840 ;
        RECT 897.070 265.780 897.390 265.840 ;
        RECT 896.150 265.640 897.390 265.780 ;
        RECT 896.150 265.580 896.470 265.640 ;
        RECT 897.070 265.580 897.390 265.640 ;
        RECT 896.150 234.500 896.470 234.560 ;
        RECT 897.070 234.500 897.390 234.560 ;
        RECT 896.150 234.360 897.390 234.500 ;
        RECT 896.150 234.300 896.470 234.360 ;
        RECT 897.070 234.300 897.390 234.360 ;
        RECT 896.150 186.560 896.470 186.620 ;
        RECT 897.530 186.560 897.850 186.620 ;
        RECT 896.150 186.420 897.850 186.560 ;
        RECT 896.150 186.360 896.470 186.420 ;
        RECT 897.530 186.360 897.850 186.420 ;
        RECT 897.530 96.460 897.850 96.520 ;
        RECT 898.450 96.460 898.770 96.520 ;
        RECT 897.530 96.320 898.770 96.460 ;
        RECT 897.530 96.260 897.850 96.320 ;
        RECT 898.450 96.260 898.770 96.320 ;
        RECT 897.530 48.520 897.850 48.580 ;
        RECT 898.910 48.520 899.230 48.580 ;
        RECT 897.530 48.380 899.230 48.520 ;
        RECT 897.530 48.320 897.850 48.380 ;
        RECT 898.910 48.320 899.230 48.380 ;
        RECT 448.570 16.220 448.890 16.280 ;
        RECT 898.910 16.220 899.230 16.280 ;
        RECT 448.570 16.080 899.230 16.220 ;
        RECT 448.570 16.020 448.890 16.080 ;
        RECT 898.910 16.020 899.230 16.080 ;
      LAYER via ;
        RECT 897.560 531.120 897.820 531.380 ;
        RECT 898.020 531.120 898.280 531.380 ;
        RECT 898.020 496.780 898.280 497.040 ;
        RECT 897.560 496.440 897.820 496.700 ;
        RECT 897.100 448.500 897.360 448.760 ;
        RECT 898.020 448.500 898.280 448.760 ;
        RECT 898.480 352.280 898.740 352.540 ;
        RECT 898.020 351.600 898.280 351.860 ;
        RECT 896.180 265.580 896.440 265.840 ;
        RECT 897.100 265.580 897.360 265.840 ;
        RECT 896.180 234.300 896.440 234.560 ;
        RECT 897.100 234.300 897.360 234.560 ;
        RECT 896.180 186.360 896.440 186.620 ;
        RECT 897.560 186.360 897.820 186.620 ;
        RECT 897.560 96.260 897.820 96.520 ;
        RECT 898.480 96.260 898.740 96.520 ;
        RECT 897.560 48.320 897.820 48.580 ;
        RECT 898.940 48.320 899.200 48.580 ;
        RECT 448.600 16.020 448.860 16.280 ;
        RECT 898.940 16.020 899.200 16.280 ;
      LAYER met2 ;
        RECT 901.010 600.170 901.290 604.000 ;
        RECT 899.460 600.030 901.290 600.170 ;
        RECT 899.460 596.770 899.600 600.030 ;
        RECT 901.010 600.000 901.290 600.030 ;
        RECT 897.620 596.630 899.600 596.770 ;
        RECT 897.620 569.400 897.760 596.630 ;
        RECT 897.160 569.260 897.760 569.400 ;
        RECT 897.160 545.090 897.300 569.260 ;
        RECT 897.160 544.950 897.760 545.090 ;
        RECT 897.620 531.410 897.760 544.950 ;
        RECT 897.560 531.090 897.820 531.410 ;
        RECT 898.020 531.090 898.280 531.410 ;
        RECT 898.080 497.070 898.220 531.090 ;
        RECT 898.020 496.750 898.280 497.070 ;
        RECT 897.560 496.410 897.820 496.730 ;
        RECT 897.620 483.210 897.760 496.410 ;
        RECT 897.620 483.070 898.220 483.210 ;
        RECT 898.080 448.790 898.220 483.070 ;
        RECT 897.100 448.530 897.360 448.790 ;
        RECT 897.100 448.470 897.760 448.530 ;
        RECT 898.020 448.470 898.280 448.790 ;
        RECT 897.160 448.390 897.760 448.470 ;
        RECT 897.620 447.850 897.760 448.390 ;
        RECT 897.620 447.710 898.680 447.850 ;
        RECT 898.540 387.330 898.680 447.710 ;
        RECT 898.080 387.190 898.680 387.330 ;
        RECT 898.080 386.650 898.220 387.190 ;
        RECT 898.080 386.510 898.680 386.650 ;
        RECT 898.540 352.570 898.680 386.510 ;
        RECT 898.480 352.250 898.740 352.570 ;
        RECT 898.020 351.570 898.280 351.890 ;
        RECT 898.080 303.690 898.220 351.570 ;
        RECT 897.160 303.550 898.220 303.690 ;
        RECT 897.160 265.870 897.300 303.550 ;
        RECT 896.180 265.550 896.440 265.870 ;
        RECT 897.100 265.550 897.360 265.870 ;
        RECT 896.240 241.925 896.380 265.550 ;
        RECT 896.170 241.555 896.450 241.925 ;
        RECT 897.090 241.555 897.370 241.925 ;
        RECT 897.160 234.590 897.300 241.555 ;
        RECT 896.180 234.270 896.440 234.590 ;
        RECT 897.100 234.270 897.360 234.590 ;
        RECT 896.240 186.650 896.380 234.270 ;
        RECT 896.180 186.330 896.440 186.650 ;
        RECT 897.560 186.330 897.820 186.650 ;
        RECT 897.620 110.570 897.760 186.330 ;
        RECT 897.620 110.430 898.680 110.570 ;
        RECT 898.540 96.550 898.680 110.430 ;
        RECT 897.560 96.230 897.820 96.550 ;
        RECT 898.480 96.230 898.740 96.550 ;
        RECT 897.620 48.610 897.760 96.230 ;
        RECT 897.560 48.290 897.820 48.610 ;
        RECT 898.940 48.290 899.200 48.610 ;
        RECT 899.000 16.310 899.140 48.290 ;
        RECT 448.600 15.990 448.860 16.310 ;
        RECT 898.940 15.990 899.200 16.310 ;
        RECT 448.660 2.400 448.800 15.990 ;
        RECT 448.450 -4.800 449.010 2.400 ;
      LAYER via2 ;
        RECT 896.170 241.600 896.450 241.880 ;
        RECT 897.090 241.600 897.370 241.880 ;
      LAYER met3 ;
        RECT 896.145 241.890 896.475 241.905 ;
        RECT 897.065 241.890 897.395 241.905 ;
        RECT 896.145 241.590 897.395 241.890 ;
        RECT 896.145 241.575 896.475 241.590 ;
        RECT 897.065 241.575 897.395 241.590 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 33.900 466.830 33.960 ;
        RECT 904.890 33.900 905.210 33.960 ;
        RECT 466.510 33.760 905.210 33.900 ;
        RECT 466.510 33.700 466.830 33.760 ;
        RECT 904.890 33.700 905.210 33.760 ;
      LAYER via ;
        RECT 466.540 33.700 466.800 33.960 ;
        RECT 904.920 33.700 905.180 33.960 ;
      LAYER met2 ;
        RECT 910.210 600.170 910.490 604.000 ;
        RECT 907.740 600.030 910.490 600.170 ;
        RECT 907.740 596.770 907.880 600.030 ;
        RECT 910.210 600.000 910.490 600.030 ;
        RECT 905.900 596.630 907.880 596.770 ;
        RECT 905.900 569.400 906.040 596.630 ;
        RECT 904.980 569.260 906.040 569.400 ;
        RECT 904.980 33.990 905.120 569.260 ;
        RECT 466.540 33.670 466.800 33.990 ;
        RECT 904.920 33.670 905.180 33.990 ;
        RECT 466.600 2.400 466.740 33.670 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 917.770 15.880 918.090 15.940 ;
        RECT 496.960 15.740 918.090 15.880 ;
        RECT 484.450 15.540 484.770 15.600 ;
        RECT 496.960 15.540 497.100 15.740 ;
        RECT 917.770 15.680 918.090 15.740 ;
        RECT 484.450 15.400 497.100 15.540 ;
        RECT 484.450 15.340 484.770 15.400 ;
      LAYER via ;
        RECT 484.480 15.340 484.740 15.600 ;
        RECT 917.800 15.680 918.060 15.940 ;
      LAYER met2 ;
        RECT 919.410 600.170 919.690 604.000 ;
        RECT 917.860 600.030 919.690 600.170 ;
        RECT 917.860 15.970 918.000 600.030 ;
        RECT 919.410 600.000 919.690 600.030 ;
        RECT 917.800 15.650 918.060 15.970 ;
        RECT 484.480 15.310 484.740 15.630 ;
        RECT 484.540 2.400 484.680 15.310 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 502.390 40.360 502.710 40.420 ;
        RECT 924.670 40.360 924.990 40.420 ;
        RECT 502.390 40.220 924.990 40.360 ;
        RECT 502.390 40.160 502.710 40.220 ;
        RECT 924.670 40.160 924.990 40.220 ;
      LAYER via ;
        RECT 502.420 40.160 502.680 40.420 ;
        RECT 924.700 40.160 924.960 40.420 ;
      LAYER met2 ;
        RECT 928.610 600.170 928.890 604.000 ;
        RECT 927.060 600.030 928.890 600.170 ;
        RECT 927.060 596.770 927.200 600.030 ;
        RECT 928.610 600.000 928.890 600.030 ;
        RECT 925.220 596.630 927.200 596.770 ;
        RECT 925.220 569.400 925.360 596.630 ;
        RECT 924.760 569.260 925.360 569.400 ;
        RECT 924.760 40.450 924.900 569.260 ;
        RECT 502.420 40.130 502.680 40.450 ;
        RECT 924.700 40.130 924.960 40.450 ;
        RECT 502.480 2.400 502.620 40.130 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 15.540 520.190 15.600 ;
        RECT 932.950 15.540 933.270 15.600 ;
        RECT 519.870 15.400 933.270 15.540 ;
        RECT 519.870 15.340 520.190 15.400 ;
        RECT 932.950 15.340 933.270 15.400 ;
      LAYER via ;
        RECT 519.900 15.340 520.160 15.600 ;
        RECT 932.980 15.340 933.240 15.600 ;
      LAYER met2 ;
        RECT 937.350 600.170 937.630 604.000 ;
        RECT 935.340 600.030 937.630 600.170 ;
        RECT 935.340 596.770 935.480 600.030 ;
        RECT 937.350 600.000 937.630 600.030 ;
        RECT 933.500 596.630 935.480 596.770 ;
        RECT 933.500 568.890 933.640 596.630 ;
        RECT 933.040 568.750 933.640 568.890 ;
        RECT 933.040 15.630 933.180 568.750 ;
        RECT 519.900 15.310 520.160 15.630 ;
        RECT 932.980 15.310 933.240 15.630 ;
        RECT 519.960 2.400 520.100 15.310 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 40.700 538.130 40.760 ;
        RECT 945.830 40.700 946.150 40.760 ;
        RECT 537.810 40.560 946.150 40.700 ;
        RECT 537.810 40.500 538.130 40.560 ;
        RECT 945.830 40.500 946.150 40.560 ;
      LAYER via ;
        RECT 537.840 40.500 538.100 40.760 ;
        RECT 945.860 40.500 946.120 40.760 ;
      LAYER met2 ;
        RECT 946.550 600.170 946.830 604.000 ;
        RECT 945.920 600.030 946.830 600.170 ;
        RECT 945.920 40.790 946.060 600.030 ;
        RECT 946.550 600.000 946.830 600.030 ;
        RECT 537.840 40.470 538.100 40.790 ;
        RECT 945.860 40.470 946.120 40.790 ;
        RECT 537.900 2.400 538.040 40.470 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 953.650 579.940 953.970 580.000 ;
        RECT 955.030 579.940 955.350 580.000 ;
        RECT 953.650 579.800 955.350 579.940 ;
        RECT 953.650 579.740 953.970 579.800 ;
        RECT 955.030 579.740 955.350 579.800 ;
        RECT 953.190 496.980 953.510 497.040 ;
        RECT 954.110 496.980 954.430 497.040 ;
        RECT 953.190 496.840 954.430 496.980 ;
        RECT 953.190 496.780 953.510 496.840 ;
        RECT 954.110 496.780 954.430 496.840 ;
        RECT 952.730 379.680 953.050 379.740 ;
        RECT 954.110 379.680 954.430 379.740 ;
        RECT 952.730 379.540 954.430 379.680 ;
        RECT 952.730 379.480 953.050 379.540 ;
        RECT 954.110 379.480 954.430 379.540 ;
        RECT 952.730 379.000 953.050 379.060 ;
        RECT 953.650 379.000 953.970 379.060 ;
        RECT 952.730 378.860 953.970 379.000 ;
        RECT 952.730 378.800 953.050 378.860 ;
        RECT 953.650 378.800 953.970 378.860 ;
        RECT 953.650 351.940 953.970 352.200 ;
        RECT 953.190 351.800 953.510 351.860 ;
        RECT 953.740 351.800 953.880 351.940 ;
        RECT 953.190 351.660 953.880 351.800 ;
        RECT 953.190 351.600 953.510 351.660 ;
        RECT 953.190 303.520 953.510 303.580 ;
        RECT 954.110 303.520 954.430 303.580 ;
        RECT 953.190 303.380 954.430 303.520 ;
        RECT 953.190 303.320 953.510 303.380 ;
        RECT 954.110 303.320 954.430 303.380 ;
        RECT 952.730 186.560 953.050 186.620 ;
        RECT 953.650 186.560 953.970 186.620 ;
        RECT 952.730 186.420 953.970 186.560 ;
        RECT 952.730 186.360 953.050 186.420 ;
        RECT 953.650 186.360 953.970 186.420 ;
        RECT 953.190 137.740 953.510 138.000 ;
        RECT 953.280 137.320 953.420 137.740 ;
        RECT 953.190 137.060 953.510 137.320 ;
        RECT 555.750 15.200 556.070 15.260 ;
        RECT 953.190 15.200 953.510 15.260 ;
        RECT 555.750 15.060 953.510 15.200 ;
        RECT 555.750 15.000 556.070 15.060 ;
        RECT 953.190 15.000 953.510 15.060 ;
      LAYER via ;
        RECT 953.680 579.740 953.940 580.000 ;
        RECT 955.060 579.740 955.320 580.000 ;
        RECT 953.220 496.780 953.480 497.040 ;
        RECT 954.140 496.780 954.400 497.040 ;
        RECT 952.760 379.480 953.020 379.740 ;
        RECT 954.140 379.480 954.400 379.740 ;
        RECT 952.760 378.800 953.020 379.060 ;
        RECT 953.680 378.800 953.940 379.060 ;
        RECT 953.680 351.940 953.940 352.200 ;
        RECT 953.220 351.600 953.480 351.860 ;
        RECT 953.220 303.320 953.480 303.580 ;
        RECT 954.140 303.320 954.400 303.580 ;
        RECT 952.760 186.360 953.020 186.620 ;
        RECT 953.680 186.360 953.940 186.620 ;
        RECT 953.220 137.740 953.480 138.000 ;
        RECT 953.220 137.060 953.480 137.320 ;
        RECT 555.780 15.000 556.040 15.260 ;
        RECT 953.220 15.000 953.480 15.260 ;
      LAYER met2 ;
        RECT 955.750 600.170 956.030 604.000 ;
        RECT 955.120 600.030 956.030 600.170 ;
        RECT 955.120 580.030 955.260 600.030 ;
        RECT 955.750 600.000 956.030 600.030 ;
        RECT 953.680 579.710 953.940 580.030 ;
        RECT 955.060 579.710 955.320 580.030 ;
        RECT 953.740 555.290 953.880 579.710 ;
        RECT 953.740 555.150 954.800 555.290 ;
        RECT 954.660 544.410 954.800 555.150 ;
        RECT 954.200 544.270 954.800 544.410 ;
        RECT 954.200 497.070 954.340 544.270 ;
        RECT 953.220 496.750 953.480 497.070 ;
        RECT 954.140 496.750 954.400 497.070 ;
        RECT 953.280 434.930 953.420 496.750 ;
        RECT 953.280 434.790 953.880 434.930 ;
        RECT 953.740 400.930 953.880 434.790 ;
        RECT 953.740 400.790 954.340 400.930 ;
        RECT 954.200 379.770 954.340 400.790 ;
        RECT 952.760 379.450 953.020 379.770 ;
        RECT 954.140 379.450 954.400 379.770 ;
        RECT 952.820 379.090 952.960 379.450 ;
        RECT 952.760 378.770 953.020 379.090 ;
        RECT 953.680 378.770 953.940 379.090 ;
        RECT 953.740 352.230 953.880 378.770 ;
        RECT 953.680 351.910 953.940 352.230 ;
        RECT 953.220 351.570 953.480 351.890 ;
        RECT 953.280 303.610 953.420 351.570 ;
        RECT 953.220 303.290 953.480 303.610 ;
        RECT 954.140 303.290 954.400 303.610 ;
        RECT 954.200 255.410 954.340 303.290 ;
        RECT 953.740 255.270 954.340 255.410 ;
        RECT 953.740 186.650 953.880 255.270 ;
        RECT 952.760 186.330 953.020 186.650 ;
        RECT 953.680 186.330 953.940 186.650 ;
        RECT 952.820 158.170 952.960 186.330 ;
        RECT 952.820 158.030 953.420 158.170 ;
        RECT 953.280 138.030 953.420 158.030 ;
        RECT 953.220 137.710 953.480 138.030 ;
        RECT 953.220 137.030 953.480 137.350 ;
        RECT 953.280 15.290 953.420 137.030 ;
        RECT 555.780 14.970 556.040 15.290 ;
        RECT 953.220 14.970 953.480 15.290 ;
        RECT 555.840 2.400 555.980 14.970 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 959.630 569.400 959.950 569.460 ;
        RECT 963.310 569.400 963.630 569.460 ;
        RECT 959.630 569.260 963.630 569.400 ;
        RECT 959.630 569.200 959.950 569.260 ;
        RECT 963.310 569.200 963.630 569.260 ;
        RECT 573.690 41.040 574.010 41.100 ;
        RECT 959.630 41.040 959.950 41.100 ;
        RECT 573.690 40.900 959.950 41.040 ;
        RECT 573.690 40.840 574.010 40.900 ;
        RECT 959.630 40.840 959.950 40.900 ;
      LAYER via ;
        RECT 959.660 569.200 959.920 569.460 ;
        RECT 963.340 569.200 963.600 569.460 ;
        RECT 573.720 40.840 573.980 41.100 ;
        RECT 959.660 40.840 959.920 41.100 ;
      LAYER met2 ;
        RECT 964.950 600.170 965.230 604.000 ;
        RECT 963.400 600.030 965.230 600.170 ;
        RECT 963.400 569.490 963.540 600.030 ;
        RECT 964.950 600.000 965.230 600.030 ;
        RECT 959.660 569.170 959.920 569.490 ;
        RECT 963.340 569.170 963.600 569.490 ;
        RECT 959.720 41.130 959.860 569.170 ;
        RECT 573.720 40.810 573.980 41.130 ;
        RECT 959.660 40.810 959.920 41.130 ;
        RECT 573.780 2.400 573.920 40.810 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 591.170 14.860 591.490 14.920 ;
        RECT 973.890 14.860 974.210 14.920 ;
        RECT 591.170 14.720 974.210 14.860 ;
        RECT 591.170 14.660 591.490 14.720 ;
        RECT 973.890 14.660 974.210 14.720 ;
      LAYER via ;
        RECT 591.200 14.660 591.460 14.920 ;
        RECT 973.920 14.660 974.180 14.920 ;
      LAYER met2 ;
        RECT 974.150 600.000 974.430 604.000 ;
        RECT 974.210 598.810 974.350 600.000 ;
        RECT 973.980 598.670 974.350 598.810 ;
        RECT 973.980 14.950 974.120 598.670 ;
        RECT 591.200 14.630 591.460 14.950 ;
        RECT 973.920 14.630 974.180 14.950 ;
        RECT 591.260 2.400 591.400 14.630 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 18.600 97.910 18.660 ;
        RECT 717.670 18.600 717.990 18.660 ;
        RECT 97.590 18.460 717.990 18.600 ;
        RECT 97.590 18.400 97.910 18.460 ;
        RECT 717.670 18.400 717.990 18.460 ;
      LAYER via ;
        RECT 97.620 18.400 97.880 18.660 ;
        RECT 717.700 18.400 717.960 18.660 ;
      LAYER met2 ;
        RECT 720.230 600.170 720.510 604.000 ;
        RECT 717.760 600.030 720.510 600.170 ;
        RECT 717.760 18.690 717.900 600.030 ;
        RECT 720.230 600.000 720.510 600.030 ;
        RECT 97.620 18.370 97.880 18.690 ;
        RECT 717.700 18.370 717.960 18.690 ;
        RECT 97.680 2.400 97.820 18.370 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 37.640 609.430 37.700 ;
        RECT 980.330 37.640 980.650 37.700 ;
        RECT 609.110 37.500 980.650 37.640 ;
        RECT 609.110 37.440 609.430 37.500 ;
        RECT 980.330 37.440 980.650 37.500 ;
      LAYER via ;
        RECT 609.140 37.440 609.400 37.700 ;
        RECT 980.360 37.440 980.620 37.700 ;
      LAYER met2 ;
        RECT 983.350 600.850 983.630 604.000 ;
        RECT 981.340 600.710 983.630 600.850 ;
        RECT 981.340 583.170 981.480 600.710 ;
        RECT 983.350 600.000 983.630 600.710 ;
        RECT 980.420 583.030 981.480 583.170 ;
        RECT 980.420 37.730 980.560 583.030 ;
        RECT 609.140 37.410 609.400 37.730 ;
        RECT 980.360 37.410 980.620 37.730 ;
        RECT 609.200 2.400 609.340 37.410 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 987.230 36.960 987.550 37.020 ;
        RECT 638.640 36.820 987.550 36.960 ;
        RECT 627.050 36.620 627.370 36.680 ;
        RECT 638.640 36.620 638.780 36.820 ;
        RECT 987.230 36.760 987.550 36.820 ;
        RECT 627.050 36.480 638.780 36.620 ;
        RECT 627.050 36.420 627.370 36.480 ;
      LAYER via ;
        RECT 627.080 36.420 627.340 36.680 ;
        RECT 987.260 36.760 987.520 37.020 ;
      LAYER met2 ;
        RECT 992.550 600.850 992.830 604.000 ;
        RECT 990.540 600.710 992.830 600.850 ;
        RECT 990.540 583.170 990.680 600.710 ;
        RECT 992.550 600.000 992.830 600.710 ;
        RECT 987.320 583.030 990.680 583.170 ;
        RECT 987.320 37.050 987.460 583.030 ;
        RECT 987.260 36.730 987.520 37.050 ;
        RECT 627.080 36.390 627.340 36.710 ;
        RECT 627.140 2.400 627.280 36.390 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 18.940 121.830 19.000 ;
        RECT 731.470 18.940 731.790 19.000 ;
        RECT 121.510 18.800 731.790 18.940 ;
        RECT 121.510 18.740 121.830 18.800 ;
        RECT 731.470 18.740 731.790 18.800 ;
      LAYER via ;
        RECT 121.540 18.740 121.800 19.000 ;
        RECT 731.500 18.740 731.760 19.000 ;
      LAYER met2 ;
        RECT 732.650 600.170 732.930 604.000 ;
        RECT 731.560 600.030 732.930 600.170 ;
        RECT 731.560 19.030 731.700 600.030 ;
        RECT 732.650 600.000 732.930 600.030 ;
        RECT 121.540 18.710 121.800 19.030 ;
        RECT 731.500 18.710 731.760 19.030 ;
        RECT 121.600 2.400 121.740 18.710 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 740.670 427.620 740.990 427.680 ;
        RECT 741.590 427.620 741.910 427.680 ;
        RECT 740.670 427.480 741.910 427.620 ;
        RECT 740.670 427.420 740.990 427.480 ;
        RECT 741.590 427.420 741.910 427.480 ;
        RECT 739.750 379.680 740.070 379.740 ;
        RECT 741.590 379.680 741.910 379.740 ;
        RECT 739.750 379.540 741.910 379.680 ;
        RECT 739.750 379.480 740.070 379.540 ;
        RECT 741.590 379.480 741.910 379.540 ;
        RECT 739.750 338.200 740.070 338.260 ;
        RECT 740.210 338.200 740.530 338.260 ;
        RECT 739.750 338.060 740.530 338.200 ;
        RECT 739.750 338.000 740.070 338.060 ;
        RECT 740.210 338.000 740.530 338.060 ;
        RECT 740.210 255.580 740.530 255.640 ;
        RECT 739.840 255.440 740.530 255.580 ;
        RECT 739.840 255.300 739.980 255.440 ;
        RECT 740.210 255.380 740.530 255.440 ;
        RECT 739.750 255.040 740.070 255.300 ;
        RECT 739.750 234.500 740.070 234.560 ;
        RECT 739.380 234.360 740.070 234.500 ;
        RECT 739.380 234.220 739.520 234.360 ;
        RECT 739.750 234.300 740.070 234.360 ;
        RECT 739.290 233.960 739.610 234.220 ;
        RECT 739.290 120.940 739.610 121.000 ;
        RECT 740.210 120.940 740.530 121.000 ;
        RECT 739.290 120.800 740.530 120.940 ;
        RECT 739.290 120.740 739.610 120.800 ;
        RECT 740.210 120.740 740.530 120.800 ;
        RECT 145.430 25.400 145.750 25.460 ;
        RECT 740.210 25.400 740.530 25.460 ;
        RECT 145.430 25.260 740.530 25.400 ;
        RECT 145.430 25.200 145.750 25.260 ;
        RECT 740.210 25.200 740.530 25.260 ;
      LAYER via ;
        RECT 740.700 427.420 740.960 427.680 ;
        RECT 741.620 427.420 741.880 427.680 ;
        RECT 739.780 379.480 740.040 379.740 ;
        RECT 741.620 379.480 741.880 379.740 ;
        RECT 739.780 338.000 740.040 338.260 ;
        RECT 740.240 338.000 740.500 338.260 ;
        RECT 740.240 255.380 740.500 255.640 ;
        RECT 739.780 255.040 740.040 255.300 ;
        RECT 739.780 234.300 740.040 234.560 ;
        RECT 739.320 233.960 739.580 234.220 ;
        RECT 739.320 120.740 739.580 121.000 ;
        RECT 740.240 120.740 740.500 121.000 ;
        RECT 145.460 25.200 145.720 25.460 ;
        RECT 740.240 25.200 740.500 25.460 ;
      LAYER met2 ;
        RECT 744.610 600.170 744.890 604.000 ;
        RECT 743.060 600.030 744.890 600.170 ;
        RECT 743.060 569.570 743.200 600.030 ;
        RECT 744.610 600.000 744.890 600.030 ;
        RECT 739.840 569.430 743.200 569.570 ;
        RECT 739.840 448.530 739.980 569.430 ;
        RECT 739.840 448.390 740.900 448.530 ;
        RECT 740.760 427.710 740.900 448.390 ;
        RECT 740.700 427.390 740.960 427.710 ;
        RECT 741.620 427.390 741.880 427.710 ;
        RECT 741.680 379.770 741.820 427.390 ;
        RECT 739.780 379.450 740.040 379.770 ;
        RECT 741.620 379.450 741.880 379.770 ;
        RECT 739.840 338.290 739.980 379.450 ;
        RECT 739.780 337.970 740.040 338.290 ;
        RECT 740.240 337.970 740.500 338.290 ;
        RECT 740.300 255.670 740.440 337.970 ;
        RECT 740.240 255.350 740.500 255.670 ;
        RECT 739.780 255.010 740.040 255.330 ;
        RECT 739.840 234.590 739.980 255.010 ;
        RECT 739.780 234.270 740.040 234.590 ;
        RECT 739.320 233.930 739.580 234.250 ;
        RECT 739.380 121.030 739.520 233.930 ;
        RECT 739.320 120.710 739.580 121.030 ;
        RECT 740.240 120.710 740.500 121.030 ;
        RECT 740.300 25.490 740.440 120.710 ;
        RECT 145.460 25.170 145.720 25.490 ;
        RECT 740.240 25.170 740.500 25.490 ;
        RECT 145.520 2.400 145.660 25.170 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 19.620 163.690 19.680 ;
        RECT 753.090 19.620 753.410 19.680 ;
        RECT 163.370 19.480 753.410 19.620 ;
        RECT 163.370 19.420 163.690 19.480 ;
        RECT 753.090 19.420 753.410 19.480 ;
      LAYER via ;
        RECT 163.400 19.420 163.660 19.680 ;
        RECT 753.120 19.420 753.380 19.680 ;
      LAYER met2 ;
        RECT 753.810 600.170 754.090 604.000 ;
        RECT 752.260 600.030 754.090 600.170 ;
        RECT 752.260 28.290 752.400 600.030 ;
        RECT 753.810 600.000 754.090 600.030 ;
        RECT 752.260 28.150 753.320 28.290 ;
        RECT 753.180 19.710 753.320 28.150 ;
        RECT 163.400 19.390 163.660 19.710 ;
        RECT 753.120 19.390 753.380 19.710 ;
        RECT 163.460 2.400 163.600 19.390 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 759.070 569.400 759.390 569.460 ;
        RECT 761.370 569.400 761.690 569.460 ;
        RECT 759.070 569.260 761.690 569.400 ;
        RECT 759.070 569.200 759.390 569.260 ;
        RECT 761.370 569.200 761.690 569.260 ;
        RECT 180.850 46.140 181.170 46.200 ;
        RECT 759.070 46.140 759.390 46.200 ;
        RECT 180.850 46.000 759.390 46.140 ;
        RECT 180.850 45.940 181.170 46.000 ;
        RECT 759.070 45.940 759.390 46.000 ;
      LAYER via ;
        RECT 759.100 569.200 759.360 569.460 ;
        RECT 761.400 569.200 761.660 569.460 ;
        RECT 180.880 45.940 181.140 46.200 ;
        RECT 759.100 45.940 759.360 46.200 ;
      LAYER met2 ;
        RECT 763.010 600.170 763.290 604.000 ;
        RECT 761.460 600.030 763.290 600.170 ;
        RECT 761.460 569.490 761.600 600.030 ;
        RECT 763.010 600.000 763.290 600.030 ;
        RECT 759.100 569.170 759.360 569.490 ;
        RECT 761.400 569.170 761.660 569.490 ;
        RECT 759.160 46.230 759.300 569.170 ;
        RECT 180.880 45.910 181.140 46.230 ;
        RECT 759.100 45.910 759.360 46.230 ;
        RECT 180.940 2.400 181.080 45.910 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 765.970 569.400 766.290 569.460 ;
        RECT 770.570 569.400 770.890 569.460 ;
        RECT 765.970 569.260 770.890 569.400 ;
        RECT 765.970 569.200 766.290 569.260 ;
        RECT 770.570 569.200 770.890 569.260 ;
        RECT 198.790 20.300 199.110 20.360 ;
        RECT 743.890 20.300 744.210 20.360 ;
        RECT 198.790 20.160 744.210 20.300 ;
        RECT 198.790 20.100 199.110 20.160 ;
        RECT 743.890 20.100 744.210 20.160 ;
        RECT 743.890 19.280 744.210 19.340 ;
        RECT 765.970 19.280 766.290 19.340 ;
        RECT 743.890 19.140 766.290 19.280 ;
        RECT 743.890 19.080 744.210 19.140 ;
        RECT 765.970 19.080 766.290 19.140 ;
      LAYER via ;
        RECT 766.000 569.200 766.260 569.460 ;
        RECT 770.600 569.200 770.860 569.460 ;
        RECT 198.820 20.100 199.080 20.360 ;
        RECT 743.920 20.100 744.180 20.360 ;
        RECT 743.920 19.080 744.180 19.340 ;
        RECT 766.000 19.080 766.260 19.340 ;
      LAYER met2 ;
        RECT 772.210 600.170 772.490 604.000 ;
        RECT 770.660 600.030 772.490 600.170 ;
        RECT 770.660 569.490 770.800 600.030 ;
        RECT 772.210 600.000 772.490 600.030 ;
        RECT 766.000 569.170 766.260 569.490 ;
        RECT 770.600 569.170 770.860 569.490 ;
        RECT 198.820 20.070 199.080 20.390 ;
        RECT 743.920 20.070 744.180 20.390 ;
        RECT 198.880 2.400 199.020 20.070 ;
        RECT 743.980 19.370 744.120 20.070 ;
        RECT 766.060 19.370 766.200 569.170 ;
        RECT 743.920 19.050 744.180 19.370 ;
        RECT 766.000 19.050 766.260 19.370 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 46.820 217.050 46.880 ;
        RECT 780.230 46.820 780.550 46.880 ;
        RECT 216.730 46.680 780.550 46.820 ;
        RECT 216.730 46.620 217.050 46.680 ;
        RECT 780.230 46.620 780.550 46.680 ;
      LAYER via ;
        RECT 216.760 46.620 217.020 46.880 ;
        RECT 780.260 46.620 780.520 46.880 ;
      LAYER met2 ;
        RECT 781.410 600.170 781.690 604.000 ;
        RECT 780.320 600.030 781.690 600.170 ;
        RECT 780.320 46.910 780.460 600.030 ;
        RECT 781.410 600.000 781.690 600.030 ;
        RECT 216.760 46.590 217.020 46.910 ;
        RECT 780.260 46.590 780.520 46.910 ;
        RECT 216.820 2.400 216.960 46.590 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 787.130 531.320 787.450 531.380 ;
        RECT 787.590 531.320 787.910 531.380 ;
        RECT 787.130 531.180 787.910 531.320 ;
        RECT 787.130 531.120 787.450 531.180 ;
        RECT 787.590 531.120 787.910 531.180 ;
        RECT 787.130 496.640 787.450 496.700 ;
        RECT 788.050 496.640 788.370 496.700 ;
        RECT 787.130 496.500 788.370 496.640 ;
        RECT 787.130 496.440 787.450 496.500 ;
        RECT 788.050 496.440 788.370 496.500 ;
        RECT 785.750 420.820 786.070 420.880 ;
        RECT 788.510 420.820 788.830 420.880 ;
        RECT 785.750 420.680 788.830 420.820 ;
        RECT 785.750 420.620 786.070 420.680 ;
        RECT 788.510 420.620 788.830 420.680 ;
        RECT 785.750 414.020 786.070 414.080 ;
        RECT 787.130 414.020 787.450 414.080 ;
        RECT 785.750 413.880 787.450 414.020 ;
        RECT 785.750 413.820 786.070 413.880 ;
        RECT 787.130 413.820 787.450 413.880 ;
        RECT 787.130 282.920 787.450 283.180 ;
        RECT 786.670 282.780 786.990 282.840 ;
        RECT 787.220 282.780 787.360 282.920 ;
        RECT 786.670 282.640 787.360 282.780 ;
        RECT 786.670 282.580 786.990 282.640 ;
        RECT 786.670 276.320 786.990 276.380 ;
        RECT 787.590 276.320 787.910 276.380 ;
        RECT 786.670 276.180 787.910 276.320 ;
        RECT 786.670 276.120 786.990 276.180 ;
        RECT 787.590 276.120 787.910 276.180 ;
        RECT 787.130 193.360 787.450 193.420 ;
        RECT 788.050 193.360 788.370 193.420 ;
        RECT 787.130 193.220 788.370 193.360 ;
        RECT 787.130 193.160 787.450 193.220 ;
        RECT 788.050 193.160 788.370 193.220 ;
        RECT 737.910 20.980 738.230 21.040 ;
        RECT 737.910 20.840 745.500 20.980 ;
        RECT 737.910 20.780 738.230 20.840 ;
        RECT 234.670 20.640 234.990 20.700 ;
        RECT 372.670 20.640 372.990 20.700 ;
        RECT 234.670 20.500 372.990 20.640 ;
        RECT 234.670 20.440 234.990 20.500 ;
        RECT 372.670 20.440 372.990 20.500 ;
        RECT 420.510 20.640 420.830 20.700 ;
        RECT 469.270 20.640 469.590 20.700 ;
        RECT 420.510 20.500 469.590 20.640 ;
        RECT 420.510 20.440 420.830 20.500 ;
        RECT 469.270 20.440 469.590 20.500 ;
        RECT 517.110 20.640 517.430 20.700 ;
        RECT 565.870 20.640 566.190 20.700 ;
        RECT 517.110 20.500 566.190 20.640 ;
        RECT 517.110 20.440 517.430 20.500 ;
        RECT 565.870 20.440 566.190 20.500 ;
        RECT 617.390 20.640 617.710 20.700 ;
        RECT 665.690 20.640 666.010 20.700 ;
        RECT 617.390 20.500 666.010 20.640 ;
        RECT 617.390 20.440 617.710 20.500 ;
        RECT 665.690 20.440 666.010 20.500 ;
        RECT 745.360 20.300 745.500 20.840 ;
        RECT 786.670 20.300 786.990 20.360 ;
        RECT 745.360 20.160 786.990 20.300 ;
        RECT 786.670 20.100 786.990 20.160 ;
        RECT 372.670 15.880 372.990 15.940 ;
        RECT 420.510 15.880 420.830 15.940 ;
        RECT 372.670 15.740 420.830 15.880 ;
        RECT 372.670 15.680 372.990 15.740 ;
        RECT 420.510 15.680 420.830 15.740 ;
        RECT 469.270 14.860 469.590 14.920 ;
        RECT 517.110 14.860 517.430 14.920 ;
        RECT 469.270 14.720 517.430 14.860 ;
        RECT 469.270 14.660 469.590 14.720 ;
        RECT 517.110 14.660 517.430 14.720 ;
        RECT 565.870 14.520 566.190 14.580 ;
        RECT 617.390 14.520 617.710 14.580 ;
        RECT 565.870 14.380 617.710 14.520 ;
        RECT 565.870 14.320 566.190 14.380 ;
        RECT 617.390 14.320 617.710 14.380 ;
        RECT 665.690 14.520 666.010 14.580 ;
        RECT 737.910 14.520 738.230 14.580 ;
        RECT 665.690 14.380 738.230 14.520 ;
        RECT 665.690 14.320 666.010 14.380 ;
        RECT 737.910 14.320 738.230 14.380 ;
      LAYER via ;
        RECT 787.160 531.120 787.420 531.380 ;
        RECT 787.620 531.120 787.880 531.380 ;
        RECT 787.160 496.440 787.420 496.700 ;
        RECT 788.080 496.440 788.340 496.700 ;
        RECT 785.780 420.620 786.040 420.880 ;
        RECT 788.540 420.620 788.800 420.880 ;
        RECT 785.780 413.820 786.040 414.080 ;
        RECT 787.160 413.820 787.420 414.080 ;
        RECT 787.160 282.920 787.420 283.180 ;
        RECT 786.700 282.580 786.960 282.840 ;
        RECT 786.700 276.120 786.960 276.380 ;
        RECT 787.620 276.120 787.880 276.380 ;
        RECT 787.160 193.160 787.420 193.420 ;
        RECT 788.080 193.160 788.340 193.420 ;
        RECT 737.940 20.780 738.200 21.040 ;
        RECT 234.700 20.440 234.960 20.700 ;
        RECT 372.700 20.440 372.960 20.700 ;
        RECT 420.540 20.440 420.800 20.700 ;
        RECT 469.300 20.440 469.560 20.700 ;
        RECT 517.140 20.440 517.400 20.700 ;
        RECT 565.900 20.440 566.160 20.700 ;
        RECT 617.420 20.440 617.680 20.700 ;
        RECT 665.720 20.440 665.980 20.700 ;
        RECT 786.700 20.100 786.960 20.360 ;
        RECT 372.700 15.680 372.960 15.940 ;
        RECT 420.540 15.680 420.800 15.940 ;
        RECT 469.300 14.660 469.560 14.920 ;
        RECT 517.140 14.660 517.400 14.920 ;
        RECT 565.900 14.320 566.160 14.580 ;
        RECT 617.420 14.320 617.680 14.580 ;
        RECT 665.720 14.320 665.980 14.580 ;
        RECT 737.940 14.320 738.200 14.580 ;
      LAYER met2 ;
        RECT 790.610 600.170 790.890 604.000 ;
        RECT 789.520 600.030 790.890 600.170 ;
        RECT 789.520 579.885 789.660 600.030 ;
        RECT 790.610 600.000 790.890 600.030 ;
        RECT 787.610 579.515 787.890 579.885 ;
        RECT 789.450 579.515 789.730 579.885 ;
        RECT 787.680 531.410 787.820 579.515 ;
        RECT 787.160 531.090 787.420 531.410 ;
        RECT 787.620 531.090 787.880 531.410 ;
        RECT 787.220 496.730 787.360 531.090 ;
        RECT 787.160 496.410 787.420 496.730 ;
        RECT 788.080 496.410 788.340 496.730 ;
        RECT 788.140 483.210 788.280 496.410 ;
        RECT 788.140 483.070 788.740 483.210 ;
        RECT 788.600 420.910 788.740 483.070 ;
        RECT 785.780 420.590 786.040 420.910 ;
        RECT 788.540 420.590 788.800 420.910 ;
        RECT 785.840 414.110 785.980 420.590 ;
        RECT 785.780 413.790 786.040 414.110 ;
        RECT 787.160 413.790 787.420 414.110 ;
        RECT 787.220 283.210 787.360 413.790 ;
        RECT 787.160 282.890 787.420 283.210 ;
        RECT 786.700 282.550 786.960 282.870 ;
        RECT 786.760 276.410 786.900 282.550 ;
        RECT 786.700 276.090 786.960 276.410 ;
        RECT 787.620 276.090 787.880 276.410 ;
        RECT 787.680 254.730 787.820 276.090 ;
        RECT 787.220 254.590 787.820 254.730 ;
        RECT 787.220 193.450 787.360 254.590 ;
        RECT 787.160 193.130 787.420 193.450 ;
        RECT 788.080 193.130 788.340 193.450 ;
        RECT 788.140 110.570 788.280 193.130 ;
        RECT 787.680 110.430 788.280 110.570 ;
        RECT 787.680 62.290 787.820 110.430 ;
        RECT 786.760 62.150 787.820 62.290 ;
        RECT 737.940 20.750 738.200 21.070 ;
        RECT 234.700 20.410 234.960 20.730 ;
        RECT 372.700 20.410 372.960 20.730 ;
        RECT 420.540 20.410 420.800 20.730 ;
        RECT 469.300 20.410 469.560 20.730 ;
        RECT 517.140 20.410 517.400 20.730 ;
        RECT 565.900 20.410 566.160 20.730 ;
        RECT 617.420 20.410 617.680 20.730 ;
        RECT 665.720 20.410 665.980 20.730 ;
        RECT 234.760 2.400 234.900 20.410 ;
        RECT 372.760 15.970 372.900 20.410 ;
        RECT 420.600 15.970 420.740 20.410 ;
        RECT 372.700 15.650 372.960 15.970 ;
        RECT 420.540 15.650 420.800 15.970 ;
        RECT 469.360 14.950 469.500 20.410 ;
        RECT 517.200 14.950 517.340 20.410 ;
        RECT 469.300 14.630 469.560 14.950 ;
        RECT 517.140 14.630 517.400 14.950 ;
        RECT 565.960 14.610 566.100 20.410 ;
        RECT 617.480 14.610 617.620 20.410 ;
        RECT 665.780 14.610 665.920 20.410 ;
        RECT 738.000 14.610 738.140 20.750 ;
        RECT 786.760 20.390 786.900 62.150 ;
        RECT 786.700 20.070 786.960 20.390 ;
        RECT 565.900 14.290 566.160 14.610 ;
        RECT 617.420 14.290 617.680 14.610 ;
        RECT 665.720 14.290 665.980 14.610 ;
        RECT 737.940 14.290 738.200 14.610 ;
        RECT 234.550 -4.800 235.110 2.400 ;
      LAYER via2 ;
        RECT 787.610 579.560 787.890 579.840 ;
        RECT 789.450 579.560 789.730 579.840 ;
      LAYER met3 ;
        RECT 787.585 579.850 787.915 579.865 ;
        RECT 789.425 579.850 789.755 579.865 ;
        RECT 787.585 579.550 789.755 579.850 ;
        RECT 787.585 579.535 787.915 579.550 ;
        RECT 789.425 579.535 789.755 579.550 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 56.190 45.120 56.510 45.180 ;
        RECT 697.430 45.120 697.750 45.180 ;
        RECT 56.190 44.980 697.750 45.120 ;
        RECT 56.190 44.920 56.510 44.980 ;
        RECT 697.430 44.920 697.750 44.980 ;
      LAYER via ;
        RECT 56.220 44.920 56.480 45.180 ;
        RECT 697.460 44.920 697.720 45.180 ;
      LAYER met2 ;
        RECT 698.610 600.170 698.890 604.000 ;
        RECT 697.520 600.030 698.890 600.170 ;
        RECT 697.520 45.210 697.660 600.030 ;
        RECT 698.610 600.000 698.890 600.030 ;
        RECT 56.220 44.890 56.480 45.210 ;
        RECT 697.460 44.890 697.720 45.210 ;
        RECT 56.280 2.400 56.420 44.890 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 80.110 17.920 80.430 17.980 ;
        RECT 711.690 17.920 712.010 17.980 ;
        RECT 80.110 17.780 712.010 17.920 ;
        RECT 80.110 17.720 80.430 17.780 ;
        RECT 711.690 17.720 712.010 17.780 ;
      LAYER via ;
        RECT 80.140 17.720 80.400 17.980 ;
        RECT 711.720 17.720 711.980 17.980 ;
      LAYER met2 ;
        RECT 711.030 600.170 711.310 604.000 ;
        RECT 711.030 600.030 711.920 600.170 ;
        RECT 711.030 600.000 711.310 600.030 ;
        RECT 711.780 18.010 711.920 600.030 ;
        RECT 80.140 17.690 80.400 18.010 ;
        RECT 711.720 17.690 711.980 18.010 ;
        RECT 80.200 2.400 80.340 17.690 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 718.130 545.260 718.450 545.320 ;
        RECT 720.890 545.260 721.210 545.320 ;
        RECT 718.130 545.120 721.210 545.260 ;
        RECT 718.130 545.060 718.450 545.120 ;
        RECT 720.890 545.060 721.210 545.120 ;
        RECT 103.570 45.460 103.890 45.520 ;
        RECT 718.130 45.460 718.450 45.520 ;
        RECT 103.570 45.320 718.450 45.460 ;
        RECT 103.570 45.260 103.890 45.320 ;
        RECT 718.130 45.260 718.450 45.320 ;
      LAYER via ;
        RECT 718.160 545.060 718.420 545.320 ;
        RECT 720.920 545.060 721.180 545.320 ;
        RECT 103.600 45.260 103.860 45.520 ;
        RECT 718.160 45.260 718.420 45.520 ;
      LAYER met2 ;
        RECT 723.450 600.170 723.730 604.000 ;
        RECT 720.980 600.030 723.730 600.170 ;
        RECT 720.980 545.350 721.120 600.030 ;
        RECT 723.450 600.000 723.730 600.030 ;
        RECT 718.160 545.030 718.420 545.350 ;
        RECT 720.920 545.030 721.180 545.350 ;
        RECT 718.220 45.550 718.360 545.030 ;
        RECT 103.600 45.230 103.860 45.550 ;
        RECT 718.160 45.230 718.420 45.550 ;
        RECT 103.660 2.400 103.800 45.230 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 19.280 127.810 19.340 ;
        RECT 731.930 19.280 732.250 19.340 ;
        RECT 127.490 19.140 732.250 19.280 ;
        RECT 127.490 19.080 127.810 19.140 ;
        RECT 731.930 19.080 732.250 19.140 ;
      LAYER via ;
        RECT 127.520 19.080 127.780 19.340 ;
        RECT 731.960 19.080 732.220 19.340 ;
      LAYER met2 ;
        RECT 735.410 600.170 735.690 604.000 ;
        RECT 733.860 600.030 735.690 600.170 ;
        RECT 733.860 596.770 734.000 600.030 ;
        RECT 735.410 600.000 735.690 600.030 ;
        RECT 732.020 596.630 734.000 596.770 ;
        RECT 732.020 19.370 732.160 596.630 ;
        RECT 127.520 19.050 127.780 19.370 ;
        RECT 731.960 19.050 732.220 19.370 ;
        RECT 127.580 2.400 127.720 19.050 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 44.780 26.610 44.840 ;
        RECT 684.090 44.780 684.410 44.840 ;
        RECT 26.290 44.640 684.410 44.780 ;
        RECT 26.290 44.580 26.610 44.640 ;
        RECT 684.090 44.580 684.410 44.640 ;
      LAYER via ;
        RECT 26.320 44.580 26.580 44.840 ;
        RECT 684.120 44.580 684.380 44.840 ;
      LAYER met2 ;
        RECT 683.430 600.170 683.710 604.000 ;
        RECT 683.430 600.030 684.320 600.170 ;
        RECT 683.430 600.000 683.710 600.030 ;
        RECT 684.180 44.870 684.320 600.030 ;
        RECT 26.320 44.550 26.580 44.870 ;
        RECT 684.120 44.550 684.380 44.870 ;
        RECT 26.380 2.400 26.520 44.550 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 17.240 32.590 17.300 ;
        RECT 684.550 17.240 684.870 17.300 ;
        RECT 32.270 17.100 684.870 17.240 ;
        RECT 32.270 17.040 32.590 17.100 ;
        RECT 684.550 17.040 684.870 17.100 ;
      LAYER via ;
        RECT 32.300 17.040 32.560 17.300 ;
        RECT 684.580 17.040 684.840 17.300 ;
      LAYER met2 ;
        RECT 686.650 600.170 686.930 604.000 ;
        RECT 684.640 600.030 686.930 600.170 ;
        RECT 684.640 17.330 684.780 600.030 ;
        RECT 686.650 600.000 686.930 600.030 ;
        RECT 32.300 17.010 32.560 17.330 ;
        RECT 684.580 17.010 684.840 17.330 ;
        RECT 32.360 2.400 32.500 17.010 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 1982.750 367.020 3529.000 ;
        RECT 544.020 2760.520 547.020 3529.000 ;
        RECT 457.645 2610.640 459.245 2747.120 ;
        RECT 544.020 1982.750 547.020 2599.000 ;
        RECT 381.040 1710.640 382.640 1969.520 ;
        RECT 364.020 -9.320 367.020 1699.000 ;
        RECT 544.020 -9.320 547.020 1699.000 ;
        RECT 724.020 1001.000 727.020 3529.000 ;
        RECT 904.020 1001.000 907.020 3529.000 ;
        RECT 1084.020 2801.000 1087.020 3529.000 ;
        RECT 1019.545 2610.640 1021.145 2787.920 ;
        RECT 1084.020 2045.110 1087.020 2599.000 ;
        RECT 1264.020 2045.110 1267.020 3529.000 ;
        RECT 1021.040 1710.640 1022.640 2032.080 ;
        RECT 1084.020 1001.000 1087.020 1699.000 ;
        RECT 1264.020 1001.000 1267.020 1699.000 ;
        RECT 1444.020 1001.000 1447.020 3529.000 ;
        RECT 1624.020 2901.055 1627.020 3529.000 ;
        RECT 1804.020 2901.055 1807.020 3529.000 ;
        RECT 1521.040 2510.640 1522.640 2889.200 ;
        RECT 1624.020 1001.000 1627.020 2499.000 ;
        RECT 1804.020 1001.000 1807.020 2499.000 ;
        RECT 1984.020 1918.095 1987.020 3529.000 ;
        RECT 1948.870 1760.640 1950.470 1905.280 ;
        RECT 1984.020 1001.000 1987.020 1749.000 ;
        RECT 2164.020 1001.000 2167.020 3529.000 ;
        RECT 2344.020 1938.745 2347.020 3529.000 ;
        RECT 2524.020 2774.820 2527.020 3529.000 ;
        RECT 2427.190 2610.640 2428.790 2760.720 ;
        RECT 2524.020 1938.745 2527.020 2599.000 ;
        RECT 2321.040 1710.640 2322.640 1926.000 ;
        RECT 691.040 610.640 692.640 989.200 ;
        RECT 724.020 -9.320 727.020 599.000 ;
        RECT 904.020 -9.320 907.020 599.000 ;
        RECT 1084.020 -9.320 1087.020 599.000 ;
        RECT 1264.020 -9.320 1267.020 599.000 ;
        RECT 1444.020 -9.320 1447.020 599.000 ;
        RECT 1624.020 -9.320 1627.020 599.000 ;
        RECT 1804.020 -9.320 1807.020 599.000 ;
        RECT 1984.020 -9.320 1987.020 599.000 ;
        RECT 2164.020 -9.320 2167.020 599.000 ;
        RECT 2344.020 -9.320 2347.020 1699.000 ;
        RECT 2524.020 -9.320 2527.020 1699.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 457.855 2711.090 459.035 2712.270 ;
        RECT 457.855 2709.490 459.035 2710.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 381.250 1811.090 382.430 1812.270 ;
        RECT 381.250 1809.490 382.430 1810.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 1019.755 2711.090 1020.935 2712.270 ;
        RECT 1019.755 2709.490 1020.935 2710.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1521.250 2711.090 1522.430 2712.270 ;
        RECT 1521.250 2709.490 1522.430 2710.670 ;
        RECT 1521.250 2531.090 1522.430 2532.270 ;
        RECT 1521.250 2529.490 1522.430 2530.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 1021.250 1991.090 1022.430 1992.270 ;
        RECT 1021.250 1989.490 1022.430 1990.670 ;
        RECT 1021.250 1811.090 1022.430 1812.270 ;
        RECT 1021.250 1809.490 1022.430 1810.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1949.080 1811.090 1950.260 1812.270 ;
        RECT 1949.080 1809.490 1950.260 1810.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2427.400 2711.090 2428.580 2712.270 ;
        RECT 2427.400 2709.490 2428.580 2710.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 2321.250 1811.090 2322.430 1812.270 ;
        RECT 2321.250 1809.490 2322.430 1810.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 691.250 911.090 692.430 912.270 ;
        RECT 691.250 909.490 692.430 910.670 ;
        RECT 691.250 731.090 692.430 732.270 ;
        RECT 691.250 729.490 692.430 730.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 457.645 2712.380 459.245 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1019.545 2712.380 1021.145 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1521.040 2712.380 1522.640 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2427.190 2712.380 2428.790 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 457.645 2709.370 459.245 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1019.545 2709.370 1021.145 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1521.040 2709.370 1522.640 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2427.190 2709.370 2428.790 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1521.040 2532.380 1522.640 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1521.040 2529.370 1522.640 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1021.040 1992.380 1022.640 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1021.040 1989.370 1022.640 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 381.040 1812.380 382.640 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1021.040 1812.380 1022.640 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1948.870 1812.380 1950.470 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2321.040 1812.380 2322.640 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 381.040 1809.370 382.640 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1021.040 1809.370 1022.640 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1948.870 1809.370 1950.470 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2321.040 1809.370 2322.640 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 691.040 912.380 692.640 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 691.040 909.370 692.640 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 691.040 732.380 692.640 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 691.040 729.370 692.640 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 2760.520 457.020 3529.000 ;
        RECT 480.565 2610.640 482.165 2747.120 ;
        RECT 454.020 1982.750 457.020 2599.000 ;
        RECT 457.840 1710.640 459.440 1969.520 ;
        RECT 454.020 -9.320 457.020 1699.000 ;
        RECT 634.020 -9.320 637.020 3529.000 ;
        RECT 814.020 1001.000 817.020 3529.000 ;
        RECT 994.020 1001.000 997.020 3529.000 ;
        RECT 1034.375 2610.640 1035.975 2787.920 ;
        RECT 1174.020 2045.110 1177.020 3529.000 ;
        RECT 1097.840 1710.640 1099.440 2032.080 ;
        RECT 1174.020 1001.000 1177.020 1699.000 ;
        RECT 1354.020 1001.000 1357.020 3529.000 ;
        RECT 1534.020 2901.055 1537.020 3529.000 ;
        RECT 1714.020 2901.055 1717.020 3529.000 ;
        RECT 1597.840 2510.640 1599.440 2889.200 ;
        RECT 1534.020 1001.000 1537.020 2499.000 ;
        RECT 1714.020 1001.000 1717.020 2499.000 ;
        RECT 1894.020 1001.000 1897.020 3529.000 ;
        RECT 2074.020 1918.095 2077.020 3529.000 ;
        RECT 1973.020 1760.640 1974.620 1905.280 ;
        RECT 2074.020 1001.000 2077.020 1749.000 ;
        RECT 767.840 610.640 769.440 989.200 ;
        RECT 814.020 -9.320 817.020 599.000 ;
        RECT 994.020 -9.320 997.020 599.000 ;
        RECT 1174.020 -9.320 1177.020 599.000 ;
        RECT 1354.020 -9.320 1357.020 599.000 ;
        RECT 1534.020 -9.320 1537.020 599.000 ;
        RECT 1714.020 -9.320 1717.020 599.000 ;
        RECT 1894.020 -9.320 1897.020 599.000 ;
        RECT 2074.020 -9.320 2077.020 599.000 ;
        RECT 2254.020 -9.320 2257.020 3529.000 ;
        RECT 2434.020 2774.820 2437.020 3529.000 ;
        RECT 2452.490 2610.640 2454.090 2760.720 ;
        RECT 2434.020 1938.745 2437.020 2599.000 ;
        RECT 2397.840 1710.640 2399.440 1926.000 ;
        RECT 2434.020 -9.320 2437.020 1699.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 480.775 2621.090 481.955 2622.270 ;
        RECT 480.775 2619.490 481.955 2620.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 458.050 1901.090 459.230 1902.270 ;
        RECT 458.050 1899.490 459.230 1900.670 ;
        RECT 458.050 1721.090 459.230 1722.270 ;
        RECT 458.050 1719.490 459.230 1720.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 1034.585 2621.090 1035.765 2622.270 ;
        RECT 1034.585 2619.490 1035.765 2620.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1598.050 2801.090 1599.230 2802.270 ;
        RECT 1598.050 2799.490 1599.230 2800.670 ;
        RECT 1598.050 2621.090 1599.230 2622.270 ;
        RECT 1598.050 2619.490 1599.230 2620.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 1098.050 1901.090 1099.230 1902.270 ;
        RECT 1098.050 1899.490 1099.230 1900.670 ;
        RECT 1098.050 1721.090 1099.230 1722.270 ;
        RECT 1098.050 1719.490 1099.230 1720.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2452.700 2621.090 2453.880 2622.270 ;
        RECT 2452.700 2619.490 2453.880 2620.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1973.230 1901.090 1974.410 1902.270 ;
        RECT 1973.230 1899.490 1974.410 1900.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2398.050 1901.090 2399.230 1902.270 ;
        RECT 2398.050 1899.490 2399.230 1900.670 ;
        RECT 2398.050 1721.090 2399.230 1722.270 ;
        RECT 2398.050 1719.490 2399.230 1720.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 768.050 821.090 769.230 822.270 ;
        RECT 768.050 819.490 769.230 820.670 ;
        RECT 768.050 641.090 769.230 642.270 ;
        RECT 768.050 639.490 769.230 640.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1597.840 2802.380 1599.440 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1597.840 2799.370 1599.440 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 480.565 2622.380 482.165 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1034.375 2622.380 1035.975 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1597.840 2622.380 1599.440 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2452.490 2622.380 2454.090 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 480.565 2619.370 482.165 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1034.375 2619.370 1035.975 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1597.840 2619.370 1599.440 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2452.490 2619.370 2454.090 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 457.840 1902.380 459.440 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1097.840 1902.380 1099.440 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 1973.020 1902.380 1974.620 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2397.840 1902.380 2399.440 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 457.840 1899.370 459.440 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1097.840 1899.370 1099.440 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 1973.020 1899.370 1974.620 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2397.840 1899.370 2399.440 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 457.840 1722.380 459.440 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1097.840 1722.380 1099.440 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2397.840 1722.380 2399.440 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 457.840 1719.370 459.440 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1097.840 1719.370 1099.440 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2397.840 1719.370 2399.440 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 767.840 822.380 769.440 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 767.840 819.370 769.440 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 767.840 642.380 769.440 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 767.840 639.370 769.440 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 382.020 1982.750 385.020 3538.400 ;
        RECT 562.020 2760.520 565.020 3538.400 ;
        RECT 562.020 1982.750 565.020 2599.000 ;
        RECT 382.020 -18.720 385.020 1699.000 ;
        RECT 562.020 -18.720 565.020 1699.000 ;
        RECT 742.020 1001.000 745.020 3538.400 ;
        RECT 922.020 1001.000 925.020 3538.400 ;
        RECT 1102.020 2045.110 1105.020 3538.400 ;
        RECT 1282.020 2045.110 1285.020 3538.400 ;
        RECT 1102.020 1001.000 1105.020 1699.000 ;
        RECT 1282.020 1001.000 1285.020 1699.000 ;
        RECT 1462.020 1001.000 1465.020 3538.400 ;
        RECT 1642.020 2901.055 1645.020 3538.400 ;
        RECT 1822.020 2901.055 1825.020 3538.400 ;
        RECT 1642.020 1001.000 1645.020 2499.000 ;
        RECT 1822.020 1001.000 1825.020 2499.000 ;
        RECT 2002.020 1918.095 2005.020 3538.400 ;
        RECT 2002.020 1001.000 2005.020 1749.000 ;
        RECT 742.020 -18.720 745.020 599.000 ;
        RECT 922.020 -18.720 925.020 599.000 ;
        RECT 1102.020 -18.720 1105.020 599.000 ;
        RECT 1282.020 -18.720 1285.020 599.000 ;
        RECT 1462.020 -18.720 1465.020 599.000 ;
        RECT 1642.020 -18.720 1645.020 599.000 ;
        RECT 1822.020 -18.720 1825.020 599.000 ;
        RECT 2002.020 -18.720 2005.020 599.000 ;
        RECT 2182.020 -18.720 2185.020 3538.400 ;
        RECT 2362.020 1938.745 2365.020 3538.400 ;
        RECT 2542.020 2774.820 2545.020 3538.400 ;
        RECT 2362.020 -18.720 2365.020 1699.000 ;
        RECT 2542.020 -18.720 2545.020 2599.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 292.020 -18.720 295.020 3538.400 ;
        RECT 472.020 2760.520 475.020 3538.400 ;
        RECT 472.020 1982.750 475.020 2599.000 ;
        RECT 472.020 -18.720 475.020 1699.000 ;
        RECT 652.020 -18.720 655.020 3538.400 ;
        RECT 832.020 1001.000 835.020 3538.400 ;
        RECT 1012.020 2801.000 1015.020 3538.400 ;
        RECT 1012.020 2045.110 1015.020 2599.000 ;
        RECT 1192.020 2045.110 1195.020 3538.400 ;
        RECT 1012.020 1001.000 1015.020 1699.000 ;
        RECT 1192.020 1001.000 1195.020 1699.000 ;
        RECT 1372.020 1001.000 1375.020 3538.400 ;
        RECT 1552.020 2901.055 1555.020 3538.400 ;
        RECT 1732.020 2901.055 1735.020 3538.400 ;
        RECT 1552.020 1001.000 1555.020 2499.000 ;
        RECT 1732.020 1001.000 1735.020 2499.000 ;
        RECT 1912.020 1001.000 1915.020 3538.400 ;
        RECT 2092.020 1001.000 2095.020 3538.400 ;
        RECT 832.020 -18.720 835.020 599.000 ;
        RECT 1012.020 -18.720 1015.020 599.000 ;
        RECT 1192.020 -18.720 1195.020 599.000 ;
        RECT 1372.020 -18.720 1375.020 599.000 ;
        RECT 1552.020 -18.720 1555.020 599.000 ;
        RECT 1732.020 -18.720 1735.020 599.000 ;
        RECT 1912.020 -18.720 1915.020 599.000 ;
        RECT 2092.020 -18.720 2095.020 599.000 ;
        RECT 2272.020 -18.720 2275.020 3538.400 ;
        RECT 2452.020 2774.820 2455.020 3538.400 ;
        RECT 2452.020 1938.745 2455.020 2599.000 ;
        RECT 2452.020 -18.720 2455.020 1699.000 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 400.020 1982.750 403.020 3547.800 ;
        RECT 580.020 1982.750 583.020 3547.800 ;
        RECT 400.020 -28.120 403.020 1699.000 ;
        RECT 580.020 -28.120 583.020 1699.000 ;
        RECT 760.020 1001.000 763.020 3547.800 ;
        RECT 940.020 1001.000 943.020 3547.800 ;
        RECT 1120.020 2045.110 1123.020 3547.800 ;
        RECT 1300.020 2045.110 1303.020 3547.800 ;
        RECT 1120.020 1001.000 1123.020 1699.000 ;
        RECT 1300.020 1001.000 1303.020 1699.000 ;
        RECT 1480.020 1001.000 1483.020 3547.800 ;
        RECT 1660.020 2901.055 1663.020 3547.800 ;
        RECT 1840.020 2901.055 1843.020 3547.800 ;
        RECT 1660.020 1001.000 1663.020 2499.000 ;
        RECT 1840.020 1001.000 1843.020 2499.000 ;
        RECT 2020.020 1918.095 2023.020 3547.800 ;
        RECT 2020.020 1001.000 2023.020 1749.000 ;
        RECT 760.020 -28.120 763.020 599.000 ;
        RECT 940.020 -28.120 943.020 599.000 ;
        RECT 1120.020 -28.120 1123.020 599.000 ;
        RECT 1300.020 -28.120 1303.020 599.000 ;
        RECT 1480.020 -28.120 1483.020 599.000 ;
        RECT 1660.020 -28.120 1663.020 599.000 ;
        RECT 1840.020 -28.120 1843.020 599.000 ;
        RECT 2020.020 -28.120 2023.020 599.000 ;
        RECT 2200.020 -28.120 2203.020 3547.800 ;
        RECT 2380.020 1938.745 2383.020 3547.800 ;
        RECT 2380.020 -28.120 2383.020 1699.000 ;
        RECT 2560.020 -28.120 2563.020 3547.800 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 310.020 -28.120 313.020 3547.800 ;
        RECT 490.020 2760.520 493.020 3547.800 ;
        RECT 490.020 1982.750 493.020 2599.000 ;
        RECT 490.020 -28.120 493.020 1699.000 ;
        RECT 670.020 1001.000 673.020 3547.800 ;
        RECT 850.020 1001.000 853.020 3547.800 ;
        RECT 1030.020 2801.000 1033.020 3547.800 ;
        RECT 1030.020 2045.110 1033.020 2599.000 ;
        RECT 1210.020 2045.110 1213.020 3547.800 ;
        RECT 1030.020 1001.000 1033.020 1699.000 ;
        RECT 1210.020 1001.000 1213.020 1699.000 ;
        RECT 1390.020 1001.000 1393.020 3547.800 ;
        RECT 1570.020 2901.055 1573.020 3547.800 ;
        RECT 1750.020 2901.055 1753.020 3547.800 ;
        RECT 1570.020 1001.000 1573.020 2499.000 ;
        RECT 1750.020 1001.000 1753.020 2499.000 ;
        RECT 1930.020 1918.095 1933.020 3547.800 ;
        RECT 1930.020 1001.000 1933.020 1749.000 ;
        RECT 2110.020 1001.000 2113.020 3547.800 ;
        RECT 670.020 -28.120 673.020 599.000 ;
        RECT 850.020 -28.120 853.020 599.000 ;
        RECT 1030.020 -28.120 1033.020 599.000 ;
        RECT 1210.020 -28.120 1213.020 599.000 ;
        RECT 1390.020 -28.120 1393.020 599.000 ;
        RECT 1570.020 -28.120 1573.020 599.000 ;
        RECT 1750.020 -28.120 1753.020 599.000 ;
        RECT 1930.020 -28.120 1933.020 599.000 ;
        RECT 2110.020 -28.120 2113.020 599.000 ;
        RECT 2290.020 -28.120 2293.020 3547.800 ;
        RECT 2470.020 2774.820 2473.020 3547.800 ;
        RECT 2470.020 1938.745 2473.020 2599.000 ;
        RECT 2470.020 -28.120 2473.020 1699.000 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 418.020 1982.750 421.020 3557.200 ;
        RECT 598.020 1982.750 601.020 3557.200 ;
        RECT 418.020 -37.520 421.020 1699.000 ;
        RECT 598.020 -37.520 601.020 1699.000 ;
        RECT 778.020 1001.000 781.020 3557.200 ;
        RECT 958.020 1001.000 961.020 3557.200 ;
        RECT 1138.020 2045.110 1141.020 3557.200 ;
        RECT 1318.020 2045.110 1321.020 3557.200 ;
        RECT 1498.020 2901.055 1501.020 3557.200 ;
        RECT 1678.020 2901.055 1681.020 3557.200 ;
        RECT 1858.020 2901.055 1861.020 3557.200 ;
        RECT 1138.020 1001.000 1141.020 1699.000 ;
        RECT 1318.020 1001.000 1321.020 1699.000 ;
        RECT 1498.020 1001.000 1501.020 2499.000 ;
        RECT 1678.020 1001.000 1681.020 2499.000 ;
        RECT 1858.020 1001.000 1861.020 2499.000 ;
        RECT 2038.020 1918.095 2041.020 3557.200 ;
        RECT 2038.020 1001.000 2041.020 1749.000 ;
        RECT 778.020 -37.520 781.020 599.000 ;
        RECT 958.020 -37.520 961.020 599.000 ;
        RECT 1138.020 -37.520 1141.020 599.000 ;
        RECT 1318.020 -37.520 1321.020 599.000 ;
        RECT 1498.020 -37.520 1501.020 599.000 ;
        RECT 1678.020 -37.520 1681.020 599.000 ;
        RECT 1858.020 -37.520 1861.020 599.000 ;
        RECT 2038.020 -37.520 2041.020 599.000 ;
        RECT 2218.020 -37.520 2221.020 3557.200 ;
        RECT 2398.020 2774.820 2401.020 3557.200 ;
        RECT 2398.020 1938.745 2401.020 2599.000 ;
        RECT 2398.020 -37.520 2401.020 1699.000 ;
        RECT 2578.020 -37.520 2581.020 3557.200 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 328.020 -37.520 331.020 3557.200 ;
        RECT 508.020 2760.520 511.020 3557.200 ;
        RECT 508.020 1982.750 511.020 2599.000 ;
        RECT 508.020 -37.520 511.020 1699.000 ;
        RECT 688.020 1001.000 691.020 3557.200 ;
        RECT 868.020 1001.000 871.020 3557.200 ;
        RECT 1048.020 2801.000 1051.020 3557.200 ;
        RECT 1048.020 2045.110 1051.020 2599.000 ;
        RECT 1228.020 2045.110 1231.020 3557.200 ;
        RECT 1048.020 1001.000 1051.020 1699.000 ;
        RECT 1228.020 1001.000 1231.020 1699.000 ;
        RECT 1408.020 1001.000 1411.020 3557.200 ;
        RECT 1588.020 2901.055 1591.020 3557.200 ;
        RECT 1768.020 2901.055 1771.020 3557.200 ;
        RECT 1588.020 1001.000 1591.020 2499.000 ;
        RECT 1768.020 1001.000 1771.020 2499.000 ;
        RECT 1948.020 1918.095 1951.020 3557.200 ;
        RECT 1948.020 1001.000 1951.020 1749.000 ;
        RECT 2128.020 1001.000 2131.020 3557.200 ;
        RECT 2308.020 1938.745 2311.020 3557.200 ;
        RECT 2488.020 2774.820 2491.020 3557.200 ;
        RECT 2488.020 1938.745 2491.020 2599.000 ;
        RECT 688.020 -37.520 691.020 599.000 ;
        RECT 868.020 -37.520 871.020 599.000 ;
        RECT 1048.020 -37.520 1051.020 599.000 ;
        RECT 1228.020 -37.520 1231.020 599.000 ;
        RECT 1408.020 -37.520 1411.020 599.000 ;
        RECT 1588.020 -37.520 1591.020 599.000 ;
        RECT 1768.020 -37.520 1771.020 599.000 ;
        RECT 1948.020 -37.520 1951.020 599.000 ;
        RECT 2128.020 -37.520 2131.020 599.000 ;
        RECT 2308.020 -37.520 2311.020 1699.000 ;
        RECT 2488.020 -37.520 2491.020 1699.000 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 435.520 2610.795 573.060 2746.965 ;
        RECT 1005.520 2610.795 1094.300 2787.765 ;
        RECT 1505.520 2510.795 1883.640 2889.045 ;
        RECT 2402.690 2610.795 2554.490 2760.565 ;
        RECT 365.520 1710.795 625.420 1969.365 ;
        RECT 1005.520 1710.795 1327.520 2031.925 ;
        RECT 1925.520 1760.795 2070.420 1905.125 ;
        RECT 2305.520 1710.795 2521.260 1925.845 ;
        RECT 675.520 610.795 2164.080 998.055 ;
      LAYER met1 ;
        RECT 1352.010 2918.120 1352.330 2918.180 ;
        RECT 1535.090 2918.120 1535.410 2918.180 ;
        RECT 1352.010 2917.980 1535.410 2918.120 ;
        RECT 1352.010 2917.920 1352.330 2917.980 ;
        RECT 1535.090 2917.920 1535.410 2917.980 ;
        RECT 1431.590 2917.780 1431.910 2917.840 ;
        RECT 1598.570 2917.780 1598.890 2917.840 ;
        RECT 1431.590 2917.640 1598.890 2917.780 ;
        RECT 1431.590 2917.580 1431.910 2917.640 ;
        RECT 1598.570 2917.580 1598.890 2917.640 ;
        RECT 1459.190 2916.080 1459.510 2916.140 ;
        RECT 1641.810 2916.080 1642.130 2916.140 ;
        RECT 1459.190 2915.940 1642.130 2916.080 ;
        RECT 1459.190 2915.880 1459.510 2915.940 ;
        RECT 1641.810 2915.880 1642.130 2915.940 ;
        RECT 1494.610 2915.740 1494.930 2915.800 ;
        RECT 1705.290 2915.740 1705.610 2915.800 ;
        RECT 1494.610 2915.600 1705.610 2915.740 ;
        RECT 1494.610 2915.540 1494.930 2915.600 ;
        RECT 1705.290 2915.540 1705.610 2915.600 ;
        RECT 1472.990 2915.400 1473.310 2915.460 ;
        RECT 1694.250 2915.400 1694.570 2915.460 ;
        RECT 1472.990 2915.260 1694.570 2915.400 ;
        RECT 1472.990 2915.200 1473.310 2915.260 ;
        RECT 1694.250 2915.200 1694.570 2915.260 ;
        RECT 1406.750 2915.060 1407.070 2915.120 ;
        RECT 1630.770 2915.060 1631.090 2915.120 ;
        RECT 1406.750 2914.920 1631.090 2915.060 ;
        RECT 1406.750 2914.860 1407.070 2914.920 ;
        RECT 1630.770 2914.860 1631.090 2914.920 ;
        RECT 1495.070 2914.720 1495.390 2914.780 ;
        RECT 1768.770 2914.720 1769.090 2914.780 ;
        RECT 1495.070 2914.580 1769.090 2914.720 ;
        RECT 1495.070 2914.520 1495.390 2914.580 ;
        RECT 1768.770 2914.520 1769.090 2914.580 ;
        RECT 1493.230 2914.380 1493.550 2914.440 ;
        RECT 1779.810 2914.380 1780.130 2914.440 ;
        RECT 1493.230 2914.240 1780.130 2914.380 ;
        RECT 1493.230 2914.180 1493.550 2914.240 ;
        RECT 1779.810 2914.180 1780.130 2914.240 ;
        RECT 1455.510 2914.040 1455.830 2914.100 ;
        RECT 1758.650 2914.040 1758.970 2914.100 ;
        RECT 1455.510 2913.900 1758.970 2914.040 ;
        RECT 1455.510 2913.840 1455.830 2913.900 ;
        RECT 1758.650 2913.840 1758.970 2913.900 ;
        RECT 1493.690 2913.700 1494.010 2913.760 ;
        RECT 1800.970 2913.700 1801.290 2913.760 ;
        RECT 1493.690 2913.560 1801.290 2913.700 ;
        RECT 1493.690 2913.500 1494.010 2913.560 ;
        RECT 1800.970 2913.500 1801.290 2913.560 ;
        RECT 1500.590 2913.360 1500.910 2913.420 ;
        RECT 1812.010 2913.360 1812.330 2913.420 ;
        RECT 1500.590 2913.220 1812.330 2913.360 ;
        RECT 1500.590 2913.160 1500.910 2913.220 ;
        RECT 1812.010 2913.160 1812.330 2913.220 ;
        RECT 1833.170 2913.360 1833.490 2913.420 ;
        RECT 1894.350 2913.360 1894.670 2913.420 ;
        RECT 1833.170 2913.220 1894.670 2913.360 ;
        RECT 1833.170 2913.160 1833.490 2913.220 ;
        RECT 1894.350 2913.160 1894.670 2913.220 ;
        RECT 1494.150 2913.020 1494.470 2913.080 ;
        RECT 1662.970 2913.020 1663.290 2913.080 ;
        RECT 1494.150 2912.880 1663.290 2913.020 ;
        RECT 1494.150 2912.820 1494.470 2912.880 ;
        RECT 1662.970 2912.820 1663.290 2912.880 ;
        RECT 1789.930 2913.020 1790.250 2913.080 ;
        RECT 1892.050 2913.020 1892.370 2913.080 ;
        RECT 1789.930 2912.880 1892.370 2913.020 ;
        RECT 1789.930 2912.820 1790.250 2912.880 ;
        RECT 1892.050 2912.820 1892.370 2912.880 ;
        RECT 1492.310 2912.680 1492.630 2912.740 ;
        RECT 1609.610 2912.680 1609.930 2912.740 ;
        RECT 1492.310 2912.540 1609.930 2912.680 ;
        RECT 1492.310 2912.480 1492.630 2912.540 ;
        RECT 1609.610 2912.480 1609.930 2912.540 ;
        RECT 1854.330 2912.680 1854.650 2912.740 ;
        RECT 1893.430 2912.680 1893.750 2912.740 ;
        RECT 1854.330 2912.540 1893.750 2912.680 ;
        RECT 1854.330 2912.480 1854.650 2912.540 ;
        RECT 1893.430 2912.480 1893.750 2912.540 ;
        RECT 1438.490 2912.340 1438.810 2912.400 ;
        RECT 1567.290 2912.340 1567.610 2912.400 ;
        RECT 1438.490 2912.200 1567.610 2912.340 ;
        RECT 1438.490 2912.140 1438.810 2912.200 ;
        RECT 1567.290 2912.140 1567.610 2912.200 ;
        RECT 1492.770 2912.000 1493.090 2912.060 ;
        RECT 1546.130 2912.000 1546.450 2912.060 ;
        RECT 1492.770 2911.860 1546.450 2912.000 ;
        RECT 1492.770 2911.800 1493.090 2911.860 ;
        RECT 1546.130 2911.800 1546.450 2911.860 ;
        RECT 1864.450 2912.000 1864.770 2912.060 ;
        RECT 1892.970 2912.000 1893.290 2912.060 ;
        RECT 1864.450 2911.860 1893.290 2912.000 ;
        RECT 1864.450 2911.800 1864.770 2911.860 ;
        RECT 1892.970 2911.800 1893.290 2911.860 ;
        RECT 1496.910 2898.400 1497.230 2898.460 ;
        RECT 1524.050 2898.400 1524.370 2898.460 ;
        RECT 1496.910 2898.260 1524.370 2898.400 ;
        RECT 1496.910 2898.200 1497.230 2898.260 ;
        RECT 1524.050 2898.200 1524.370 2898.260 ;
        RECT 1497.370 2896.700 1497.690 2896.760 ;
        RECT 1503.350 2896.700 1503.670 2896.760 ;
        RECT 1497.370 2896.560 1503.670 2896.700 ;
        RECT 1497.370 2896.500 1497.690 2896.560 ;
        RECT 1503.350 2896.500 1503.670 2896.560 ;
        RECT 1876.870 2896.700 1877.190 2896.760 ;
        RECT 1892.510 2896.700 1892.830 2896.760 ;
        RECT 1876.870 2896.560 1892.830 2896.700 ;
        RECT 1876.870 2896.500 1877.190 2896.560 ;
        RECT 1892.510 2896.500 1892.830 2896.560 ;
        RECT 1362.590 2849.780 1362.910 2849.840 ;
        RECT 1483.570 2849.780 1483.890 2849.840 ;
        RECT 1362.590 2849.640 1483.890 2849.780 ;
        RECT 1362.590 2849.580 1362.910 2849.640 ;
        RECT 1483.570 2849.580 1483.890 2849.640 ;
        RECT 1501.510 2842.980 1501.830 2843.040 ;
        RECT 1501.970 2842.980 1502.290 2843.040 ;
        RECT 1501.510 2842.840 1502.290 2842.980 ;
        RECT 1501.510 2842.780 1501.830 2842.840 ;
        RECT 1501.970 2842.780 1502.290 2842.840 ;
        RECT 1501.510 2815.920 1501.830 2816.180 ;
        RECT 1501.600 2815.500 1501.740 2815.920 ;
        RECT 1501.510 2815.240 1501.830 2815.500 ;
        RECT 979.410 2810.340 979.730 2810.400 ;
        RECT 979.410 2810.200 1044.500 2810.340 ;
        RECT 979.410 2810.140 979.730 2810.200 ;
        RECT 985.390 2809.660 985.710 2809.720 ;
        RECT 1043.350 2809.660 1043.670 2809.720 ;
        RECT 985.390 2809.520 1043.670 2809.660 ;
        RECT 1044.360 2809.660 1044.500 2810.200 ;
        RECT 1089.350 2809.660 1089.670 2809.720 ;
        RECT 1044.360 2809.520 1089.670 2809.660 ;
        RECT 985.390 2809.460 985.710 2809.520 ;
        RECT 1043.350 2809.460 1043.670 2809.520 ;
        RECT 1089.350 2809.460 1089.670 2809.520 ;
        RECT 984.930 2809.320 985.250 2809.380 ;
        RECT 1027.710 2809.320 1028.030 2809.380 ;
        RECT 984.930 2809.180 1028.030 2809.320 ;
        RECT 984.930 2809.120 985.250 2809.180 ;
        RECT 1027.710 2809.120 1028.030 2809.180 ;
        RECT 986.310 2808.980 986.630 2809.040 ;
        RECT 1073.710 2808.980 1074.030 2809.040 ;
        RECT 986.310 2808.840 1074.030 2808.980 ;
        RECT 986.310 2808.780 986.630 2808.840 ;
        RECT 1073.710 2808.780 1074.030 2808.840 ;
        RECT 985.850 2808.640 986.170 2808.700 ;
        RECT 1012.070 2808.640 1012.390 2808.700 ;
        RECT 985.850 2808.500 1012.390 2808.640 ;
        RECT 985.850 2808.440 986.170 2808.500 ;
        RECT 1012.070 2808.440 1012.390 2808.500 ;
        RECT 1501.510 2794.700 1501.830 2794.760 ;
        RECT 1501.970 2794.700 1502.290 2794.760 ;
        RECT 1501.510 2794.560 1502.290 2794.700 ;
        RECT 1501.510 2794.500 1501.830 2794.560 ;
        RECT 1501.970 2794.500 1502.290 2794.560 ;
        RECT 445.810 2769.540 446.130 2769.600 ;
        RECT 810.590 2769.540 810.910 2769.600 ;
        RECT 445.810 2769.400 810.910 2769.540 ;
        RECT 445.810 2769.340 446.130 2769.400 ;
        RECT 810.590 2769.340 810.910 2769.400 ;
        RECT 532.290 2768.180 532.610 2768.240 ;
        RECT 700.190 2768.180 700.510 2768.240 ;
        RECT 532.290 2768.040 700.510 2768.180 ;
        RECT 532.290 2767.980 532.610 2768.040 ;
        RECT 700.190 2767.980 700.510 2768.040 ;
        RECT 518.490 2767.840 518.810 2767.900 ;
        RECT 755.390 2767.840 755.710 2767.900 ;
        RECT 518.490 2767.700 755.710 2767.840 ;
        RECT 518.490 2767.640 518.810 2767.700 ;
        RECT 755.390 2767.640 755.710 2767.700 ;
        RECT 489.050 2767.500 489.370 2767.560 ;
        RECT 789.890 2767.500 790.210 2767.560 ;
        RECT 489.050 2767.360 790.210 2767.500 ;
        RECT 489.050 2767.300 489.370 2767.360 ;
        RECT 789.890 2767.300 790.210 2767.360 ;
      LAYER met1 ;
        RECT 432.830 2606.500 575.750 2747.120 ;
      LAYER met1 ;
        RECT 586.570 2684.200 586.890 2684.260 ;
        RECT 734.690 2684.200 735.010 2684.260 ;
        RECT 586.570 2684.060 735.010 2684.200 ;
        RECT 586.570 2684.000 586.890 2684.060 ;
        RECT 734.690 2684.000 735.010 2684.060 ;
        RECT 586.570 2663.800 586.890 2663.860 ;
        RECT 803.690 2663.800 804.010 2663.860 ;
        RECT 586.570 2663.660 804.010 2663.800 ;
        RECT 586.570 2663.600 586.890 2663.660 ;
        RECT 803.690 2663.600 804.010 2663.660 ;
      LAYER met1 ;
        RECT 1002.830 2610.640 1095.150 2787.920 ;
      LAYER met1 ;
        RECT 1365.810 2781.100 1366.130 2781.160 ;
        RECT 1485.410 2781.100 1485.730 2781.160 ;
        RECT 1365.810 2780.960 1485.730 2781.100 ;
        RECT 1365.810 2780.900 1366.130 2780.960 ;
        RECT 1485.410 2780.900 1485.730 2780.960 ;
        RECT 1501.970 2766.960 1502.290 2767.220 ;
        RECT 1502.060 2766.540 1502.200 2766.960 ;
        RECT 1501.970 2766.280 1502.290 2766.540 ;
        RECT 1501.510 2753.220 1501.830 2753.280 ;
        RECT 1501.970 2753.220 1502.290 2753.280 ;
        RECT 1501.510 2753.080 1502.290 2753.220 ;
        RECT 1501.510 2753.020 1501.830 2753.080 ;
        RECT 1501.970 2753.020 1502.290 2753.080 ;
        RECT 1501.510 2719.020 1501.830 2719.280 ;
        RECT 1501.600 2718.600 1501.740 2719.020 ;
        RECT 1501.510 2718.340 1501.830 2718.600 ;
        RECT 1434.350 2691.340 1434.670 2691.400 ;
        RECT 1488.630 2691.340 1488.950 2691.400 ;
        RECT 1434.350 2691.200 1488.950 2691.340 ;
        RECT 1434.350 2691.140 1434.670 2691.200 ;
        RECT 1488.630 2691.140 1488.950 2691.200 ;
        RECT 1501.510 2670.600 1501.830 2670.660 ;
        RECT 1501.510 2670.460 1502.200 2670.600 ;
        RECT 1501.510 2670.400 1501.830 2670.460 ;
        RECT 1502.060 2670.320 1502.200 2670.460 ;
        RECT 1501.970 2670.060 1502.290 2670.320 ;
        RECT 1501.510 2656.660 1501.830 2656.720 ;
        RECT 1501.970 2656.660 1502.290 2656.720 ;
        RECT 1501.510 2656.520 1502.290 2656.660 ;
        RECT 1501.510 2656.460 1501.830 2656.520 ;
        RECT 1501.970 2656.460 1502.290 2656.520 ;
        RECT 1501.510 2622.460 1501.830 2622.720 ;
        RECT 1501.600 2622.040 1501.740 2622.460 ;
        RECT 1501.510 2621.780 1501.830 2622.040 ;
        RECT 1400.310 2608.380 1400.630 2608.440 ;
        RECT 1485.410 2608.380 1485.730 2608.440 ;
        RECT 1400.310 2608.240 1485.730 2608.380 ;
        RECT 1400.310 2608.180 1400.630 2608.240 ;
        RECT 1485.410 2608.180 1485.730 2608.240 ;
        RECT 996.890 2605.660 997.210 2605.720 ;
        RECT 1111.890 2605.660 1112.210 2605.720 ;
        RECT 996.890 2605.520 1112.210 2605.660 ;
        RECT 996.890 2605.460 997.210 2605.520 ;
        RECT 1111.890 2605.460 1112.210 2605.520 ;
        RECT 997.350 2605.320 997.670 2605.380 ;
        RECT 1112.810 2605.320 1113.130 2605.380 ;
        RECT 997.350 2605.180 1113.130 2605.320 ;
        RECT 997.350 2605.120 997.670 2605.180 ;
        RECT 1112.810 2605.120 1113.130 2605.180 ;
        RECT 991.370 2604.980 991.690 2605.040 ;
        RECT 1113.270 2604.980 1113.590 2605.040 ;
        RECT 991.370 2604.840 1113.590 2604.980 ;
        RECT 991.370 2604.780 991.690 2604.840 ;
        RECT 1113.270 2604.780 1113.590 2604.840 ;
        RECT 990.910 2604.640 991.230 2604.700 ;
        RECT 1112.350 2604.640 1112.670 2604.700 ;
        RECT 990.910 2604.500 1112.670 2604.640 ;
        RECT 990.910 2604.440 991.230 2604.500 ;
        RECT 1112.350 2604.440 1112.670 2604.500 ;
        RECT 1397.090 2594.780 1397.410 2594.840 ;
        RECT 1488.630 2594.780 1488.950 2594.840 ;
        RECT 1397.090 2594.640 1488.950 2594.780 ;
        RECT 1397.090 2594.580 1397.410 2594.640 ;
        RECT 1488.630 2594.580 1488.950 2594.640 ;
        RECT 533.210 2591.720 533.530 2591.780 ;
        RECT 769.190 2591.720 769.510 2591.780 ;
        RECT 533.210 2591.580 769.510 2591.720 ;
        RECT 533.210 2591.520 533.530 2591.580 ;
        RECT 769.190 2591.520 769.510 2591.580 ;
        RECT 504.690 2591.380 505.010 2591.440 ;
        RECT 796.790 2591.380 797.110 2591.440 ;
        RECT 504.690 2591.240 797.110 2591.380 ;
        RECT 504.690 2591.180 505.010 2591.240 ;
        RECT 796.790 2591.180 797.110 2591.240 ;
        RECT 990.450 2591.380 990.770 2591.440 ;
        RECT 1094.870 2591.380 1095.190 2591.440 ;
        RECT 990.450 2591.240 1095.190 2591.380 ;
        RECT 990.450 2591.180 990.770 2591.240 ;
        RECT 1094.870 2591.180 1095.190 2591.240 ;
        RECT 1028.170 2587.640 1028.490 2587.700 ;
        RECT 1033.230 2587.640 1033.550 2587.700 ;
        RECT 1028.170 2587.500 1033.550 2587.640 ;
        RECT 1028.170 2587.440 1028.490 2587.500 ;
        RECT 1033.230 2587.440 1033.550 2587.500 ;
        RECT 1424.690 2580.840 1425.010 2580.900 ;
        RECT 1488.630 2580.840 1488.950 2580.900 ;
        RECT 1424.690 2580.700 1488.950 2580.840 ;
        RECT 1424.690 2580.640 1425.010 2580.700 ;
        RECT 1488.630 2580.640 1488.950 2580.700 ;
        RECT 1469.310 2546.500 1469.630 2546.560 ;
        RECT 1483.570 2546.500 1483.890 2546.560 ;
        RECT 1469.310 2546.360 1483.890 2546.500 ;
        RECT 1469.310 2546.300 1469.630 2546.360 ;
        RECT 1483.570 2546.300 1483.890 2546.360 ;
        RECT 1500.130 2512.160 1500.450 2512.220 ;
        RECT 1501.970 2512.160 1502.290 2512.220 ;
        RECT 1500.130 2512.020 1502.290 2512.160 ;
        RECT 1500.130 2511.960 1500.450 2512.020 ;
        RECT 1501.970 2511.960 1502.290 2512.020 ;
      LAYER met1 ;
        RECT 1502.830 2510.640 1885.870 2889.200 ;
      LAYER met1 ;
        RECT 2100.890 2781.440 2101.210 2781.500 ;
        RECT 2556.290 2781.440 2556.610 2781.500 ;
        RECT 2100.890 2781.300 2556.610 2781.440 ;
        RECT 2100.890 2781.240 2101.210 2781.300 ;
        RECT 2556.290 2781.240 2556.610 2781.300 ;
        RECT 1893.890 2781.100 1894.210 2781.160 ;
        RECT 2421.970 2781.100 2422.290 2781.160 ;
        RECT 1893.890 2780.960 2422.290 2781.100 ;
        RECT 1893.890 2780.900 1894.210 2780.960 ;
        RECT 2421.970 2780.900 2422.290 2780.960 ;
      LAYER met1 ;
        RECT 2400.000 2610.640 2556.720 2760.720 ;
      LAYER met1 ;
        RECT 1902.170 2504.000 1902.490 2504.060 ;
        RECT 1903.550 2504.000 1903.870 2504.060 ;
        RECT 1902.170 2503.860 1903.870 2504.000 ;
        RECT 1902.170 2503.800 1902.490 2503.860 ;
        RECT 1903.550 2503.800 1903.870 2503.860 ;
        RECT 1501.970 2495.840 1502.290 2495.900 ;
        RECT 1559.470 2495.840 1559.790 2495.900 ;
        RECT 1501.970 2495.700 1559.790 2495.840 ;
        RECT 1501.970 2495.640 1502.290 2495.700 ;
        RECT 1559.470 2495.640 1559.790 2495.700 ;
        RECT 1494.610 2495.500 1494.930 2495.560 ;
        RECT 1553.030 2495.500 1553.350 2495.560 ;
        RECT 1494.610 2495.360 1553.350 2495.500 ;
        RECT 1494.610 2495.300 1494.930 2495.360 ;
        RECT 1553.030 2495.300 1553.350 2495.360 ;
        RECT 1621.110 2495.500 1621.430 2495.560 ;
        RECT 1892.050 2495.500 1892.370 2495.560 ;
        RECT 1621.110 2495.360 1892.370 2495.500 ;
        RECT 1621.110 2495.300 1621.430 2495.360 ;
        RECT 1892.050 2495.300 1892.370 2495.360 ;
        RECT 1495.070 2495.160 1495.390 2495.220 ;
        RECT 1574.190 2495.160 1574.510 2495.220 ;
        RECT 1495.070 2495.020 1574.510 2495.160 ;
        RECT 1495.070 2494.960 1495.390 2495.020 ;
        RECT 1574.190 2494.960 1574.510 2495.020 ;
        RECT 1607.310 2495.160 1607.630 2495.220 ;
        RECT 1892.510 2495.160 1892.830 2495.220 ;
        RECT 1607.310 2495.020 1892.830 2495.160 ;
        RECT 1607.310 2494.960 1607.630 2495.020 ;
        RECT 1892.510 2494.960 1892.830 2495.020 ;
        RECT 1493.230 2494.820 1493.550 2494.880 ;
        RECT 1580.170 2494.820 1580.490 2494.880 ;
        RECT 1493.230 2494.680 1580.490 2494.820 ;
        RECT 1493.230 2494.620 1493.550 2494.680 ;
        RECT 1580.170 2494.620 1580.490 2494.680 ;
        RECT 1586.610 2494.820 1586.930 2494.880 ;
        RECT 1894.350 2494.820 1894.670 2494.880 ;
        RECT 1586.610 2494.680 1894.670 2494.820 ;
        RECT 1586.610 2494.620 1586.930 2494.680 ;
        RECT 1894.350 2494.620 1894.670 2494.680 ;
        RECT 1494.150 2494.480 1494.470 2494.540 ;
        RECT 1545.670 2494.480 1545.990 2494.540 ;
        RECT 1494.150 2494.340 1545.990 2494.480 ;
        RECT 1494.150 2494.280 1494.470 2494.340 ;
        RECT 1545.670 2494.280 1545.990 2494.340 ;
        RECT 1552.110 2494.480 1552.430 2494.540 ;
        RECT 1893.430 2494.480 1893.750 2494.540 ;
        RECT 1552.110 2494.340 1893.750 2494.480 ;
        RECT 1552.110 2494.280 1552.430 2494.340 ;
        RECT 1893.430 2494.280 1893.750 2494.340 ;
        RECT 1492.310 2494.140 1492.630 2494.200 ;
        RECT 1532.330 2494.140 1532.650 2494.200 ;
        RECT 1492.310 2494.000 1532.650 2494.140 ;
        RECT 1492.310 2493.940 1492.630 2494.000 ;
        RECT 1532.330 2493.940 1532.650 2494.000 ;
        RECT 1545.210 2494.140 1545.530 2494.200 ;
        RECT 1892.970 2494.140 1893.290 2494.200 ;
        RECT 1545.210 2494.000 1893.290 2494.140 ;
        RECT 1545.210 2493.940 1545.530 2494.000 ;
        RECT 1892.970 2493.940 1893.290 2494.000 ;
        RECT 1492.770 2491.420 1493.090 2491.480 ;
        RECT 1512.090 2491.420 1512.410 2491.480 ;
        RECT 1492.770 2491.280 1512.410 2491.420 ;
        RECT 1492.770 2491.220 1493.090 2491.280 ;
        RECT 1512.090 2491.220 1512.410 2491.280 ;
        RECT 1600.410 2489.720 1600.730 2489.780 ;
        RECT 1789.930 2489.720 1790.250 2489.780 ;
        RECT 1600.410 2489.580 1790.250 2489.720 ;
        RECT 1600.410 2489.520 1600.730 2489.580 ;
        RECT 1789.930 2489.520 1790.250 2489.580 ;
        RECT 1693.790 2489.380 1694.110 2489.440 ;
        RECT 1811.090 2489.380 1811.410 2489.440 ;
        RECT 1693.790 2489.240 1811.410 2489.380 ;
        RECT 1693.790 2489.180 1694.110 2489.240 ;
        RECT 1811.090 2489.180 1811.410 2489.240 ;
        RECT 1420.550 2489.040 1420.870 2489.100 ;
        RECT 1842.370 2489.040 1842.690 2489.100 ;
        RECT 1420.550 2488.900 1842.690 2489.040 ;
        RECT 1420.550 2488.840 1420.870 2488.900 ;
        RECT 1842.370 2488.840 1842.690 2488.900 ;
        RECT 1455.050 2488.700 1455.370 2488.760 ;
        RECT 1885.610 2488.700 1885.930 2488.760 ;
        RECT 1455.050 2488.560 1885.930 2488.700 ;
        RECT 1455.050 2488.500 1455.370 2488.560 ;
        RECT 1885.610 2488.500 1885.930 2488.560 ;
        RECT 1421.010 2488.360 1421.330 2488.420 ;
        RECT 1874.570 2488.360 1874.890 2488.420 ;
        RECT 1421.010 2488.220 1874.890 2488.360 ;
        RECT 1421.010 2488.160 1421.330 2488.220 ;
        RECT 1874.570 2488.160 1874.890 2488.220 ;
        RECT 1530.030 2488.020 1530.350 2488.080 ;
        RECT 1832.250 2488.020 1832.570 2488.080 ;
        RECT 1530.030 2487.880 1832.570 2488.020 ;
        RECT 1530.030 2487.820 1530.350 2487.880 ;
        RECT 1832.250 2487.820 1832.570 2487.880 ;
        RECT 1427.910 2487.000 1428.230 2487.060 ;
        RECT 1725.530 2487.000 1725.850 2487.060 ;
        RECT 1427.910 2486.860 1725.850 2487.000 ;
        RECT 1427.910 2486.800 1428.230 2486.860 ;
        RECT 1725.530 2486.800 1725.850 2486.860 ;
        RECT 1461.490 2486.660 1461.810 2486.720 ;
        RECT 1757.730 2486.660 1758.050 2486.720 ;
        RECT 1461.490 2486.520 1758.050 2486.660 ;
        RECT 1461.490 2486.460 1461.810 2486.520 ;
        RECT 1757.730 2486.460 1758.050 2486.520 ;
        RECT 1386.510 2486.320 1386.830 2486.380 ;
        RECT 1587.530 2486.320 1587.850 2486.380 ;
        RECT 1386.510 2486.180 1587.850 2486.320 ;
        RECT 1386.510 2486.120 1386.830 2486.180 ;
        RECT 1587.530 2486.120 1587.850 2486.180 ;
        RECT 1686.890 2486.320 1687.210 2486.380 ;
        RECT 1778.890 2486.320 1779.210 2486.380 ;
        RECT 1686.890 2486.180 1779.210 2486.320 ;
        RECT 1686.890 2486.120 1687.210 2486.180 ;
        RECT 1778.890 2486.120 1779.210 2486.180 ;
        RECT 1383.290 2485.980 1383.610 2486.040 ;
        RECT 1555.330 2485.980 1555.650 2486.040 ;
        RECT 1383.290 2485.840 1555.650 2485.980 ;
        RECT 1383.290 2485.780 1383.610 2485.840 ;
        RECT 1555.330 2485.780 1555.650 2485.840 ;
        RECT 1579.710 2485.980 1580.030 2486.040 ;
        RECT 1746.690 2485.980 1747.010 2486.040 ;
        RECT 1579.710 2485.840 1747.010 2485.980 ;
        RECT 1579.710 2485.780 1580.030 2485.840 ;
        RECT 1746.690 2485.780 1747.010 2485.840 ;
        RECT 1442.630 2485.640 1442.950 2485.700 ;
        RECT 1608.690 2485.640 1609.010 2485.700 ;
        RECT 1442.630 2485.500 1609.010 2485.640 ;
        RECT 1442.630 2485.440 1442.950 2485.500 ;
        RECT 1608.690 2485.440 1609.010 2485.500 ;
        RECT 1507.490 2485.300 1507.810 2485.360 ;
        RECT 1629.850 2485.300 1630.170 2485.360 ;
        RECT 1507.490 2485.160 1630.170 2485.300 ;
        RECT 1507.490 2485.100 1507.810 2485.160 ;
        RECT 1629.850 2485.100 1630.170 2485.160 ;
        RECT 1432.050 2484.960 1432.370 2485.020 ;
        RECT 1534.170 2484.960 1534.490 2485.020 ;
        RECT 1432.050 2484.820 1534.490 2484.960 ;
        RECT 1432.050 2484.760 1432.370 2484.820 ;
        RECT 1534.170 2484.760 1534.490 2484.820 ;
        RECT 1544.750 2484.960 1545.070 2485.020 ;
        RECT 1608.690 2484.960 1609.010 2485.020 ;
        RECT 1544.750 2484.820 1609.010 2484.960 ;
        RECT 1544.750 2484.760 1545.070 2484.820 ;
        RECT 1608.690 2484.760 1609.010 2484.820 ;
        RECT 1528.190 2484.620 1528.510 2484.680 ;
        RECT 1619.730 2484.620 1620.050 2484.680 ;
        RECT 1528.190 2484.480 1620.050 2484.620 ;
        RECT 1528.190 2484.420 1528.510 2484.480 ;
        RECT 1619.730 2484.420 1620.050 2484.480 ;
        RECT 1541.990 2484.280 1542.310 2484.340 ;
        RECT 1576.490 2484.280 1576.810 2484.340 ;
        RECT 1541.990 2484.140 1576.810 2484.280 ;
        RECT 1541.990 2484.080 1542.310 2484.140 ;
        RECT 1576.490 2484.080 1576.810 2484.140 ;
        RECT 1652.390 2484.280 1652.710 2484.340 ;
        RECT 1683.210 2484.280 1683.530 2484.340 ;
        RECT 1652.390 2484.140 1683.530 2484.280 ;
        RECT 1652.390 2484.080 1652.710 2484.140 ;
        RECT 1683.210 2484.080 1683.530 2484.140 ;
        RECT 1700.690 2484.280 1701.010 2484.340 ;
        RECT 1715.410 2484.280 1715.730 2484.340 ;
        RECT 1700.690 2484.140 1715.730 2484.280 ;
        RECT 1700.690 2484.080 1701.010 2484.140 ;
        RECT 1715.410 2484.080 1715.730 2484.140 ;
        RECT 1441.710 2429.340 1442.030 2429.600 ;
        RECT 1441.250 2428.520 1441.570 2428.580 ;
        RECT 1441.800 2428.520 1441.940 2429.340 ;
        RECT 1520.830 2429.000 1521.150 2429.260 ;
        RECT 1441.250 2428.380 1441.940 2428.520 ;
        RECT 1520.920 2428.520 1521.060 2429.000 ;
        RECT 1521.290 2428.520 1521.610 2428.580 ;
        RECT 1520.920 2428.380 1521.610 2428.520 ;
        RECT 1441.250 2428.320 1441.570 2428.380 ;
        RECT 1521.290 2428.320 1521.610 2428.380 ;
        RECT 1441.250 2414.920 1441.570 2414.980 ;
        RECT 1441.710 2414.920 1442.030 2414.980 ;
        RECT 1441.250 2414.780 1442.030 2414.920 ;
        RECT 1441.250 2414.720 1441.570 2414.780 ;
        RECT 1441.710 2414.720 1442.030 2414.780 ;
        RECT 1519.910 2414.920 1520.230 2414.980 ;
        RECT 1521.290 2414.920 1521.610 2414.980 ;
        RECT 1519.910 2414.780 1521.610 2414.920 ;
        RECT 1519.910 2414.720 1520.230 2414.780 ;
        RECT 1521.290 2414.720 1521.610 2414.780 ;
        RECT 1441.710 2380.580 1442.030 2380.640 ;
        RECT 1441.340 2380.440 1442.030 2380.580 ;
        RECT 1441.340 2380.300 1441.480 2380.440 ;
        RECT 1441.710 2380.380 1442.030 2380.440 ;
        RECT 1441.250 2380.040 1441.570 2380.300 ;
        RECT 1440.330 2342.500 1440.650 2342.560 ;
        RECT 1441.710 2342.500 1442.030 2342.560 ;
        RECT 1440.330 2342.360 1442.030 2342.500 ;
        RECT 1440.330 2342.300 1440.650 2342.360 ;
        RECT 1441.710 2342.300 1442.030 2342.360 ;
        RECT 1520.830 2332.100 1521.150 2332.360 ;
        RECT 1520.920 2331.960 1521.060 2332.100 ;
        RECT 1521.290 2331.960 1521.610 2332.020 ;
        RECT 1520.920 2331.820 1521.610 2331.960 ;
        RECT 1521.290 2331.760 1521.610 2331.820 ;
        RECT 1440.330 2319.040 1440.650 2319.100 ;
        RECT 1441.250 2319.040 1441.570 2319.100 ;
        RECT 1440.330 2318.900 1441.570 2319.040 ;
        RECT 1440.330 2318.840 1440.650 2318.900 ;
        RECT 1441.250 2318.840 1441.570 2318.900 ;
        RECT 1441.250 2318.360 1441.570 2318.420 ;
        RECT 1441.710 2318.360 1442.030 2318.420 ;
        RECT 1441.250 2318.220 1442.030 2318.360 ;
        RECT 1441.250 2318.160 1441.570 2318.220 ;
        RECT 1441.710 2318.160 1442.030 2318.220 ;
        RECT 1521.290 2284.160 1521.610 2284.420 ;
        RECT 1441.710 2284.020 1442.030 2284.080 ;
        RECT 1441.340 2283.880 1442.030 2284.020 ;
        RECT 1441.340 2283.740 1441.480 2283.880 ;
        RECT 1441.710 2283.820 1442.030 2283.880 ;
        RECT 1521.380 2283.740 1521.520 2284.160 ;
        RECT 1441.250 2283.480 1441.570 2283.740 ;
        RECT 1521.290 2283.480 1521.610 2283.740 ;
        RECT 1521.290 2270.080 1521.610 2270.140 ;
        RECT 1521.750 2270.080 1522.070 2270.140 ;
        RECT 1521.290 2269.940 1522.070 2270.080 ;
        RECT 1521.290 2269.880 1521.610 2269.940 ;
        RECT 1521.750 2269.880 1522.070 2269.940 ;
        RECT 1520.830 2262.940 1521.150 2263.000 ;
        RECT 1521.750 2262.940 1522.070 2263.000 ;
        RECT 1520.830 2262.800 1522.070 2262.940 ;
        RECT 1520.830 2262.740 1521.150 2262.800 ;
        RECT 1521.750 2262.740 1522.070 2262.800 ;
        RECT 1440.330 2245.940 1440.650 2246.000 ;
        RECT 1441.710 2245.940 1442.030 2246.000 ;
        RECT 1440.330 2245.800 1442.030 2245.940 ;
        RECT 1440.330 2245.740 1440.650 2245.800 ;
        RECT 1441.710 2245.740 1442.030 2245.800 ;
        RECT 1440.330 2222.480 1440.650 2222.540 ;
        RECT 1441.250 2222.480 1441.570 2222.540 ;
        RECT 1440.330 2222.340 1441.570 2222.480 ;
        RECT 1440.330 2222.280 1440.650 2222.340 ;
        RECT 1441.250 2222.280 1441.570 2222.340 ;
        RECT 1441.250 2221.800 1441.570 2221.860 ;
        RECT 1441.710 2221.800 1442.030 2221.860 ;
        RECT 1441.250 2221.660 1442.030 2221.800 ;
        RECT 1441.250 2221.600 1441.570 2221.660 ;
        RECT 1441.710 2221.600 1442.030 2221.660 ;
        RECT 1520.370 2215.000 1520.690 2215.060 ;
        RECT 1520.830 2215.000 1521.150 2215.060 ;
        RECT 1520.370 2214.860 1521.150 2215.000 ;
        RECT 1520.370 2214.800 1520.690 2214.860 ;
        RECT 1520.830 2214.800 1521.150 2214.860 ;
        RECT 1441.710 2187.460 1442.030 2187.520 ;
        RECT 1441.340 2187.320 1442.030 2187.460 ;
        RECT 1441.340 2187.180 1441.480 2187.320 ;
        RECT 1441.710 2187.260 1442.030 2187.320 ;
        RECT 1441.250 2186.920 1441.570 2187.180 ;
        RECT 1520.370 2173.860 1520.690 2173.920 ;
        RECT 1520.830 2173.860 1521.150 2173.920 ;
        RECT 1520.370 2173.720 1521.150 2173.860 ;
        RECT 1520.370 2173.660 1520.690 2173.720 ;
        RECT 1520.830 2173.660 1521.150 2173.720 ;
        RECT 1520.830 2162.980 1521.150 2163.040 ;
        RECT 1521.750 2162.980 1522.070 2163.040 ;
        RECT 1520.830 2162.840 1522.070 2162.980 ;
        RECT 1520.830 2162.780 1521.150 2162.840 ;
        RECT 1521.750 2162.780 1522.070 2162.840 ;
        RECT 1440.330 2149.380 1440.650 2149.440 ;
        RECT 1441.710 2149.380 1442.030 2149.440 ;
        RECT 1440.330 2149.240 1442.030 2149.380 ;
        RECT 1440.330 2149.180 1440.650 2149.240 ;
        RECT 1441.710 2149.180 1442.030 2149.240 ;
        RECT 1440.330 2125.920 1440.650 2125.980 ;
        RECT 1441.250 2125.920 1441.570 2125.980 ;
        RECT 1440.330 2125.780 1441.570 2125.920 ;
        RECT 1440.330 2125.720 1440.650 2125.780 ;
        RECT 1441.250 2125.720 1441.570 2125.780 ;
        RECT 1440.330 2125.240 1440.650 2125.300 ;
        RECT 1441.250 2125.240 1441.570 2125.300 ;
        RECT 1440.330 2125.100 1441.570 2125.240 ;
        RECT 1440.330 2125.040 1440.650 2125.100 ;
        RECT 1441.250 2125.040 1441.570 2125.100 ;
        RECT 1519.910 2076.960 1520.230 2077.020 ;
        RECT 1520.370 2076.960 1520.690 2077.020 ;
        RECT 1519.910 2076.820 1520.690 2076.960 ;
        RECT 1519.910 2076.760 1520.230 2076.820 ;
        RECT 1520.370 2076.760 1520.690 2076.820 ;
        RECT 1518.990 2069.820 1519.310 2069.880 ;
        RECT 1519.910 2069.820 1520.230 2069.880 ;
        RECT 1518.990 2069.680 1520.230 2069.820 ;
        RECT 1518.990 2069.620 1519.310 2069.680 ;
        RECT 1519.910 2069.620 1520.230 2069.680 ;
        RECT 1244.830 2054.180 1245.150 2054.240 ;
        RECT 1332.690 2054.180 1333.010 2054.240 ;
        RECT 1244.830 2054.040 1333.010 2054.180 ;
        RECT 1244.830 2053.980 1245.150 2054.040 ;
        RECT 1332.690 2053.980 1333.010 2054.040 ;
        RECT 1230.110 2053.840 1230.430 2053.900 ;
        RECT 1338.670 2053.840 1338.990 2053.900 ;
        RECT 1230.110 2053.700 1338.990 2053.840 ;
        RECT 1230.110 2053.640 1230.430 2053.700 ;
        RECT 1338.670 2053.640 1338.990 2053.700 ;
        RECT 1173.070 2053.500 1173.390 2053.560 ;
        RECT 1333.150 2053.500 1333.470 2053.560 ;
        RECT 1173.070 2053.360 1333.470 2053.500 ;
        RECT 1173.070 2053.300 1173.390 2053.360 ;
        RECT 1333.150 2053.300 1333.470 2053.360 ;
        RECT 1144.550 2053.160 1144.870 2053.220 ;
        RECT 1334.990 2053.160 1335.310 2053.220 ;
        RECT 1144.550 2053.020 1335.310 2053.160 ;
        RECT 1144.550 2052.960 1144.870 2053.020 ;
        RECT 1334.990 2052.960 1335.310 2053.020 ;
        RECT 1116.950 2052.820 1117.270 2052.880 ;
        RECT 1334.530 2052.820 1334.850 2052.880 ;
        RECT 1116.950 2052.680 1334.850 2052.820 ;
        RECT 1116.950 2052.620 1117.270 2052.680 ;
        RECT 1334.530 2052.620 1334.850 2052.680 ;
        RECT 1059.910 2052.480 1060.230 2052.540 ;
        RECT 1335.450 2052.480 1335.770 2052.540 ;
        RECT 1059.910 2052.340 1335.770 2052.480 ;
        RECT 1059.910 2052.280 1060.230 2052.340 ;
        RECT 1335.450 2052.280 1335.770 2052.340 ;
        RECT 1031.390 2052.140 1031.710 2052.200 ;
        RECT 1331.770 2052.140 1332.090 2052.200 ;
        RECT 1031.390 2052.000 1332.090 2052.140 ;
        RECT 1031.390 2051.940 1031.710 2052.000 ;
        RECT 1331.770 2051.940 1332.090 2052.000 ;
        RECT 1216.310 2051.800 1216.630 2051.860 ;
        RECT 1334.070 2051.800 1334.390 2051.860 ;
        RECT 1216.310 2051.660 1334.390 2051.800 ;
        RECT 1216.310 2051.600 1216.630 2051.660 ;
        RECT 1334.070 2051.600 1334.390 2051.660 ;
        RECT 1201.590 2051.460 1201.910 2051.520 ;
        RECT 1333.610 2051.460 1333.930 2051.520 ;
        RECT 1201.590 2051.320 1333.930 2051.460 ;
        RECT 1201.590 2051.260 1201.910 2051.320 ;
        RECT 1333.610 2051.260 1333.930 2051.320 ;
        RECT 1187.790 2051.120 1188.110 2051.180 ;
        RECT 1338.210 2051.120 1338.530 2051.180 ;
        RECT 1187.790 2050.980 1338.530 2051.120 ;
        RECT 1187.790 2050.920 1188.110 2050.980 ;
        RECT 1338.210 2050.920 1338.530 2050.980 ;
        RECT 984.470 2050.780 984.790 2050.840 ;
        RECT 1002.870 2050.780 1003.190 2050.840 ;
        RECT 984.470 2050.640 1003.190 2050.780 ;
        RECT 984.470 2050.580 984.790 2050.640 ;
        RECT 1002.870 2050.580 1003.190 2050.640 ;
        RECT 1287.150 2050.780 1287.470 2050.840 ;
        RECT 1343.730 2050.780 1344.050 2050.840 ;
        RECT 1287.150 2050.640 1344.050 2050.780 ;
        RECT 1287.150 2050.580 1287.470 2050.640 ;
        RECT 1343.730 2050.580 1344.050 2050.640 ;
        RECT 998.730 2050.440 999.050 2050.500 ;
        RECT 1088.430 2050.440 1088.750 2050.500 ;
        RECT 998.730 2050.300 1088.750 2050.440 ;
        RECT 998.730 2050.240 999.050 2050.300 ;
        RECT 1088.430 2050.240 1088.750 2050.300 ;
        RECT 1273.350 2050.440 1273.670 2050.500 ;
        RECT 1344.190 2050.440 1344.510 2050.500 ;
        RECT 1273.350 2050.300 1344.510 2050.440 ;
        RECT 1273.350 2050.240 1273.670 2050.300 ;
        RECT 1344.190 2050.240 1344.510 2050.300 ;
        RECT 999.650 2050.100 999.970 2050.160 ;
        RECT 1102.230 2050.100 1102.550 2050.160 ;
        RECT 999.650 2049.960 1102.550 2050.100 ;
        RECT 999.650 2049.900 999.970 2049.960 ;
        RECT 1102.230 2049.900 1102.550 2049.960 ;
        RECT 1258.630 2050.100 1258.950 2050.160 ;
        RECT 1332.230 2050.100 1332.550 2050.160 ;
        RECT 1258.630 2049.960 1332.550 2050.100 ;
        RECT 1258.630 2049.900 1258.950 2049.960 ;
        RECT 1332.230 2049.900 1332.550 2049.960 ;
        RECT 1000.110 2049.760 1000.430 2049.820 ;
        RECT 1073.710 2049.760 1074.030 2049.820 ;
        RECT 1000.110 2049.620 1074.030 2049.760 ;
        RECT 1000.110 2049.560 1000.430 2049.620 ;
        RECT 1073.710 2049.560 1074.030 2049.620 ;
        RECT 1301.870 2049.760 1302.190 2049.820 ;
        RECT 1337.750 2049.760 1338.070 2049.820 ;
        RECT 1301.870 2049.620 1338.070 2049.760 ;
        RECT 1301.870 2049.560 1302.190 2049.620 ;
        RECT 1337.750 2049.560 1338.070 2049.620 ;
        RECT 999.190 2049.420 999.510 2049.480 ;
        RECT 1045.190 2049.420 1045.510 2049.480 ;
        RECT 999.190 2049.280 1045.510 2049.420 ;
        RECT 999.190 2049.220 999.510 2049.280 ;
        RECT 1045.190 2049.220 1045.510 2049.280 ;
        RECT 1329.470 2049.420 1329.790 2049.480 ;
        RECT 1344.650 2049.420 1344.970 2049.480 ;
        RECT 1329.470 2049.280 1344.970 2049.420 ;
        RECT 1329.470 2049.220 1329.790 2049.280 ;
        RECT 1344.650 2049.220 1344.970 2049.280 ;
        RECT 997.810 2048.400 998.130 2048.460 ;
        RECT 1014.370 2048.400 1014.690 2048.460 ;
        RECT 997.810 2048.260 1014.690 2048.400 ;
        RECT 997.810 2048.200 998.130 2048.260 ;
        RECT 1014.370 2048.200 1014.690 2048.260 ;
        RECT 998.270 2048.060 998.590 2048.120 ;
        RECT 1028.170 2048.060 1028.490 2048.120 ;
        RECT 998.270 2047.920 1028.490 2048.060 ;
        RECT 998.270 2047.860 998.590 2047.920 ;
        RECT 1028.170 2047.860 1028.490 2047.920 ;
        RECT 984.010 2047.720 984.330 2047.780 ;
        RECT 1048.870 2047.720 1049.190 2047.780 ;
        RECT 984.010 2047.580 1049.190 2047.720 ;
        RECT 984.010 2047.520 984.330 2047.580 ;
        RECT 1048.870 2047.520 1049.190 2047.580 ;
        RECT 978.490 2047.380 978.810 2047.440 ;
        RECT 1062.670 2047.380 1062.990 2047.440 ;
        RECT 978.490 2047.240 1062.990 2047.380 ;
        RECT 978.490 2047.180 978.810 2047.240 ;
        RECT 1062.670 2047.180 1062.990 2047.240 ;
        RECT 978.950 2047.040 979.270 2047.100 ;
        RECT 1076.470 2047.040 1076.790 2047.100 ;
        RECT 978.950 2046.900 1076.790 2047.040 ;
        RECT 978.950 2046.840 979.270 2046.900 ;
        RECT 1076.470 2046.840 1076.790 2046.900 ;
        RECT 983.550 2046.700 983.870 2046.760 ;
        RECT 1113.730 2046.700 1114.050 2046.760 ;
        RECT 983.550 2046.560 1114.050 2046.700 ;
        RECT 983.550 2046.500 983.870 2046.560 ;
        RECT 1113.730 2046.500 1114.050 2046.560 ;
        RECT 983.090 2046.360 983.410 2046.420 ;
        RECT 1114.190 2046.360 1114.510 2046.420 ;
        RECT 983.090 2046.220 1114.510 2046.360 ;
        RECT 983.090 2046.160 983.410 2046.220 ;
        RECT 1114.190 2046.160 1114.510 2046.220 ;
        RECT 978.030 2046.020 978.350 2046.080 ;
        RECT 1110.970 2046.020 1111.290 2046.080 ;
        RECT 978.030 2045.880 1111.290 2046.020 ;
        RECT 978.030 2045.820 978.350 2045.880 ;
        RECT 1110.970 2045.820 1111.290 2045.880 ;
        RECT 977.570 2045.680 977.890 2045.740 ;
        RECT 1111.430 2045.680 1111.750 2045.740 ;
        RECT 977.570 2045.540 1111.750 2045.680 ;
        RECT 977.570 2045.480 977.890 2045.540 ;
        RECT 1111.430 2045.480 1111.750 2045.540 ;
        RECT 1439.410 2042.620 1439.730 2042.680 ;
        RECT 1439.870 2042.620 1440.190 2042.680 ;
        RECT 1439.410 2042.480 1440.190 2042.620 ;
        RECT 1439.410 2042.420 1439.730 2042.480 ;
        RECT 1439.870 2042.420 1440.190 2042.480 ;
        RECT 579.210 1988.900 579.530 1988.960 ;
        RECT 632.110 1988.900 632.430 1988.960 ;
        RECT 579.210 1988.760 632.430 1988.900 ;
        RECT 579.210 1988.700 579.530 1988.760 ;
        RECT 632.110 1988.700 632.430 1988.760 ;
        RECT 529.990 1988.220 530.310 1988.280 ;
        RECT 638.090 1988.220 638.410 1988.280 ;
        RECT 529.990 1988.080 638.410 1988.220 ;
        RECT 529.990 1988.020 530.310 1988.080 ;
        RECT 638.090 1988.020 638.410 1988.080 ;
        RECT 419.590 1980.060 419.910 1980.120 ;
        RECT 420.510 1980.060 420.830 1980.120 ;
        RECT 419.590 1979.920 420.830 1980.060 ;
        RECT 419.590 1979.860 419.910 1979.920 ;
        RECT 420.510 1979.860 420.830 1979.920 ;
        RECT 420.050 1978.700 420.370 1978.760 ;
        RECT 420.050 1978.560 420.740 1978.700 ;
        RECT 420.050 1978.500 420.370 1978.560 ;
        RECT 419.590 1978.160 419.910 1978.420 ;
        RECT 419.680 1977.680 419.820 1978.160 ;
        RECT 420.600 1978.020 420.740 1978.560 ;
        RECT 843.250 1978.020 843.570 1978.080 ;
        RECT 420.600 1977.880 843.570 1978.020 ;
        RECT 843.250 1977.820 843.570 1977.880 ;
        RECT 897.530 1977.680 897.850 1977.740 ;
        RECT 419.680 1977.540 897.850 1977.680 ;
        RECT 897.530 1977.480 897.850 1977.540 ;
      LAYER met1 ;
        RECT 362.830 1704.460 628.110 1977.400 ;
      LAYER met1 ;
        RECT 996.430 1714.520 996.750 1714.580 ;
        RECT 1001.030 1714.520 1001.350 1714.580 ;
        RECT 996.430 1714.380 1001.350 1714.520 ;
        RECT 996.430 1714.320 996.750 1714.380 ;
        RECT 1001.030 1714.320 1001.350 1714.380 ;
      LAYER met1 ;
        RECT 1002.830 1710.640 1329.750 2032.080 ;
      LAYER met1 ;
        RECT 1441.710 1994.000 1442.030 1994.060 ;
        RECT 1442.630 1994.000 1442.950 1994.060 ;
        RECT 1441.710 1993.860 1442.950 1994.000 ;
        RECT 1441.710 1993.800 1442.030 1993.860 ;
        RECT 1442.630 1993.800 1442.950 1993.860 ;
        RECT 1519.910 1994.000 1520.230 1994.060 ;
        RECT 1521.290 1994.000 1521.610 1994.060 ;
        RECT 1519.910 1993.860 1521.610 1994.000 ;
        RECT 1519.910 1993.800 1520.230 1993.860 ;
        RECT 1521.290 1993.800 1521.610 1993.860 ;
        RECT 2082.950 1947.080 2083.270 1947.140 ;
        RECT 2321.230 1947.080 2321.550 1947.140 ;
        RECT 2082.950 1946.940 2321.550 1947.080 ;
        RECT 2082.950 1946.880 2083.270 1946.940 ;
        RECT 2321.230 1946.880 2321.550 1946.940 ;
        RECT 2073.290 1946.740 2073.610 1946.800 ;
        RECT 2379.190 1946.740 2379.510 1946.800 ;
        RECT 2073.290 1946.600 2379.510 1946.740 ;
        RECT 2073.290 1946.540 2073.610 1946.600 ;
        RECT 2379.190 1946.540 2379.510 1946.600 ;
        RECT 2090.310 1946.400 2090.630 1946.460 ;
        RECT 2437.150 1946.400 2437.470 1946.460 ;
        RECT 2090.310 1946.260 2437.470 1946.400 ;
        RECT 2090.310 1946.200 2090.630 1946.260 ;
        RECT 2437.150 1946.200 2437.470 1946.260 ;
        RECT 1521.290 1946.060 1521.610 1946.120 ;
        RECT 1520.920 1945.920 1521.610 1946.060 ;
        RECT 1520.920 1945.780 1521.060 1945.920 ;
        RECT 1521.290 1945.860 1521.610 1945.920 ;
        RECT 2083.410 1946.060 2083.730 1946.120 ;
        RECT 2495.110 1946.060 2495.430 1946.120 ;
        RECT 2083.410 1945.920 2495.430 1946.060 ;
        RECT 2083.410 1945.860 2083.730 1945.920 ;
        RECT 2495.110 1945.860 2495.430 1945.920 ;
        RECT 1520.830 1945.520 1521.150 1945.780 ;
        RECT 1876.410 1935.520 1876.730 1935.580 ;
        RECT 2394.370 1935.520 2394.690 1935.580 ;
        RECT 1876.410 1935.380 2394.690 1935.520 ;
        RECT 1876.410 1935.320 1876.730 1935.380 ;
        RECT 2394.370 1935.320 2394.690 1935.380 ;
        RECT 1521.290 1931.780 1521.610 1931.840 ;
        RECT 1522.210 1931.780 1522.530 1931.840 ;
        RECT 1521.290 1931.640 1522.530 1931.780 ;
        RECT 1521.290 1931.580 1521.610 1931.640 ;
        RECT 1522.210 1931.580 1522.530 1931.640 ;
        RECT 1724.610 1929.060 1724.930 1929.120 ;
        RECT 2044.310 1929.060 2044.630 1929.120 ;
        RECT 1724.610 1928.920 2044.630 1929.060 ;
        RECT 1724.610 1928.860 1724.930 1928.920 ;
        RECT 2044.310 1928.860 2044.630 1928.920 ;
        RECT 1845.590 1928.040 1845.910 1928.100 ;
        RECT 1964.270 1928.040 1964.590 1928.100 ;
        RECT 1845.590 1927.900 1964.590 1928.040 ;
        RECT 1845.590 1927.840 1845.910 1927.900 ;
        RECT 1964.270 1927.840 1964.590 1927.900 ;
        RECT 1745.310 1927.700 1745.630 1927.760 ;
        RECT 1929.310 1927.700 1929.630 1927.760 ;
        RECT 1745.310 1927.560 1929.630 1927.700 ;
        RECT 1745.310 1927.500 1745.630 1927.560 ;
        RECT 1929.310 1927.500 1929.630 1927.560 ;
        RECT 1779.350 1927.360 1779.670 1927.420 ;
        RECT 1998.310 1927.360 1998.630 1927.420 ;
        RECT 1779.350 1927.220 1998.630 1927.360 ;
        RECT 1779.350 1927.160 1779.670 1927.220 ;
        RECT 1998.310 1927.160 1998.630 1927.220 ;
        RECT 1786.710 1927.020 1787.030 1927.080 ;
        RECT 2033.270 1927.020 2033.590 1927.080 ;
        RECT 1786.710 1926.880 2033.590 1927.020 ;
        RECT 1786.710 1926.820 1787.030 1926.880 ;
        RECT 2033.270 1926.820 2033.590 1926.880 ;
        RECT 1766.010 1926.680 1766.330 1926.740 ;
        RECT 2010.270 1926.680 2010.590 1926.740 ;
        RECT 1766.010 1926.540 2010.590 1926.680 ;
        RECT 1766.010 1926.480 1766.330 1926.540 ;
        RECT 2010.270 1926.480 2010.590 1926.540 ;
        RECT 1738.410 1926.340 1738.730 1926.400 ;
        RECT 1987.270 1926.340 1987.590 1926.400 ;
        RECT 1738.410 1926.200 1987.590 1926.340 ;
        RECT 1738.410 1926.140 1738.730 1926.200 ;
        RECT 1987.270 1926.140 1987.590 1926.200 ;
        RECT 1717.710 1926.000 1718.030 1926.060 ;
        RECT 1975.310 1926.000 1975.630 1926.060 ;
        RECT 1717.710 1925.860 1975.630 1926.000 ;
        RECT 1717.710 1925.800 1718.030 1925.860 ;
        RECT 1975.310 1925.800 1975.630 1925.860 ;
        RECT 1779.810 1925.660 1780.130 1925.720 ;
        RECT 2067.310 1925.660 2067.630 1925.720 ;
        RECT 1779.810 1925.520 2067.630 1925.660 ;
        RECT 1779.810 1925.460 1780.130 1925.520 ;
        RECT 2067.310 1925.460 2067.630 1925.520 ;
        RECT 1835.010 1925.320 1835.330 1925.380 ;
        RECT 1952.310 1925.320 1952.630 1925.380 ;
        RECT 1835.010 1925.180 1952.630 1925.320 ;
        RECT 1835.010 1925.120 1835.330 1925.180 ;
        RECT 1952.310 1925.120 1952.630 1925.180 ;
        RECT 1441.710 1897.440 1442.030 1897.500 ;
        RECT 1442.630 1897.440 1442.950 1897.500 ;
        RECT 1441.710 1897.300 1442.950 1897.440 ;
        RECT 1441.710 1897.240 1442.030 1897.300 ;
        RECT 1442.630 1897.240 1442.950 1897.300 ;
        RECT 1759.110 1883.840 1759.430 1883.900 ;
        RECT 1904.470 1883.840 1904.790 1883.900 ;
        RECT 1759.110 1883.700 1904.790 1883.840 ;
        RECT 1759.110 1883.640 1759.430 1883.700 ;
        RECT 1904.470 1883.640 1904.790 1883.700 ;
        RECT 1821.210 1870.240 1821.530 1870.300 ;
        RECT 1904.470 1870.240 1904.790 1870.300 ;
        RECT 1821.210 1870.100 1904.790 1870.240 ;
        RECT 1821.210 1870.040 1821.530 1870.100 ;
        RECT 1904.470 1870.040 1904.790 1870.100 ;
        RECT 1521.290 1859.700 1521.610 1859.760 ;
        RECT 1522.210 1859.700 1522.530 1859.760 ;
        RECT 1521.290 1859.560 1522.530 1859.700 ;
        RECT 1521.290 1859.500 1521.610 1859.560 ;
        RECT 1522.210 1859.500 1522.530 1859.560 ;
        RECT 1737.950 1849.500 1738.270 1849.560 ;
        RECT 1904.470 1849.500 1904.790 1849.560 ;
        RECT 1737.950 1849.360 1904.790 1849.500 ;
        RECT 1737.950 1849.300 1738.270 1849.360 ;
        RECT 1904.470 1849.300 1904.790 1849.360 ;
        RECT 1669.410 1814.820 1669.730 1814.880 ;
        RECT 1904.470 1814.820 1904.790 1814.880 ;
        RECT 1669.410 1814.680 1904.790 1814.820 ;
        RECT 1669.410 1814.620 1669.730 1814.680 ;
        RECT 1904.470 1814.620 1904.790 1814.680 ;
        RECT 1772.910 1766.540 1773.230 1766.600 ;
        RECT 1904.470 1766.540 1904.790 1766.600 ;
        RECT 1772.910 1766.400 1904.790 1766.540 ;
        RECT 1772.910 1766.340 1773.230 1766.400 ;
        RECT 1904.470 1766.340 1904.790 1766.400 ;
        RECT 1521.290 1763.140 1521.610 1763.200 ;
        RECT 1522.210 1763.140 1522.530 1763.200 ;
        RECT 1521.290 1763.000 1522.530 1763.140 ;
        RECT 1521.290 1762.940 1521.610 1763.000 ;
        RECT 1522.210 1762.940 1522.530 1763.000 ;
      LAYER met1 ;
        RECT 1922.830 1760.240 2072.190 1905.280 ;
      LAYER met1 ;
        RECT 2080.190 1870.240 2080.510 1870.300 ;
        RECT 2283.970 1870.240 2284.290 1870.300 ;
        RECT 2080.190 1870.100 2284.290 1870.240 ;
        RECT 2080.190 1870.040 2080.510 1870.100 ;
        RECT 2283.970 1870.040 2284.290 1870.100 ;
        RECT 1907.690 1738.660 1908.010 1738.720 ;
        RECT 1933.910 1738.660 1934.230 1738.720 ;
        RECT 1907.690 1738.520 1934.230 1738.660 ;
        RECT 1907.690 1738.460 1908.010 1738.520 ;
        RECT 1933.910 1738.460 1934.230 1738.520 ;
        RECT 1800.510 1738.320 1800.830 1738.380 ;
        RECT 1956.910 1738.320 1957.230 1738.380 ;
        RECT 1800.510 1738.180 1957.230 1738.320 ;
        RECT 1800.510 1738.120 1800.830 1738.180 ;
        RECT 1956.910 1738.120 1957.230 1738.180 ;
        RECT 1814.310 1737.980 1814.630 1738.040 ;
        RECT 1990.950 1737.980 1991.270 1738.040 ;
        RECT 1814.310 1737.840 1991.270 1737.980 ;
        RECT 1814.310 1737.780 1814.630 1737.840 ;
        RECT 1990.950 1737.780 1991.270 1737.840 ;
        RECT 1793.610 1737.640 1793.930 1737.700 ;
        RECT 1967.950 1737.640 1968.270 1737.700 ;
        RECT 1793.610 1737.500 1968.270 1737.640 ;
        RECT 1793.610 1737.440 1793.930 1737.500 ;
        RECT 1967.950 1737.440 1968.270 1737.500 ;
        RECT 1813.850 1737.300 1814.170 1737.360 ;
        RECT 2013.950 1737.300 2014.270 1737.360 ;
        RECT 1813.850 1737.160 2014.270 1737.300 ;
        RECT 1813.850 1737.100 1814.170 1737.160 ;
        RECT 2013.950 1737.100 2014.270 1737.160 ;
        RECT 1752.210 1736.960 1752.530 1737.020 ;
        RECT 1979.910 1736.960 1980.230 1737.020 ;
        RECT 1752.210 1736.820 1980.230 1736.960 ;
        RECT 1752.210 1736.760 1752.530 1736.820 ;
        RECT 1979.910 1736.760 1980.230 1736.820 ;
        RECT 1710.810 1736.620 1711.130 1736.680 ;
        RECT 1944.950 1736.620 1945.270 1736.680 ;
        RECT 1710.810 1736.480 1945.270 1736.620 ;
        RECT 1710.810 1736.420 1711.130 1736.480 ;
        RECT 1944.950 1736.420 1945.270 1736.480 ;
        RECT 1807.410 1736.280 1807.730 1736.340 ;
        RECT 2036.950 1736.280 2037.270 1736.340 ;
        RECT 1807.410 1736.140 2037.270 1736.280 ;
        RECT 1807.410 1736.080 1807.730 1736.140 ;
        RECT 2036.950 1736.080 2037.270 1736.140 ;
        RECT 1772.450 1735.940 1772.770 1736.000 ;
        RECT 2002.910 1735.940 2003.230 1736.000 ;
        RECT 1772.450 1735.800 2003.230 1735.940 ;
        RECT 1772.450 1735.740 1772.770 1735.800 ;
        RECT 2002.910 1735.740 2003.230 1735.800 ;
        RECT 1806.950 1735.600 1807.270 1735.660 ;
        RECT 2071.910 1735.600 2072.230 1735.660 ;
        RECT 1806.950 1735.460 2072.230 1735.600 ;
        RECT 1806.950 1735.400 1807.270 1735.460 ;
        RECT 2071.910 1735.400 2072.230 1735.460 ;
        RECT 1668.950 1735.260 1669.270 1735.320 ;
        RECT 2059.950 1735.260 2060.270 1735.320 ;
        RECT 1668.950 1735.120 2060.270 1735.260 ;
        RECT 1668.950 1735.060 1669.270 1735.120 ;
        RECT 2059.950 1735.060 2060.270 1735.120 ;
      LAYER met1 ;
        RECT 2302.830 1710.640 2521.260 1926.000 ;
      LAYER met1 ;
        RECT 2519.030 1710.100 2519.350 1710.160 ;
        RECT 2520.870 1710.100 2521.190 1710.160 ;
        RECT 2519.030 1709.960 2521.190 1710.100 ;
        RECT 2519.030 1709.900 2519.350 1709.960 ;
        RECT 2520.870 1709.900 2521.190 1709.960 ;
        RECT 2523.630 1704.320 2523.950 1704.380 ;
        RECT 2520.500 1704.180 2523.950 1704.320 ;
        RECT 2519.490 1703.980 2519.810 1704.040 ;
        RECT 2520.500 1703.980 2520.640 1704.180 ;
        RECT 2523.630 1704.120 2523.950 1704.180 ;
        RECT 2519.490 1703.840 2520.640 1703.980 ;
        RECT 2519.490 1703.780 2519.810 1703.840 ;
        RECT 1310.610 1695.820 1310.930 1695.880 ;
        RECT 1344.650 1695.820 1344.970 1695.880 ;
        RECT 1310.610 1695.680 1344.970 1695.820 ;
        RECT 1310.610 1695.620 1310.930 1695.680 ;
        RECT 1344.650 1695.620 1344.970 1695.680 ;
        RECT 990.450 1695.140 990.770 1695.200 ;
        RECT 1048.870 1695.140 1049.190 1695.200 ;
        RECT 990.450 1695.000 1049.190 1695.140 ;
        RECT 990.450 1694.940 990.770 1695.000 ;
        RECT 1048.870 1694.940 1049.190 1695.000 ;
        RECT 997.350 1694.800 997.670 1694.860 ;
        RECT 1069.570 1694.800 1069.890 1694.860 ;
        RECT 997.350 1694.660 1069.890 1694.800 ;
        RECT 997.350 1694.600 997.670 1694.660 ;
        RECT 1069.570 1694.600 1069.890 1694.660 ;
        RECT 1288.530 1694.800 1288.850 1694.860 ;
        RECT 1337.750 1694.800 1338.070 1694.860 ;
        RECT 1288.530 1694.660 1338.070 1694.800 ;
        RECT 1288.530 1694.600 1288.850 1694.660 ;
        RECT 1337.750 1694.600 1338.070 1694.660 ;
        RECT 996.890 1694.460 997.210 1694.520 ;
        RECT 1076.470 1694.460 1076.790 1694.520 ;
        RECT 996.890 1694.320 1076.790 1694.460 ;
        RECT 996.890 1694.260 997.210 1694.320 ;
        RECT 1076.470 1694.260 1076.790 1694.320 ;
        RECT 1268.290 1694.460 1268.610 1694.520 ;
        RECT 1344.190 1694.460 1344.510 1694.520 ;
        RECT 1268.290 1694.320 1344.510 1694.460 ;
        RECT 1268.290 1694.260 1268.610 1694.320 ;
        RECT 1344.190 1694.260 1344.510 1694.320 ;
        RECT 991.370 1694.120 991.690 1694.180 ;
        RECT 1104.070 1694.120 1104.390 1694.180 ;
        RECT 991.370 1693.980 1104.390 1694.120 ;
        RECT 991.370 1693.920 991.690 1693.980 ;
        RECT 1104.070 1693.920 1104.390 1693.980 ;
        RECT 1220.910 1694.120 1221.230 1694.180 ;
        RECT 1343.730 1694.120 1344.050 1694.180 ;
        RECT 1220.910 1693.980 1344.050 1694.120 ;
        RECT 1220.910 1693.920 1221.230 1693.980 ;
        RECT 1343.730 1693.920 1344.050 1693.980 ;
        RECT 990.910 1693.780 991.230 1693.840 ;
        RECT 1110.970 1693.780 1111.290 1693.840 ;
        RECT 990.910 1693.640 1111.290 1693.780 ;
        RECT 990.910 1693.580 991.230 1693.640 ;
        RECT 1110.970 1693.580 1111.290 1693.640 ;
        RECT 1186.410 1693.780 1186.730 1693.840 ;
        RECT 1338.210 1693.780 1338.530 1693.840 ;
        RECT 1186.410 1693.640 1338.530 1693.780 ;
        RECT 1186.410 1693.580 1186.730 1693.640 ;
        RECT 1338.210 1693.580 1338.530 1693.640 ;
        RECT 1520.830 1690.720 1521.150 1690.780 ;
        RECT 1522.210 1690.720 1522.530 1690.780 ;
        RECT 1520.830 1690.580 1522.530 1690.720 ;
        RECT 1520.830 1690.520 1521.150 1690.580 ;
        RECT 1522.210 1690.520 1522.530 1690.580 ;
        RECT 1102.230 1690.040 1102.550 1690.100 ;
        RECT 1190.550 1690.040 1190.870 1690.100 ;
        RECT 1102.230 1689.900 1190.870 1690.040 ;
        RECT 1102.230 1689.840 1102.550 1689.900 ;
        RECT 1190.550 1689.840 1190.870 1689.900 ;
        RECT 1045.190 1689.700 1045.510 1689.760 ;
        RECT 1100.390 1689.700 1100.710 1689.760 ;
        RECT 1045.190 1689.560 1100.710 1689.700 ;
        RECT 1045.190 1689.500 1045.510 1689.560 ;
        RECT 1100.390 1689.500 1100.710 1689.560 ;
        RECT 1130.750 1689.700 1131.070 1689.760 ;
        RECT 1243.450 1689.700 1243.770 1689.760 ;
        RECT 1130.750 1689.560 1243.770 1689.700 ;
        RECT 1130.750 1689.500 1131.070 1689.560 ;
        RECT 1243.450 1689.500 1243.770 1689.560 ;
        RECT 1254.950 1689.700 1255.270 1689.760 ;
        RECT 1300.950 1689.700 1301.270 1689.760 ;
        RECT 1254.950 1689.560 1301.270 1689.700 ;
        RECT 1254.950 1689.500 1255.270 1689.560 ;
        RECT 1300.950 1689.500 1301.270 1689.560 ;
        RECT 1016.670 1689.360 1016.990 1689.420 ;
        RECT 1079.690 1689.360 1080.010 1689.420 ;
        RECT 1016.670 1689.220 1080.010 1689.360 ;
        RECT 1016.670 1689.160 1016.990 1689.220 ;
        RECT 1079.690 1689.160 1080.010 1689.220 ;
        RECT 1087.510 1689.360 1087.830 1689.420 ;
        RECT 1195.150 1689.360 1195.470 1689.420 ;
        RECT 1087.510 1689.220 1195.470 1689.360 ;
        RECT 1087.510 1689.160 1087.830 1689.220 ;
        RECT 1195.150 1689.160 1195.470 1689.220 ;
        RECT 1207.110 1689.360 1207.430 1689.420 ;
        RECT 1230.110 1689.360 1230.430 1689.420 ;
        RECT 1207.110 1689.220 1230.430 1689.360 ;
        RECT 1207.110 1689.160 1207.430 1689.220 ;
        RECT 1230.110 1689.160 1230.430 1689.220 ;
        RECT 1268.750 1689.360 1269.070 1689.420 ;
        RECT 1315.670 1689.360 1315.990 1689.420 ;
        RECT 1268.750 1689.220 1315.990 1689.360 ;
        RECT 1268.750 1689.160 1269.070 1689.220 ;
        RECT 1315.670 1689.160 1315.990 1689.220 ;
        RECT 1002.870 1689.020 1003.190 1689.080 ;
        RECT 1167.550 1689.020 1167.870 1689.080 ;
        RECT 1002.870 1688.880 1167.870 1689.020 ;
        RECT 1002.870 1688.820 1003.190 1688.880 ;
        RECT 1167.550 1688.820 1167.870 1688.880 ;
        RECT 1173.070 1689.020 1173.390 1689.080 ;
        RECT 1188.710 1689.020 1189.030 1689.080 ;
        RECT 1173.070 1688.880 1189.030 1689.020 ;
        RECT 1173.070 1688.820 1173.390 1688.880 ;
        RECT 1188.710 1688.820 1189.030 1688.880 ;
        RECT 1200.210 1689.020 1200.530 1689.080 ;
        RECT 1215.390 1689.020 1215.710 1689.080 ;
        RECT 1200.210 1688.880 1215.710 1689.020 ;
        RECT 1200.210 1688.820 1200.530 1688.880 ;
        RECT 1215.390 1688.820 1215.710 1688.880 ;
        RECT 1238.390 1689.020 1238.710 1689.080 ;
        RECT 1287.150 1689.020 1287.470 1689.080 ;
        RECT 1238.390 1688.880 1287.470 1689.020 ;
        RECT 1238.390 1688.820 1238.710 1688.880 ;
        RECT 1287.150 1688.820 1287.470 1688.880 ;
        RECT 463.750 1688.680 464.070 1688.740 ;
        RECT 468.810 1688.680 469.130 1688.740 ;
        RECT 463.750 1688.540 469.130 1688.680 ;
        RECT 463.750 1688.480 464.070 1688.540 ;
        RECT 468.810 1688.480 469.130 1688.540 ;
        RECT 514.350 1688.680 514.670 1688.740 ;
        RECT 517.110 1688.680 517.430 1688.740 ;
        RECT 514.350 1688.540 517.430 1688.680 ;
        RECT 514.350 1688.480 514.670 1688.540 ;
        RECT 517.110 1688.480 517.430 1688.540 ;
        RECT 1073.710 1688.680 1074.030 1688.740 ;
        RECT 1293.590 1688.680 1293.910 1688.740 ;
        RECT 1073.710 1688.540 1293.910 1688.680 ;
        RECT 1073.710 1688.480 1074.030 1688.540 ;
        RECT 1293.590 1688.480 1293.910 1688.540 ;
        RECT 1030.470 1688.340 1030.790 1688.400 ;
        RECT 1258.170 1688.340 1258.490 1688.400 ;
        RECT 1030.470 1688.200 1258.490 1688.340 ;
        RECT 1030.470 1688.140 1030.790 1688.200 ;
        RECT 1258.170 1688.140 1258.490 1688.200 ;
        RECT 1258.630 1688.340 1258.950 1688.400 ;
        RECT 1262.310 1688.340 1262.630 1688.400 ;
        RECT 1258.630 1688.200 1262.630 1688.340 ;
        RECT 1258.630 1688.140 1258.950 1688.200 ;
        RECT 1262.310 1688.140 1262.630 1688.200 ;
        RECT 2007.510 1688.000 2007.830 1688.060 ;
        RECT 2302.830 1688.000 2303.150 1688.060 ;
        RECT 2007.510 1687.860 2303.150 1688.000 ;
        RECT 2007.510 1687.800 2007.830 1687.860 ;
        RECT 2302.830 1687.800 2303.150 1687.860 ;
        RECT 2055.810 1687.660 2056.130 1687.720 ;
        RECT 2360.790 1687.660 2361.110 1687.720 ;
        RECT 2055.810 1687.520 2361.110 1687.660 ;
        RECT 2055.810 1687.460 2056.130 1687.520 ;
        RECT 2360.790 1687.460 2361.110 1687.520 ;
        RECT 2042.010 1687.320 2042.330 1687.380 ;
        RECT 2418.750 1687.320 2419.070 1687.380 ;
        RECT 2042.010 1687.180 2419.070 1687.320 ;
        RECT 2042.010 1687.120 2042.330 1687.180 ;
        RECT 2418.750 1687.120 2419.070 1687.180 ;
        RECT 2069.610 1686.980 2069.930 1687.040 ;
        RECT 2476.710 1686.980 2477.030 1687.040 ;
        RECT 2069.610 1686.840 2477.030 1686.980 ;
        RECT 2069.610 1686.780 2069.930 1686.840 ;
        RECT 2476.710 1686.780 2477.030 1686.840 ;
        RECT 1159.270 1686.640 1159.590 1686.700 ;
        RECT 1243.910 1686.640 1244.230 1686.700 ;
        RECT 1159.270 1686.500 1244.230 1686.640 ;
        RECT 1159.270 1686.440 1159.590 1686.500 ;
        RECT 1243.910 1686.440 1244.230 1686.500 ;
        RECT 1258.170 1686.640 1258.490 1686.700 ;
        RECT 1276.570 1686.640 1276.890 1686.700 ;
        RECT 1258.170 1686.500 1276.890 1686.640 ;
        RECT 1258.170 1686.440 1258.490 1686.500 ;
        RECT 1276.570 1686.440 1276.890 1686.500 ;
        RECT 1144.550 1686.300 1144.870 1686.360 ;
        RECT 1162.490 1686.300 1162.810 1686.360 ;
        RECT 1144.550 1686.160 1162.810 1686.300 ;
        RECT 1144.550 1686.100 1144.870 1686.160 ;
        RECT 1162.490 1686.100 1162.810 1686.160 ;
        RECT 1187.790 1686.300 1188.110 1686.360 ;
        RECT 1215.390 1686.300 1215.710 1686.360 ;
        RECT 1187.790 1686.160 1215.710 1686.300 ;
        RECT 1187.790 1686.100 1188.110 1686.160 ;
        RECT 1215.390 1686.100 1215.710 1686.160 ;
        RECT 1167.550 1685.960 1167.870 1686.020 ;
        RECT 1190.090 1685.960 1190.410 1686.020 ;
        RECT 1167.550 1685.820 1190.410 1685.960 ;
        RECT 1167.550 1685.760 1167.870 1685.820 ;
        RECT 1190.090 1685.760 1190.410 1685.820 ;
        RECT 1195.150 1685.960 1195.470 1686.020 ;
        RECT 1224.590 1685.960 1224.910 1686.020 ;
        RECT 1195.150 1685.820 1224.910 1685.960 ;
        RECT 1195.150 1685.760 1195.470 1685.820 ;
        RECT 1224.590 1685.760 1224.910 1685.820 ;
        RECT 1116.030 1684.260 1116.350 1684.320 ;
        RECT 1148.690 1684.260 1149.010 1684.320 ;
        RECT 1116.030 1684.120 1149.010 1684.260 ;
        RECT 1116.030 1684.060 1116.350 1684.120 ;
        RECT 1148.690 1684.060 1149.010 1684.120 ;
        RECT 1220.450 1684.260 1220.770 1684.320 ;
        RECT 1242.990 1684.260 1243.310 1684.320 ;
        RECT 1220.450 1684.120 1243.310 1684.260 ;
        RECT 1220.450 1684.060 1220.770 1684.120 ;
        RECT 1242.990 1684.060 1243.310 1684.120 ;
        RECT 1272.430 1684.260 1272.750 1684.320 ;
        RECT 1291.290 1684.260 1291.610 1684.320 ;
        RECT 1272.430 1684.120 1291.610 1684.260 ;
        RECT 1272.430 1684.060 1272.750 1684.120 ;
        RECT 1291.290 1684.060 1291.610 1684.120 ;
        RECT 1288.530 1656.180 1288.850 1656.440 ;
        RECT 1521.290 1656.380 1521.610 1656.440 ;
        RECT 1520.920 1656.240 1521.610 1656.380 ;
        RECT 1288.620 1655.700 1288.760 1656.180 ;
        RECT 1520.920 1656.100 1521.060 1656.240 ;
        RECT 1521.290 1656.180 1521.610 1656.240 ;
        RECT 1520.830 1655.840 1521.150 1656.100 ;
        RECT 2518.110 1656.040 2518.430 1656.100 ;
        RECT 2519.950 1656.040 2520.270 1656.100 ;
        RECT 2518.110 1655.900 2520.270 1656.040 ;
        RECT 2518.110 1655.840 2518.430 1655.900 ;
        RECT 2519.950 1655.840 2520.270 1655.900 ;
        RECT 1288.990 1655.700 1289.310 1655.760 ;
        RECT 1288.620 1655.560 1289.310 1655.700 ;
        RECT 1288.990 1655.500 1289.310 1655.560 ;
        RECT 1441.710 1642.440 1442.030 1642.500 ;
        RECT 1443.090 1642.440 1443.410 1642.500 ;
        RECT 1441.710 1642.300 1443.410 1642.440 ;
        RECT 1441.710 1642.240 1442.030 1642.300 ;
        RECT 1443.090 1642.240 1443.410 1642.300 ;
        RECT 2517.650 1642.100 2517.970 1642.160 ;
        RECT 2518.570 1642.100 2518.890 1642.160 ;
        RECT 2517.650 1641.960 2518.890 1642.100 ;
        RECT 2517.650 1641.900 2517.970 1641.960 ;
        RECT 2518.570 1641.900 2518.890 1641.960 ;
        RECT 1441.710 1617.960 1442.030 1618.020 ;
        RECT 1442.630 1617.960 1442.950 1618.020 ;
        RECT 1441.710 1617.820 1442.950 1617.960 ;
        RECT 1441.710 1617.760 1442.030 1617.820 ;
        RECT 1442.630 1617.760 1442.950 1617.820 ;
        RECT 2519.950 1617.960 2520.270 1618.020 ;
        RECT 2520.870 1617.960 2521.190 1618.020 ;
        RECT 2519.950 1617.820 2521.190 1617.960 ;
        RECT 2519.950 1617.760 2520.270 1617.820 ;
        RECT 2520.870 1617.760 2521.190 1617.820 ;
        RECT 1520.830 1607.760 1521.150 1607.820 ;
        RECT 1521.290 1607.760 1521.610 1607.820 ;
        RECT 1520.830 1607.620 1521.610 1607.760 ;
        RECT 1520.830 1607.560 1521.150 1607.620 ;
        RECT 1521.290 1607.560 1521.610 1607.620 ;
        RECT 1288.990 1594.980 1289.310 1595.240 ;
        RECT 1289.080 1593.880 1289.220 1594.980 ;
        RECT 1441.710 1594.160 1442.030 1594.220 ;
        RECT 1442.630 1594.160 1442.950 1594.220 ;
        RECT 1441.710 1594.020 1442.950 1594.160 ;
        RECT 1441.710 1593.960 1442.030 1594.020 ;
        RECT 1442.630 1593.960 1442.950 1594.020 ;
        RECT 2517.650 1594.160 2517.970 1594.220 ;
        RECT 2518.570 1594.160 2518.890 1594.220 ;
        RECT 2517.650 1594.020 2518.890 1594.160 ;
        RECT 2517.650 1593.960 2517.970 1594.020 ;
        RECT 2518.570 1593.960 2518.890 1594.020 ;
        RECT 2519.950 1594.160 2520.270 1594.220 ;
        RECT 2520.870 1594.160 2521.190 1594.220 ;
        RECT 2519.950 1594.020 2521.190 1594.160 ;
        RECT 2519.950 1593.960 2520.270 1594.020 ;
        RECT 2520.870 1593.960 2521.190 1594.020 ;
        RECT 1288.990 1593.620 1289.310 1593.880 ;
        RECT 1521.290 1593.820 1521.610 1593.880 ;
        RECT 1522.670 1593.820 1522.990 1593.880 ;
        RECT 1521.290 1593.680 1522.990 1593.820 ;
        RECT 1521.290 1593.620 1521.610 1593.680 ;
        RECT 1522.670 1593.620 1522.990 1593.680 ;
        RECT 1288.990 1587.020 1289.310 1587.080 ;
        RECT 1290.370 1587.020 1290.690 1587.080 ;
        RECT 1288.990 1586.880 1290.690 1587.020 ;
        RECT 1288.990 1586.820 1289.310 1586.880 ;
        RECT 1290.370 1586.820 1290.690 1586.880 ;
        RECT 1440.330 1569.680 1440.650 1569.740 ;
        RECT 1441.710 1569.680 1442.030 1569.740 ;
        RECT 1440.330 1569.540 1442.030 1569.680 ;
        RECT 1440.330 1569.480 1440.650 1569.540 ;
        RECT 1441.710 1569.480 1442.030 1569.540 ;
        RECT 2517.190 1569.680 2517.510 1569.740 ;
        RECT 2518.570 1569.680 2518.890 1569.740 ;
        RECT 2517.190 1569.540 2518.890 1569.680 ;
        RECT 2517.190 1569.480 2517.510 1569.540 ;
        RECT 2518.570 1569.480 2518.890 1569.540 ;
        RECT 2518.110 1559.480 2518.430 1559.540 ;
        RECT 2519.950 1559.480 2520.270 1559.540 ;
        RECT 2518.110 1559.340 2520.270 1559.480 ;
        RECT 2518.110 1559.280 2518.430 1559.340 ;
        RECT 2519.950 1559.280 2520.270 1559.340 ;
        RECT 1288.990 1558.800 1289.310 1558.860 ;
        RECT 1290.370 1558.800 1290.690 1558.860 ;
        RECT 1288.990 1558.660 1290.690 1558.800 ;
        RECT 1288.990 1558.600 1289.310 1558.660 ;
        RECT 1290.370 1558.600 1290.690 1558.660 ;
        RECT 2518.110 1558.800 2518.430 1558.860 ;
        RECT 2519.950 1558.800 2520.270 1558.860 ;
        RECT 2518.110 1558.660 2520.270 1558.800 ;
        RECT 2518.110 1558.600 2518.430 1558.660 ;
        RECT 2519.950 1558.600 2520.270 1558.660 ;
        RECT 1521.290 1546.220 1521.610 1546.280 ;
        RECT 1522.670 1546.220 1522.990 1546.280 ;
        RECT 1521.290 1546.080 1522.990 1546.220 ;
        RECT 1521.290 1546.020 1521.610 1546.080 ;
        RECT 1522.670 1546.020 1522.990 1546.080 ;
        RECT 1440.330 1545.880 1440.650 1545.940 ;
        RECT 1440.790 1545.880 1441.110 1545.940 ;
        RECT 1440.330 1545.740 1441.110 1545.880 ;
        RECT 1440.330 1545.680 1440.650 1545.740 ;
        RECT 1440.790 1545.680 1441.110 1545.740 ;
        RECT 2517.190 1545.880 2517.510 1545.940 ;
        RECT 2519.030 1545.880 2519.350 1545.940 ;
        RECT 2517.190 1545.740 2519.350 1545.880 ;
        RECT 2517.190 1545.680 2517.510 1545.740 ;
        RECT 2519.030 1545.680 2519.350 1545.740 ;
        RECT 1521.290 1545.540 1521.610 1545.600 ;
        RECT 1522.210 1545.540 1522.530 1545.600 ;
        RECT 1521.290 1545.400 1522.530 1545.540 ;
        RECT 1521.290 1545.340 1521.610 1545.400 ;
        RECT 1522.210 1545.340 1522.530 1545.400 ;
        RECT 1440.330 1545.200 1440.650 1545.260 ;
        RECT 1440.790 1545.200 1441.110 1545.260 ;
        RECT 1440.330 1545.060 1441.110 1545.200 ;
        RECT 1440.330 1545.000 1440.650 1545.060 ;
        RECT 1440.790 1545.000 1441.110 1545.060 ;
        RECT 1288.530 1538.740 1288.850 1538.800 ;
        RECT 1288.990 1538.740 1289.310 1538.800 ;
        RECT 1288.530 1538.600 1289.310 1538.740 ;
        RECT 1288.530 1538.540 1288.850 1538.600 ;
        RECT 1288.990 1538.540 1289.310 1538.600 ;
        RECT 1440.330 1497.600 1440.650 1497.660 ;
        RECT 1441.710 1497.600 1442.030 1497.660 ;
        RECT 1440.330 1497.460 1442.030 1497.600 ;
        RECT 1440.330 1497.400 1440.650 1497.460 ;
        RECT 1441.710 1497.400 1442.030 1497.460 ;
        RECT 1521.290 1497.260 1521.610 1497.320 ;
        RECT 1522.670 1497.260 1522.990 1497.320 ;
        RECT 1521.290 1497.120 1522.990 1497.260 ;
        RECT 1521.290 1497.060 1521.610 1497.120 ;
        RECT 1522.670 1497.060 1522.990 1497.120 ;
        RECT 1288.530 1490.800 1288.850 1490.860 ;
        RECT 1289.450 1490.800 1289.770 1490.860 ;
        RECT 1288.530 1490.660 1289.770 1490.800 ;
        RECT 1288.530 1490.600 1288.850 1490.660 ;
        RECT 1289.450 1490.600 1289.770 1490.660 ;
        RECT 1440.330 1473.120 1440.650 1473.180 ;
        RECT 1441.710 1473.120 1442.030 1473.180 ;
        RECT 1440.330 1472.980 1442.030 1473.120 ;
        RECT 1440.330 1472.920 1440.650 1472.980 ;
        RECT 1441.710 1472.920 1442.030 1472.980 ;
        RECT 1521.290 1449.660 1521.610 1449.720 ;
        RECT 1522.670 1449.660 1522.990 1449.720 ;
        RECT 1521.290 1449.520 1522.990 1449.660 ;
        RECT 1521.290 1449.460 1521.610 1449.520 ;
        RECT 1522.670 1449.460 1522.990 1449.520 ;
        RECT 1440.330 1449.320 1440.650 1449.380 ;
        RECT 1440.790 1449.320 1441.110 1449.380 ;
        RECT 1440.330 1449.180 1441.110 1449.320 ;
        RECT 1440.330 1449.120 1440.650 1449.180 ;
        RECT 1440.790 1449.120 1441.110 1449.180 ;
        RECT 1521.290 1448.980 1521.610 1449.040 ;
        RECT 1522.210 1448.980 1522.530 1449.040 ;
        RECT 1521.290 1448.840 1522.530 1448.980 ;
        RECT 1521.290 1448.780 1521.610 1448.840 ;
        RECT 1522.210 1448.780 1522.530 1448.840 ;
        RECT 1440.790 1448.640 1441.110 1448.700 ;
        RECT 1442.630 1448.640 1442.950 1448.700 ;
        RECT 1440.790 1448.500 1442.950 1448.640 ;
        RECT 1440.790 1448.440 1441.110 1448.500 ;
        RECT 1442.630 1448.440 1442.950 1448.500 ;
        RECT 1288.990 1442.180 1289.310 1442.240 ;
        RECT 1289.450 1442.180 1289.770 1442.240 ;
        RECT 1288.990 1442.040 1289.770 1442.180 ;
        RECT 1288.990 1441.980 1289.310 1442.040 ;
        RECT 1289.450 1441.980 1289.770 1442.040 ;
        RECT 2518.570 1415.320 2518.890 1415.380 ;
        RECT 2518.570 1415.180 2519.260 1415.320 ;
        RECT 2518.570 1415.120 2518.890 1415.180 ;
        RECT 2519.120 1415.040 2519.260 1415.180 ;
        RECT 2519.030 1414.780 2519.350 1415.040 ;
        RECT 1288.990 1414.640 1289.310 1414.700 ;
        RECT 1289.910 1414.640 1290.230 1414.700 ;
        RECT 1288.990 1414.500 1290.230 1414.640 ;
        RECT 1288.990 1414.440 1289.310 1414.500 ;
        RECT 1289.910 1414.440 1290.230 1414.500 ;
        RECT 1521.290 1400.700 1521.610 1400.760 ;
        RECT 1522.670 1400.700 1522.990 1400.760 ;
        RECT 1521.290 1400.560 1522.990 1400.700 ;
        RECT 1521.290 1400.500 1521.610 1400.560 ;
        RECT 1522.670 1400.500 1522.990 1400.560 ;
        RECT 1441.710 1387.100 1442.030 1387.160 ;
        RECT 1442.630 1387.100 1442.950 1387.160 ;
        RECT 1441.710 1386.960 1442.950 1387.100 ;
        RECT 1441.710 1386.900 1442.030 1386.960 ;
        RECT 1442.630 1386.900 1442.950 1386.960 ;
        RECT 2518.110 1366.700 2518.430 1366.760 ;
        RECT 2519.950 1366.700 2520.270 1366.760 ;
        RECT 2518.110 1366.560 2520.270 1366.700 ;
        RECT 2518.110 1366.500 2518.430 1366.560 ;
        RECT 2519.950 1366.500 2520.270 1366.560 ;
        RECT 2518.110 1366.020 2518.430 1366.080 ;
        RECT 2519.950 1366.020 2520.270 1366.080 ;
        RECT 2518.110 1365.880 2520.270 1366.020 ;
        RECT 2518.110 1365.820 2518.430 1365.880 ;
        RECT 2519.950 1365.820 2520.270 1365.880 ;
        RECT 1521.290 1353.100 1521.610 1353.160 ;
        RECT 1522.670 1353.100 1522.990 1353.160 ;
        RECT 1521.290 1352.960 1522.990 1353.100 ;
        RECT 1521.290 1352.900 1521.610 1352.960 ;
        RECT 1522.670 1352.900 1522.990 1352.960 ;
        RECT 1288.990 1352.420 1289.310 1352.480 ;
        RECT 1289.910 1352.420 1290.230 1352.480 ;
        RECT 1288.990 1352.280 1290.230 1352.420 ;
        RECT 1288.990 1352.220 1289.310 1352.280 ;
        RECT 1289.910 1352.220 1290.230 1352.280 ;
        RECT 1521.290 1352.420 1521.610 1352.480 ;
        RECT 1522.670 1352.420 1522.990 1352.480 ;
        RECT 1521.290 1352.280 1522.990 1352.420 ;
        RECT 1521.290 1352.220 1521.610 1352.280 ;
        RECT 1522.670 1352.220 1522.990 1352.280 ;
        RECT 2518.570 1318.420 2518.890 1318.480 ;
        RECT 2519.950 1318.420 2520.270 1318.480 ;
        RECT 2518.570 1318.280 2520.270 1318.420 ;
        RECT 2518.570 1318.220 2518.890 1318.280 ;
        RECT 2519.950 1318.220 2520.270 1318.280 ;
        RECT 1288.990 1317.740 1289.310 1317.800 ;
        RECT 1289.910 1317.740 1290.230 1317.800 ;
        RECT 1288.990 1317.600 1290.230 1317.740 ;
        RECT 1288.990 1317.540 1289.310 1317.600 ;
        RECT 1289.910 1317.540 1290.230 1317.600 ;
        RECT 2518.570 1317.740 2518.890 1317.800 ;
        RECT 2519.950 1317.740 2520.270 1317.800 ;
        RECT 2518.570 1317.600 2520.270 1317.740 ;
        RECT 2518.570 1317.540 2518.890 1317.600 ;
        RECT 2519.950 1317.540 2520.270 1317.600 ;
        RECT 1521.290 1317.400 1521.610 1317.460 ;
        RECT 1522.670 1317.400 1522.990 1317.460 ;
        RECT 1521.290 1317.260 1522.990 1317.400 ;
        RECT 1521.290 1317.200 1521.610 1317.260 ;
        RECT 1522.670 1317.200 1522.990 1317.260 ;
        RECT 1288.990 1304.140 1289.310 1304.200 ;
        RECT 1290.370 1304.140 1290.690 1304.200 ;
        RECT 1288.990 1304.000 1290.690 1304.140 ;
        RECT 1288.990 1303.940 1289.310 1304.000 ;
        RECT 1290.370 1303.940 1290.690 1304.000 ;
        RECT 1521.290 1304.140 1521.610 1304.200 ;
        RECT 1522.670 1304.140 1522.990 1304.200 ;
        RECT 1521.290 1304.000 1522.990 1304.140 ;
        RECT 1521.290 1303.940 1521.610 1304.000 ;
        RECT 1522.670 1303.940 1522.990 1304.000 ;
        RECT 1440.790 1290.200 1441.110 1290.260 ;
        RECT 1441.710 1290.200 1442.030 1290.260 ;
        RECT 1440.790 1290.060 1442.030 1290.200 ;
        RECT 1440.790 1290.000 1441.110 1290.060 ;
        RECT 1441.710 1290.000 1442.030 1290.060 ;
        RECT 2518.110 1270.140 2518.430 1270.200 ;
        RECT 2519.950 1270.140 2520.270 1270.200 ;
        RECT 2518.110 1270.000 2520.270 1270.140 ;
        RECT 2518.110 1269.940 2518.430 1270.000 ;
        RECT 2519.950 1269.940 2520.270 1270.000 ;
        RECT 2518.110 1269.460 2518.430 1269.520 ;
        RECT 2519.950 1269.460 2520.270 1269.520 ;
        RECT 2518.110 1269.320 2520.270 1269.460 ;
        RECT 2518.110 1269.260 2518.430 1269.320 ;
        RECT 2519.950 1269.260 2520.270 1269.320 ;
        RECT 1288.990 1269.120 1289.310 1269.180 ;
        RECT 1290.370 1269.120 1290.690 1269.180 ;
        RECT 1288.990 1268.980 1290.690 1269.120 ;
        RECT 1288.990 1268.920 1289.310 1268.980 ;
        RECT 1290.370 1268.920 1290.690 1268.980 ;
        RECT 1287.610 1255.860 1287.930 1255.920 ;
        RECT 1288.990 1255.860 1289.310 1255.920 ;
        RECT 1287.610 1255.720 1289.310 1255.860 ;
        RECT 1287.610 1255.660 1287.930 1255.720 ;
        RECT 1288.990 1255.660 1289.310 1255.720 ;
        RECT 1440.330 1242.260 1440.650 1242.320 ;
        RECT 1440.790 1242.260 1441.110 1242.320 ;
        RECT 1440.330 1242.120 1441.110 1242.260 ;
        RECT 1440.330 1242.060 1440.650 1242.120 ;
        RECT 1440.790 1242.060 1441.110 1242.120 ;
        RECT 2518.570 1222.200 2518.890 1222.260 ;
        RECT 2518.570 1222.060 2519.260 1222.200 ;
        RECT 2518.570 1222.000 2518.890 1222.060 ;
        RECT 2519.120 1221.920 2519.260 1222.060 ;
        RECT 2519.030 1221.660 2519.350 1221.920 ;
        RECT 1440.330 1220.840 1440.650 1220.900 ;
        RECT 1441.710 1220.840 1442.030 1220.900 ;
        RECT 1440.330 1220.700 1442.030 1220.840 ;
        RECT 1440.330 1220.640 1440.650 1220.700 ;
        RECT 1441.710 1220.640 1442.030 1220.700 ;
        RECT 1287.610 1207.580 1287.930 1207.640 ;
        RECT 1288.530 1207.580 1288.850 1207.640 ;
        RECT 1287.610 1207.440 1288.850 1207.580 ;
        RECT 1287.610 1207.380 1287.930 1207.440 ;
        RECT 1288.530 1207.380 1288.850 1207.440 ;
        RECT 1520.830 1207.580 1521.150 1207.640 ;
        RECT 1521.750 1207.580 1522.070 1207.640 ;
        RECT 1520.830 1207.440 1522.070 1207.580 ;
        RECT 1520.830 1207.380 1521.150 1207.440 ;
        RECT 1521.750 1207.380 1522.070 1207.440 ;
        RECT 1519.450 1206.900 1519.770 1206.960 ;
        RECT 1520.830 1206.900 1521.150 1206.960 ;
        RECT 1519.450 1206.760 1521.150 1206.900 ;
        RECT 1519.450 1206.700 1519.770 1206.760 ;
        RECT 1520.830 1206.700 1521.150 1206.760 ;
        RECT 2518.110 1173.580 2518.430 1173.640 ;
        RECT 2519.950 1173.580 2520.270 1173.640 ;
        RECT 2518.110 1173.440 2520.270 1173.580 ;
        RECT 2518.110 1173.380 2518.430 1173.440 ;
        RECT 2519.950 1173.380 2520.270 1173.440 ;
        RECT 1288.530 1173.040 1288.850 1173.300 ;
        RECT 1288.620 1172.560 1288.760 1173.040 ;
        RECT 2518.110 1172.900 2518.430 1172.960 ;
        RECT 2519.950 1172.900 2520.270 1172.960 ;
        RECT 2518.110 1172.760 2520.270 1172.900 ;
        RECT 2518.110 1172.700 2518.430 1172.760 ;
        RECT 2519.950 1172.700 2520.270 1172.760 ;
        RECT 1288.990 1172.560 1289.310 1172.620 ;
        RECT 1288.620 1172.420 1289.310 1172.560 ;
        RECT 1288.990 1172.360 1289.310 1172.420 ;
        RECT 1519.450 1159.300 1519.770 1159.360 ;
        RECT 1520.830 1159.300 1521.150 1159.360 ;
        RECT 1519.450 1159.160 1521.150 1159.300 ;
        RECT 1519.450 1159.100 1519.770 1159.160 ;
        RECT 1520.830 1159.100 1521.150 1159.160 ;
        RECT 2518.570 1125.640 2518.890 1125.700 ;
        RECT 2518.570 1125.500 2519.260 1125.640 ;
        RECT 2518.570 1125.440 2518.890 1125.500 ;
        RECT 2519.120 1125.360 2519.260 1125.500 ;
        RECT 2519.030 1125.100 2519.350 1125.360 ;
        RECT 1288.530 1124.960 1288.850 1125.020 ;
        RECT 1521.290 1124.960 1521.610 1125.020 ;
        RECT 1288.530 1124.820 1289.220 1124.960 ;
        RECT 1288.530 1124.760 1288.850 1124.820 ;
        RECT 1289.080 1124.680 1289.220 1124.820 ;
        RECT 1521.290 1124.820 1521.980 1124.960 ;
        RECT 1521.290 1124.760 1521.610 1124.820 ;
        RECT 1288.990 1124.420 1289.310 1124.680 ;
        RECT 1521.840 1124.340 1521.980 1124.820 ;
        RECT 1521.750 1124.080 1522.070 1124.340 ;
        RECT 1288.530 1111.020 1288.850 1111.080 ;
        RECT 1288.990 1111.020 1289.310 1111.080 ;
        RECT 1288.530 1110.880 1289.310 1111.020 ;
        RECT 1288.530 1110.820 1288.850 1110.880 ;
        RECT 1288.990 1110.820 1289.310 1110.880 ;
        RECT 1441.710 1111.020 1442.030 1111.080 ;
        RECT 1442.630 1111.020 1442.950 1111.080 ;
        RECT 1441.710 1110.880 1442.950 1111.020 ;
        RECT 1441.710 1110.820 1442.030 1110.880 ;
        RECT 1442.630 1110.820 1442.950 1110.880 ;
        RECT 1520.370 1080.080 1520.690 1080.140 ;
        RECT 1521.290 1080.080 1521.610 1080.140 ;
        RECT 1520.370 1079.940 1521.610 1080.080 ;
        RECT 1520.370 1079.880 1520.690 1079.940 ;
        RECT 1521.290 1079.880 1521.610 1079.940 ;
        RECT 2518.110 1077.020 2518.430 1077.080 ;
        RECT 2519.950 1077.020 2520.270 1077.080 ;
        RECT 2518.110 1076.880 2520.270 1077.020 ;
        RECT 2518.110 1076.820 2518.430 1076.880 ;
        RECT 2519.950 1076.820 2520.270 1076.880 ;
        RECT 1288.530 1076.480 1288.850 1076.740 ;
        RECT 1288.620 1076.000 1288.760 1076.480 ;
        RECT 2518.110 1076.340 2518.430 1076.400 ;
        RECT 2519.950 1076.340 2520.270 1076.400 ;
        RECT 2518.110 1076.200 2520.270 1076.340 ;
        RECT 2518.110 1076.140 2518.430 1076.200 ;
        RECT 2519.950 1076.140 2520.270 1076.200 ;
        RECT 1288.990 1076.000 1289.310 1076.060 ;
        RECT 1288.620 1075.860 1289.310 1076.000 ;
        RECT 1288.990 1075.800 1289.310 1075.860 ;
        RECT 1440.330 1062.740 1440.650 1062.800 ;
        RECT 1440.790 1062.740 1441.110 1062.800 ;
        RECT 1440.330 1062.600 1441.110 1062.740 ;
        RECT 1440.330 1062.540 1440.650 1062.600 ;
        RECT 1440.790 1062.540 1441.110 1062.600 ;
        RECT 2082.030 1062.740 2082.350 1062.800 ;
        RECT 2083.410 1062.740 2083.730 1062.800 ;
        RECT 2082.030 1062.600 2083.730 1062.740 ;
        RECT 2082.030 1062.540 2082.350 1062.600 ;
        RECT 2083.410 1062.540 2083.730 1062.600 ;
        RECT 1454.590 1052.200 1454.910 1052.260 ;
        RECT 1455.510 1052.200 1455.830 1052.260 ;
        RECT 1454.590 1052.060 1455.830 1052.200 ;
        RECT 1454.590 1052.000 1454.910 1052.060 ;
        RECT 1455.510 1052.000 1455.830 1052.060 ;
        RECT 1062.210 1051.860 1062.530 1051.920 ;
        RECT 1098.550 1051.860 1098.870 1051.920 ;
        RECT 1062.210 1051.720 1098.870 1051.860 ;
        RECT 1062.210 1051.660 1062.530 1051.720 ;
        RECT 1098.550 1051.660 1098.870 1051.720 ;
        RECT 1219.990 1048.800 1220.310 1048.860 ;
        RECT 1220.910 1048.800 1221.230 1048.860 ;
        RECT 1219.990 1048.660 1221.230 1048.800 ;
        RECT 1219.990 1048.600 1220.310 1048.660 ;
        RECT 1220.910 1048.600 1221.230 1048.660 ;
        RECT 2518.570 1029.080 2518.890 1029.140 ;
        RECT 2518.570 1028.940 2519.260 1029.080 ;
        RECT 2518.570 1028.880 2518.890 1028.940 ;
        RECT 2519.120 1028.800 2519.260 1028.940 ;
        RECT 2519.030 1028.540 2519.350 1028.800 ;
        RECT 632.110 1028.400 632.430 1028.460 ;
        RECT 1288.530 1028.400 1288.850 1028.460 ;
        RECT 2518.570 1028.400 2518.890 1028.460 ;
        RECT 2519.950 1028.400 2520.270 1028.460 ;
        RECT 632.110 1028.260 633.260 1028.400 ;
        RECT 632.110 1028.200 632.430 1028.260 ;
        RECT 632.110 1027.720 632.430 1027.780 ;
        RECT 633.120 1027.720 633.260 1028.260 ;
        RECT 1288.530 1028.260 1289.220 1028.400 ;
        RECT 1288.530 1028.200 1288.850 1028.260 ;
        RECT 1289.080 1028.120 1289.220 1028.260 ;
        RECT 2518.570 1028.260 2520.270 1028.400 ;
        RECT 2518.570 1028.200 2518.890 1028.260 ;
        RECT 2519.950 1028.200 2520.270 1028.260 ;
        RECT 1288.990 1027.860 1289.310 1028.120 ;
        RECT 632.110 1027.580 633.260 1027.720 ;
        RECT 632.110 1027.520 632.430 1027.580 ;
        RECT 983.550 1026.700 983.870 1026.760 ;
        RECT 1134.430 1026.700 1134.750 1026.760 ;
        RECT 983.550 1026.560 1134.750 1026.700 ;
        RECT 983.550 1026.500 983.870 1026.560 ;
        RECT 1134.430 1026.500 1134.750 1026.560 ;
        RECT 983.090 1026.360 983.410 1026.420 ;
        RECT 1139.490 1026.360 1139.810 1026.420 ;
        RECT 983.090 1026.220 1139.810 1026.360 ;
        RECT 983.090 1026.160 983.410 1026.220 ;
        RECT 1139.490 1026.160 1139.810 1026.220 ;
        RECT 979.410 1026.020 979.730 1026.080 ;
        RECT 1143.170 1026.020 1143.490 1026.080 ;
        RECT 979.410 1025.880 1143.490 1026.020 ;
        RECT 979.410 1025.820 979.730 1025.880 ;
        RECT 1143.170 1025.820 1143.490 1025.880 ;
        RECT 978.490 1025.680 978.810 1025.740 ;
        RECT 1147.770 1025.680 1148.090 1025.740 ;
        RECT 978.490 1025.540 1148.090 1025.680 ;
        RECT 978.490 1025.480 978.810 1025.540 ;
        RECT 1147.770 1025.480 1148.090 1025.540 ;
        RECT 978.950 1025.340 979.270 1025.400 ;
        RECT 1152.370 1025.340 1152.690 1025.400 ;
        RECT 978.950 1025.200 1152.690 1025.340 ;
        RECT 978.950 1025.140 979.270 1025.200 ;
        RECT 1152.370 1025.140 1152.690 1025.200 ;
        RECT 1196.070 1025.340 1196.390 1025.400 ;
        RECT 1200.210 1025.340 1200.530 1025.400 ;
        RECT 1196.070 1025.200 1200.530 1025.340 ;
        RECT 1196.070 1025.140 1196.390 1025.200 ;
        RECT 1200.210 1025.140 1200.530 1025.200 ;
        RECT 977.570 1025.000 977.890 1025.060 ;
        RECT 1156.050 1025.000 1156.370 1025.060 ;
        RECT 977.570 1024.860 1156.370 1025.000 ;
        RECT 977.570 1024.800 977.890 1024.860 ;
        RECT 1156.050 1024.800 1156.370 1024.860 ;
        RECT 978.030 1024.660 978.350 1024.720 ;
        RECT 1166.170 1024.660 1166.490 1024.720 ;
        RECT 978.030 1024.520 1166.490 1024.660 ;
        RECT 978.030 1024.460 978.350 1024.520 ;
        RECT 1166.170 1024.460 1166.490 1024.520 ;
        RECT 1472.070 1021.260 1472.390 1021.320 ;
        RECT 1704.370 1021.260 1704.690 1021.320 ;
        RECT 1472.070 1021.120 1704.690 1021.260 ;
        RECT 1472.070 1021.060 1472.390 1021.120 ;
        RECT 1704.370 1021.060 1704.690 1021.120 ;
        RECT 1728.750 1021.260 1729.070 1021.320 ;
        RECT 2085.250 1021.260 2085.570 1021.320 ;
        RECT 1728.750 1021.120 2085.570 1021.260 ;
        RECT 1728.750 1021.060 1729.070 1021.120 ;
        RECT 2085.250 1021.060 2085.570 1021.120 ;
        RECT 1278.870 1020.920 1279.190 1020.980 ;
        RECT 1340.970 1020.920 1341.290 1020.980 ;
        RECT 1278.870 1020.780 1341.290 1020.920 ;
        RECT 1278.870 1020.720 1279.190 1020.780 ;
        RECT 1340.970 1020.720 1341.290 1020.780 ;
        RECT 1489.550 1020.920 1489.870 1020.980 ;
        RECT 1521.290 1020.920 1521.610 1020.980 ;
        RECT 1489.550 1020.780 1521.610 1020.920 ;
        RECT 1489.550 1020.720 1489.870 1020.780 ;
        RECT 1521.290 1020.720 1521.610 1020.780 ;
        RECT 1533.250 1020.920 1533.570 1020.980 ;
        RECT 1902.170 1020.920 1902.490 1020.980 ;
        RECT 1533.250 1020.780 1902.490 1020.920 ;
        RECT 1533.250 1020.720 1533.570 1020.780 ;
        RECT 1902.170 1020.720 1902.490 1020.780 ;
        RECT 1267.830 1020.580 1268.150 1020.640 ;
        RECT 1345.110 1020.580 1345.430 1020.640 ;
        RECT 1267.830 1020.440 1345.430 1020.580 ;
        RECT 1267.830 1020.380 1268.150 1020.440 ;
        RECT 1345.110 1020.380 1345.430 1020.440 ;
        RECT 1507.030 1020.580 1507.350 1020.640 ;
        RECT 1898.030 1020.580 1898.350 1020.640 ;
        RECT 1507.030 1020.440 1898.350 1020.580 ;
        RECT 1507.030 1020.380 1507.350 1020.440 ;
        RECT 1898.030 1020.380 1898.350 1020.440 ;
        RECT 1252.650 1020.240 1252.970 1020.300 ;
        RECT 1339.590 1020.240 1339.910 1020.300 ;
        RECT 1252.650 1020.100 1339.910 1020.240 ;
        RECT 1252.650 1020.040 1252.970 1020.100 ;
        RECT 1339.590 1020.040 1339.910 1020.100 ;
        RECT 1495.070 1020.240 1495.390 1020.300 ;
        RECT 1901.710 1020.240 1902.030 1020.300 ;
        RECT 1495.070 1020.100 1902.030 1020.240 ;
        RECT 1495.070 1020.040 1495.390 1020.100 ;
        RECT 1901.710 1020.040 1902.030 1020.100 ;
        RECT 995.050 1019.900 995.370 1019.960 ;
        RECT 1193.770 1019.900 1194.090 1019.960 ;
        RECT 995.050 1019.760 1194.090 1019.900 ;
        RECT 995.050 1019.700 995.370 1019.760 ;
        RECT 1193.770 1019.700 1194.090 1019.760 ;
        RECT 1237.930 1019.900 1238.250 1019.960 ;
        RECT 1340.510 1019.900 1340.830 1019.960 ;
        RECT 1237.930 1019.760 1340.830 1019.900 ;
        RECT 1237.930 1019.700 1238.250 1019.760 ;
        RECT 1340.510 1019.700 1340.830 1019.760 ;
        RECT 1474.370 1019.900 1474.690 1019.960 ;
        RECT 1886.990 1019.900 1887.310 1019.960 ;
        RECT 1474.370 1019.760 1887.310 1019.900 ;
        RECT 1474.370 1019.700 1474.690 1019.760 ;
        RECT 1886.990 1019.700 1887.310 1019.760 ;
        RECT 988.610 1019.560 988.930 1019.620 ;
        RECT 1285.770 1019.560 1286.090 1019.620 ;
        RECT 988.610 1019.420 1286.090 1019.560 ;
        RECT 988.610 1019.360 988.930 1019.420 ;
        RECT 1285.770 1019.360 1286.090 1019.420 ;
        RECT 1461.030 1019.560 1461.350 1019.620 ;
        RECT 1898.950 1019.560 1899.270 1019.620 ;
        RECT 1461.030 1019.420 1899.270 1019.560 ;
        RECT 1461.030 1019.360 1461.350 1019.420 ;
        RECT 1898.950 1019.360 1899.270 1019.420 ;
        RECT 989.990 1019.220 990.310 1019.280 ;
        RECT 1301.870 1019.220 1302.190 1019.280 ;
        RECT 989.990 1019.080 1302.190 1019.220 ;
        RECT 989.990 1019.020 990.310 1019.080 ;
        RECT 1301.870 1019.020 1302.190 1019.080 ;
        RECT 1462.410 1019.220 1462.730 1019.280 ;
        RECT 1899.410 1019.220 1899.730 1019.280 ;
        RECT 1462.410 1019.080 1899.730 1019.220 ;
        RECT 1462.410 1019.020 1462.730 1019.080 ;
        RECT 1899.410 1019.020 1899.730 1019.080 ;
        RECT 992.290 1018.880 992.610 1018.940 ;
        RECT 1313.830 1018.880 1314.150 1018.940 ;
        RECT 992.290 1018.740 1314.150 1018.880 ;
        RECT 992.290 1018.680 992.610 1018.740 ;
        RECT 1313.830 1018.680 1314.150 1018.740 ;
        RECT 1434.810 1018.880 1435.130 1018.940 ;
        RECT 1886.530 1018.880 1886.850 1018.940 ;
        RECT 1434.810 1018.740 1886.850 1018.880 ;
        RECT 1434.810 1018.680 1435.130 1018.740 ;
        RECT 1886.530 1018.680 1886.850 1018.740 ;
        RECT 987.230 1018.540 987.550 1018.600 ;
        RECT 1314.750 1018.540 1315.070 1018.600 ;
        RECT 987.230 1018.400 1315.070 1018.540 ;
        RECT 987.230 1018.340 987.550 1018.400 ;
        RECT 1314.750 1018.340 1315.070 1018.400 ;
        RECT 1437.570 1018.540 1437.890 1018.600 ;
        RECT 1898.490 1018.540 1898.810 1018.600 ;
        RECT 1437.570 1018.400 1898.810 1018.540 ;
        RECT 1437.570 1018.340 1437.890 1018.400 ;
        RECT 1898.490 1018.340 1898.810 1018.400 ;
        RECT 989.070 1018.200 989.390 1018.260 ;
        RECT 1326.250 1018.200 1326.570 1018.260 ;
        RECT 989.070 1018.060 1326.570 1018.200 ;
        RECT 989.070 1018.000 989.390 1018.060 ;
        RECT 1326.250 1018.000 1326.570 1018.060 ;
        RECT 1358.910 1018.200 1359.230 1018.260 ;
        RECT 1849.270 1018.200 1849.590 1018.260 ;
        RECT 1358.910 1018.060 1849.590 1018.200 ;
        RECT 1358.910 1018.000 1359.230 1018.060 ;
        RECT 1849.270 1018.000 1849.590 1018.060 ;
        RECT 991.830 1017.860 992.150 1017.920 ;
        RECT 1337.750 1017.860 1338.070 1017.920 ;
        RECT 991.830 1017.720 1338.070 1017.860 ;
        RECT 991.830 1017.660 992.150 1017.720 ;
        RECT 1337.750 1017.660 1338.070 1017.720 ;
        RECT 1402.610 1017.860 1402.930 1017.920 ;
        RECT 1899.870 1017.860 1900.190 1017.920 ;
        RECT 1402.610 1017.720 1900.190 1017.860 ;
        RECT 1402.610 1017.660 1402.930 1017.720 ;
        RECT 1899.870 1017.660 1900.190 1017.720 ;
        RECT 1567.750 1017.520 1568.070 1017.580 ;
        RECT 1897.570 1017.520 1897.890 1017.580 ;
        RECT 1567.750 1017.380 1897.890 1017.520 ;
        RECT 1567.750 1017.320 1568.070 1017.380 ;
        RECT 1897.570 1017.320 1897.890 1017.380 ;
        RECT 1480.810 1017.180 1481.130 1017.240 ;
        RECT 1766.470 1017.180 1766.790 1017.240 ;
        RECT 1480.810 1017.040 1766.790 1017.180 ;
        RECT 1480.810 1016.980 1481.130 1017.040 ;
        RECT 1766.470 1016.980 1766.790 1017.040 ;
        RECT 1614.670 1016.840 1614.990 1016.900 ;
        RECT 1900.790 1016.840 1901.110 1016.900 ;
        RECT 1614.670 1016.700 1901.110 1016.840 ;
        RECT 1614.670 1016.640 1614.990 1016.700 ;
        RECT 1900.790 1016.640 1901.110 1016.700 ;
        RECT 1514.390 1016.500 1514.710 1016.560 ;
        RECT 1656.070 1016.500 1656.390 1016.560 ;
        RECT 1514.390 1016.360 1656.390 1016.500 ;
        RECT 1514.390 1016.300 1514.710 1016.360 ;
        RECT 1656.070 1016.300 1656.390 1016.360 ;
        RECT 1490.010 1016.160 1490.330 1016.220 ;
        RECT 1625.710 1016.160 1626.030 1016.220 ;
        RECT 1490.010 1016.020 1626.030 1016.160 ;
        RECT 1490.010 1015.960 1490.330 1016.020 ;
        RECT 1625.710 1015.960 1626.030 1016.020 ;
        RECT 1288.530 1014.460 1288.850 1014.520 ;
        RECT 1288.990 1014.460 1289.310 1014.520 ;
        RECT 1300.950 1014.460 1301.270 1014.520 ;
        RECT 1288.530 1014.320 1289.310 1014.460 ;
        RECT 1288.530 1014.260 1288.850 1014.320 ;
        RECT 1288.990 1014.260 1289.310 1014.320 ;
        RECT 1293.680 1014.320 1301.270 1014.460 ;
        RECT 810.590 1014.120 810.910 1014.180 ;
        RECT 845.550 1014.120 845.870 1014.180 ;
        RECT 810.590 1013.980 845.870 1014.120 ;
        RECT 810.590 1013.920 810.910 1013.980 ;
        RECT 845.550 1013.920 845.870 1013.980 ;
        RECT 994.590 1014.120 994.910 1014.180 ;
        RECT 997.350 1014.120 997.670 1014.180 ;
        RECT 994.590 1013.980 997.670 1014.120 ;
        RECT 994.590 1013.920 994.910 1013.980 ;
        RECT 997.350 1013.920 997.670 1013.980 ;
        RECT 1000.110 1014.120 1000.430 1014.180 ;
        RECT 1197.910 1014.120 1198.230 1014.180 ;
        RECT 1000.110 1013.980 1198.230 1014.120 ;
        RECT 1000.110 1013.920 1000.430 1013.980 ;
        RECT 1197.910 1013.920 1198.230 1013.980 ;
        RECT 1198.370 1014.120 1198.690 1014.180 ;
        RECT 1200.670 1014.120 1200.990 1014.180 ;
        RECT 1198.370 1013.980 1200.990 1014.120 ;
        RECT 1198.370 1013.920 1198.690 1013.980 ;
        RECT 1200.670 1013.920 1200.990 1013.980 ;
        RECT 1202.510 1014.120 1202.830 1014.180 ;
        RECT 1207.110 1014.120 1207.430 1014.180 ;
        RECT 1202.510 1013.980 1207.430 1014.120 ;
        RECT 1202.510 1013.920 1202.830 1013.980 ;
        RECT 1207.110 1013.920 1207.430 1013.980 ;
        RECT 1214.930 1014.120 1215.250 1014.180 ;
        RECT 1220.450 1014.120 1220.770 1014.180 ;
        RECT 1214.930 1013.980 1220.770 1014.120 ;
        RECT 1214.930 1013.920 1215.250 1013.980 ;
        RECT 1220.450 1013.920 1220.770 1013.980 ;
        RECT 1259.090 1014.120 1259.410 1014.180 ;
        RECT 1284.850 1014.120 1285.170 1014.180 ;
        RECT 1293.680 1014.120 1293.820 1014.320 ;
        RECT 1300.950 1014.260 1301.270 1014.320 ;
        RECT 1494.240 1014.320 1508.180 1014.460 ;
        RECT 1259.090 1013.980 1276.340 1014.120 ;
        RECT 1259.090 1013.920 1259.410 1013.980 ;
        RECT 984.470 1013.780 984.790 1013.840 ;
        RECT 1208.950 1013.780 1209.270 1013.840 ;
        RECT 984.470 1013.640 1209.270 1013.780 ;
        RECT 984.470 1013.580 984.790 1013.640 ;
        RECT 1208.950 1013.580 1209.270 1013.640 ;
        RECT 1262.310 1013.780 1262.630 1013.840 ;
        RECT 1269.210 1013.780 1269.530 1013.840 ;
        RECT 1262.310 1013.640 1269.530 1013.780 ;
        RECT 1276.200 1013.780 1276.340 1013.980 ;
        RECT 1284.850 1013.980 1293.820 1014.120 ;
        RECT 1294.050 1014.120 1294.370 1014.180 ;
        RECT 1333.610 1014.120 1333.930 1014.180 ;
        RECT 1294.050 1013.980 1333.930 1014.120 ;
        RECT 1284.850 1013.920 1285.170 1013.980 ;
        RECT 1294.050 1013.920 1294.370 1013.980 ;
        RECT 1333.610 1013.920 1333.930 1013.980 ;
        RECT 1361.210 1014.120 1361.530 1014.180 ;
        RECT 1365.810 1014.120 1366.130 1014.180 ;
        RECT 1361.210 1013.980 1366.130 1014.120 ;
        RECT 1361.210 1013.920 1361.530 1013.980 ;
        RECT 1365.810 1013.920 1366.130 1013.980 ;
        RECT 1452.750 1014.120 1453.070 1014.180 ;
        RECT 1455.050 1014.120 1455.370 1014.180 ;
        RECT 1452.750 1013.980 1455.370 1014.120 ;
        RECT 1452.750 1013.920 1453.070 1013.980 ;
        RECT 1455.050 1013.920 1455.370 1013.980 ;
        RECT 1456.890 1014.120 1457.210 1014.180 ;
        RECT 1461.490 1014.120 1461.810 1014.180 ;
        RECT 1456.890 1013.980 1461.810 1014.120 ;
        RECT 1456.890 1013.920 1457.210 1013.980 ;
        RECT 1461.490 1013.920 1461.810 1013.980 ;
        RECT 1465.630 1014.120 1465.950 1014.180 ;
        RECT 1472.990 1014.120 1473.310 1014.180 ;
        RECT 1465.630 1013.980 1473.310 1014.120 ;
        RECT 1465.630 1013.920 1465.950 1013.980 ;
        RECT 1472.990 1013.920 1473.310 1013.980 ;
        RECT 1478.970 1014.120 1479.290 1014.180 ;
        RECT 1482.190 1014.120 1482.510 1014.180 ;
        RECT 1489.550 1014.120 1489.870 1014.180 ;
        RECT 1493.690 1014.120 1494.010 1014.180 ;
        RECT 1478.970 1013.980 1482.510 1014.120 ;
        RECT 1478.970 1013.920 1479.290 1013.980 ;
        RECT 1482.190 1013.920 1482.510 1013.980 ;
        RECT 1482.740 1013.980 1489.320 1014.120 ;
        RECT 1339.130 1013.780 1339.450 1013.840 ;
        RECT 1276.200 1013.640 1339.450 1013.780 ;
        RECT 1262.310 1013.580 1262.630 1013.640 ;
        RECT 1269.210 1013.580 1269.530 1013.640 ;
        RECT 1339.130 1013.580 1339.450 1013.640 ;
        RECT 1446.310 1013.780 1446.630 1013.840 ;
        RECT 1459.190 1013.780 1459.510 1013.840 ;
        RECT 1446.310 1013.640 1459.510 1013.780 ;
        RECT 1446.310 1013.580 1446.630 1013.640 ;
        RECT 1459.190 1013.580 1459.510 1013.640 ;
        RECT 999.190 1013.440 999.510 1013.500 ;
        RECT 1197.450 1013.440 1197.770 1013.500 ;
        RECT 999.190 1013.300 1197.770 1013.440 ;
        RECT 999.190 1013.240 999.510 1013.300 ;
        RECT 1197.450 1013.240 1197.770 1013.300 ;
        RECT 1197.910 1013.440 1198.230 1013.500 ;
        RECT 1225.970 1013.440 1226.290 1013.500 ;
        RECT 1197.910 1013.300 1226.290 1013.440 ;
        RECT 1197.910 1013.240 1198.230 1013.300 ;
        RECT 1225.970 1013.240 1226.290 1013.300 ;
        RECT 1244.830 1013.440 1245.150 1013.500 ;
        RECT 1292.670 1013.440 1292.990 1013.500 ;
        RECT 1333.150 1013.440 1333.470 1013.500 ;
        RECT 1244.830 1013.300 1292.440 1013.440 ;
        RECT 1244.830 1013.240 1245.150 1013.300 ;
        RECT 988.150 1013.100 988.470 1013.160 ;
        RECT 1223.670 1013.100 1223.990 1013.160 ;
        RECT 988.150 1012.960 1223.990 1013.100 ;
        RECT 988.150 1012.900 988.470 1012.960 ;
        RECT 1223.670 1012.900 1223.990 1012.960 ;
        RECT 1224.130 1013.100 1224.450 1013.160 ;
        RECT 1259.550 1013.100 1259.870 1013.160 ;
        RECT 1224.130 1012.960 1259.870 1013.100 ;
        RECT 1224.130 1012.900 1224.450 1012.960 ;
        RECT 1259.550 1012.900 1259.870 1012.960 ;
        RECT 1265.530 1013.100 1265.850 1013.160 ;
        RECT 1268.750 1013.100 1269.070 1013.160 ;
        RECT 1265.530 1012.960 1269.070 1013.100 ;
        RECT 1292.300 1013.100 1292.440 1013.300 ;
        RECT 1292.670 1013.300 1333.470 1013.440 ;
        RECT 1292.670 1013.240 1292.990 1013.300 ;
        RECT 1333.150 1013.240 1333.470 1013.300 ;
        RECT 1341.430 1013.100 1341.750 1013.160 ;
        RECT 1292.300 1012.960 1341.750 1013.100 ;
        RECT 1265.530 1012.900 1265.850 1012.960 ;
        RECT 1268.750 1012.900 1269.070 1012.960 ;
        RECT 1341.430 1012.900 1341.750 1012.960 ;
        RECT 1444.010 1013.100 1444.330 1013.160 ;
        RECT 1482.740 1013.100 1482.880 1013.980 ;
        RECT 1489.180 1013.780 1489.320 1013.980 ;
        RECT 1489.550 1013.980 1494.010 1014.120 ;
        RECT 1489.550 1013.920 1489.870 1013.980 ;
        RECT 1493.690 1013.920 1494.010 1013.980 ;
        RECT 1494.240 1013.780 1494.380 1014.320 ;
        RECT 1494.610 1014.120 1494.930 1014.180 ;
        RECT 1507.490 1014.120 1507.810 1014.180 ;
        RECT 1494.610 1013.980 1507.810 1014.120 ;
        RECT 1508.040 1014.120 1508.180 1014.320 ;
        RECT 1528.190 1014.120 1528.510 1014.180 ;
        RECT 1508.040 1013.980 1528.510 1014.120 ;
        RECT 1494.610 1013.920 1494.930 1013.980 ;
        RECT 1507.490 1013.920 1507.810 1013.980 ;
        RECT 1528.190 1013.920 1528.510 1013.980 ;
        RECT 1545.670 1014.120 1545.990 1014.180 ;
        RECT 1547.970 1014.120 1548.290 1014.180 ;
        RECT 1545.670 1013.980 1548.290 1014.120 ;
        RECT 1545.670 1013.920 1545.990 1013.980 ;
        RECT 1547.970 1013.920 1548.290 1013.980 ;
        RECT 1559.470 1014.120 1559.790 1014.180 ;
        RECT 1562.690 1014.120 1563.010 1014.180 ;
        RECT 1559.470 1013.980 1563.010 1014.120 ;
        RECT 1559.470 1013.920 1559.790 1013.980 ;
        RECT 1562.690 1013.920 1563.010 1013.980 ;
        RECT 1574.190 1014.120 1574.510 1014.180 ;
        RECT 1577.870 1014.120 1578.190 1014.180 ;
        RECT 1574.190 1013.980 1578.190 1014.120 ;
        RECT 1574.190 1013.920 1574.510 1013.980 ;
        RECT 1577.870 1013.920 1578.190 1013.980 ;
        RECT 1578.330 1014.120 1578.650 1014.180 ;
        RECT 1886.070 1014.120 1886.390 1014.180 ;
        RECT 1578.330 1013.980 1886.390 1014.120 ;
        RECT 1578.330 1013.920 1578.650 1013.980 ;
        RECT 1886.070 1013.920 1886.390 1013.980 ;
        RECT 2002.910 1014.120 2003.230 1014.180 ;
        RECT 2007.510 1014.120 2007.830 1014.180 ;
        RECT 2002.910 1013.980 2007.830 1014.120 ;
        RECT 2002.910 1013.920 2003.230 1013.980 ;
        RECT 2007.510 1013.920 2007.830 1013.980 ;
        RECT 1489.180 1013.640 1494.380 1013.780 ;
        RECT 1495.530 1013.780 1495.850 1013.840 ;
        RECT 1511.630 1013.780 1511.950 1013.840 ;
        RECT 1495.530 1013.640 1511.950 1013.780 ;
        RECT 1495.530 1013.580 1495.850 1013.640 ;
        RECT 1511.630 1013.580 1511.950 1013.640 ;
        RECT 1517.150 1013.780 1517.470 1013.840 ;
        RECT 1591.670 1013.780 1591.990 1013.840 ;
        RECT 1517.150 1013.640 1591.990 1013.780 ;
        RECT 1517.150 1013.580 1517.470 1013.640 ;
        RECT 1591.670 1013.580 1591.990 1013.640 ;
        RECT 1596.270 1013.780 1596.590 1013.840 ;
        RECT 1600.410 1013.780 1600.730 1013.840 ;
        RECT 1596.270 1013.640 1600.730 1013.780 ;
        RECT 1596.270 1013.580 1596.590 1013.640 ;
        RECT 1600.410 1013.580 1600.730 1013.640 ;
        RECT 1665.730 1013.780 1666.050 1013.840 ;
        RECT 1669.410 1013.780 1669.730 1013.840 ;
        RECT 1665.730 1013.640 1669.730 1013.780 ;
        RECT 1665.730 1013.580 1666.050 1013.640 ;
        RECT 1669.410 1013.580 1669.730 1013.640 ;
        RECT 1754.970 1013.780 1755.290 1013.840 ;
        RECT 1759.110 1013.780 1759.430 1013.840 ;
        RECT 1754.970 1013.640 1759.430 1013.780 ;
        RECT 1754.970 1013.580 1755.290 1013.640 ;
        RECT 1759.110 1013.580 1759.430 1013.640 ;
        RECT 1759.570 1013.780 1759.890 1013.840 ;
        RECT 2085.710 1013.780 2086.030 1013.840 ;
        RECT 1759.570 1013.640 2086.030 1013.780 ;
        RECT 1759.570 1013.580 1759.890 1013.640 ;
        RECT 2085.710 1013.580 2086.030 1013.640 ;
        RECT 1495.990 1013.440 1496.310 1013.500 ;
        RECT 1518.530 1013.440 1518.850 1013.500 ;
        RECT 1628.470 1013.440 1628.790 1013.500 ;
        RECT 1495.990 1013.300 1518.850 1013.440 ;
        RECT 1495.990 1013.240 1496.310 1013.300 ;
        RECT 1518.530 1013.240 1518.850 1013.300 ;
        RECT 1523.680 1013.300 1628.790 1013.440 ;
        RECT 1444.010 1012.960 1482.880 1013.100 ;
        RECT 1498.290 1013.100 1498.610 1013.160 ;
        RECT 1523.680 1013.100 1523.820 1013.300 ;
        RECT 1628.470 1013.240 1628.790 1013.300 ;
        RECT 1720.010 1013.440 1720.330 1013.500 ;
        RECT 2084.330 1013.440 2084.650 1013.500 ;
        RECT 1720.010 1013.300 2084.650 1013.440 ;
        RECT 1720.010 1013.240 1720.330 1013.300 ;
        RECT 2084.330 1013.240 2084.650 1013.300 ;
        RECT 1498.290 1012.960 1523.820 1013.100 ;
        RECT 1524.050 1013.100 1524.370 1013.160 ;
        RECT 1693.790 1013.100 1694.110 1013.160 ;
        RECT 1524.050 1012.960 1694.110 1013.100 ;
        RECT 1444.010 1012.900 1444.330 1012.960 ;
        RECT 1498.290 1012.900 1498.610 1012.960 ;
        RECT 1524.050 1012.900 1524.370 1012.960 ;
        RECT 1693.790 1012.900 1694.110 1012.960 ;
        RECT 1707.130 1013.100 1707.450 1013.160 ;
        RECT 1710.810 1013.100 1711.130 1013.160 ;
        RECT 1707.130 1012.960 1711.130 1013.100 ;
        RECT 1707.130 1012.900 1707.450 1012.960 ;
        RECT 1710.810 1012.900 1711.130 1012.960 ;
        RECT 1715.410 1013.100 1715.730 1013.160 ;
        RECT 1717.710 1013.100 1718.030 1013.160 ;
        RECT 1715.410 1012.960 1718.030 1013.100 ;
        RECT 1715.410 1012.900 1715.730 1012.960 ;
        RECT 1717.710 1012.900 1718.030 1012.960 ;
        RECT 1733.350 1013.100 1733.670 1013.160 ;
        RECT 1737.950 1013.100 1738.270 1013.160 ;
        RECT 1733.350 1012.960 1738.270 1013.100 ;
        RECT 1733.350 1012.900 1733.670 1012.960 ;
        RECT 1737.950 1012.900 1738.270 1012.960 ;
        RECT 1738.870 1013.100 1739.190 1013.160 ;
        RECT 2076.970 1013.100 2077.290 1013.160 ;
        RECT 1738.870 1012.960 2077.290 1013.100 ;
        RECT 1738.870 1012.900 1739.190 1012.960 ;
        RECT 2076.970 1012.900 2077.290 1012.960 ;
        RECT 796.790 1012.760 797.110 1012.820 ;
        RECT 884.650 1012.760 884.970 1012.820 ;
        RECT 796.790 1012.620 884.970 1012.760 ;
        RECT 796.790 1012.560 797.110 1012.620 ;
        RECT 884.650 1012.560 884.970 1012.620 ;
        RECT 987.690 1012.760 988.010 1012.820 ;
        RECT 1228.270 1012.760 1228.590 1012.820 ;
        RECT 987.690 1012.620 1228.590 1012.760 ;
        RECT 987.690 1012.560 988.010 1012.620 ;
        RECT 1228.270 1012.560 1228.590 1012.620 ;
        RECT 1237.470 1012.760 1237.790 1012.820 ;
        RECT 1338.670 1012.760 1338.990 1012.820 ;
        RECT 1237.470 1012.620 1338.990 1012.760 ;
        RECT 1237.470 1012.560 1237.790 1012.620 ;
        RECT 1338.670 1012.560 1338.990 1012.620 ;
        RECT 1357.070 1012.760 1357.390 1012.820 ;
        RECT 1362.590 1012.760 1362.910 1012.820 ;
        RECT 1357.070 1012.620 1362.910 1012.760 ;
        RECT 1357.070 1012.560 1357.390 1012.620 ;
        RECT 1362.590 1012.560 1362.910 1012.620 ;
        RECT 1496.910 1012.760 1497.230 1012.820 ;
        RECT 1517.150 1012.760 1517.470 1012.820 ;
        RECT 1866.290 1012.760 1866.610 1012.820 ;
        RECT 1887.450 1012.760 1887.770 1012.820 ;
        RECT 1496.910 1012.620 1517.470 1012.760 ;
        RECT 1496.910 1012.560 1497.230 1012.620 ;
        RECT 1517.150 1012.560 1517.470 1012.620 ;
        RECT 1518.160 1012.620 1866.610 1012.760 ;
        RECT 803.690 1012.420 804.010 1012.480 ;
        RECT 890.170 1012.420 890.490 1012.480 ;
        RECT 803.690 1012.280 890.490 1012.420 ;
        RECT 803.690 1012.220 804.010 1012.280 ;
        RECT 890.170 1012.220 890.490 1012.280 ;
        RECT 986.770 1012.420 987.090 1012.480 ;
        RECT 1224.130 1012.420 1224.450 1012.480 ;
        RECT 986.770 1012.280 1224.450 1012.420 ;
        RECT 986.770 1012.220 987.090 1012.280 ;
        RECT 1224.130 1012.220 1224.450 1012.280 ;
        RECT 1224.590 1012.420 1224.910 1012.480 ;
        RECT 1230.110 1012.420 1230.430 1012.480 ;
        RECT 1224.590 1012.280 1230.430 1012.420 ;
        RECT 1224.590 1012.220 1224.910 1012.280 ;
        RECT 1230.110 1012.220 1230.430 1012.280 ;
        RECT 1243.910 1012.420 1244.230 1012.480 ;
        RECT 1284.850 1012.420 1285.170 1012.480 ;
        RECT 1294.510 1012.420 1294.830 1012.480 ;
        RECT 1341.890 1012.420 1342.210 1012.480 ;
        RECT 1243.910 1012.280 1285.170 1012.420 ;
        RECT 1243.910 1012.220 1244.230 1012.280 ;
        RECT 1284.850 1012.220 1285.170 1012.280 ;
        RECT 1285.860 1012.280 1294.830 1012.420 ;
        RECT 789.890 1012.080 790.210 1012.140 ;
        RECT 910.870 1012.080 911.190 1012.140 ;
        RECT 789.890 1011.940 911.190 1012.080 ;
        RECT 789.890 1011.880 790.210 1011.940 ;
        RECT 910.870 1011.880 911.190 1011.940 ;
        RECT 995.970 1012.080 996.290 1012.140 ;
        RECT 1270.130 1012.080 1270.450 1012.140 ;
        RECT 995.970 1011.940 1270.450 1012.080 ;
        RECT 995.970 1011.880 996.290 1011.940 ;
        RECT 1270.130 1011.880 1270.450 1011.940 ;
        RECT 1276.110 1012.080 1276.430 1012.140 ;
        RECT 1285.860 1012.080 1286.000 1012.280 ;
        RECT 1294.510 1012.220 1294.830 1012.280 ;
        RECT 1295.520 1012.280 1342.210 1012.420 ;
        RECT 1276.110 1011.940 1286.000 1012.080 ;
        RECT 1276.110 1011.880 1276.430 1011.940 ;
        RECT 769.190 1011.740 769.510 1011.800 ;
        RECT 906.270 1011.740 906.590 1011.800 ;
        RECT 769.190 1011.600 906.590 1011.740 ;
        RECT 769.190 1011.540 769.510 1011.600 ;
        RECT 906.270 1011.540 906.590 1011.600 ;
        RECT 1000.110 1011.740 1000.430 1011.800 ;
        RECT 1075.550 1011.740 1075.870 1011.800 ;
        RECT 1000.110 1011.600 1075.870 1011.740 ;
        RECT 1000.110 1011.540 1000.430 1011.600 ;
        RECT 1075.550 1011.540 1075.870 1011.600 ;
        RECT 1079.690 1011.740 1080.010 1011.800 ;
        RECT 1081.070 1011.740 1081.390 1011.800 ;
        RECT 1079.690 1011.600 1081.390 1011.740 ;
        RECT 1079.690 1011.540 1080.010 1011.600 ;
        RECT 1081.070 1011.540 1081.390 1011.600 ;
        RECT 1104.070 1011.740 1104.390 1011.800 ;
        RECT 1106.370 1011.740 1106.690 1011.800 ;
        RECT 1104.070 1011.600 1106.690 1011.740 ;
        RECT 1104.070 1011.540 1104.390 1011.600 ;
        RECT 1106.370 1011.540 1106.690 1011.600 ;
        RECT 1106.830 1011.740 1107.150 1011.800 ;
        RECT 1145.470 1011.740 1145.790 1011.800 ;
        RECT 1106.830 1011.600 1145.790 1011.740 ;
        RECT 1106.830 1011.540 1107.150 1011.600 ;
        RECT 1145.470 1011.540 1145.790 1011.600 ;
        RECT 1169.390 1011.740 1169.710 1011.800 ;
        RECT 1262.310 1011.740 1262.630 1011.800 ;
        RECT 1295.520 1011.740 1295.660 1012.280 ;
        RECT 1341.890 1012.220 1342.210 1012.280 ;
        RECT 1369.950 1012.420 1370.270 1012.480 ;
        RECT 1372.710 1012.420 1373.030 1012.480 ;
        RECT 1369.950 1012.280 1373.030 1012.420 ;
        RECT 1369.950 1012.220 1370.270 1012.280 ;
        RECT 1372.710 1012.220 1373.030 1012.280 ;
        RECT 1384.670 1012.420 1384.990 1012.480 ;
        RECT 1386.510 1012.420 1386.830 1012.480 ;
        RECT 1384.670 1012.280 1386.830 1012.420 ;
        RECT 1384.670 1012.220 1384.990 1012.280 ;
        RECT 1386.510 1012.220 1386.830 1012.280 ;
        RECT 1393.410 1012.420 1393.730 1012.480 ;
        RECT 1397.090 1012.420 1397.410 1012.480 ;
        RECT 1393.410 1012.280 1397.410 1012.420 ;
        RECT 1393.410 1012.220 1393.730 1012.280 ;
        RECT 1397.090 1012.220 1397.410 1012.280 ;
        RECT 1404.910 1012.420 1405.230 1012.480 ;
        RECT 1406.750 1012.420 1407.070 1012.480 ;
        RECT 1404.910 1012.280 1407.070 1012.420 ;
        RECT 1404.910 1012.220 1405.230 1012.280 ;
        RECT 1406.750 1012.220 1407.070 1012.280 ;
        RECT 1488.630 1012.420 1488.950 1012.480 ;
        RECT 1516.690 1012.420 1517.010 1012.480 ;
        RECT 1488.630 1012.280 1517.010 1012.420 ;
        RECT 1488.630 1012.220 1488.950 1012.280 ;
        RECT 1516.690 1012.220 1517.010 1012.280 ;
        RECT 1295.890 1012.080 1296.210 1012.140 ;
        RECT 1342.350 1012.080 1342.670 1012.140 ;
        RECT 1295.890 1011.940 1342.670 1012.080 ;
        RECT 1295.890 1011.880 1296.210 1011.940 ;
        RECT 1342.350 1011.880 1342.670 1011.940 ;
        RECT 1376.390 1012.080 1376.710 1012.140 ;
        RECT 1432.050 1012.080 1432.370 1012.140 ;
        RECT 1376.390 1011.940 1432.370 1012.080 ;
        RECT 1376.390 1011.880 1376.710 1011.940 ;
        RECT 1432.050 1011.880 1432.370 1011.940 ;
        RECT 1509.330 1012.080 1509.650 1012.140 ;
        RECT 1518.160 1012.080 1518.300 1012.620 ;
        RECT 1866.290 1012.560 1866.610 1012.620 ;
        RECT 1868.220 1012.620 1887.770 1012.760 ;
        RECT 1524.510 1012.420 1524.830 1012.480 ;
        RECT 1545.670 1012.420 1545.990 1012.480 ;
        RECT 1524.510 1012.280 1545.990 1012.420 ;
        RECT 1524.510 1012.220 1524.830 1012.280 ;
        RECT 1545.670 1012.220 1545.990 1012.280 ;
        RECT 1553.030 1012.420 1553.350 1012.480 ;
        RECT 1556.250 1012.420 1556.570 1012.480 ;
        RECT 1553.030 1012.280 1556.570 1012.420 ;
        RECT 1553.030 1012.220 1553.350 1012.280 ;
        RECT 1556.250 1012.220 1556.570 1012.280 ;
        RECT 1556.710 1012.420 1557.030 1012.480 ;
        RECT 1868.220 1012.420 1868.360 1012.620 ;
        RECT 1887.450 1012.560 1887.770 1012.620 ;
        RECT 2004.750 1012.760 2005.070 1012.820 ;
        RECT 2073.290 1012.760 2073.610 1012.820 ;
        RECT 2004.750 1012.620 2073.610 1012.760 ;
        RECT 2004.750 1012.560 2005.070 1012.620 ;
        RECT 2073.290 1012.560 2073.610 1012.620 ;
        RECT 2073.840 1012.620 2080.880 1012.760 ;
        RECT 1556.710 1012.280 1868.360 1012.420 ;
        RECT 1872.270 1012.420 1872.590 1012.480 ;
        RECT 1876.410 1012.420 1876.730 1012.480 ;
        RECT 1872.270 1012.280 1876.730 1012.420 ;
        RECT 1556.710 1012.220 1557.030 1012.280 ;
        RECT 1872.270 1012.220 1872.590 1012.280 ;
        RECT 1876.410 1012.220 1876.730 1012.280 ;
        RECT 1509.330 1011.940 1518.300 1012.080 ;
        RECT 1518.530 1012.080 1518.850 1012.140 ;
        RECT 1525.430 1012.080 1525.750 1012.140 ;
        RECT 1518.530 1011.940 1525.750 1012.080 ;
        RECT 1509.330 1011.880 1509.650 1011.940 ;
        RECT 1518.530 1011.880 1518.850 1011.940 ;
        RECT 1525.430 1011.880 1525.750 1011.940 ;
        RECT 1535.090 1012.080 1535.410 1012.140 ;
        RECT 1541.990 1012.080 1542.310 1012.140 ;
        RECT 1535.090 1011.940 1542.310 1012.080 ;
        RECT 1535.090 1011.880 1535.410 1011.940 ;
        RECT 1541.990 1011.880 1542.310 1011.940 ;
        RECT 1542.450 1012.080 1542.770 1012.140 ;
        RECT 1614.670 1012.080 1614.990 1012.140 ;
        RECT 1542.450 1011.940 1614.990 1012.080 ;
        RECT 1542.450 1011.880 1542.770 1011.940 ;
        RECT 1614.670 1011.880 1614.990 1011.940 ;
        RECT 1662.510 1012.080 1662.830 1012.140 ;
        RECT 2061.330 1012.080 2061.650 1012.140 ;
        RECT 2073.840 1012.080 2073.980 1012.620 ;
        RECT 2080.740 1012.420 2080.880 1012.620 ;
        RECT 2287.190 1012.420 2287.510 1012.480 ;
        RECT 2080.740 1012.280 2287.510 1012.420 ;
        RECT 2287.190 1012.220 2287.510 1012.280 ;
        RECT 1662.510 1011.940 2053.740 1012.080 ;
        RECT 1662.510 1011.880 1662.830 1011.940 ;
        RECT 1334.070 1011.740 1334.390 1011.800 ;
        RECT 1169.390 1011.600 1244.600 1011.740 ;
        RECT 1169.390 1011.540 1169.710 1011.600 ;
        RECT 700.190 1011.400 700.510 1011.460 ;
        RECT 841.870 1011.400 842.190 1011.460 ;
        RECT 700.190 1011.260 842.190 1011.400 ;
        RECT 700.190 1011.200 700.510 1011.260 ;
        RECT 841.870 1011.200 842.190 1011.260 ;
        RECT 997.350 1011.400 997.670 1011.460 ;
        RECT 1076.010 1011.400 1076.330 1011.460 ;
        RECT 997.350 1011.260 1076.330 1011.400 ;
        RECT 997.350 1011.200 997.670 1011.260 ;
        RECT 1076.010 1011.200 1076.330 1011.260 ;
        RECT 1076.930 1011.400 1077.250 1011.460 ;
        RECT 1145.930 1011.400 1146.250 1011.460 ;
        RECT 1076.930 1011.260 1146.250 1011.400 ;
        RECT 1076.930 1011.200 1077.250 1011.260 ;
        RECT 1145.930 1011.200 1146.250 1011.260 ;
        RECT 1166.630 1011.400 1166.950 1011.460 ;
        RECT 1243.910 1011.400 1244.230 1011.460 ;
        RECT 1166.630 1011.260 1244.230 1011.400 ;
        RECT 1244.460 1011.400 1244.600 1011.600 ;
        RECT 1262.310 1011.600 1295.660 1011.740 ;
        RECT 1310.240 1011.600 1334.390 1011.740 ;
        RECT 1262.310 1011.540 1262.630 1011.600 ;
        RECT 1289.450 1011.400 1289.770 1011.460 ;
        RECT 1309.690 1011.400 1310.010 1011.460 ;
        RECT 1244.460 1011.260 1289.770 1011.400 ;
        RECT 1166.630 1011.200 1166.950 1011.260 ;
        RECT 1243.910 1011.200 1244.230 1011.260 ;
        RECT 1289.450 1011.200 1289.770 1011.260 ;
        RECT 1290.000 1011.260 1310.010 1011.400 ;
        RECT 517.110 1011.060 517.430 1011.120 ;
        RECT 712.610 1011.060 712.930 1011.120 ;
        RECT 517.110 1010.920 712.930 1011.060 ;
        RECT 517.110 1010.860 517.430 1010.920 ;
        RECT 712.610 1010.860 712.930 1010.920 ;
        RECT 755.390 1011.060 755.710 1011.120 ;
        RECT 901.670 1011.060 901.990 1011.120 ;
        RECT 755.390 1010.920 901.990 1011.060 ;
        RECT 755.390 1010.860 755.710 1010.920 ;
        RECT 901.670 1010.860 901.990 1010.920 ;
        RECT 994.130 1011.060 994.450 1011.120 ;
        RECT 1290.000 1011.060 1290.140 1011.260 ;
        RECT 1309.690 1011.200 1310.010 1011.260 ;
        RECT 994.130 1010.920 1290.140 1011.060 ;
        RECT 1290.370 1011.060 1290.690 1011.120 ;
        RECT 1310.240 1011.060 1310.380 1011.600 ;
        RECT 1334.070 1011.540 1334.390 1011.600 ;
        RECT 1378.690 1011.740 1379.010 1011.800 ;
        RECT 1431.590 1011.740 1431.910 1011.800 ;
        RECT 1378.690 1011.600 1431.910 1011.740 ;
        RECT 1378.690 1011.540 1379.010 1011.600 ;
        RECT 1431.590 1011.540 1431.910 1011.600 ;
        RECT 1500.590 1011.740 1500.910 1011.800 ;
        RECT 1865.830 1011.740 1866.150 1011.800 ;
        RECT 1500.590 1011.600 1866.150 1011.740 ;
        RECT 1500.590 1011.540 1500.910 1011.600 ;
        RECT 1865.830 1011.540 1866.150 1011.600 ;
        RECT 1866.290 1011.740 1866.610 1011.800 ;
        RECT 1894.810 1011.740 1895.130 1011.800 ;
        RECT 1866.290 1011.600 1895.130 1011.740 ;
        RECT 2053.600 1011.740 2053.740 1011.940 ;
        RECT 2061.330 1011.940 2073.980 1012.080 ;
        RECT 2078.810 1012.080 2079.130 1012.140 ;
        RECT 2082.950 1012.080 2083.270 1012.140 ;
        RECT 2078.810 1011.940 2083.270 1012.080 ;
        RECT 2061.330 1011.880 2061.650 1011.940 ;
        RECT 2078.810 1011.880 2079.130 1011.940 ;
        RECT 2082.950 1011.880 2083.270 1011.940 ;
        RECT 2087.550 1012.080 2087.870 1012.140 ;
        RECT 2090.310 1012.080 2090.630 1012.140 ;
        RECT 2087.550 1011.940 2090.630 1012.080 ;
        RECT 2087.550 1011.880 2087.870 1011.940 ;
        RECT 2090.310 1011.880 2090.630 1011.940 ;
        RECT 2083.870 1011.740 2084.190 1011.800 ;
        RECT 2519.490 1011.740 2519.810 1011.800 ;
        RECT 2053.600 1011.600 2084.190 1011.740 ;
        RECT 1866.290 1011.540 1866.610 1011.600 ;
        RECT 1894.810 1011.540 1895.130 1011.600 ;
        RECT 2083.870 1011.540 2084.190 1011.600 ;
        RECT 2084.420 1011.600 2519.810 1011.740 ;
        RECT 1386.510 1011.400 1386.830 1011.460 ;
        RECT 1890.670 1011.400 1890.990 1011.460 ;
        RECT 1386.510 1011.260 1890.990 1011.400 ;
        RECT 1386.510 1011.200 1386.830 1011.260 ;
        RECT 1890.670 1011.200 1890.990 1011.260 ;
        RECT 2074.670 1011.400 2074.990 1011.460 ;
        RECT 2084.420 1011.400 2084.560 1011.600 ;
        RECT 2519.490 1011.540 2519.810 1011.600 ;
        RECT 2519.030 1011.400 2519.350 1011.460 ;
        RECT 2074.670 1011.260 2084.560 1011.400 ;
        RECT 2084.880 1011.260 2519.350 1011.400 ;
        RECT 2074.670 1011.200 2074.990 1011.260 ;
        RECT 1290.370 1010.920 1310.380 1011.060 ;
        RECT 1320.270 1011.060 1320.590 1011.120 ;
        RECT 1342.810 1011.060 1343.130 1011.120 ;
        RECT 1320.270 1010.920 1343.130 1011.060 ;
        RECT 994.130 1010.860 994.450 1010.920 ;
        RECT 1290.370 1010.860 1290.690 1010.920 ;
        RECT 1320.270 1010.860 1320.590 1010.920 ;
        RECT 1342.810 1010.860 1343.130 1010.920 ;
        RECT 1354.770 1011.060 1355.090 1011.120 ;
        RECT 1873.190 1011.060 1873.510 1011.120 ;
        RECT 1891.590 1011.060 1891.910 1011.120 ;
        RECT 1354.770 1010.920 1873.510 1011.060 ;
        RECT 1354.770 1010.860 1355.090 1010.920 ;
        RECT 1873.190 1010.860 1873.510 1010.920 ;
        RECT 1873.740 1010.920 1891.910 1011.060 ;
        RECT 468.810 1010.720 469.130 1010.780 ;
        RECT 673.510 1010.720 673.830 1010.780 ;
        RECT 468.810 1010.580 673.830 1010.720 ;
        RECT 468.810 1010.520 469.130 1010.580 ;
        RECT 673.510 1010.520 673.830 1010.580 ;
        RECT 734.690 1010.720 735.010 1010.780 ;
        RECT 893.390 1010.720 893.710 1010.780 ;
        RECT 734.690 1010.580 893.710 1010.720 ;
        RECT 734.690 1010.520 735.010 1010.580 ;
        RECT 893.390 1010.520 893.710 1010.580 ;
        RECT 989.530 1010.720 989.850 1010.780 ;
        RECT 1347.410 1010.720 1347.730 1010.780 ;
        RECT 989.530 1010.580 1347.730 1010.720 ;
        RECT 989.530 1010.520 989.850 1010.580 ;
        RECT 1347.410 1010.520 1347.730 1010.580 ;
        RECT 1417.790 1010.720 1418.110 1010.780 ;
        RECT 1700.690 1010.720 1701.010 1010.780 ;
        RECT 1417.790 1010.580 1701.010 1010.720 ;
        RECT 1417.790 1010.520 1418.110 1010.580 ;
        RECT 1700.690 1010.520 1701.010 1010.580 ;
        RECT 1710.810 1010.720 1711.130 1010.780 ;
        RECT 1738.870 1010.720 1739.190 1010.780 ;
        RECT 1710.810 1010.580 1739.190 1010.720 ;
        RECT 1710.810 1010.520 1711.130 1010.580 ;
        RECT 1738.870 1010.520 1739.190 1010.580 ;
        RECT 1741.630 1010.720 1741.950 1010.780 ;
        RECT 1759.570 1010.720 1759.890 1010.780 ;
        RECT 1741.630 1010.580 1759.890 1010.720 ;
        RECT 1741.630 1010.520 1741.950 1010.580 ;
        RECT 1759.570 1010.520 1759.890 1010.580 ;
        RECT 1767.850 1010.720 1768.170 1010.780 ;
        RECT 1772.910 1010.720 1773.230 1010.780 ;
        RECT 1767.850 1010.580 1773.230 1010.720 ;
        RECT 1767.850 1010.520 1768.170 1010.580 ;
        RECT 1772.910 1010.520 1773.230 1010.580 ;
        RECT 1830.870 1010.720 1831.190 1010.780 ;
        RECT 1835.010 1010.720 1835.330 1010.780 ;
        RECT 1830.870 1010.580 1835.330 1010.720 ;
        RECT 1830.870 1010.520 1831.190 1010.580 ;
        RECT 1835.010 1010.520 1835.330 1010.580 ;
        RECT 1865.830 1010.720 1866.150 1010.780 ;
        RECT 1873.740 1010.720 1873.880 1010.920 ;
        RECT 1891.590 1010.860 1891.910 1010.920 ;
        RECT 2055.350 1011.060 2055.670 1011.120 ;
        RECT 2084.880 1011.060 2085.020 1011.260 ;
        RECT 2519.030 1011.200 2519.350 1011.260 ;
        RECT 2055.350 1010.920 2085.020 1011.060 ;
        RECT 2085.250 1011.060 2085.570 1011.120 ;
        RECT 2518.570 1011.060 2518.890 1011.120 ;
        RECT 2085.250 1010.920 2518.890 1011.060 ;
        RECT 2055.350 1010.860 2055.670 1010.920 ;
        RECT 2085.250 1010.860 2085.570 1010.920 ;
        RECT 2518.570 1010.860 2518.890 1010.920 ;
        RECT 1865.830 1010.580 1873.880 1010.720 ;
        RECT 1883.310 1010.720 1883.630 1010.780 ;
        RECT 2532.370 1010.720 2532.690 1010.780 ;
        RECT 1883.310 1010.580 2532.690 1010.720 ;
        RECT 1865.830 1010.520 1866.150 1010.580 ;
        RECT 1883.310 1010.520 1883.630 1010.580 ;
        RECT 2532.370 1010.520 2532.690 1010.580 ;
        RECT 995.510 1010.380 995.830 1010.440 ;
        RECT 999.190 1010.380 999.510 1010.440 ;
        RECT 995.510 1010.240 999.510 1010.380 ;
        RECT 995.510 1010.180 995.830 1010.240 ;
        RECT 999.190 1010.180 999.510 1010.240 ;
        RECT 999.650 1010.380 999.970 1010.440 ;
        RECT 1146.390 1010.380 1146.710 1010.440 ;
        RECT 999.650 1010.240 1146.710 1010.380 ;
        RECT 999.650 1010.180 999.970 1010.240 ;
        RECT 1146.390 1010.180 1146.710 1010.240 ;
        RECT 1204.810 1010.380 1205.130 1010.440 ;
        RECT 1336.830 1010.380 1337.150 1010.440 ;
        RECT 1204.810 1010.240 1337.150 1010.380 ;
        RECT 1204.810 1010.180 1205.130 1010.240 ;
        RECT 1336.830 1010.180 1337.150 1010.240 ;
        RECT 1447.690 1010.380 1448.010 1010.440 ;
        RECT 1520.830 1010.380 1521.150 1010.440 ;
        RECT 1556.710 1010.380 1557.030 1010.440 ;
        RECT 1447.690 1010.240 1521.150 1010.380 ;
        RECT 1447.690 1010.180 1448.010 1010.240 ;
        RECT 1520.830 1010.180 1521.150 1010.240 ;
        RECT 1525.060 1010.240 1557.030 1010.380 ;
        RECT 998.730 1010.040 999.050 1010.100 ;
        RECT 1150.990 1010.040 1151.310 1010.100 ;
        RECT 1160.190 1010.040 1160.510 1010.100 ;
        RECT 998.730 1009.900 1151.310 1010.040 ;
        RECT 998.730 1009.840 999.050 1009.900 ;
        RECT 1150.990 1009.840 1151.310 1009.900 ;
        RECT 1159.820 1009.900 1160.510 1010.040 ;
        RECT 993.210 1009.700 993.530 1009.760 ;
        RECT 1080.150 1009.700 1080.470 1009.760 ;
        RECT 993.210 1009.560 1080.470 1009.700 ;
        RECT 993.210 1009.500 993.530 1009.560 ;
        RECT 1080.150 1009.500 1080.470 1009.560 ;
        RECT 1081.070 1009.700 1081.390 1009.760 ;
        RECT 1159.820 1009.700 1159.960 1009.900 ;
        RECT 1160.190 1009.840 1160.510 1009.900 ;
        RECT 1183.190 1010.040 1183.510 1010.100 ;
        RECT 1186.410 1010.040 1186.730 1010.100 ;
        RECT 1183.190 1009.900 1186.730 1010.040 ;
        RECT 1183.190 1009.840 1183.510 1009.900 ;
        RECT 1186.410 1009.840 1186.730 1009.900 ;
        RECT 1223.210 1010.040 1223.530 1010.100 ;
        RECT 1340.050 1010.040 1340.370 1010.100 ;
        RECT 1223.210 1009.900 1340.370 1010.040 ;
        RECT 1223.210 1009.840 1223.530 1009.900 ;
        RECT 1340.050 1009.840 1340.370 1009.900 ;
        RECT 1503.810 1010.040 1504.130 1010.100 ;
        RECT 1525.060 1010.040 1525.200 1010.240 ;
        RECT 1556.710 1010.180 1557.030 1010.240 ;
        RECT 1576.490 1010.380 1576.810 1010.440 ;
        RECT 1579.710 1010.380 1580.030 1010.440 ;
        RECT 1576.490 1010.240 1580.030 1010.380 ;
        RECT 1576.490 1010.180 1576.810 1010.240 ;
        RECT 1579.710 1010.180 1580.030 1010.240 ;
        RECT 1580.170 1010.380 1580.490 1010.440 ;
        RECT 1585.690 1010.380 1586.010 1010.440 ;
        RECT 1580.170 1010.240 1586.010 1010.380 ;
        RECT 1580.170 1010.180 1580.490 1010.240 ;
        RECT 1585.690 1010.180 1586.010 1010.240 ;
        RECT 1593.050 1010.380 1593.370 1010.440 ;
        RECT 1686.890 1010.380 1687.210 1010.440 ;
        RECT 1593.050 1010.240 1687.210 1010.380 ;
        RECT 1593.050 1010.180 1593.370 1010.240 ;
        RECT 1686.890 1010.180 1687.210 1010.240 ;
        RECT 1749.910 1010.380 1750.230 1010.440 ;
        RECT 1752.210 1010.380 1752.530 1010.440 ;
        RECT 1749.910 1010.240 1752.530 1010.380 ;
        RECT 1749.910 1010.180 1750.230 1010.240 ;
        RECT 1752.210 1010.180 1752.530 1010.240 ;
        RECT 1763.710 1010.380 1764.030 1010.440 ;
        RECT 1766.010 1010.380 1766.330 1010.440 ;
        RECT 2086.170 1010.380 2086.490 1010.440 ;
        RECT 1763.710 1010.240 1766.330 1010.380 ;
        RECT 1763.710 1010.180 1764.030 1010.240 ;
        RECT 1766.010 1010.180 1766.330 1010.240 ;
        RECT 1766.560 1010.240 2086.490 1010.380 ;
        RECT 1576.950 1010.040 1577.270 1010.100 ;
        RECT 1503.810 1009.900 1525.200 1010.040 ;
        RECT 1531.500 1009.900 1577.270 1010.040 ;
        RECT 1503.810 1009.840 1504.130 1009.900 ;
        RECT 1081.070 1009.560 1159.960 1009.700 ;
        RECT 1176.290 1009.700 1176.610 1009.760 ;
        RECT 1205.270 1009.700 1205.590 1009.760 ;
        RECT 1210.330 1009.700 1210.650 1009.760 ;
        RECT 1238.390 1009.700 1238.710 1009.760 ;
        RECT 1176.290 1009.560 1205.590 1009.700 ;
        RECT 1081.070 1009.500 1081.390 1009.560 ;
        RECT 1176.290 1009.500 1176.610 1009.560 ;
        RECT 1205.270 1009.500 1205.590 1009.560 ;
        RECT 1207.890 1009.560 1208.720 1009.700 ;
        RECT 993.670 1009.360 993.990 1009.420 ;
        RECT 1058.530 1009.360 1058.850 1009.420 ;
        RECT 993.670 1009.220 1058.850 1009.360 ;
        RECT 993.670 1009.160 993.990 1009.220 ;
        RECT 1058.530 1009.160 1058.850 1009.220 ;
        RECT 1069.570 1009.360 1069.890 1009.420 ;
        RECT 1071.870 1009.360 1072.190 1009.420 ;
        RECT 1069.570 1009.220 1072.190 1009.360 ;
        RECT 1069.570 1009.160 1069.890 1009.220 ;
        RECT 1071.870 1009.160 1072.190 1009.220 ;
        RECT 1077.390 1009.360 1077.710 1009.420 ;
        RECT 1106.830 1009.360 1107.150 1009.420 ;
        RECT 1077.390 1009.220 1107.150 1009.360 ;
        RECT 1077.390 1009.160 1077.710 1009.220 ;
        RECT 1106.830 1009.160 1107.150 1009.220 ;
        RECT 1200.210 1009.360 1200.530 1009.420 ;
        RECT 1207.890 1009.360 1208.030 1009.560 ;
        RECT 1200.210 1009.220 1208.030 1009.360 ;
        RECT 1208.580 1009.360 1208.720 1009.560 ;
        RECT 1210.330 1009.560 1238.710 1009.700 ;
        RECT 1210.330 1009.500 1210.650 1009.560 ;
        RECT 1238.390 1009.500 1238.710 1009.560 ;
        RECT 1274.270 1009.700 1274.590 1009.760 ;
        RECT 1334.530 1009.700 1334.850 1009.760 ;
        RECT 1274.270 1009.560 1334.850 1009.700 ;
        RECT 1274.270 1009.500 1274.590 1009.560 ;
        RECT 1334.530 1009.500 1334.850 1009.560 ;
        RECT 1489.090 1009.700 1489.410 1009.760 ;
        RECT 1524.510 1009.700 1524.830 1009.760 ;
        RECT 1489.090 1009.560 1524.830 1009.700 ;
        RECT 1489.090 1009.500 1489.410 1009.560 ;
        RECT 1524.510 1009.500 1524.830 1009.560 ;
        RECT 1210.790 1009.360 1211.110 1009.420 ;
        RECT 1208.580 1009.220 1211.110 1009.360 ;
        RECT 1200.210 1009.160 1200.530 1009.220 ;
        RECT 1210.790 1009.160 1211.110 1009.220 ;
        RECT 1279.790 1009.360 1280.110 1009.420 ;
        RECT 1320.270 1009.360 1320.590 1009.420 ;
        RECT 1337.290 1009.360 1337.610 1009.420 ;
        RECT 1279.790 1009.220 1320.590 1009.360 ;
        RECT 1279.790 1009.160 1280.110 1009.220 ;
        RECT 1320.270 1009.160 1320.590 1009.220 ;
        RECT 1320.820 1009.220 1337.610 1009.360 ;
        RECT 984.010 1009.020 984.330 1009.080 ;
        RECT 1079.690 1009.020 1080.010 1009.080 ;
        RECT 984.010 1008.880 1080.010 1009.020 ;
        RECT 984.010 1008.820 984.330 1008.880 ;
        RECT 1079.690 1008.820 1080.010 1008.880 ;
        RECT 1098.550 1009.020 1098.870 1009.080 ;
        RECT 1111.430 1009.020 1111.750 1009.080 ;
        RECT 1098.550 1008.880 1111.750 1009.020 ;
        RECT 1098.550 1008.820 1098.870 1008.880 ;
        RECT 1111.430 1008.820 1111.750 1008.880 ;
        RECT 1145.930 1009.020 1146.250 1009.080 ;
        RECT 1159.730 1009.020 1160.050 1009.080 ;
        RECT 1145.930 1008.880 1160.050 1009.020 ;
        RECT 1145.930 1008.820 1146.250 1008.880 ;
        RECT 1159.730 1008.820 1160.050 1008.880 ;
        RECT 1162.490 1009.020 1162.810 1009.080 ;
        RECT 1183.650 1009.020 1183.970 1009.080 ;
        RECT 1162.490 1008.880 1183.970 1009.020 ;
        RECT 1162.490 1008.820 1162.810 1008.880 ;
        RECT 1183.650 1008.820 1183.970 1008.880 ;
        RECT 1190.550 1009.020 1190.870 1009.080 ;
        RECT 1207.570 1009.020 1207.890 1009.080 ;
        RECT 1190.550 1008.880 1207.890 1009.020 ;
        RECT 1190.550 1008.820 1190.870 1008.880 ;
        RECT 1207.570 1008.820 1207.890 1008.880 ;
        RECT 1209.410 1009.020 1209.730 1009.080 ;
        RECT 1304.170 1009.020 1304.490 1009.080 ;
        RECT 1209.410 1008.880 1304.490 1009.020 ;
        RECT 1209.410 1008.820 1209.730 1008.880 ;
        RECT 1304.170 1008.820 1304.490 1008.880 ;
        RECT 996.430 1008.680 996.750 1008.740 ;
        RECT 1097.630 1008.680 1097.950 1008.740 ;
        RECT 996.430 1008.540 1097.950 1008.680 ;
        RECT 996.430 1008.480 996.750 1008.540 ;
        RECT 1097.630 1008.480 1097.950 1008.540 ;
        RECT 1100.850 1008.680 1101.170 1008.740 ;
        RECT 1159.270 1008.680 1159.590 1008.740 ;
        RECT 1100.850 1008.540 1159.590 1008.680 ;
        RECT 1100.850 1008.480 1101.170 1008.540 ;
        RECT 1159.270 1008.480 1159.590 1008.540 ;
        RECT 1161.110 1008.680 1161.430 1008.740 ;
        RECT 1269.210 1008.680 1269.530 1008.740 ;
        RECT 1317.970 1008.680 1318.290 1008.740 ;
        RECT 1161.110 1008.540 1208.260 1008.680 ;
        RECT 1161.110 1008.480 1161.430 1008.540 ;
        RECT 1208.120 1008.400 1208.260 1008.540 ;
        RECT 1269.210 1008.540 1318.290 1008.680 ;
        RECT 1269.210 1008.480 1269.530 1008.540 ;
        RECT 1317.970 1008.480 1318.290 1008.540 ;
        RECT 997.810 1008.340 998.130 1008.400 ;
        RECT 1093.030 1008.340 1093.350 1008.400 ;
        RECT 997.810 1008.200 1093.350 1008.340 ;
        RECT 997.810 1008.140 998.130 1008.200 ;
        RECT 1093.030 1008.140 1093.350 1008.200 ;
        RECT 1148.690 1008.340 1149.010 1008.400 ;
        RECT 1186.870 1008.340 1187.190 1008.400 ;
        RECT 1148.690 1008.200 1187.190 1008.340 ;
        RECT 1148.690 1008.140 1149.010 1008.200 ;
        RECT 1186.870 1008.140 1187.190 1008.200 ;
        RECT 1190.090 1008.340 1190.410 1008.400 ;
        RECT 1207.570 1008.340 1207.890 1008.400 ;
        RECT 1190.090 1008.200 1207.890 1008.340 ;
        RECT 1190.090 1008.140 1190.410 1008.200 ;
        RECT 1207.570 1008.140 1207.890 1008.200 ;
        RECT 1208.030 1008.140 1208.350 1008.400 ;
        RECT 1209.410 1008.340 1209.730 1008.400 ;
        RECT 1297.270 1008.340 1297.590 1008.400 ;
        RECT 1209.410 1008.200 1297.590 1008.340 ;
        RECT 1209.410 1008.140 1209.730 1008.200 ;
        RECT 1297.270 1008.140 1297.590 1008.200 ;
        RECT 1300.490 1008.340 1300.810 1008.400 ;
        RECT 1320.820 1008.340 1320.960 1009.220 ;
        RECT 1337.290 1009.160 1337.610 1009.220 ;
        RECT 1487.710 1009.360 1488.030 1009.420 ;
        RECT 1530.950 1009.360 1531.270 1009.420 ;
        RECT 1487.710 1009.220 1531.270 1009.360 ;
        RECT 1487.710 1009.160 1488.030 1009.220 ;
        RECT 1530.950 1009.160 1531.270 1009.220 ;
        RECT 1331.310 1009.020 1331.630 1009.080 ;
        RECT 1345.570 1009.020 1345.890 1009.080 ;
        RECT 1331.310 1008.880 1345.890 1009.020 ;
        RECT 1331.310 1008.820 1331.630 1008.880 ;
        RECT 1345.570 1008.820 1345.890 1008.880 ;
        RECT 1497.830 1009.020 1498.150 1009.080 ;
        RECT 1531.500 1009.020 1531.640 1009.900 ;
        RECT 1576.950 1009.840 1577.270 1009.900 ;
        RECT 1591.670 1010.040 1591.990 1010.100 ;
        RECT 1603.170 1010.040 1603.490 1010.100 ;
        RECT 1591.670 1009.900 1603.490 1010.040 ;
        RECT 1591.670 1009.840 1591.990 1009.900 ;
        RECT 1603.170 1009.840 1603.490 1009.900 ;
        RECT 1758.650 1010.040 1758.970 1010.100 ;
        RECT 1766.560 1010.040 1766.700 1010.240 ;
        RECT 2086.170 1010.180 2086.490 1010.240 ;
        RECT 1758.650 1009.900 1766.700 1010.040 ;
        RECT 1826.730 1010.040 1827.050 1010.100 ;
        RECT 1845.590 1010.040 1845.910 1010.100 ;
        RECT 1826.730 1009.900 1845.910 1010.040 ;
        RECT 1758.650 1009.840 1758.970 1009.900 ;
        RECT 1826.730 1009.840 1827.050 1009.900 ;
        RECT 1845.590 1009.840 1845.910 1009.900 ;
        RECT 1878.710 1010.040 1879.030 1010.100 ;
        RECT 1893.890 1010.040 1894.210 1010.100 ;
        RECT 1878.710 1009.900 1894.210 1010.040 ;
        RECT 1878.710 1009.840 1879.030 1009.900 ;
        RECT 1893.890 1009.840 1894.210 1009.900 ;
        RECT 1531.870 1009.700 1532.190 1009.760 ;
        RECT 1542.450 1009.700 1542.770 1009.760 ;
        RECT 1531.870 1009.560 1542.770 1009.700 ;
        RECT 1531.870 1009.500 1532.190 1009.560 ;
        RECT 1542.450 1009.500 1542.770 1009.560 ;
        RECT 1555.790 1009.700 1556.110 1009.760 ;
        RECT 1652.390 1009.700 1652.710 1009.760 ;
        RECT 1555.790 1009.560 1652.710 1009.700 ;
        RECT 1555.790 1009.500 1556.110 1009.560 ;
        RECT 1652.390 1009.500 1652.710 1009.560 ;
        RECT 1789.470 1009.700 1789.790 1009.760 ;
        RECT 2084.790 1009.700 2085.110 1009.760 ;
        RECT 1789.470 1009.560 2085.110 1009.700 ;
        RECT 1789.470 1009.500 1789.790 1009.560 ;
        RECT 2084.790 1009.500 2085.110 1009.560 ;
        RECT 1568.210 1009.360 1568.530 1009.420 ;
        RECT 1497.830 1008.880 1531.640 1009.020 ;
        RECT 1531.960 1009.220 1568.530 1009.360 ;
        RECT 1497.830 1008.820 1498.150 1008.880 ;
        RECT 1325.790 1008.680 1326.110 1008.740 ;
        RECT 1335.910 1008.680 1336.230 1008.740 ;
        RECT 1325.790 1008.540 1336.230 1008.680 ;
        RECT 1325.790 1008.480 1326.110 1008.540 ;
        RECT 1335.910 1008.480 1336.230 1008.540 ;
        RECT 1491.850 1008.680 1492.170 1008.740 ;
        RECT 1524.050 1008.680 1524.370 1008.740 ;
        RECT 1491.850 1008.540 1524.370 1008.680 ;
        RECT 1491.850 1008.480 1492.170 1008.540 ;
        RECT 1524.050 1008.480 1524.370 1008.540 ;
        RECT 1524.970 1008.680 1525.290 1008.740 ;
        RECT 1528.190 1008.680 1528.510 1008.740 ;
        RECT 1524.970 1008.540 1528.510 1008.680 ;
        RECT 1524.970 1008.480 1525.290 1008.540 ;
        RECT 1528.190 1008.480 1528.510 1008.540 ;
        RECT 1300.490 1008.200 1320.960 1008.340 ;
        RECT 1335.450 1008.340 1335.770 1008.400 ;
        RECT 1340.970 1008.340 1341.290 1008.400 ;
        RECT 1335.450 1008.200 1341.290 1008.340 ;
        RECT 1300.490 1008.140 1300.810 1008.200 ;
        RECT 1335.450 1008.140 1335.770 1008.200 ;
        RECT 1340.970 1008.140 1341.290 1008.200 ;
        RECT 1368.110 1008.340 1368.430 1008.400 ;
        RECT 1383.290 1008.340 1383.610 1008.400 ;
        RECT 1368.110 1008.200 1383.610 1008.340 ;
        RECT 1368.110 1008.140 1368.430 1008.200 ;
        RECT 1383.290 1008.140 1383.610 1008.200 ;
        RECT 1497.370 1008.340 1497.690 1008.400 ;
        RECT 1531.960 1008.340 1532.100 1009.220 ;
        RECT 1568.210 1009.160 1568.530 1009.220 ;
        RECT 1602.710 1009.360 1603.030 1009.420 ;
        RECT 1607.310 1009.360 1607.630 1009.420 ;
        RECT 1602.710 1009.220 1607.630 1009.360 ;
        RECT 1602.710 1009.160 1603.030 1009.220 ;
        RECT 1607.310 1009.160 1607.630 1009.220 ;
        RECT 1613.750 1009.360 1614.070 1009.420 ;
        RECT 1891.130 1009.360 1891.450 1009.420 ;
        RECT 1613.750 1009.220 1891.450 1009.360 ;
        RECT 1613.750 1009.160 1614.070 1009.220 ;
        RECT 1891.130 1009.160 1891.450 1009.220 ;
        RECT 2046.150 1009.360 2046.470 1009.420 ;
        RECT 2085.250 1009.360 2085.570 1009.420 ;
        RECT 2046.150 1009.220 2085.570 1009.360 ;
        RECT 2046.150 1009.160 2046.470 1009.220 ;
        RECT 2085.250 1009.160 2085.570 1009.220 ;
        RECT 1559.930 1009.020 1560.250 1009.080 ;
        RECT 1537.020 1008.880 1560.250 1009.020 ;
        RECT 1532.330 1008.680 1532.650 1008.740 ;
        RECT 1536.470 1008.680 1536.790 1008.740 ;
        RECT 1532.330 1008.540 1536.790 1008.680 ;
        RECT 1532.330 1008.480 1532.650 1008.540 ;
        RECT 1536.470 1008.480 1536.790 1008.540 ;
        RECT 1497.370 1008.200 1532.100 1008.340 ;
        RECT 1497.370 1008.140 1497.690 1008.200 ;
        RECT 632.110 1008.000 632.430 1008.060 ;
        RECT 670.750 1008.000 671.070 1008.060 ;
        RECT 632.110 1007.860 671.070 1008.000 ;
        RECT 632.110 1007.800 632.430 1007.860 ;
        RECT 670.750 1007.800 671.070 1007.860 ;
        RECT 998.270 1008.000 998.590 1008.060 ;
        RECT 1084.290 1008.000 1084.610 1008.060 ;
        RECT 998.270 1007.860 1084.610 1008.000 ;
        RECT 998.270 1007.800 998.590 1007.860 ;
        RECT 1084.290 1007.800 1084.610 1007.860 ;
        RECT 1150.990 1008.000 1151.310 1008.060 ;
        RECT 1191.010 1008.000 1191.330 1008.060 ;
        RECT 1150.990 1007.860 1191.330 1008.000 ;
        RECT 1150.990 1007.800 1151.310 1007.860 ;
        RECT 1191.010 1007.800 1191.330 1007.860 ;
        RECT 1191.470 1008.000 1191.790 1008.060 ;
        RECT 1238.850 1008.000 1239.170 1008.060 ;
        RECT 1191.470 1007.860 1239.170 1008.000 ;
        RECT 1191.470 1007.800 1191.790 1007.860 ;
        RECT 1238.850 1007.800 1239.170 1007.860 ;
        RECT 1250.350 1008.000 1250.670 1008.060 ;
        RECT 1254.950 1008.000 1255.270 1008.060 ;
        RECT 1292.670 1008.000 1292.990 1008.060 ;
        RECT 1250.350 1007.860 1255.270 1008.000 ;
        RECT 1250.350 1007.800 1250.670 1007.860 ;
        RECT 1254.950 1007.800 1255.270 1007.860 ;
        RECT 1255.500 1007.860 1292.990 1008.000 ;
        RECT 638.090 1007.660 638.410 1007.720 ;
        RECT 671.670 1007.660 671.990 1007.720 ;
        RECT 638.090 1007.520 671.990 1007.660 ;
        RECT 638.090 1007.460 638.410 1007.520 ;
        RECT 671.670 1007.460 671.990 1007.520 ;
        RECT 992.750 1007.660 993.070 1007.720 ;
        RECT 1014.370 1007.660 1014.690 1007.720 ;
        RECT 992.750 1007.520 1014.690 1007.660 ;
        RECT 992.750 1007.460 993.070 1007.520 ;
        RECT 1014.370 1007.460 1014.690 1007.520 ;
        RECT 1079.690 1007.660 1080.010 1007.720 ;
        RECT 1115.110 1007.660 1115.430 1007.720 ;
        RECT 1079.690 1007.520 1115.430 1007.660 ;
        RECT 1079.690 1007.460 1080.010 1007.520 ;
        RECT 1115.110 1007.460 1115.430 1007.520 ;
        RECT 1145.470 1007.660 1145.790 1007.720 ;
        RECT 1169.390 1007.660 1169.710 1007.720 ;
        RECT 1145.470 1007.520 1169.710 1007.660 ;
        RECT 1145.470 1007.460 1145.790 1007.520 ;
        RECT 1169.390 1007.460 1169.710 1007.520 ;
        RECT 1197.450 1007.660 1197.770 1007.720 ;
        RECT 1232.410 1007.660 1232.730 1007.720 ;
        RECT 1197.450 1007.520 1232.730 1007.660 ;
        RECT 1197.450 1007.460 1197.770 1007.520 ;
        RECT 1232.410 1007.460 1232.730 1007.520 ;
        RECT 1254.490 1007.660 1254.810 1007.720 ;
        RECT 1255.500 1007.660 1255.640 1007.860 ;
        RECT 1292.670 1007.800 1292.990 1007.860 ;
        RECT 1293.590 1008.000 1293.910 1008.060 ;
        RECT 1319.350 1008.000 1319.670 1008.060 ;
        RECT 1293.590 1007.860 1319.670 1008.000 ;
        RECT 1293.590 1007.800 1293.910 1007.860 ;
        RECT 1319.350 1007.800 1319.670 1007.860 ;
        RECT 1334.990 1008.000 1335.310 1008.060 ;
        RECT 1338.670 1008.000 1338.990 1008.060 ;
        RECT 1334.990 1007.860 1338.990 1008.000 ;
        RECT 1334.990 1007.800 1335.310 1007.860 ;
        RECT 1338.670 1007.800 1338.990 1007.860 ;
        RECT 1396.170 1008.000 1396.490 1008.060 ;
        RECT 1400.310 1008.000 1400.630 1008.060 ;
        RECT 1396.170 1007.860 1400.630 1008.000 ;
        RECT 1396.170 1007.800 1396.490 1007.860 ;
        RECT 1400.310 1007.800 1400.630 1007.860 ;
        RECT 1413.190 1008.000 1413.510 1008.060 ;
        RECT 1438.490 1008.000 1438.810 1008.060 ;
        RECT 1413.190 1007.860 1438.810 1008.000 ;
        RECT 1413.190 1007.800 1413.510 1007.860 ;
        RECT 1438.490 1007.800 1438.810 1007.860 ;
        RECT 1496.450 1008.000 1496.770 1008.060 ;
        RECT 1537.020 1008.000 1537.160 1008.880 ;
        RECT 1559.930 1008.820 1560.250 1008.880 ;
        RECT 1834.550 1009.020 1834.870 1009.080 ;
        RECT 2100.890 1009.020 2101.210 1009.080 ;
        RECT 1834.550 1008.880 2101.210 1009.020 ;
        RECT 1834.550 1008.820 1834.870 1008.880 ;
        RECT 2100.890 1008.820 2101.210 1008.880 ;
        RECT 1541.990 1008.680 1542.310 1008.740 ;
        RECT 1578.330 1008.680 1578.650 1008.740 ;
        RECT 1541.990 1008.540 1578.650 1008.680 ;
        RECT 1541.990 1008.480 1542.310 1008.540 ;
        RECT 1578.330 1008.480 1578.650 1008.540 ;
        RECT 1824.430 1008.680 1824.750 1008.740 ;
        RECT 1907.690 1008.680 1908.010 1008.740 ;
        RECT 1824.430 1008.540 1908.010 1008.680 ;
        RECT 1824.430 1008.480 1824.750 1008.540 ;
        RECT 1907.690 1008.480 1908.010 1008.540 ;
        RECT 2050.750 1008.680 2051.070 1008.740 ;
        RECT 2055.810 1008.680 2056.130 1008.740 ;
        RECT 2050.750 1008.540 2056.130 1008.680 ;
        RECT 2050.750 1008.480 2051.070 1008.540 ;
        RECT 2055.810 1008.480 2056.130 1008.540 ;
        RECT 2065.930 1008.680 2066.250 1008.740 ;
        RECT 2080.190 1008.680 2080.510 1008.740 ;
        RECT 2065.930 1008.540 2080.510 1008.680 ;
        RECT 2065.930 1008.480 2066.250 1008.540 ;
        RECT 2080.190 1008.480 2080.510 1008.540 ;
        RECT 1873.190 1008.340 1873.510 1008.400 ;
        RECT 1900.330 1008.340 1900.650 1008.400 ;
        RECT 1873.190 1008.200 1900.650 1008.340 ;
        RECT 1873.190 1008.140 1873.510 1008.200 ;
        RECT 1900.330 1008.140 1900.650 1008.200 ;
        RECT 1496.450 1007.860 1537.160 1008.000 ;
        RECT 1574.650 1008.000 1574.970 1008.060 ;
        RECT 1901.250 1008.000 1901.570 1008.060 ;
        RECT 1574.650 1007.860 1901.570 1008.000 ;
        RECT 1496.450 1007.800 1496.770 1007.860 ;
        RECT 1574.650 1007.800 1574.970 1007.860 ;
        RECT 1901.250 1007.800 1901.570 1007.860 ;
        RECT 1254.490 1007.520 1255.640 1007.660 ;
        RECT 1257.250 1007.660 1257.570 1007.720 ;
        RECT 1294.050 1007.660 1294.370 1007.720 ;
        RECT 1257.250 1007.520 1294.370 1007.660 ;
        RECT 1254.490 1007.460 1254.810 1007.520 ;
        RECT 1257.250 1007.460 1257.570 1007.520 ;
        RECT 1294.050 1007.460 1294.370 1007.520 ;
        RECT 1324.410 1007.660 1324.730 1007.720 ;
        RECT 1332.690 1007.660 1333.010 1007.720 ;
        RECT 1324.410 1007.520 1333.010 1007.660 ;
        RECT 1324.410 1007.460 1324.730 1007.520 ;
        RECT 1332.690 1007.460 1333.010 1007.520 ;
        RECT 1333.150 1007.660 1333.470 1007.720 ;
        RECT 1336.370 1007.660 1336.690 1007.720 ;
        RECT 1333.150 1007.520 1336.690 1007.660 ;
        RECT 1333.150 1007.460 1333.470 1007.520 ;
        RECT 1336.370 1007.460 1336.690 1007.520 ;
        RECT 1411.350 1007.660 1411.670 1007.720 ;
        RECT 1424.690 1007.660 1425.010 1007.720 ;
        RECT 1411.350 1007.520 1425.010 1007.660 ;
        RECT 1411.350 1007.460 1411.670 1007.520 ;
        RECT 1424.690 1007.460 1425.010 1007.520 ;
        RECT 1431.130 1007.660 1431.450 1007.720 ;
        RECT 1434.810 1007.660 1435.130 1007.720 ;
        RECT 1431.130 1007.520 1435.130 1007.660 ;
        RECT 1431.130 1007.460 1431.450 1007.520 ;
        RECT 1434.810 1007.460 1435.130 1007.520 ;
        RECT 1511.630 1007.660 1511.950 1007.720 ;
        RECT 1514.850 1007.660 1515.170 1007.720 ;
        RECT 1511.630 1007.520 1515.170 1007.660 ;
        RECT 1511.630 1007.460 1511.950 1007.520 ;
        RECT 1514.850 1007.460 1515.170 1007.520 ;
        RECT 1620.190 1007.660 1620.510 1007.720 ;
        RECT 1635.370 1007.660 1635.690 1007.720 ;
        RECT 1620.190 1007.520 1635.690 1007.660 ;
        RECT 1620.190 1007.460 1620.510 1007.520 ;
        RECT 1635.370 1007.460 1635.690 1007.520 ;
        RECT 1776.590 1007.660 1776.910 1007.720 ;
        RECT 1779.810 1007.660 1780.130 1007.720 ;
        RECT 1776.590 1007.520 1780.130 1007.660 ;
        RECT 1776.590 1007.460 1776.910 1007.520 ;
        RECT 1779.810 1007.460 1780.130 1007.520 ;
        RECT 1798.210 1007.660 1798.530 1007.720 ;
        RECT 1800.510 1007.660 1800.830 1007.720 ;
        RECT 1798.210 1007.520 1800.830 1007.660 ;
        RECT 1798.210 1007.460 1798.530 1007.520 ;
        RECT 1800.510 1007.460 1800.830 1007.520 ;
        RECT 1802.810 1007.660 1803.130 1007.720 ;
        RECT 1806.950 1007.660 1807.270 1007.720 ;
        RECT 1802.810 1007.520 1807.270 1007.660 ;
        RECT 1802.810 1007.460 1803.130 1007.520 ;
        RECT 1806.950 1007.460 1807.270 1007.520 ;
        RECT 1811.550 1007.660 1811.870 1007.720 ;
        RECT 1813.850 1007.660 1814.170 1007.720 ;
        RECT 1811.550 1007.520 1814.170 1007.660 ;
        RECT 1811.550 1007.460 1811.870 1007.520 ;
        RECT 1813.850 1007.460 1814.170 1007.520 ;
        RECT 1075.550 1007.320 1075.870 1007.380 ;
        RECT 1077.390 1007.320 1077.710 1007.380 ;
        RECT 1075.550 1007.180 1077.710 1007.320 ;
        RECT 1075.550 1007.120 1075.870 1007.180 ;
        RECT 1077.390 1007.120 1077.710 1007.180 ;
        RECT 1076.010 1006.980 1076.330 1007.040 ;
        RECT 1076.930 1006.980 1077.250 1007.040 ;
        RECT 1076.010 1006.840 1077.250 1006.980 ;
        RECT 1076.010 1006.780 1076.330 1006.840 ;
        RECT 1076.930 1006.780 1077.250 1006.840 ;
        RECT 1332.230 1005.960 1332.550 1006.020 ;
        RECT 1338.210 1005.960 1338.530 1006.020 ;
        RECT 1332.230 1005.820 1338.530 1005.960 ;
        RECT 1332.230 1005.760 1332.550 1005.820 ;
        RECT 1338.210 1005.760 1338.530 1005.820 ;
        RECT 1208.030 1001.200 1208.350 1001.260 ;
        RECT 1216.540 1001.200 1216.860 1001.260 ;
        RECT 1208.030 1001.060 1216.860 1001.200 ;
        RECT 1208.030 1001.000 1208.350 1001.060 ;
        RECT 1216.540 1001.000 1216.860 1001.060 ;
        RECT 1332.230 1000.520 1332.550 1000.580 ;
        RECT 1333.610 1000.520 1333.930 1000.580 ;
        RECT 1332.230 1000.380 1333.930 1000.520 ;
        RECT 1332.230 1000.320 1332.550 1000.380 ;
        RECT 1333.610 1000.320 1333.930 1000.380 ;
        RECT 1193.770 999.500 1194.090 999.560 ;
        RECT 1197.450 999.500 1197.770 999.560 ;
        RECT 1193.770 999.360 1197.770 999.500 ;
        RECT 1193.770 999.300 1194.090 999.360 ;
        RECT 1197.450 999.300 1197.770 999.360 ;
        RECT 1215.390 999.500 1215.710 999.560 ;
        RECT 1219.070 999.500 1219.390 999.560 ;
        RECT 1215.390 999.360 1219.390 999.500 ;
        RECT 1215.390 999.300 1215.710 999.360 ;
        RECT 1219.070 999.300 1219.390 999.360 ;
      LAYER met1 ;
        RECT 670.990 604.460 2169.070 998.780 ;
      LAYER via ;
        RECT 1352.040 2917.920 1352.300 2918.180 ;
        RECT 1535.120 2917.920 1535.380 2918.180 ;
        RECT 1431.620 2917.580 1431.880 2917.840 ;
        RECT 1598.600 2917.580 1598.860 2917.840 ;
        RECT 1459.220 2915.880 1459.480 2916.140 ;
        RECT 1641.840 2915.880 1642.100 2916.140 ;
        RECT 1494.640 2915.540 1494.900 2915.800 ;
        RECT 1705.320 2915.540 1705.580 2915.800 ;
        RECT 1473.020 2915.200 1473.280 2915.460 ;
        RECT 1694.280 2915.200 1694.540 2915.460 ;
        RECT 1406.780 2914.860 1407.040 2915.120 ;
        RECT 1630.800 2914.860 1631.060 2915.120 ;
        RECT 1495.100 2914.520 1495.360 2914.780 ;
        RECT 1768.800 2914.520 1769.060 2914.780 ;
        RECT 1493.260 2914.180 1493.520 2914.440 ;
        RECT 1779.840 2914.180 1780.100 2914.440 ;
        RECT 1455.540 2913.840 1455.800 2914.100 ;
        RECT 1758.680 2913.840 1758.940 2914.100 ;
        RECT 1493.720 2913.500 1493.980 2913.760 ;
        RECT 1801.000 2913.500 1801.260 2913.760 ;
        RECT 1500.620 2913.160 1500.880 2913.420 ;
        RECT 1812.040 2913.160 1812.300 2913.420 ;
        RECT 1833.200 2913.160 1833.460 2913.420 ;
        RECT 1894.380 2913.160 1894.640 2913.420 ;
        RECT 1494.180 2912.820 1494.440 2913.080 ;
        RECT 1663.000 2912.820 1663.260 2913.080 ;
        RECT 1789.960 2912.820 1790.220 2913.080 ;
        RECT 1892.080 2912.820 1892.340 2913.080 ;
        RECT 1492.340 2912.480 1492.600 2912.740 ;
        RECT 1609.640 2912.480 1609.900 2912.740 ;
        RECT 1854.360 2912.480 1854.620 2912.740 ;
        RECT 1893.460 2912.480 1893.720 2912.740 ;
        RECT 1438.520 2912.140 1438.780 2912.400 ;
        RECT 1567.320 2912.140 1567.580 2912.400 ;
        RECT 1492.800 2911.800 1493.060 2912.060 ;
        RECT 1546.160 2911.800 1546.420 2912.060 ;
        RECT 1864.480 2911.800 1864.740 2912.060 ;
        RECT 1893.000 2911.800 1893.260 2912.060 ;
        RECT 1496.940 2898.200 1497.200 2898.460 ;
        RECT 1524.080 2898.200 1524.340 2898.460 ;
        RECT 1497.400 2896.500 1497.660 2896.760 ;
        RECT 1503.380 2896.500 1503.640 2896.760 ;
        RECT 1876.900 2896.500 1877.160 2896.760 ;
        RECT 1892.540 2896.500 1892.800 2896.760 ;
        RECT 1362.620 2849.580 1362.880 2849.840 ;
        RECT 1483.600 2849.580 1483.860 2849.840 ;
        RECT 1501.540 2842.780 1501.800 2843.040 ;
        RECT 1502.000 2842.780 1502.260 2843.040 ;
        RECT 1501.540 2815.920 1501.800 2816.180 ;
        RECT 1501.540 2815.240 1501.800 2815.500 ;
        RECT 979.440 2810.140 979.700 2810.400 ;
        RECT 985.420 2809.460 985.680 2809.720 ;
        RECT 1043.380 2809.460 1043.640 2809.720 ;
        RECT 1089.380 2809.460 1089.640 2809.720 ;
        RECT 984.960 2809.120 985.220 2809.380 ;
        RECT 1027.740 2809.120 1028.000 2809.380 ;
        RECT 986.340 2808.780 986.600 2809.040 ;
        RECT 1073.740 2808.780 1074.000 2809.040 ;
        RECT 985.880 2808.440 986.140 2808.700 ;
        RECT 1012.100 2808.440 1012.360 2808.700 ;
        RECT 1501.540 2794.500 1501.800 2794.760 ;
        RECT 1502.000 2794.500 1502.260 2794.760 ;
        RECT 445.840 2769.340 446.100 2769.600 ;
        RECT 810.620 2769.340 810.880 2769.600 ;
        RECT 532.320 2767.980 532.580 2768.240 ;
        RECT 700.220 2767.980 700.480 2768.240 ;
        RECT 518.520 2767.640 518.780 2767.900 ;
        RECT 755.420 2767.640 755.680 2767.900 ;
        RECT 489.080 2767.300 489.340 2767.560 ;
        RECT 789.920 2767.300 790.180 2767.560 ;
        RECT 586.600 2684.000 586.860 2684.260 ;
        RECT 734.720 2684.000 734.980 2684.260 ;
        RECT 586.600 2663.600 586.860 2663.860 ;
        RECT 803.720 2663.600 803.980 2663.860 ;
        RECT 1365.840 2780.900 1366.100 2781.160 ;
        RECT 1485.440 2780.900 1485.700 2781.160 ;
        RECT 1502.000 2766.960 1502.260 2767.220 ;
        RECT 1502.000 2766.280 1502.260 2766.540 ;
        RECT 1501.540 2753.020 1501.800 2753.280 ;
        RECT 1502.000 2753.020 1502.260 2753.280 ;
        RECT 1501.540 2719.020 1501.800 2719.280 ;
        RECT 1501.540 2718.340 1501.800 2718.600 ;
        RECT 1434.380 2691.140 1434.640 2691.400 ;
        RECT 1488.660 2691.140 1488.920 2691.400 ;
        RECT 1501.540 2670.400 1501.800 2670.660 ;
        RECT 1502.000 2670.060 1502.260 2670.320 ;
        RECT 1501.540 2656.460 1501.800 2656.720 ;
        RECT 1502.000 2656.460 1502.260 2656.720 ;
        RECT 1501.540 2622.460 1501.800 2622.720 ;
        RECT 1501.540 2621.780 1501.800 2622.040 ;
        RECT 1400.340 2608.180 1400.600 2608.440 ;
        RECT 1485.440 2608.180 1485.700 2608.440 ;
        RECT 996.920 2605.460 997.180 2605.720 ;
        RECT 1111.920 2605.460 1112.180 2605.720 ;
        RECT 997.380 2605.120 997.640 2605.380 ;
        RECT 1112.840 2605.120 1113.100 2605.380 ;
        RECT 991.400 2604.780 991.660 2605.040 ;
        RECT 1113.300 2604.780 1113.560 2605.040 ;
        RECT 990.940 2604.440 991.200 2604.700 ;
        RECT 1112.380 2604.440 1112.640 2604.700 ;
        RECT 1397.120 2594.580 1397.380 2594.840 ;
        RECT 1488.660 2594.580 1488.920 2594.840 ;
        RECT 533.240 2591.520 533.500 2591.780 ;
        RECT 769.220 2591.520 769.480 2591.780 ;
        RECT 504.720 2591.180 504.980 2591.440 ;
        RECT 796.820 2591.180 797.080 2591.440 ;
        RECT 990.480 2591.180 990.740 2591.440 ;
        RECT 1094.900 2591.180 1095.160 2591.440 ;
        RECT 1028.200 2587.440 1028.460 2587.700 ;
        RECT 1033.260 2587.440 1033.520 2587.700 ;
        RECT 1424.720 2580.640 1424.980 2580.900 ;
        RECT 1488.660 2580.640 1488.920 2580.900 ;
        RECT 1469.340 2546.300 1469.600 2546.560 ;
        RECT 1483.600 2546.300 1483.860 2546.560 ;
        RECT 1500.160 2511.960 1500.420 2512.220 ;
        RECT 1502.000 2511.960 1502.260 2512.220 ;
        RECT 2100.920 2781.240 2101.180 2781.500 ;
        RECT 2556.320 2781.240 2556.580 2781.500 ;
        RECT 1893.920 2780.900 1894.180 2781.160 ;
        RECT 2422.000 2780.900 2422.260 2781.160 ;
        RECT 1902.200 2503.800 1902.460 2504.060 ;
        RECT 1903.580 2503.800 1903.840 2504.060 ;
        RECT 1502.000 2495.640 1502.260 2495.900 ;
        RECT 1559.500 2495.640 1559.760 2495.900 ;
        RECT 1494.640 2495.300 1494.900 2495.560 ;
        RECT 1553.060 2495.300 1553.320 2495.560 ;
        RECT 1621.140 2495.300 1621.400 2495.560 ;
        RECT 1892.080 2495.300 1892.340 2495.560 ;
        RECT 1495.100 2494.960 1495.360 2495.220 ;
        RECT 1574.220 2494.960 1574.480 2495.220 ;
        RECT 1607.340 2494.960 1607.600 2495.220 ;
        RECT 1892.540 2494.960 1892.800 2495.220 ;
        RECT 1493.260 2494.620 1493.520 2494.880 ;
        RECT 1580.200 2494.620 1580.460 2494.880 ;
        RECT 1586.640 2494.620 1586.900 2494.880 ;
        RECT 1894.380 2494.620 1894.640 2494.880 ;
        RECT 1494.180 2494.280 1494.440 2494.540 ;
        RECT 1545.700 2494.280 1545.960 2494.540 ;
        RECT 1552.140 2494.280 1552.400 2494.540 ;
        RECT 1893.460 2494.280 1893.720 2494.540 ;
        RECT 1492.340 2493.940 1492.600 2494.200 ;
        RECT 1532.360 2493.940 1532.620 2494.200 ;
        RECT 1545.240 2493.940 1545.500 2494.200 ;
        RECT 1893.000 2493.940 1893.260 2494.200 ;
        RECT 1492.800 2491.220 1493.060 2491.480 ;
        RECT 1512.120 2491.220 1512.380 2491.480 ;
        RECT 1600.440 2489.520 1600.700 2489.780 ;
        RECT 1789.960 2489.520 1790.220 2489.780 ;
        RECT 1693.820 2489.180 1694.080 2489.440 ;
        RECT 1811.120 2489.180 1811.380 2489.440 ;
        RECT 1420.580 2488.840 1420.840 2489.100 ;
        RECT 1842.400 2488.840 1842.660 2489.100 ;
        RECT 1455.080 2488.500 1455.340 2488.760 ;
        RECT 1885.640 2488.500 1885.900 2488.760 ;
        RECT 1421.040 2488.160 1421.300 2488.420 ;
        RECT 1874.600 2488.160 1874.860 2488.420 ;
        RECT 1530.060 2487.820 1530.320 2488.080 ;
        RECT 1832.280 2487.820 1832.540 2488.080 ;
        RECT 1427.940 2486.800 1428.200 2487.060 ;
        RECT 1725.560 2486.800 1725.820 2487.060 ;
        RECT 1461.520 2486.460 1461.780 2486.720 ;
        RECT 1757.760 2486.460 1758.020 2486.720 ;
        RECT 1386.540 2486.120 1386.800 2486.380 ;
        RECT 1587.560 2486.120 1587.820 2486.380 ;
        RECT 1686.920 2486.120 1687.180 2486.380 ;
        RECT 1778.920 2486.120 1779.180 2486.380 ;
        RECT 1383.320 2485.780 1383.580 2486.040 ;
        RECT 1555.360 2485.780 1555.620 2486.040 ;
        RECT 1579.740 2485.780 1580.000 2486.040 ;
        RECT 1746.720 2485.780 1746.980 2486.040 ;
        RECT 1442.660 2485.440 1442.920 2485.700 ;
        RECT 1608.720 2485.440 1608.980 2485.700 ;
        RECT 1507.520 2485.100 1507.780 2485.360 ;
        RECT 1629.880 2485.100 1630.140 2485.360 ;
        RECT 1432.080 2484.760 1432.340 2485.020 ;
        RECT 1534.200 2484.760 1534.460 2485.020 ;
        RECT 1544.780 2484.760 1545.040 2485.020 ;
        RECT 1608.720 2484.760 1608.980 2485.020 ;
        RECT 1528.220 2484.420 1528.480 2484.680 ;
        RECT 1619.760 2484.420 1620.020 2484.680 ;
        RECT 1542.020 2484.080 1542.280 2484.340 ;
        RECT 1576.520 2484.080 1576.780 2484.340 ;
        RECT 1652.420 2484.080 1652.680 2484.340 ;
        RECT 1683.240 2484.080 1683.500 2484.340 ;
        RECT 1700.720 2484.080 1700.980 2484.340 ;
        RECT 1715.440 2484.080 1715.700 2484.340 ;
        RECT 1441.740 2429.340 1442.000 2429.600 ;
        RECT 1441.280 2428.320 1441.540 2428.580 ;
        RECT 1520.860 2429.000 1521.120 2429.260 ;
        RECT 1521.320 2428.320 1521.580 2428.580 ;
        RECT 1441.280 2414.720 1441.540 2414.980 ;
        RECT 1441.740 2414.720 1442.000 2414.980 ;
        RECT 1519.940 2414.720 1520.200 2414.980 ;
        RECT 1521.320 2414.720 1521.580 2414.980 ;
        RECT 1441.740 2380.380 1442.000 2380.640 ;
        RECT 1441.280 2380.040 1441.540 2380.300 ;
        RECT 1440.360 2342.300 1440.620 2342.560 ;
        RECT 1441.740 2342.300 1442.000 2342.560 ;
        RECT 1520.860 2332.100 1521.120 2332.360 ;
        RECT 1521.320 2331.760 1521.580 2332.020 ;
        RECT 1440.360 2318.840 1440.620 2319.100 ;
        RECT 1441.280 2318.840 1441.540 2319.100 ;
        RECT 1441.280 2318.160 1441.540 2318.420 ;
        RECT 1441.740 2318.160 1442.000 2318.420 ;
        RECT 1521.320 2284.160 1521.580 2284.420 ;
        RECT 1441.740 2283.820 1442.000 2284.080 ;
        RECT 1441.280 2283.480 1441.540 2283.740 ;
        RECT 1521.320 2283.480 1521.580 2283.740 ;
        RECT 1521.320 2269.880 1521.580 2270.140 ;
        RECT 1521.780 2269.880 1522.040 2270.140 ;
        RECT 1520.860 2262.740 1521.120 2263.000 ;
        RECT 1521.780 2262.740 1522.040 2263.000 ;
        RECT 1440.360 2245.740 1440.620 2246.000 ;
        RECT 1441.740 2245.740 1442.000 2246.000 ;
        RECT 1440.360 2222.280 1440.620 2222.540 ;
        RECT 1441.280 2222.280 1441.540 2222.540 ;
        RECT 1441.280 2221.600 1441.540 2221.860 ;
        RECT 1441.740 2221.600 1442.000 2221.860 ;
        RECT 1520.400 2214.800 1520.660 2215.060 ;
        RECT 1520.860 2214.800 1521.120 2215.060 ;
        RECT 1441.740 2187.260 1442.000 2187.520 ;
        RECT 1441.280 2186.920 1441.540 2187.180 ;
        RECT 1520.400 2173.660 1520.660 2173.920 ;
        RECT 1520.860 2173.660 1521.120 2173.920 ;
        RECT 1520.860 2162.780 1521.120 2163.040 ;
        RECT 1521.780 2162.780 1522.040 2163.040 ;
        RECT 1440.360 2149.180 1440.620 2149.440 ;
        RECT 1441.740 2149.180 1442.000 2149.440 ;
        RECT 1440.360 2125.720 1440.620 2125.980 ;
        RECT 1441.280 2125.720 1441.540 2125.980 ;
        RECT 1440.360 2125.040 1440.620 2125.300 ;
        RECT 1441.280 2125.040 1441.540 2125.300 ;
        RECT 1519.940 2076.760 1520.200 2077.020 ;
        RECT 1520.400 2076.760 1520.660 2077.020 ;
        RECT 1519.020 2069.620 1519.280 2069.880 ;
        RECT 1519.940 2069.620 1520.200 2069.880 ;
        RECT 1244.860 2053.980 1245.120 2054.240 ;
        RECT 1332.720 2053.980 1332.980 2054.240 ;
        RECT 1230.140 2053.640 1230.400 2053.900 ;
        RECT 1338.700 2053.640 1338.960 2053.900 ;
        RECT 1173.100 2053.300 1173.360 2053.560 ;
        RECT 1333.180 2053.300 1333.440 2053.560 ;
        RECT 1144.580 2052.960 1144.840 2053.220 ;
        RECT 1335.020 2052.960 1335.280 2053.220 ;
        RECT 1116.980 2052.620 1117.240 2052.880 ;
        RECT 1334.560 2052.620 1334.820 2052.880 ;
        RECT 1059.940 2052.280 1060.200 2052.540 ;
        RECT 1335.480 2052.280 1335.740 2052.540 ;
        RECT 1031.420 2051.940 1031.680 2052.200 ;
        RECT 1331.800 2051.940 1332.060 2052.200 ;
        RECT 1216.340 2051.600 1216.600 2051.860 ;
        RECT 1334.100 2051.600 1334.360 2051.860 ;
        RECT 1201.620 2051.260 1201.880 2051.520 ;
        RECT 1333.640 2051.260 1333.900 2051.520 ;
        RECT 1187.820 2050.920 1188.080 2051.180 ;
        RECT 1338.240 2050.920 1338.500 2051.180 ;
        RECT 984.500 2050.580 984.760 2050.840 ;
        RECT 1002.900 2050.580 1003.160 2050.840 ;
        RECT 1287.180 2050.580 1287.440 2050.840 ;
        RECT 1343.760 2050.580 1344.020 2050.840 ;
        RECT 998.760 2050.240 999.020 2050.500 ;
        RECT 1088.460 2050.240 1088.720 2050.500 ;
        RECT 1273.380 2050.240 1273.640 2050.500 ;
        RECT 1344.220 2050.240 1344.480 2050.500 ;
        RECT 999.680 2049.900 999.940 2050.160 ;
        RECT 1102.260 2049.900 1102.520 2050.160 ;
        RECT 1258.660 2049.900 1258.920 2050.160 ;
        RECT 1332.260 2049.900 1332.520 2050.160 ;
        RECT 1000.140 2049.560 1000.400 2049.820 ;
        RECT 1073.740 2049.560 1074.000 2049.820 ;
        RECT 1301.900 2049.560 1302.160 2049.820 ;
        RECT 1337.780 2049.560 1338.040 2049.820 ;
        RECT 999.220 2049.220 999.480 2049.480 ;
        RECT 1045.220 2049.220 1045.480 2049.480 ;
        RECT 1329.500 2049.220 1329.760 2049.480 ;
        RECT 1344.680 2049.220 1344.940 2049.480 ;
        RECT 997.840 2048.200 998.100 2048.460 ;
        RECT 1014.400 2048.200 1014.660 2048.460 ;
        RECT 998.300 2047.860 998.560 2048.120 ;
        RECT 1028.200 2047.860 1028.460 2048.120 ;
        RECT 984.040 2047.520 984.300 2047.780 ;
        RECT 1048.900 2047.520 1049.160 2047.780 ;
        RECT 978.520 2047.180 978.780 2047.440 ;
        RECT 1062.700 2047.180 1062.960 2047.440 ;
        RECT 978.980 2046.840 979.240 2047.100 ;
        RECT 1076.500 2046.840 1076.760 2047.100 ;
        RECT 983.580 2046.500 983.840 2046.760 ;
        RECT 1113.760 2046.500 1114.020 2046.760 ;
        RECT 983.120 2046.160 983.380 2046.420 ;
        RECT 1114.220 2046.160 1114.480 2046.420 ;
        RECT 978.060 2045.820 978.320 2046.080 ;
        RECT 1111.000 2045.820 1111.260 2046.080 ;
        RECT 977.600 2045.480 977.860 2045.740 ;
        RECT 1111.460 2045.480 1111.720 2045.740 ;
        RECT 1439.440 2042.420 1439.700 2042.680 ;
        RECT 1439.900 2042.420 1440.160 2042.680 ;
        RECT 579.240 1988.700 579.500 1988.960 ;
        RECT 632.140 1988.700 632.400 1988.960 ;
        RECT 530.020 1988.020 530.280 1988.280 ;
        RECT 638.120 1988.020 638.380 1988.280 ;
        RECT 419.620 1979.860 419.880 1980.120 ;
        RECT 420.540 1979.860 420.800 1980.120 ;
        RECT 420.080 1978.500 420.340 1978.760 ;
        RECT 419.620 1978.160 419.880 1978.420 ;
        RECT 843.280 1977.820 843.540 1978.080 ;
        RECT 897.560 1977.480 897.820 1977.740 ;
        RECT 996.460 1714.320 996.720 1714.580 ;
        RECT 1001.060 1714.320 1001.320 1714.580 ;
        RECT 1441.740 1993.800 1442.000 1994.060 ;
        RECT 1442.660 1993.800 1442.920 1994.060 ;
        RECT 1519.940 1993.800 1520.200 1994.060 ;
        RECT 1521.320 1993.800 1521.580 1994.060 ;
        RECT 2082.980 1946.880 2083.240 1947.140 ;
        RECT 2321.260 1946.880 2321.520 1947.140 ;
        RECT 2073.320 1946.540 2073.580 1946.800 ;
        RECT 2379.220 1946.540 2379.480 1946.800 ;
        RECT 2090.340 1946.200 2090.600 1946.460 ;
        RECT 2437.180 1946.200 2437.440 1946.460 ;
        RECT 1521.320 1945.860 1521.580 1946.120 ;
        RECT 2083.440 1945.860 2083.700 1946.120 ;
        RECT 2495.140 1945.860 2495.400 1946.120 ;
        RECT 1520.860 1945.520 1521.120 1945.780 ;
        RECT 1876.440 1935.320 1876.700 1935.580 ;
        RECT 2394.400 1935.320 2394.660 1935.580 ;
        RECT 1521.320 1931.580 1521.580 1931.840 ;
        RECT 1522.240 1931.580 1522.500 1931.840 ;
        RECT 1724.640 1928.860 1724.900 1929.120 ;
        RECT 2044.340 1928.860 2044.600 1929.120 ;
        RECT 1845.620 1927.840 1845.880 1928.100 ;
        RECT 1964.300 1927.840 1964.560 1928.100 ;
        RECT 1745.340 1927.500 1745.600 1927.760 ;
        RECT 1929.340 1927.500 1929.600 1927.760 ;
        RECT 1779.380 1927.160 1779.640 1927.420 ;
        RECT 1998.340 1927.160 1998.600 1927.420 ;
        RECT 1786.740 1926.820 1787.000 1927.080 ;
        RECT 2033.300 1926.820 2033.560 1927.080 ;
        RECT 1766.040 1926.480 1766.300 1926.740 ;
        RECT 2010.300 1926.480 2010.560 1926.740 ;
        RECT 1738.440 1926.140 1738.700 1926.400 ;
        RECT 1987.300 1926.140 1987.560 1926.400 ;
        RECT 1717.740 1925.800 1718.000 1926.060 ;
        RECT 1975.340 1925.800 1975.600 1926.060 ;
        RECT 1779.840 1925.460 1780.100 1925.720 ;
        RECT 2067.340 1925.460 2067.600 1925.720 ;
        RECT 1835.040 1925.120 1835.300 1925.380 ;
        RECT 1952.340 1925.120 1952.600 1925.380 ;
        RECT 1441.740 1897.240 1442.000 1897.500 ;
        RECT 1442.660 1897.240 1442.920 1897.500 ;
        RECT 1759.140 1883.640 1759.400 1883.900 ;
        RECT 1904.500 1883.640 1904.760 1883.900 ;
        RECT 1821.240 1870.040 1821.500 1870.300 ;
        RECT 1904.500 1870.040 1904.760 1870.300 ;
        RECT 1521.320 1859.500 1521.580 1859.760 ;
        RECT 1522.240 1859.500 1522.500 1859.760 ;
        RECT 1737.980 1849.300 1738.240 1849.560 ;
        RECT 1904.500 1849.300 1904.760 1849.560 ;
        RECT 1669.440 1814.620 1669.700 1814.880 ;
        RECT 1904.500 1814.620 1904.760 1814.880 ;
        RECT 1772.940 1766.340 1773.200 1766.600 ;
        RECT 1904.500 1766.340 1904.760 1766.600 ;
        RECT 1521.320 1762.940 1521.580 1763.200 ;
        RECT 1522.240 1762.940 1522.500 1763.200 ;
        RECT 2080.220 1870.040 2080.480 1870.300 ;
        RECT 2284.000 1870.040 2284.260 1870.300 ;
        RECT 1907.720 1738.460 1907.980 1738.720 ;
        RECT 1933.940 1738.460 1934.200 1738.720 ;
        RECT 1800.540 1738.120 1800.800 1738.380 ;
        RECT 1956.940 1738.120 1957.200 1738.380 ;
        RECT 1814.340 1737.780 1814.600 1738.040 ;
        RECT 1990.980 1737.780 1991.240 1738.040 ;
        RECT 1793.640 1737.440 1793.900 1737.700 ;
        RECT 1967.980 1737.440 1968.240 1737.700 ;
        RECT 1813.880 1737.100 1814.140 1737.360 ;
        RECT 2013.980 1737.100 2014.240 1737.360 ;
        RECT 1752.240 1736.760 1752.500 1737.020 ;
        RECT 1979.940 1736.760 1980.200 1737.020 ;
        RECT 1710.840 1736.420 1711.100 1736.680 ;
        RECT 1944.980 1736.420 1945.240 1736.680 ;
        RECT 1807.440 1736.080 1807.700 1736.340 ;
        RECT 2036.980 1736.080 2037.240 1736.340 ;
        RECT 1772.480 1735.740 1772.740 1736.000 ;
        RECT 2002.940 1735.740 2003.200 1736.000 ;
        RECT 1806.980 1735.400 1807.240 1735.660 ;
        RECT 2071.940 1735.400 2072.200 1735.660 ;
        RECT 1668.980 1735.060 1669.240 1735.320 ;
        RECT 2059.980 1735.060 2060.240 1735.320 ;
        RECT 2519.060 1709.900 2519.320 1710.160 ;
        RECT 2520.900 1709.900 2521.160 1710.160 ;
        RECT 2519.520 1703.780 2519.780 1704.040 ;
        RECT 2523.660 1704.120 2523.920 1704.380 ;
        RECT 1310.640 1695.620 1310.900 1695.880 ;
        RECT 1344.680 1695.620 1344.940 1695.880 ;
        RECT 990.480 1694.940 990.740 1695.200 ;
        RECT 1048.900 1694.940 1049.160 1695.200 ;
        RECT 997.380 1694.600 997.640 1694.860 ;
        RECT 1069.600 1694.600 1069.860 1694.860 ;
        RECT 1288.560 1694.600 1288.820 1694.860 ;
        RECT 1337.780 1694.600 1338.040 1694.860 ;
        RECT 996.920 1694.260 997.180 1694.520 ;
        RECT 1076.500 1694.260 1076.760 1694.520 ;
        RECT 1268.320 1694.260 1268.580 1694.520 ;
        RECT 1344.220 1694.260 1344.480 1694.520 ;
        RECT 991.400 1693.920 991.660 1694.180 ;
        RECT 1104.100 1693.920 1104.360 1694.180 ;
        RECT 1220.940 1693.920 1221.200 1694.180 ;
        RECT 1343.760 1693.920 1344.020 1694.180 ;
        RECT 990.940 1693.580 991.200 1693.840 ;
        RECT 1111.000 1693.580 1111.260 1693.840 ;
        RECT 1186.440 1693.580 1186.700 1693.840 ;
        RECT 1338.240 1693.580 1338.500 1693.840 ;
        RECT 1520.860 1690.520 1521.120 1690.780 ;
        RECT 1522.240 1690.520 1522.500 1690.780 ;
        RECT 1102.260 1689.840 1102.520 1690.100 ;
        RECT 1190.580 1689.840 1190.840 1690.100 ;
        RECT 1045.220 1689.500 1045.480 1689.760 ;
        RECT 1100.420 1689.500 1100.680 1689.760 ;
        RECT 1130.780 1689.500 1131.040 1689.760 ;
        RECT 1243.480 1689.500 1243.740 1689.760 ;
        RECT 1254.980 1689.500 1255.240 1689.760 ;
        RECT 1300.980 1689.500 1301.240 1689.760 ;
        RECT 1016.700 1689.160 1016.960 1689.420 ;
        RECT 1079.720 1689.160 1079.980 1689.420 ;
        RECT 1087.540 1689.160 1087.800 1689.420 ;
        RECT 1195.180 1689.160 1195.440 1689.420 ;
        RECT 1207.140 1689.160 1207.400 1689.420 ;
        RECT 1230.140 1689.160 1230.400 1689.420 ;
        RECT 1268.780 1689.160 1269.040 1689.420 ;
        RECT 1315.700 1689.160 1315.960 1689.420 ;
        RECT 1002.900 1688.820 1003.160 1689.080 ;
        RECT 1167.580 1688.820 1167.840 1689.080 ;
        RECT 1173.100 1688.820 1173.360 1689.080 ;
        RECT 1188.740 1688.820 1189.000 1689.080 ;
        RECT 1200.240 1688.820 1200.500 1689.080 ;
        RECT 1215.420 1688.820 1215.680 1689.080 ;
        RECT 1238.420 1688.820 1238.680 1689.080 ;
        RECT 1287.180 1688.820 1287.440 1689.080 ;
        RECT 463.780 1688.480 464.040 1688.740 ;
        RECT 468.840 1688.480 469.100 1688.740 ;
        RECT 514.380 1688.480 514.640 1688.740 ;
        RECT 517.140 1688.480 517.400 1688.740 ;
        RECT 1073.740 1688.480 1074.000 1688.740 ;
        RECT 1293.620 1688.480 1293.880 1688.740 ;
        RECT 1030.500 1688.140 1030.760 1688.400 ;
        RECT 1258.200 1688.140 1258.460 1688.400 ;
        RECT 1258.660 1688.140 1258.920 1688.400 ;
        RECT 1262.340 1688.140 1262.600 1688.400 ;
        RECT 2007.540 1687.800 2007.800 1688.060 ;
        RECT 2302.860 1687.800 2303.120 1688.060 ;
        RECT 2055.840 1687.460 2056.100 1687.720 ;
        RECT 2360.820 1687.460 2361.080 1687.720 ;
        RECT 2042.040 1687.120 2042.300 1687.380 ;
        RECT 2418.780 1687.120 2419.040 1687.380 ;
        RECT 2069.640 1686.780 2069.900 1687.040 ;
        RECT 2476.740 1686.780 2477.000 1687.040 ;
        RECT 1159.300 1686.440 1159.560 1686.700 ;
        RECT 1243.940 1686.440 1244.200 1686.700 ;
        RECT 1258.200 1686.440 1258.460 1686.700 ;
        RECT 1276.600 1686.440 1276.860 1686.700 ;
        RECT 1144.580 1686.100 1144.840 1686.360 ;
        RECT 1162.520 1686.100 1162.780 1686.360 ;
        RECT 1187.820 1686.100 1188.080 1686.360 ;
        RECT 1215.420 1686.100 1215.680 1686.360 ;
        RECT 1167.580 1685.760 1167.840 1686.020 ;
        RECT 1190.120 1685.760 1190.380 1686.020 ;
        RECT 1195.180 1685.760 1195.440 1686.020 ;
        RECT 1224.620 1685.760 1224.880 1686.020 ;
        RECT 1116.060 1684.060 1116.320 1684.320 ;
        RECT 1148.720 1684.060 1148.980 1684.320 ;
        RECT 1220.480 1684.060 1220.740 1684.320 ;
        RECT 1243.020 1684.060 1243.280 1684.320 ;
        RECT 1272.460 1684.060 1272.720 1684.320 ;
        RECT 1291.320 1684.060 1291.580 1684.320 ;
        RECT 1288.560 1656.180 1288.820 1656.440 ;
        RECT 1521.320 1656.180 1521.580 1656.440 ;
        RECT 1520.860 1655.840 1521.120 1656.100 ;
        RECT 2518.140 1655.840 2518.400 1656.100 ;
        RECT 2519.980 1655.840 2520.240 1656.100 ;
        RECT 1289.020 1655.500 1289.280 1655.760 ;
        RECT 1441.740 1642.240 1442.000 1642.500 ;
        RECT 1443.120 1642.240 1443.380 1642.500 ;
        RECT 2517.680 1641.900 2517.940 1642.160 ;
        RECT 2518.600 1641.900 2518.860 1642.160 ;
        RECT 1441.740 1617.760 1442.000 1618.020 ;
        RECT 1442.660 1617.760 1442.920 1618.020 ;
        RECT 2519.980 1617.760 2520.240 1618.020 ;
        RECT 2520.900 1617.760 2521.160 1618.020 ;
        RECT 1520.860 1607.560 1521.120 1607.820 ;
        RECT 1521.320 1607.560 1521.580 1607.820 ;
        RECT 1289.020 1594.980 1289.280 1595.240 ;
        RECT 1441.740 1593.960 1442.000 1594.220 ;
        RECT 1442.660 1593.960 1442.920 1594.220 ;
        RECT 2517.680 1593.960 2517.940 1594.220 ;
        RECT 2518.600 1593.960 2518.860 1594.220 ;
        RECT 2519.980 1593.960 2520.240 1594.220 ;
        RECT 2520.900 1593.960 2521.160 1594.220 ;
        RECT 1289.020 1593.620 1289.280 1593.880 ;
        RECT 1521.320 1593.620 1521.580 1593.880 ;
        RECT 1522.700 1593.620 1522.960 1593.880 ;
        RECT 1289.020 1586.820 1289.280 1587.080 ;
        RECT 1290.400 1586.820 1290.660 1587.080 ;
        RECT 1440.360 1569.480 1440.620 1569.740 ;
        RECT 1441.740 1569.480 1442.000 1569.740 ;
        RECT 2517.220 1569.480 2517.480 1569.740 ;
        RECT 2518.600 1569.480 2518.860 1569.740 ;
        RECT 2518.140 1559.280 2518.400 1559.540 ;
        RECT 2519.980 1559.280 2520.240 1559.540 ;
        RECT 1289.020 1558.600 1289.280 1558.860 ;
        RECT 1290.400 1558.600 1290.660 1558.860 ;
        RECT 2518.140 1558.600 2518.400 1558.860 ;
        RECT 2519.980 1558.600 2520.240 1558.860 ;
        RECT 1521.320 1546.020 1521.580 1546.280 ;
        RECT 1522.700 1546.020 1522.960 1546.280 ;
        RECT 1440.360 1545.680 1440.620 1545.940 ;
        RECT 1440.820 1545.680 1441.080 1545.940 ;
        RECT 2517.220 1545.680 2517.480 1545.940 ;
        RECT 2519.060 1545.680 2519.320 1545.940 ;
        RECT 1521.320 1545.340 1521.580 1545.600 ;
        RECT 1522.240 1545.340 1522.500 1545.600 ;
        RECT 1440.360 1545.000 1440.620 1545.260 ;
        RECT 1440.820 1545.000 1441.080 1545.260 ;
        RECT 1288.560 1538.540 1288.820 1538.800 ;
        RECT 1289.020 1538.540 1289.280 1538.800 ;
        RECT 1440.360 1497.400 1440.620 1497.660 ;
        RECT 1441.740 1497.400 1442.000 1497.660 ;
        RECT 1521.320 1497.060 1521.580 1497.320 ;
        RECT 1522.700 1497.060 1522.960 1497.320 ;
        RECT 1288.560 1490.600 1288.820 1490.860 ;
        RECT 1289.480 1490.600 1289.740 1490.860 ;
        RECT 1440.360 1472.920 1440.620 1473.180 ;
        RECT 1441.740 1472.920 1442.000 1473.180 ;
        RECT 1521.320 1449.460 1521.580 1449.720 ;
        RECT 1522.700 1449.460 1522.960 1449.720 ;
        RECT 1440.360 1449.120 1440.620 1449.380 ;
        RECT 1440.820 1449.120 1441.080 1449.380 ;
        RECT 1521.320 1448.780 1521.580 1449.040 ;
        RECT 1522.240 1448.780 1522.500 1449.040 ;
        RECT 1440.820 1448.440 1441.080 1448.700 ;
        RECT 1442.660 1448.440 1442.920 1448.700 ;
        RECT 1289.020 1441.980 1289.280 1442.240 ;
        RECT 1289.480 1441.980 1289.740 1442.240 ;
        RECT 2518.600 1415.120 2518.860 1415.380 ;
        RECT 2519.060 1414.780 2519.320 1415.040 ;
        RECT 1289.020 1414.440 1289.280 1414.700 ;
        RECT 1289.940 1414.440 1290.200 1414.700 ;
        RECT 1521.320 1400.500 1521.580 1400.760 ;
        RECT 1522.700 1400.500 1522.960 1400.760 ;
        RECT 1441.740 1386.900 1442.000 1387.160 ;
        RECT 1442.660 1386.900 1442.920 1387.160 ;
        RECT 2518.140 1366.500 2518.400 1366.760 ;
        RECT 2519.980 1366.500 2520.240 1366.760 ;
        RECT 2518.140 1365.820 2518.400 1366.080 ;
        RECT 2519.980 1365.820 2520.240 1366.080 ;
        RECT 1521.320 1352.900 1521.580 1353.160 ;
        RECT 1522.700 1352.900 1522.960 1353.160 ;
        RECT 1289.020 1352.220 1289.280 1352.480 ;
        RECT 1289.940 1352.220 1290.200 1352.480 ;
        RECT 1521.320 1352.220 1521.580 1352.480 ;
        RECT 1522.700 1352.220 1522.960 1352.480 ;
        RECT 2518.600 1318.220 2518.860 1318.480 ;
        RECT 2519.980 1318.220 2520.240 1318.480 ;
        RECT 1289.020 1317.540 1289.280 1317.800 ;
        RECT 1289.940 1317.540 1290.200 1317.800 ;
        RECT 2518.600 1317.540 2518.860 1317.800 ;
        RECT 2519.980 1317.540 2520.240 1317.800 ;
        RECT 1521.320 1317.200 1521.580 1317.460 ;
        RECT 1522.700 1317.200 1522.960 1317.460 ;
        RECT 1289.020 1303.940 1289.280 1304.200 ;
        RECT 1290.400 1303.940 1290.660 1304.200 ;
        RECT 1521.320 1303.940 1521.580 1304.200 ;
        RECT 1522.700 1303.940 1522.960 1304.200 ;
        RECT 1440.820 1290.000 1441.080 1290.260 ;
        RECT 1441.740 1290.000 1442.000 1290.260 ;
        RECT 2518.140 1269.940 2518.400 1270.200 ;
        RECT 2519.980 1269.940 2520.240 1270.200 ;
        RECT 2518.140 1269.260 2518.400 1269.520 ;
        RECT 2519.980 1269.260 2520.240 1269.520 ;
        RECT 1289.020 1268.920 1289.280 1269.180 ;
        RECT 1290.400 1268.920 1290.660 1269.180 ;
        RECT 1287.640 1255.660 1287.900 1255.920 ;
        RECT 1289.020 1255.660 1289.280 1255.920 ;
        RECT 1440.360 1242.060 1440.620 1242.320 ;
        RECT 1440.820 1242.060 1441.080 1242.320 ;
        RECT 2518.600 1222.000 2518.860 1222.260 ;
        RECT 2519.060 1221.660 2519.320 1221.920 ;
        RECT 1440.360 1220.640 1440.620 1220.900 ;
        RECT 1441.740 1220.640 1442.000 1220.900 ;
        RECT 1287.640 1207.380 1287.900 1207.640 ;
        RECT 1288.560 1207.380 1288.820 1207.640 ;
        RECT 1520.860 1207.380 1521.120 1207.640 ;
        RECT 1521.780 1207.380 1522.040 1207.640 ;
        RECT 1519.480 1206.700 1519.740 1206.960 ;
        RECT 1520.860 1206.700 1521.120 1206.960 ;
        RECT 2518.140 1173.380 2518.400 1173.640 ;
        RECT 2519.980 1173.380 2520.240 1173.640 ;
        RECT 1288.560 1173.040 1288.820 1173.300 ;
        RECT 2518.140 1172.700 2518.400 1172.960 ;
        RECT 2519.980 1172.700 2520.240 1172.960 ;
        RECT 1289.020 1172.360 1289.280 1172.620 ;
        RECT 1519.480 1159.100 1519.740 1159.360 ;
        RECT 1520.860 1159.100 1521.120 1159.360 ;
        RECT 2518.600 1125.440 2518.860 1125.700 ;
        RECT 2519.060 1125.100 2519.320 1125.360 ;
        RECT 1288.560 1124.760 1288.820 1125.020 ;
        RECT 1521.320 1124.760 1521.580 1125.020 ;
        RECT 1289.020 1124.420 1289.280 1124.680 ;
        RECT 1521.780 1124.080 1522.040 1124.340 ;
        RECT 1288.560 1110.820 1288.820 1111.080 ;
        RECT 1289.020 1110.820 1289.280 1111.080 ;
        RECT 1441.740 1110.820 1442.000 1111.080 ;
        RECT 1442.660 1110.820 1442.920 1111.080 ;
        RECT 1520.400 1079.880 1520.660 1080.140 ;
        RECT 1521.320 1079.880 1521.580 1080.140 ;
        RECT 2518.140 1076.820 2518.400 1077.080 ;
        RECT 2519.980 1076.820 2520.240 1077.080 ;
        RECT 1288.560 1076.480 1288.820 1076.740 ;
        RECT 2518.140 1076.140 2518.400 1076.400 ;
        RECT 2519.980 1076.140 2520.240 1076.400 ;
        RECT 1289.020 1075.800 1289.280 1076.060 ;
        RECT 1440.360 1062.540 1440.620 1062.800 ;
        RECT 1440.820 1062.540 1441.080 1062.800 ;
        RECT 2082.060 1062.540 2082.320 1062.800 ;
        RECT 2083.440 1062.540 2083.700 1062.800 ;
        RECT 1454.620 1052.000 1454.880 1052.260 ;
        RECT 1455.540 1052.000 1455.800 1052.260 ;
        RECT 1062.240 1051.660 1062.500 1051.920 ;
        RECT 1098.580 1051.660 1098.840 1051.920 ;
        RECT 1220.020 1048.600 1220.280 1048.860 ;
        RECT 1220.940 1048.600 1221.200 1048.860 ;
        RECT 2518.600 1028.880 2518.860 1029.140 ;
        RECT 2519.060 1028.540 2519.320 1028.800 ;
        RECT 632.140 1028.200 632.400 1028.460 ;
        RECT 632.140 1027.520 632.400 1027.780 ;
        RECT 1288.560 1028.200 1288.820 1028.460 ;
        RECT 2518.600 1028.200 2518.860 1028.460 ;
        RECT 2519.980 1028.200 2520.240 1028.460 ;
        RECT 1289.020 1027.860 1289.280 1028.120 ;
        RECT 983.580 1026.500 983.840 1026.760 ;
        RECT 1134.460 1026.500 1134.720 1026.760 ;
        RECT 983.120 1026.160 983.380 1026.420 ;
        RECT 1139.520 1026.160 1139.780 1026.420 ;
        RECT 979.440 1025.820 979.700 1026.080 ;
        RECT 1143.200 1025.820 1143.460 1026.080 ;
        RECT 978.520 1025.480 978.780 1025.740 ;
        RECT 1147.800 1025.480 1148.060 1025.740 ;
        RECT 978.980 1025.140 979.240 1025.400 ;
        RECT 1152.400 1025.140 1152.660 1025.400 ;
        RECT 1196.100 1025.140 1196.360 1025.400 ;
        RECT 1200.240 1025.140 1200.500 1025.400 ;
        RECT 977.600 1024.800 977.860 1025.060 ;
        RECT 1156.080 1024.800 1156.340 1025.060 ;
        RECT 978.060 1024.460 978.320 1024.720 ;
        RECT 1166.200 1024.460 1166.460 1024.720 ;
        RECT 1472.100 1021.060 1472.360 1021.320 ;
        RECT 1704.400 1021.060 1704.660 1021.320 ;
        RECT 1728.780 1021.060 1729.040 1021.320 ;
        RECT 2085.280 1021.060 2085.540 1021.320 ;
        RECT 1278.900 1020.720 1279.160 1020.980 ;
        RECT 1341.000 1020.720 1341.260 1020.980 ;
        RECT 1489.580 1020.720 1489.840 1020.980 ;
        RECT 1521.320 1020.720 1521.580 1020.980 ;
        RECT 1533.280 1020.720 1533.540 1020.980 ;
        RECT 1902.200 1020.720 1902.460 1020.980 ;
        RECT 1267.860 1020.380 1268.120 1020.640 ;
        RECT 1345.140 1020.380 1345.400 1020.640 ;
        RECT 1507.060 1020.380 1507.320 1020.640 ;
        RECT 1898.060 1020.380 1898.320 1020.640 ;
        RECT 1252.680 1020.040 1252.940 1020.300 ;
        RECT 1339.620 1020.040 1339.880 1020.300 ;
        RECT 1495.100 1020.040 1495.360 1020.300 ;
        RECT 1901.740 1020.040 1902.000 1020.300 ;
        RECT 995.080 1019.700 995.340 1019.960 ;
        RECT 1193.800 1019.700 1194.060 1019.960 ;
        RECT 1237.960 1019.700 1238.220 1019.960 ;
        RECT 1340.540 1019.700 1340.800 1019.960 ;
        RECT 1474.400 1019.700 1474.660 1019.960 ;
        RECT 1887.020 1019.700 1887.280 1019.960 ;
        RECT 988.640 1019.360 988.900 1019.620 ;
        RECT 1285.800 1019.360 1286.060 1019.620 ;
        RECT 1461.060 1019.360 1461.320 1019.620 ;
        RECT 1898.980 1019.360 1899.240 1019.620 ;
        RECT 990.020 1019.020 990.280 1019.280 ;
        RECT 1301.900 1019.020 1302.160 1019.280 ;
        RECT 1462.440 1019.020 1462.700 1019.280 ;
        RECT 1899.440 1019.020 1899.700 1019.280 ;
        RECT 992.320 1018.680 992.580 1018.940 ;
        RECT 1313.860 1018.680 1314.120 1018.940 ;
        RECT 1434.840 1018.680 1435.100 1018.940 ;
        RECT 1886.560 1018.680 1886.820 1018.940 ;
        RECT 987.260 1018.340 987.520 1018.600 ;
        RECT 1314.780 1018.340 1315.040 1018.600 ;
        RECT 1437.600 1018.340 1437.860 1018.600 ;
        RECT 1898.520 1018.340 1898.780 1018.600 ;
        RECT 989.100 1018.000 989.360 1018.260 ;
        RECT 1326.280 1018.000 1326.540 1018.260 ;
        RECT 1358.940 1018.000 1359.200 1018.260 ;
        RECT 1849.300 1018.000 1849.560 1018.260 ;
        RECT 991.860 1017.660 992.120 1017.920 ;
        RECT 1337.780 1017.660 1338.040 1017.920 ;
        RECT 1402.640 1017.660 1402.900 1017.920 ;
        RECT 1899.900 1017.660 1900.160 1017.920 ;
        RECT 1567.780 1017.320 1568.040 1017.580 ;
        RECT 1897.600 1017.320 1897.860 1017.580 ;
        RECT 1480.840 1016.980 1481.100 1017.240 ;
        RECT 1766.500 1016.980 1766.760 1017.240 ;
        RECT 1614.700 1016.640 1614.960 1016.900 ;
        RECT 1900.820 1016.640 1901.080 1016.900 ;
        RECT 1514.420 1016.300 1514.680 1016.560 ;
        RECT 1656.100 1016.300 1656.360 1016.560 ;
        RECT 1490.040 1015.960 1490.300 1016.220 ;
        RECT 1625.740 1015.960 1626.000 1016.220 ;
        RECT 1288.560 1014.260 1288.820 1014.520 ;
        RECT 1289.020 1014.260 1289.280 1014.520 ;
        RECT 810.620 1013.920 810.880 1014.180 ;
        RECT 845.580 1013.920 845.840 1014.180 ;
        RECT 994.620 1013.920 994.880 1014.180 ;
        RECT 997.380 1013.920 997.640 1014.180 ;
        RECT 1000.140 1013.920 1000.400 1014.180 ;
        RECT 1197.940 1013.920 1198.200 1014.180 ;
        RECT 1198.400 1013.920 1198.660 1014.180 ;
        RECT 1200.700 1013.920 1200.960 1014.180 ;
        RECT 1202.540 1013.920 1202.800 1014.180 ;
        RECT 1207.140 1013.920 1207.400 1014.180 ;
        RECT 1214.960 1013.920 1215.220 1014.180 ;
        RECT 1220.480 1013.920 1220.740 1014.180 ;
        RECT 1259.120 1013.920 1259.380 1014.180 ;
        RECT 984.500 1013.580 984.760 1013.840 ;
        RECT 1208.980 1013.580 1209.240 1013.840 ;
        RECT 1262.340 1013.580 1262.600 1013.840 ;
        RECT 1269.240 1013.580 1269.500 1013.840 ;
        RECT 1284.880 1013.920 1285.140 1014.180 ;
        RECT 1300.980 1014.260 1301.240 1014.520 ;
        RECT 1294.080 1013.920 1294.340 1014.180 ;
        RECT 1333.640 1013.920 1333.900 1014.180 ;
        RECT 1361.240 1013.920 1361.500 1014.180 ;
        RECT 1365.840 1013.920 1366.100 1014.180 ;
        RECT 1452.780 1013.920 1453.040 1014.180 ;
        RECT 1455.080 1013.920 1455.340 1014.180 ;
        RECT 1456.920 1013.920 1457.180 1014.180 ;
        RECT 1461.520 1013.920 1461.780 1014.180 ;
        RECT 1465.660 1013.920 1465.920 1014.180 ;
        RECT 1473.020 1013.920 1473.280 1014.180 ;
        RECT 1479.000 1013.920 1479.260 1014.180 ;
        RECT 1482.220 1013.920 1482.480 1014.180 ;
        RECT 1339.160 1013.580 1339.420 1013.840 ;
        RECT 1446.340 1013.580 1446.600 1013.840 ;
        RECT 1459.220 1013.580 1459.480 1013.840 ;
        RECT 999.220 1013.240 999.480 1013.500 ;
        RECT 1197.480 1013.240 1197.740 1013.500 ;
        RECT 1197.940 1013.240 1198.200 1013.500 ;
        RECT 1226.000 1013.240 1226.260 1013.500 ;
        RECT 1244.860 1013.240 1245.120 1013.500 ;
        RECT 988.180 1012.900 988.440 1013.160 ;
        RECT 1223.700 1012.900 1223.960 1013.160 ;
        RECT 1224.160 1012.900 1224.420 1013.160 ;
        RECT 1259.580 1012.900 1259.840 1013.160 ;
        RECT 1265.560 1012.900 1265.820 1013.160 ;
        RECT 1268.780 1012.900 1269.040 1013.160 ;
        RECT 1292.700 1013.240 1292.960 1013.500 ;
        RECT 1333.180 1013.240 1333.440 1013.500 ;
        RECT 1341.460 1012.900 1341.720 1013.160 ;
        RECT 1444.040 1012.900 1444.300 1013.160 ;
        RECT 1489.580 1013.920 1489.840 1014.180 ;
        RECT 1493.720 1013.920 1493.980 1014.180 ;
        RECT 1494.640 1013.920 1494.900 1014.180 ;
        RECT 1507.520 1013.920 1507.780 1014.180 ;
        RECT 1528.220 1013.920 1528.480 1014.180 ;
        RECT 1545.700 1013.920 1545.960 1014.180 ;
        RECT 1548.000 1013.920 1548.260 1014.180 ;
        RECT 1559.500 1013.920 1559.760 1014.180 ;
        RECT 1562.720 1013.920 1562.980 1014.180 ;
        RECT 1574.220 1013.920 1574.480 1014.180 ;
        RECT 1577.900 1013.920 1578.160 1014.180 ;
        RECT 1578.360 1013.920 1578.620 1014.180 ;
        RECT 1886.100 1013.920 1886.360 1014.180 ;
        RECT 2002.940 1013.920 2003.200 1014.180 ;
        RECT 2007.540 1013.920 2007.800 1014.180 ;
        RECT 1495.560 1013.580 1495.820 1013.840 ;
        RECT 1511.660 1013.580 1511.920 1013.840 ;
        RECT 1517.180 1013.580 1517.440 1013.840 ;
        RECT 1591.700 1013.580 1591.960 1013.840 ;
        RECT 1596.300 1013.580 1596.560 1013.840 ;
        RECT 1600.440 1013.580 1600.700 1013.840 ;
        RECT 1665.760 1013.580 1666.020 1013.840 ;
        RECT 1669.440 1013.580 1669.700 1013.840 ;
        RECT 1755.000 1013.580 1755.260 1013.840 ;
        RECT 1759.140 1013.580 1759.400 1013.840 ;
        RECT 1759.600 1013.580 1759.860 1013.840 ;
        RECT 2085.740 1013.580 2086.000 1013.840 ;
        RECT 1496.020 1013.240 1496.280 1013.500 ;
        RECT 1518.560 1013.240 1518.820 1013.500 ;
        RECT 1498.320 1012.900 1498.580 1013.160 ;
        RECT 1628.500 1013.240 1628.760 1013.500 ;
        RECT 1720.040 1013.240 1720.300 1013.500 ;
        RECT 2084.360 1013.240 2084.620 1013.500 ;
        RECT 1524.080 1012.900 1524.340 1013.160 ;
        RECT 1693.820 1012.900 1694.080 1013.160 ;
        RECT 1707.160 1012.900 1707.420 1013.160 ;
        RECT 1710.840 1012.900 1711.100 1013.160 ;
        RECT 1715.440 1012.900 1715.700 1013.160 ;
        RECT 1717.740 1012.900 1718.000 1013.160 ;
        RECT 1733.380 1012.900 1733.640 1013.160 ;
        RECT 1737.980 1012.900 1738.240 1013.160 ;
        RECT 1738.900 1012.900 1739.160 1013.160 ;
        RECT 2077.000 1012.900 2077.260 1013.160 ;
        RECT 796.820 1012.560 797.080 1012.820 ;
        RECT 884.680 1012.560 884.940 1012.820 ;
        RECT 987.720 1012.560 987.980 1012.820 ;
        RECT 1228.300 1012.560 1228.560 1012.820 ;
        RECT 1237.500 1012.560 1237.760 1012.820 ;
        RECT 1338.700 1012.560 1338.960 1012.820 ;
        RECT 1357.100 1012.560 1357.360 1012.820 ;
        RECT 1362.620 1012.560 1362.880 1012.820 ;
        RECT 1496.940 1012.560 1497.200 1012.820 ;
        RECT 1517.180 1012.560 1517.440 1012.820 ;
        RECT 803.720 1012.220 803.980 1012.480 ;
        RECT 890.200 1012.220 890.460 1012.480 ;
        RECT 986.800 1012.220 987.060 1012.480 ;
        RECT 1224.160 1012.220 1224.420 1012.480 ;
        RECT 1224.620 1012.220 1224.880 1012.480 ;
        RECT 1230.140 1012.220 1230.400 1012.480 ;
        RECT 1243.940 1012.220 1244.200 1012.480 ;
        RECT 1284.880 1012.220 1285.140 1012.480 ;
        RECT 789.920 1011.880 790.180 1012.140 ;
        RECT 910.900 1011.880 911.160 1012.140 ;
        RECT 996.000 1011.880 996.260 1012.140 ;
        RECT 1270.160 1011.880 1270.420 1012.140 ;
        RECT 1276.140 1011.880 1276.400 1012.140 ;
        RECT 1294.540 1012.220 1294.800 1012.480 ;
        RECT 769.220 1011.540 769.480 1011.800 ;
        RECT 906.300 1011.540 906.560 1011.800 ;
        RECT 1000.140 1011.540 1000.400 1011.800 ;
        RECT 1075.580 1011.540 1075.840 1011.800 ;
        RECT 1079.720 1011.540 1079.980 1011.800 ;
        RECT 1081.100 1011.540 1081.360 1011.800 ;
        RECT 1104.100 1011.540 1104.360 1011.800 ;
        RECT 1106.400 1011.540 1106.660 1011.800 ;
        RECT 1106.860 1011.540 1107.120 1011.800 ;
        RECT 1145.500 1011.540 1145.760 1011.800 ;
        RECT 1169.420 1011.540 1169.680 1011.800 ;
        RECT 700.220 1011.200 700.480 1011.460 ;
        RECT 841.900 1011.200 842.160 1011.460 ;
        RECT 997.380 1011.200 997.640 1011.460 ;
        RECT 1076.040 1011.200 1076.300 1011.460 ;
        RECT 1076.960 1011.200 1077.220 1011.460 ;
        RECT 1145.960 1011.200 1146.220 1011.460 ;
        RECT 1166.660 1011.200 1166.920 1011.460 ;
        RECT 1243.940 1011.200 1244.200 1011.460 ;
        RECT 1262.340 1011.540 1262.600 1011.800 ;
        RECT 1341.920 1012.220 1342.180 1012.480 ;
        RECT 1369.980 1012.220 1370.240 1012.480 ;
        RECT 1372.740 1012.220 1373.000 1012.480 ;
        RECT 1384.700 1012.220 1384.960 1012.480 ;
        RECT 1386.540 1012.220 1386.800 1012.480 ;
        RECT 1393.440 1012.220 1393.700 1012.480 ;
        RECT 1397.120 1012.220 1397.380 1012.480 ;
        RECT 1404.940 1012.220 1405.200 1012.480 ;
        RECT 1406.780 1012.220 1407.040 1012.480 ;
        RECT 1488.660 1012.220 1488.920 1012.480 ;
        RECT 1516.720 1012.220 1516.980 1012.480 ;
        RECT 1295.920 1011.880 1296.180 1012.140 ;
        RECT 1342.380 1011.880 1342.640 1012.140 ;
        RECT 1376.420 1011.880 1376.680 1012.140 ;
        RECT 1432.080 1011.880 1432.340 1012.140 ;
        RECT 1509.360 1011.880 1509.620 1012.140 ;
        RECT 1866.320 1012.560 1866.580 1012.820 ;
        RECT 1524.540 1012.220 1524.800 1012.480 ;
        RECT 1545.700 1012.220 1545.960 1012.480 ;
        RECT 1553.060 1012.220 1553.320 1012.480 ;
        RECT 1556.280 1012.220 1556.540 1012.480 ;
        RECT 1556.740 1012.220 1557.000 1012.480 ;
        RECT 1887.480 1012.560 1887.740 1012.820 ;
        RECT 2004.780 1012.560 2005.040 1012.820 ;
        RECT 2073.320 1012.560 2073.580 1012.820 ;
        RECT 1872.300 1012.220 1872.560 1012.480 ;
        RECT 1876.440 1012.220 1876.700 1012.480 ;
        RECT 1518.560 1011.880 1518.820 1012.140 ;
        RECT 1525.460 1011.880 1525.720 1012.140 ;
        RECT 1535.120 1011.880 1535.380 1012.140 ;
        RECT 1542.020 1011.880 1542.280 1012.140 ;
        RECT 1542.480 1011.880 1542.740 1012.140 ;
        RECT 1614.700 1011.880 1614.960 1012.140 ;
        RECT 1662.540 1011.880 1662.800 1012.140 ;
        RECT 1289.480 1011.200 1289.740 1011.460 ;
        RECT 517.140 1010.860 517.400 1011.120 ;
        RECT 712.640 1010.860 712.900 1011.120 ;
        RECT 755.420 1010.860 755.680 1011.120 ;
        RECT 901.700 1010.860 901.960 1011.120 ;
        RECT 994.160 1010.860 994.420 1011.120 ;
        RECT 1309.720 1011.200 1309.980 1011.460 ;
        RECT 1290.400 1010.860 1290.660 1011.120 ;
        RECT 1334.100 1011.540 1334.360 1011.800 ;
        RECT 1378.720 1011.540 1378.980 1011.800 ;
        RECT 1431.620 1011.540 1431.880 1011.800 ;
        RECT 1500.620 1011.540 1500.880 1011.800 ;
        RECT 1865.860 1011.540 1866.120 1011.800 ;
        RECT 1866.320 1011.540 1866.580 1011.800 ;
        RECT 1894.840 1011.540 1895.100 1011.800 ;
        RECT 2061.360 1011.880 2061.620 1012.140 ;
        RECT 2287.220 1012.220 2287.480 1012.480 ;
        RECT 2078.840 1011.880 2079.100 1012.140 ;
        RECT 2082.980 1011.880 2083.240 1012.140 ;
        RECT 2087.580 1011.880 2087.840 1012.140 ;
        RECT 2090.340 1011.880 2090.600 1012.140 ;
        RECT 2083.900 1011.540 2084.160 1011.800 ;
        RECT 1386.540 1011.200 1386.800 1011.460 ;
        RECT 1890.700 1011.200 1890.960 1011.460 ;
        RECT 2074.700 1011.200 2074.960 1011.460 ;
        RECT 2519.520 1011.540 2519.780 1011.800 ;
        RECT 1320.300 1010.860 1320.560 1011.120 ;
        RECT 1342.840 1010.860 1343.100 1011.120 ;
        RECT 1354.800 1010.860 1355.060 1011.120 ;
        RECT 1873.220 1010.860 1873.480 1011.120 ;
        RECT 468.840 1010.520 469.100 1010.780 ;
        RECT 673.540 1010.520 673.800 1010.780 ;
        RECT 734.720 1010.520 734.980 1010.780 ;
        RECT 893.420 1010.520 893.680 1010.780 ;
        RECT 989.560 1010.520 989.820 1010.780 ;
        RECT 1347.440 1010.520 1347.700 1010.780 ;
        RECT 1417.820 1010.520 1418.080 1010.780 ;
        RECT 1700.720 1010.520 1700.980 1010.780 ;
        RECT 1710.840 1010.520 1711.100 1010.780 ;
        RECT 1738.900 1010.520 1739.160 1010.780 ;
        RECT 1741.660 1010.520 1741.920 1010.780 ;
        RECT 1759.600 1010.520 1759.860 1010.780 ;
        RECT 1767.880 1010.520 1768.140 1010.780 ;
        RECT 1772.940 1010.520 1773.200 1010.780 ;
        RECT 1830.900 1010.520 1831.160 1010.780 ;
        RECT 1835.040 1010.520 1835.300 1010.780 ;
        RECT 1865.860 1010.520 1866.120 1010.780 ;
        RECT 1891.620 1010.860 1891.880 1011.120 ;
        RECT 2055.380 1010.860 2055.640 1011.120 ;
        RECT 2519.060 1011.200 2519.320 1011.460 ;
        RECT 2085.280 1010.860 2085.540 1011.120 ;
        RECT 2518.600 1010.860 2518.860 1011.120 ;
        RECT 1883.340 1010.520 1883.600 1010.780 ;
        RECT 2532.400 1010.520 2532.660 1010.780 ;
        RECT 995.540 1010.180 995.800 1010.440 ;
        RECT 999.220 1010.180 999.480 1010.440 ;
        RECT 999.680 1010.180 999.940 1010.440 ;
        RECT 1146.420 1010.180 1146.680 1010.440 ;
        RECT 1204.840 1010.180 1205.100 1010.440 ;
        RECT 1336.860 1010.180 1337.120 1010.440 ;
        RECT 1447.720 1010.180 1447.980 1010.440 ;
        RECT 1520.860 1010.180 1521.120 1010.440 ;
        RECT 998.760 1009.840 999.020 1010.100 ;
        RECT 1151.020 1009.840 1151.280 1010.100 ;
        RECT 993.240 1009.500 993.500 1009.760 ;
        RECT 1080.180 1009.500 1080.440 1009.760 ;
        RECT 1081.100 1009.500 1081.360 1009.760 ;
        RECT 1160.220 1009.840 1160.480 1010.100 ;
        RECT 1183.220 1009.840 1183.480 1010.100 ;
        RECT 1186.440 1009.840 1186.700 1010.100 ;
        RECT 1223.240 1009.840 1223.500 1010.100 ;
        RECT 1340.080 1009.840 1340.340 1010.100 ;
        RECT 1503.840 1009.840 1504.100 1010.100 ;
        RECT 1556.740 1010.180 1557.000 1010.440 ;
        RECT 1576.520 1010.180 1576.780 1010.440 ;
        RECT 1579.740 1010.180 1580.000 1010.440 ;
        RECT 1580.200 1010.180 1580.460 1010.440 ;
        RECT 1585.720 1010.180 1585.980 1010.440 ;
        RECT 1593.080 1010.180 1593.340 1010.440 ;
        RECT 1686.920 1010.180 1687.180 1010.440 ;
        RECT 1749.940 1010.180 1750.200 1010.440 ;
        RECT 1752.240 1010.180 1752.500 1010.440 ;
        RECT 1763.740 1010.180 1764.000 1010.440 ;
        RECT 1766.040 1010.180 1766.300 1010.440 ;
        RECT 1176.320 1009.500 1176.580 1009.760 ;
        RECT 1205.300 1009.500 1205.560 1009.760 ;
        RECT 993.700 1009.160 993.960 1009.420 ;
        RECT 1058.560 1009.160 1058.820 1009.420 ;
        RECT 1069.600 1009.160 1069.860 1009.420 ;
        RECT 1071.900 1009.160 1072.160 1009.420 ;
        RECT 1077.420 1009.160 1077.680 1009.420 ;
        RECT 1106.860 1009.160 1107.120 1009.420 ;
        RECT 1200.240 1009.160 1200.500 1009.420 ;
        RECT 1210.360 1009.500 1210.620 1009.760 ;
        RECT 1238.420 1009.500 1238.680 1009.760 ;
        RECT 1274.300 1009.500 1274.560 1009.760 ;
        RECT 1334.560 1009.500 1334.820 1009.760 ;
        RECT 1489.120 1009.500 1489.380 1009.760 ;
        RECT 1524.540 1009.500 1524.800 1009.760 ;
        RECT 1210.820 1009.160 1211.080 1009.420 ;
        RECT 1279.820 1009.160 1280.080 1009.420 ;
        RECT 1320.300 1009.160 1320.560 1009.420 ;
        RECT 984.040 1008.820 984.300 1009.080 ;
        RECT 1079.720 1008.820 1079.980 1009.080 ;
        RECT 1098.580 1008.820 1098.840 1009.080 ;
        RECT 1111.460 1008.820 1111.720 1009.080 ;
        RECT 1145.960 1008.820 1146.220 1009.080 ;
        RECT 1159.760 1008.820 1160.020 1009.080 ;
        RECT 1162.520 1008.820 1162.780 1009.080 ;
        RECT 1183.680 1008.820 1183.940 1009.080 ;
        RECT 1190.580 1008.820 1190.840 1009.080 ;
        RECT 1207.600 1008.820 1207.860 1009.080 ;
        RECT 1209.440 1008.820 1209.700 1009.080 ;
        RECT 1304.200 1008.820 1304.460 1009.080 ;
        RECT 996.460 1008.480 996.720 1008.740 ;
        RECT 1097.660 1008.480 1097.920 1008.740 ;
        RECT 1100.880 1008.480 1101.140 1008.740 ;
        RECT 1159.300 1008.480 1159.560 1008.740 ;
        RECT 1161.140 1008.480 1161.400 1008.740 ;
        RECT 1269.240 1008.480 1269.500 1008.740 ;
        RECT 1318.000 1008.480 1318.260 1008.740 ;
        RECT 997.840 1008.140 998.100 1008.400 ;
        RECT 1093.060 1008.140 1093.320 1008.400 ;
        RECT 1148.720 1008.140 1148.980 1008.400 ;
        RECT 1186.900 1008.140 1187.160 1008.400 ;
        RECT 1190.120 1008.140 1190.380 1008.400 ;
        RECT 1207.600 1008.140 1207.860 1008.400 ;
        RECT 1208.060 1008.140 1208.320 1008.400 ;
        RECT 1209.440 1008.140 1209.700 1008.400 ;
        RECT 1297.300 1008.140 1297.560 1008.400 ;
        RECT 1300.520 1008.140 1300.780 1008.400 ;
        RECT 1337.320 1009.160 1337.580 1009.420 ;
        RECT 1487.740 1009.160 1488.000 1009.420 ;
        RECT 1530.980 1009.160 1531.240 1009.420 ;
        RECT 1331.340 1008.820 1331.600 1009.080 ;
        RECT 1345.600 1008.820 1345.860 1009.080 ;
        RECT 1497.860 1008.820 1498.120 1009.080 ;
        RECT 1576.980 1009.840 1577.240 1010.100 ;
        RECT 1591.700 1009.840 1591.960 1010.100 ;
        RECT 1603.200 1009.840 1603.460 1010.100 ;
        RECT 1758.680 1009.840 1758.940 1010.100 ;
        RECT 2086.200 1010.180 2086.460 1010.440 ;
        RECT 1826.760 1009.840 1827.020 1010.100 ;
        RECT 1845.620 1009.840 1845.880 1010.100 ;
        RECT 1878.740 1009.840 1879.000 1010.100 ;
        RECT 1893.920 1009.840 1894.180 1010.100 ;
        RECT 1531.900 1009.500 1532.160 1009.760 ;
        RECT 1542.480 1009.500 1542.740 1009.760 ;
        RECT 1555.820 1009.500 1556.080 1009.760 ;
        RECT 1652.420 1009.500 1652.680 1009.760 ;
        RECT 1789.500 1009.500 1789.760 1009.760 ;
        RECT 2084.820 1009.500 2085.080 1009.760 ;
        RECT 1325.820 1008.480 1326.080 1008.740 ;
        RECT 1335.940 1008.480 1336.200 1008.740 ;
        RECT 1491.880 1008.480 1492.140 1008.740 ;
        RECT 1524.080 1008.480 1524.340 1008.740 ;
        RECT 1525.000 1008.480 1525.260 1008.740 ;
        RECT 1528.220 1008.480 1528.480 1008.740 ;
        RECT 1335.480 1008.140 1335.740 1008.400 ;
        RECT 1341.000 1008.140 1341.260 1008.400 ;
        RECT 1368.140 1008.140 1368.400 1008.400 ;
        RECT 1383.320 1008.140 1383.580 1008.400 ;
        RECT 1497.400 1008.140 1497.660 1008.400 ;
        RECT 1568.240 1009.160 1568.500 1009.420 ;
        RECT 1602.740 1009.160 1603.000 1009.420 ;
        RECT 1607.340 1009.160 1607.600 1009.420 ;
        RECT 1613.780 1009.160 1614.040 1009.420 ;
        RECT 1891.160 1009.160 1891.420 1009.420 ;
        RECT 2046.180 1009.160 2046.440 1009.420 ;
        RECT 2085.280 1009.160 2085.540 1009.420 ;
        RECT 1532.360 1008.480 1532.620 1008.740 ;
        RECT 1536.500 1008.480 1536.760 1008.740 ;
        RECT 632.140 1007.800 632.400 1008.060 ;
        RECT 670.780 1007.800 671.040 1008.060 ;
        RECT 998.300 1007.800 998.560 1008.060 ;
        RECT 1084.320 1007.800 1084.580 1008.060 ;
        RECT 1151.020 1007.800 1151.280 1008.060 ;
        RECT 1191.040 1007.800 1191.300 1008.060 ;
        RECT 1191.500 1007.800 1191.760 1008.060 ;
        RECT 1238.880 1007.800 1239.140 1008.060 ;
        RECT 1250.380 1007.800 1250.640 1008.060 ;
        RECT 1254.980 1007.800 1255.240 1008.060 ;
        RECT 638.120 1007.460 638.380 1007.720 ;
        RECT 671.700 1007.460 671.960 1007.720 ;
        RECT 992.780 1007.460 993.040 1007.720 ;
        RECT 1014.400 1007.460 1014.660 1007.720 ;
        RECT 1079.720 1007.460 1079.980 1007.720 ;
        RECT 1115.140 1007.460 1115.400 1007.720 ;
        RECT 1145.500 1007.460 1145.760 1007.720 ;
        RECT 1169.420 1007.460 1169.680 1007.720 ;
        RECT 1197.480 1007.460 1197.740 1007.720 ;
        RECT 1232.440 1007.460 1232.700 1007.720 ;
        RECT 1254.520 1007.460 1254.780 1007.720 ;
        RECT 1292.700 1007.800 1292.960 1008.060 ;
        RECT 1293.620 1007.800 1293.880 1008.060 ;
        RECT 1319.380 1007.800 1319.640 1008.060 ;
        RECT 1335.020 1007.800 1335.280 1008.060 ;
        RECT 1338.700 1007.800 1338.960 1008.060 ;
        RECT 1396.200 1007.800 1396.460 1008.060 ;
        RECT 1400.340 1007.800 1400.600 1008.060 ;
        RECT 1413.220 1007.800 1413.480 1008.060 ;
        RECT 1438.520 1007.800 1438.780 1008.060 ;
        RECT 1496.480 1007.800 1496.740 1008.060 ;
        RECT 1559.960 1008.820 1560.220 1009.080 ;
        RECT 1834.580 1008.820 1834.840 1009.080 ;
        RECT 2100.920 1008.820 2101.180 1009.080 ;
        RECT 1542.020 1008.480 1542.280 1008.740 ;
        RECT 1578.360 1008.480 1578.620 1008.740 ;
        RECT 1824.460 1008.480 1824.720 1008.740 ;
        RECT 1907.720 1008.480 1907.980 1008.740 ;
        RECT 2050.780 1008.480 2051.040 1008.740 ;
        RECT 2055.840 1008.480 2056.100 1008.740 ;
        RECT 2065.960 1008.480 2066.220 1008.740 ;
        RECT 2080.220 1008.480 2080.480 1008.740 ;
        RECT 1873.220 1008.140 1873.480 1008.400 ;
        RECT 1900.360 1008.140 1900.620 1008.400 ;
        RECT 1574.680 1007.800 1574.940 1008.060 ;
        RECT 1901.280 1007.800 1901.540 1008.060 ;
        RECT 1257.280 1007.460 1257.540 1007.720 ;
        RECT 1294.080 1007.460 1294.340 1007.720 ;
        RECT 1324.440 1007.460 1324.700 1007.720 ;
        RECT 1332.720 1007.460 1332.980 1007.720 ;
        RECT 1333.180 1007.460 1333.440 1007.720 ;
        RECT 1336.400 1007.460 1336.660 1007.720 ;
        RECT 1411.380 1007.460 1411.640 1007.720 ;
        RECT 1424.720 1007.460 1424.980 1007.720 ;
        RECT 1431.160 1007.460 1431.420 1007.720 ;
        RECT 1434.840 1007.460 1435.100 1007.720 ;
        RECT 1511.660 1007.460 1511.920 1007.720 ;
        RECT 1514.880 1007.460 1515.140 1007.720 ;
        RECT 1620.220 1007.460 1620.480 1007.720 ;
        RECT 1635.400 1007.460 1635.660 1007.720 ;
        RECT 1776.620 1007.460 1776.880 1007.720 ;
        RECT 1779.840 1007.460 1780.100 1007.720 ;
        RECT 1798.240 1007.460 1798.500 1007.720 ;
        RECT 1800.540 1007.460 1800.800 1007.720 ;
        RECT 1802.840 1007.460 1803.100 1007.720 ;
        RECT 1806.980 1007.460 1807.240 1007.720 ;
        RECT 1811.580 1007.460 1811.840 1007.720 ;
        RECT 1813.880 1007.460 1814.140 1007.720 ;
        RECT 1075.580 1007.120 1075.840 1007.380 ;
        RECT 1077.420 1007.120 1077.680 1007.380 ;
        RECT 1076.040 1006.780 1076.300 1007.040 ;
        RECT 1076.960 1006.780 1077.220 1007.040 ;
        RECT 1332.260 1005.760 1332.520 1006.020 ;
        RECT 1338.240 1005.760 1338.500 1006.020 ;
        RECT 1208.060 1001.000 1208.320 1001.260 ;
        RECT 1216.570 1001.000 1216.830 1001.260 ;
        RECT 1332.260 1000.320 1332.520 1000.580 ;
        RECT 1333.640 1000.320 1333.900 1000.580 ;
        RECT 1193.800 999.300 1194.060 999.560 ;
        RECT 1197.480 999.300 1197.740 999.560 ;
        RECT 1215.420 999.300 1215.680 999.560 ;
        RECT 1219.100 999.300 1219.360 999.560 ;
      LAYER met2 ;
        RECT 1352.040 2917.890 1352.300 2918.210 ;
        RECT 1535.120 2917.890 1535.380 2918.210 ;
        RECT 979.440 2810.110 979.700 2810.430 ;
        RECT 445.840 2769.310 446.100 2769.630 ;
        RECT 810.620 2769.310 810.880 2769.630 ;
        RECT 445.900 2759.520 446.040 2769.310 ;
        RECT 532.320 2767.950 532.580 2768.270 ;
        RECT 700.220 2767.950 700.480 2768.270 ;
        RECT 518.520 2767.610 518.780 2767.930 ;
        RECT 489.080 2767.270 489.340 2767.590 ;
        RECT 489.140 2759.520 489.280 2767.270 ;
        RECT 518.580 2759.520 518.720 2767.610 ;
        RECT 532.380 2759.520 532.520 2767.950 ;
        RECT 445.730 2759.100 446.040 2759.520 ;
        RECT 488.970 2759.100 489.280 2759.520 ;
        RECT 518.410 2759.100 518.720 2759.520 ;
        RECT 532.210 2759.100 532.520 2759.520 ;
        RECT 445.730 2755.520 446.010 2759.100 ;
        RECT 488.970 2755.520 489.250 2759.100 ;
        RECT 518.410 2755.520 518.690 2759.100 ;
        RECT 532.210 2755.520 532.490 2759.100 ;
      LAYER met2 ;
        RECT 432.860 2755.240 445.450 2755.520 ;
        RECT 446.290 2755.240 460.170 2755.520 ;
        RECT 461.010 2755.240 474.890 2755.520 ;
        RECT 475.730 2755.240 488.690 2755.520 ;
        RECT 489.530 2755.240 503.410 2755.520 ;
        RECT 504.250 2755.240 518.130 2755.520 ;
        RECT 518.970 2755.240 531.930 2755.520 ;
        RECT 532.770 2755.240 546.650 2755.520 ;
        RECT 547.490 2755.240 561.370 2755.520 ;
        RECT 562.210 2755.240 575.170 2755.520 ;
      LAYER met2 ;
        RECT 420.530 2728.995 420.810 2729.365 ;
        RECT 420.070 2707.235 420.350 2707.605 ;
        RECT 419.620 1979.830 419.880 1980.150 ;
        RECT 419.680 1978.450 419.820 1979.830 ;
        RECT 420.140 1978.790 420.280 2707.235 ;
        RECT 420.600 1980.150 420.740 2728.995 ;
      LAYER met2 ;
        RECT 432.860 2604.280 575.720 2755.240 ;
      LAYER met2 ;
        RECT 586.590 2686.835 586.870 2687.205 ;
        RECT 586.660 2684.290 586.800 2686.835 ;
        RECT 586.600 2683.970 586.860 2684.290 ;
        RECT 586.590 2666.435 586.870 2666.805 ;
        RECT 586.660 2663.890 586.800 2666.435 ;
        RECT 586.600 2663.570 586.860 2663.890 ;
      LAYER met2 ;
        RECT 433.410 2604.000 446.370 2604.280 ;
        RECT 447.210 2604.000 461.090 2604.280 ;
        RECT 461.930 2604.000 475.810 2604.280 ;
        RECT 476.650 2604.000 489.610 2604.280 ;
        RECT 490.450 2604.000 504.330 2604.280 ;
        RECT 505.170 2604.000 519.050 2604.280 ;
        RECT 519.890 2604.000 532.850 2604.280 ;
        RECT 533.690 2604.000 547.570 2604.280 ;
        RECT 548.410 2604.000 562.290 2604.280 ;
        RECT 563.130 2604.000 575.720 2604.280 ;
      LAYER met2 ;
        RECT 504.610 2600.660 504.890 2604.000 ;
        RECT 533.130 2600.660 533.410 2604.000 ;
        RECT 504.610 2600.000 504.920 2600.660 ;
        RECT 533.130 2600.000 533.440 2600.660 ;
        RECT 504.780 2591.470 504.920 2600.000 ;
        RECT 533.300 2591.810 533.440 2600.000 ;
        RECT 533.240 2591.490 533.500 2591.810 ;
        RECT 504.720 2591.150 504.980 2591.470 ;
        RECT 579.240 1988.670 579.500 1988.990 ;
        RECT 632.140 1988.670 632.400 1988.990 ;
        RECT 530.020 1987.990 530.280 1988.310 ;
        RECT 528.450 1981.250 528.730 1981.750 ;
        RECT 530.080 1981.250 530.220 1987.990 ;
        RECT 528.450 1981.110 530.220 1981.250 ;
        RECT 578.130 1981.250 578.410 1981.750 ;
        RECT 579.300 1981.250 579.440 1988.670 ;
        RECT 578.130 1981.110 579.440 1981.250 ;
        RECT 420.540 1979.830 420.800 1980.150 ;
        RECT 420.080 1978.470 420.340 1978.790 ;
        RECT 419.620 1978.130 419.880 1978.450 ;
        RECT 528.450 1977.750 528.730 1981.110 ;
        RECT 578.130 1977.750 578.410 1981.110 ;
      LAYER met2 ;
        RECT 362.860 1977.470 377.290 1977.750 ;
        RECT 378.130 1977.470 402.130 1977.750 ;
        RECT 402.970 1977.470 427.890 1977.750 ;
        RECT 428.730 1977.470 452.730 1977.750 ;
        RECT 453.570 1977.470 477.570 1977.750 ;
        RECT 478.410 1977.470 502.410 1977.750 ;
        RECT 503.250 1977.470 528.170 1977.750 ;
        RECT 529.010 1977.470 553.010 1977.750 ;
        RECT 553.850 1977.470 577.850 1977.750 ;
        RECT 578.690 1977.470 602.690 1977.750 ;
        RECT 603.530 1977.470 627.530 1977.750 ;
        RECT 362.860 1704.280 628.080 1977.470 ;
        RECT 363.410 1704.000 387.410 1704.280 ;
        RECT 388.250 1704.000 412.250 1704.280 ;
        RECT 413.090 1704.000 437.090 1704.280 ;
        RECT 437.930 1704.000 461.930 1704.280 ;
        RECT 462.770 1704.000 487.690 1704.280 ;
        RECT 488.530 1704.000 512.530 1704.280 ;
        RECT 513.370 1704.000 537.370 1704.280 ;
        RECT 538.210 1704.000 562.210 1704.280 ;
        RECT 563.050 1704.000 587.970 1704.280 ;
        RECT 588.810 1704.000 612.810 1704.280 ;
        RECT 613.650 1704.000 628.080 1704.280 ;
      LAYER met2 ;
        RECT 462.210 1700.410 462.490 1704.000 ;
        RECT 512.810 1700.410 513.090 1704.000 ;
        RECT 462.210 1700.270 463.980 1700.410 ;
        RECT 462.210 1700.000 462.490 1700.270 ;
        RECT 463.840 1688.770 463.980 1700.270 ;
        RECT 512.810 1700.270 514.580 1700.410 ;
        RECT 512.810 1700.000 513.090 1700.270 ;
        RECT 514.440 1688.770 514.580 1700.270 ;
        RECT 463.780 1688.450 464.040 1688.770 ;
        RECT 468.840 1688.450 469.100 1688.770 ;
        RECT 514.380 1688.450 514.640 1688.770 ;
        RECT 517.140 1688.450 517.400 1688.770 ;
        RECT 468.900 1010.810 469.040 1688.450 ;
        RECT 517.200 1011.150 517.340 1688.450 ;
        RECT 632.200 1028.490 632.340 1988.670 ;
        RECT 638.120 1987.990 638.380 1988.310 ;
        RECT 632.140 1028.170 632.400 1028.490 ;
        RECT 632.140 1027.490 632.400 1027.810 ;
        RECT 517.140 1010.830 517.400 1011.150 ;
        RECT 468.840 1010.490 469.100 1010.810 ;
        RECT 632.200 1008.090 632.340 1027.490 ;
        RECT 632.140 1007.770 632.400 1008.090 ;
        RECT 638.180 1007.750 638.320 1987.990 ;
        RECT 700.280 1011.490 700.420 2767.950 ;
        RECT 755.420 2767.610 755.680 2767.930 ;
        RECT 734.720 2683.970 734.980 2684.290 ;
        RECT 700.220 1011.170 700.480 1011.490 ;
        RECT 712.640 1010.830 712.900 1011.150 ;
        RECT 673.540 1010.490 673.800 1010.810 ;
        RECT 670.780 1007.770 671.040 1008.090 ;
        RECT 638.120 1007.430 638.380 1007.750 ;
        RECT 670.840 1000.010 670.980 1007.770 ;
        RECT 671.700 1007.430 671.960 1007.750 ;
        RECT 671.760 1000.010 671.900 1007.430 ;
        RECT 673.600 1000.010 673.740 1010.490 ;
        RECT 712.700 1000.010 712.840 1010.830 ;
        RECT 734.780 1010.810 734.920 2683.970 ;
        RECT 755.480 1011.150 755.620 2767.610 ;
        RECT 789.920 2767.270 790.180 2767.590 ;
        RECT 769.220 2591.490 769.480 2591.810 ;
        RECT 769.280 1011.830 769.420 2591.490 ;
        RECT 789.980 1012.170 790.120 2767.270 ;
        RECT 803.720 2663.570 803.980 2663.890 ;
        RECT 796.820 2591.150 797.080 2591.470 ;
        RECT 796.880 1012.850 797.020 2591.150 ;
        RECT 796.820 1012.530 797.080 1012.850 ;
        RECT 803.780 1012.510 803.920 2663.570 ;
        RECT 810.680 1014.210 810.820 2769.310 ;
        RECT 978.520 2047.150 978.780 2047.470 ;
        RECT 978.060 2045.790 978.320 2046.110 ;
        RECT 977.600 2045.450 977.860 2045.770 ;
        RECT 843.280 1977.790 843.540 1978.110 ;
        RECT 810.620 1013.890 810.880 1014.210 ;
        RECT 803.720 1012.190 803.980 1012.510 ;
        RECT 789.920 1011.850 790.180 1012.170 ;
        RECT 769.220 1011.510 769.480 1011.830 ;
        RECT 841.900 1011.170 842.160 1011.490 ;
        RECT 755.420 1010.830 755.680 1011.150 ;
        RECT 734.720 1010.490 734.980 1010.810 ;
        RECT 841.960 1000.010 842.100 1011.170 ;
        RECT 843.340 1000.010 843.480 1977.790 ;
        RECT 897.560 1977.450 897.820 1977.770 ;
        RECT 845.580 1013.890 845.840 1014.210 ;
        RECT 845.640 1000.010 845.780 1013.890 ;
        RECT 884.680 1012.530 884.940 1012.850 ;
        RECT 884.740 1000.010 884.880 1012.530 ;
        RECT 890.200 1012.190 890.460 1012.510 ;
        RECT 890.260 1000.010 890.400 1012.190 ;
        RECT 893.420 1010.490 893.680 1010.810 ;
        RECT 893.480 1000.010 893.620 1010.490 ;
        RECT 897.620 1000.010 897.760 1977.450 ;
        RECT 977.660 1025.090 977.800 2045.450 ;
        RECT 977.600 1024.770 977.860 1025.090 ;
        RECT 978.120 1024.750 978.260 2045.790 ;
        RECT 978.580 1025.770 978.720 2047.150 ;
        RECT 978.980 2046.810 979.240 2047.130 ;
        RECT 978.520 1025.450 978.780 1025.770 ;
        RECT 979.040 1025.430 979.180 2046.810 ;
        RECT 979.500 1026.110 979.640 2810.110 ;
        RECT 985.420 2809.430 985.680 2809.750 ;
        RECT 1043.380 2809.430 1043.640 2809.750 ;
        RECT 1089.380 2809.430 1089.640 2809.750 ;
        RECT 984.960 2809.090 985.220 2809.410 ;
        RECT 984.500 2050.550 984.760 2050.870 ;
        RECT 984.040 2047.490 984.300 2047.810 ;
        RECT 983.580 2046.470 983.840 2046.790 ;
        RECT 983.120 2046.130 983.380 2046.450 ;
        RECT 983.180 1026.450 983.320 2046.130 ;
        RECT 983.640 1026.790 983.780 2046.470 ;
        RECT 983.580 1026.470 983.840 1026.790 ;
        RECT 983.120 1026.130 983.380 1026.450 ;
        RECT 979.440 1025.790 979.700 1026.110 ;
        RECT 978.980 1025.110 979.240 1025.430 ;
        RECT 978.060 1024.430 978.320 1024.750 ;
        RECT 910.900 1011.850 911.160 1012.170 ;
        RECT 906.300 1011.510 906.560 1011.830 ;
        RECT 901.700 1010.830 901.960 1011.150 ;
        RECT 901.760 1000.010 901.900 1010.830 ;
        RECT 906.360 1000.010 906.500 1011.510 ;
        RECT 910.960 1000.010 911.100 1011.850 ;
        RECT 984.100 1009.110 984.240 2047.490 ;
        RECT 984.560 1013.870 984.700 2050.550 ;
        RECT 984.500 1013.550 984.760 1013.870 ;
        RECT 985.020 1013.725 985.160 2809.090 ;
        RECT 985.480 1014.405 985.620 2809.430 ;
        RECT 1027.740 2809.090 1028.000 2809.410 ;
        RECT 986.340 2808.750 986.600 2809.070 ;
        RECT 985.880 2808.410 986.140 2808.730 ;
        RECT 985.410 1014.035 985.690 1014.405 ;
        RECT 984.950 1013.355 985.230 1013.725 ;
        RECT 985.940 1011.005 986.080 2808.410 ;
        RECT 986.400 1012.365 986.540 2808.750 ;
        RECT 1012.100 2808.410 1012.360 2808.730 ;
        RECT 1012.160 2800.000 1012.300 2808.410 ;
        RECT 1027.800 2800.000 1027.940 2809.090 ;
        RECT 1043.440 2800.000 1043.580 2809.430 ;
        RECT 1058.090 2808.555 1058.370 2808.925 ;
        RECT 1073.740 2808.750 1074.000 2809.070 ;
        RECT 1058.160 2800.000 1058.300 2808.555 ;
        RECT 1073.800 2800.000 1073.940 2808.750 ;
        RECT 1089.440 2800.000 1089.580 2809.430 ;
        RECT 1012.050 2796.000 1012.330 2800.000 ;
        RECT 1027.690 2796.000 1027.970 2800.000 ;
        RECT 1043.330 2796.000 1043.610 2800.000 ;
        RECT 1058.050 2796.000 1058.330 2800.000 ;
        RECT 1073.690 2796.000 1073.970 2800.000 ;
        RECT 1089.330 2796.000 1089.610 2800.000 ;
      LAYER met2 ;
        RECT 1002.860 2795.720 1011.770 2796.000 ;
        RECT 1012.610 2795.720 1027.410 2796.000 ;
        RECT 1028.250 2795.720 1043.050 2796.000 ;
        RECT 1043.890 2795.720 1057.770 2796.000 ;
        RECT 1058.610 2795.720 1073.410 2796.000 ;
        RECT 1074.250 2795.720 1089.050 2796.000 ;
        RECT 1089.890 2795.720 1095.120 2796.000 ;
      LAYER met2 ;
        RECT 993.230 2670.515 993.510 2670.885 ;
        RECT 992.770 2622.915 993.050 2623.285 ;
        RECT 991.400 2604.750 991.660 2605.070 ;
        RECT 990.940 2604.410 991.200 2604.730 ;
        RECT 990.480 2591.150 990.740 2591.470 ;
        RECT 990.010 1893.275 990.290 1893.645 ;
        RECT 989.550 1871.515 989.830 1871.885 ;
        RECT 989.090 1851.115 989.370 1851.485 ;
        RECT 988.630 1808.955 988.910 1809.325 ;
        RECT 987.710 1787.195 987.990 1787.565 ;
        RECT 987.250 1766.795 987.530 1767.165 ;
        RECT 986.790 1745.035 987.070 1745.405 ;
        RECT 986.860 1012.510 987.000 1745.035 ;
        RECT 987.320 1018.630 987.460 1766.795 ;
        RECT 987.260 1018.310 987.520 1018.630 ;
        RECT 987.780 1012.850 987.920 1787.195 ;
        RECT 988.170 1724.635 988.450 1725.005 ;
        RECT 988.240 1013.190 988.380 1724.635 ;
        RECT 988.700 1019.650 988.840 1808.955 ;
        RECT 988.640 1019.330 988.900 1019.650 ;
        RECT 989.160 1018.290 989.300 1851.115 ;
        RECT 989.100 1017.970 989.360 1018.290 ;
        RECT 988.180 1012.870 988.440 1013.190 ;
        RECT 987.720 1012.530 987.980 1012.850 ;
        RECT 986.330 1011.995 986.610 1012.365 ;
        RECT 986.800 1012.190 987.060 1012.510 ;
        RECT 985.870 1010.635 986.150 1011.005 ;
        RECT 989.620 1010.810 989.760 1871.515 ;
        RECT 990.080 1019.310 990.220 1893.275 ;
        RECT 990.540 1695.230 990.680 2591.150 ;
        RECT 990.480 1694.910 990.740 1695.230 ;
        RECT 991.000 1693.870 991.140 2604.410 ;
        RECT 991.460 1694.210 991.600 2604.750 ;
        RECT 992.310 1997.995 992.590 1998.365 ;
        RECT 991.850 1935.435 992.130 1935.805 ;
        RECT 991.400 1693.890 991.660 1694.210 ;
        RECT 990.940 1693.550 991.200 1693.870 ;
        RECT 990.020 1018.990 990.280 1019.310 ;
        RECT 991.920 1017.950 992.060 1935.435 ;
        RECT 992.380 1018.970 992.520 1997.995 ;
        RECT 992.320 1018.650 992.580 1018.970 ;
        RECT 991.860 1017.630 992.120 1017.950 ;
        RECT 989.560 1010.490 989.820 1010.810 ;
        RECT 984.040 1008.790 984.300 1009.110 ;
        RECT 992.840 1007.750 992.980 2622.915 ;
        RECT 993.300 1009.790 993.440 2670.515 ;
        RECT 993.690 2646.035 993.970 2646.405 ;
        RECT 993.240 1009.470 993.500 1009.790 ;
        RECT 993.760 1009.450 993.900 2646.035 ;
        RECT 996.920 2605.430 997.180 2605.750 ;
        RECT 994.150 2018.395 994.430 2018.765 ;
        RECT 994.220 1011.150 994.360 2018.395 ;
        RECT 994.610 1976.235 994.890 1976.605 ;
        RECT 994.680 1014.210 994.820 1976.235 ;
        RECT 995.070 1955.835 995.350 1956.205 ;
        RECT 995.140 1019.990 995.280 1955.835 ;
        RECT 995.530 1913.675 995.810 1914.045 ;
        RECT 995.080 1019.670 995.340 1019.990 ;
        RECT 994.620 1013.890 994.880 1014.210 ;
        RECT 994.160 1010.830 994.420 1011.150 ;
        RECT 995.600 1010.470 995.740 1913.675 ;
        RECT 995.990 1829.355 996.270 1829.725 ;
        RECT 996.060 1012.170 996.200 1829.355 ;
        RECT 996.460 1714.290 996.720 1714.610 ;
        RECT 996.000 1011.850 996.260 1012.170 ;
        RECT 995.540 1010.150 995.800 1010.470 ;
        RECT 993.700 1009.130 993.960 1009.450 ;
        RECT 996.520 1008.770 996.660 1714.290 ;
        RECT 996.980 1694.550 997.120 2605.430 ;
        RECT 997.380 2605.090 997.640 2605.410 ;
        RECT 997.440 1694.890 997.580 2605.090 ;
      LAYER met2 ;
        RECT 1002.860 2604.280 1095.120 2795.720 ;
      LAYER met2 ;
        RECT 1110.990 2780.675 1111.270 2781.045 ;
      LAYER met2 ;
        RECT 1003.410 2604.000 1017.290 2604.280 ;
        RECT 1018.130 2604.000 1032.930 2604.280 ;
        RECT 1033.770 2604.000 1048.570 2604.280 ;
        RECT 1049.410 2604.000 1064.210 2604.280 ;
        RECT 1065.050 2604.000 1079.850 2604.280 ;
        RECT 1080.690 2604.000 1094.570 2604.280 ;
      LAYER met2 ;
        RECT 1002.850 2600.730 1003.130 2604.000 ;
        RECT 1017.570 2600.730 1017.850 2604.000 ;
        RECT 1001.120 2600.590 1003.130 2600.730 ;
        RECT 998.760 2050.210 999.020 2050.530 ;
        RECT 997.840 2048.170 998.100 2048.490 ;
        RECT 997.380 1694.570 997.640 1694.890 ;
        RECT 996.920 1694.230 997.180 1694.550 ;
        RECT 997.380 1013.890 997.640 1014.210 ;
        RECT 997.440 1011.490 997.580 1013.890 ;
        RECT 997.380 1011.170 997.640 1011.490 ;
        RECT 996.460 1008.450 996.720 1008.770 ;
        RECT 997.900 1008.430 998.040 2048.170 ;
        RECT 998.300 2047.830 998.560 2048.150 ;
        RECT 997.840 1008.110 998.100 1008.430 ;
        RECT 998.360 1008.090 998.500 2047.830 ;
        RECT 998.820 1010.130 998.960 2050.210 ;
        RECT 999.680 2049.870 999.940 2050.190 ;
        RECT 999.220 2049.190 999.480 2049.510 ;
        RECT 999.280 1013.530 999.420 2049.190 ;
        RECT 999.220 1013.210 999.480 1013.530 ;
        RECT 999.740 1010.470 999.880 2049.870 ;
        RECT 1000.140 2049.530 1000.400 2049.850 ;
        RECT 1000.200 1014.210 1000.340 2049.530 ;
        RECT 1001.120 1714.610 1001.260 2600.590 ;
        RECT 1002.850 2600.000 1003.130 2600.590 ;
        RECT 1014.460 2600.590 1017.850 2600.730 ;
        RECT 1002.900 2050.550 1003.160 2050.870 ;
        RECT 1002.960 2044.110 1003.100 2050.550 ;
        RECT 1014.460 2048.490 1014.600 2600.590 ;
        RECT 1017.570 2600.000 1017.850 2600.590 ;
        RECT 1033.210 2600.000 1033.490 2604.000 ;
        RECT 1048.850 2600.000 1049.130 2604.000 ;
        RECT 1064.490 2600.730 1064.770 2604.000 ;
        RECT 1080.130 2600.730 1080.410 2604.000 ;
        RECT 1062.760 2600.590 1064.770 2600.730 ;
        RECT 1033.320 2587.730 1033.460 2600.000 ;
        RECT 1028.200 2587.410 1028.460 2587.730 ;
        RECT 1033.260 2587.410 1033.520 2587.730 ;
        RECT 1016.690 2051.715 1016.970 2052.085 ;
        RECT 1014.400 2048.170 1014.660 2048.490 ;
        RECT 1016.760 2044.110 1016.900 2051.715 ;
        RECT 1028.260 2048.150 1028.400 2587.410 ;
        RECT 1031.420 2051.910 1031.680 2052.230 ;
        RECT 1028.200 2047.830 1028.460 2048.150 ;
        RECT 1031.480 2044.110 1031.620 2051.910 ;
        RECT 1045.220 2049.190 1045.480 2049.510 ;
        RECT 1045.280 2044.110 1045.420 2049.190 ;
        RECT 1048.960 2047.810 1049.100 2600.000 ;
        RECT 1059.940 2052.250 1060.200 2052.570 ;
        RECT 1048.900 2047.490 1049.160 2047.810 ;
        RECT 1060.000 2044.110 1060.140 2052.250 ;
        RECT 1062.760 2047.470 1062.900 2600.590 ;
        RECT 1064.490 2600.000 1064.770 2600.590 ;
        RECT 1076.560 2600.590 1080.410 2600.730 ;
        RECT 1073.740 2049.530 1074.000 2049.850 ;
        RECT 1062.700 2047.150 1062.960 2047.470 ;
        RECT 1073.800 2044.110 1073.940 2049.530 ;
        RECT 1076.560 2047.130 1076.700 2600.590 ;
        RECT 1080.130 2600.000 1080.410 2600.590 ;
        RECT 1094.850 2600.000 1095.130 2604.000 ;
        RECT 1094.960 2591.470 1095.100 2600.000 ;
        RECT 1094.900 2591.150 1095.160 2591.470 ;
        RECT 1088.460 2050.210 1088.720 2050.530 ;
        RECT 1076.500 2046.810 1076.760 2047.130 ;
        RECT 1088.520 2044.110 1088.660 2050.210 ;
        RECT 1102.260 2049.870 1102.520 2050.190 ;
        RECT 1102.320 2044.110 1102.460 2049.870 ;
        RECT 1111.060 2046.110 1111.200 2780.675 ;
        RECT 1111.450 2760.275 1111.730 2760.645 ;
        RECT 1111.000 2045.790 1111.260 2046.110 ;
        RECT 1111.520 2045.770 1111.660 2760.275 ;
        RECT 1112.830 2734.435 1113.110 2734.805 ;
        RECT 1112.370 2712.675 1112.650 2713.045 ;
        RECT 1111.910 2691.595 1112.190 2691.965 ;
        RECT 1111.980 2605.750 1112.120 2691.595 ;
        RECT 1111.920 2605.430 1112.180 2605.750 ;
        RECT 1112.440 2604.730 1112.580 2712.675 ;
        RECT 1112.900 2605.410 1113.040 2734.435 ;
        RECT 1113.290 2666.435 1113.570 2666.805 ;
        RECT 1112.840 2605.090 1113.100 2605.410 ;
        RECT 1113.360 2605.070 1113.500 2666.435 ;
        RECT 1113.750 2644.675 1114.030 2645.045 ;
        RECT 1113.300 2604.750 1113.560 2605.070 ;
        RECT 1112.380 2604.410 1112.640 2604.730 ;
        RECT 1113.820 2046.790 1113.960 2644.675 ;
        RECT 1114.210 2622.235 1114.490 2622.605 ;
        RECT 1113.760 2046.470 1114.020 2046.790 ;
        RECT 1114.280 2046.450 1114.420 2622.235 ;
        RECT 1244.860 2053.950 1245.120 2054.270 ;
        RECT 1332.720 2053.950 1332.980 2054.270 ;
        RECT 1230.140 2053.610 1230.400 2053.930 ;
        RECT 1173.100 2053.270 1173.360 2053.590 ;
        RECT 1144.580 2052.930 1144.840 2053.250 ;
        RECT 1116.980 2052.590 1117.240 2052.910 ;
        RECT 1114.220 2046.130 1114.480 2046.450 ;
        RECT 1111.460 2045.450 1111.720 2045.770 ;
        RECT 1117.040 2044.110 1117.180 2052.590 ;
        RECT 1130.770 2050.355 1131.050 2050.725 ;
        RECT 1130.840 2044.110 1130.980 2050.355 ;
        RECT 1144.640 2044.110 1144.780 2052.930 ;
        RECT 1159.290 2051.035 1159.570 2051.405 ;
        RECT 1159.360 2044.110 1159.500 2051.035 ;
        RECT 1173.160 2044.110 1173.300 2053.270 ;
        RECT 1216.340 2051.570 1216.600 2051.890 ;
        RECT 1201.620 2051.230 1201.880 2051.550 ;
        RECT 1187.820 2050.890 1188.080 2051.210 ;
        RECT 1187.880 2044.110 1188.020 2050.890 ;
        RECT 1201.680 2044.110 1201.820 2051.230 ;
        RECT 1216.400 2044.110 1216.540 2051.570 ;
        RECT 1230.200 2044.110 1230.340 2053.610 ;
        RECT 1244.920 2044.110 1245.060 2053.950 ;
        RECT 1331.800 2051.910 1332.060 2052.230 ;
        RECT 1287.180 2050.550 1287.440 2050.870 ;
        RECT 1273.380 2050.210 1273.640 2050.530 ;
        RECT 1258.660 2049.870 1258.920 2050.190 ;
        RECT 1258.720 2044.110 1258.860 2049.870 ;
        RECT 1273.440 2044.110 1273.580 2050.210 ;
        RECT 1287.240 2044.110 1287.380 2050.550 ;
        RECT 1301.900 2049.530 1302.160 2049.850 ;
        RECT 1315.690 2049.675 1315.970 2050.045 ;
        RECT 1301.960 2044.110 1302.100 2049.530 ;
        RECT 1315.760 2044.110 1315.900 2049.675 ;
        RECT 1329.500 2049.190 1329.760 2049.510 ;
        RECT 1329.560 2044.110 1329.700 2049.190 ;
        RECT 1002.850 2040.110 1003.130 2044.110 ;
        RECT 1016.650 2040.110 1016.930 2044.110 ;
        RECT 1031.370 2040.110 1031.650 2044.110 ;
        RECT 1045.170 2040.110 1045.450 2044.110 ;
        RECT 1059.890 2040.110 1060.170 2044.110 ;
        RECT 1073.690 2040.110 1073.970 2044.110 ;
        RECT 1088.410 2040.110 1088.690 2044.110 ;
        RECT 1102.210 2040.110 1102.490 2044.110 ;
        RECT 1116.930 2040.110 1117.210 2044.110 ;
        RECT 1130.730 2040.110 1131.010 2044.110 ;
        RECT 1144.530 2040.110 1144.810 2044.110 ;
        RECT 1159.250 2040.110 1159.530 2044.110 ;
        RECT 1173.050 2040.110 1173.330 2044.110 ;
        RECT 1187.770 2040.110 1188.050 2044.110 ;
        RECT 1201.570 2040.110 1201.850 2044.110 ;
        RECT 1216.290 2040.110 1216.570 2044.110 ;
        RECT 1230.090 2040.110 1230.370 2044.110 ;
        RECT 1244.810 2040.110 1245.090 2044.110 ;
        RECT 1258.610 2040.110 1258.890 2044.110 ;
        RECT 1273.330 2040.110 1273.610 2044.110 ;
        RECT 1287.130 2040.110 1287.410 2044.110 ;
        RECT 1301.850 2040.110 1302.130 2044.110 ;
        RECT 1315.650 2040.110 1315.930 2044.110 ;
        RECT 1329.450 2040.110 1329.730 2044.110 ;
      LAYER met2 ;
        RECT 1003.410 2039.830 1016.370 2040.110 ;
        RECT 1017.210 2039.830 1031.090 2040.110 ;
        RECT 1031.930 2039.830 1044.890 2040.110 ;
        RECT 1045.730 2039.830 1059.610 2040.110 ;
        RECT 1060.450 2039.830 1073.410 2040.110 ;
        RECT 1074.250 2039.830 1088.130 2040.110 ;
        RECT 1088.970 2039.830 1101.930 2040.110 ;
        RECT 1102.770 2039.830 1116.650 2040.110 ;
        RECT 1117.490 2039.830 1130.450 2040.110 ;
        RECT 1131.290 2039.830 1144.250 2040.110 ;
        RECT 1145.090 2039.830 1158.970 2040.110 ;
        RECT 1159.810 2039.830 1172.770 2040.110 ;
        RECT 1173.610 2039.830 1187.490 2040.110 ;
        RECT 1188.330 2039.830 1201.290 2040.110 ;
        RECT 1202.130 2039.830 1216.010 2040.110 ;
        RECT 1216.850 2039.830 1229.810 2040.110 ;
        RECT 1230.650 2039.830 1244.530 2040.110 ;
        RECT 1245.370 2039.830 1258.330 2040.110 ;
        RECT 1259.170 2039.830 1273.050 2040.110 ;
        RECT 1273.890 2039.830 1286.850 2040.110 ;
        RECT 1287.690 2039.830 1301.570 2040.110 ;
        RECT 1302.410 2039.830 1315.370 2040.110 ;
        RECT 1316.210 2039.830 1329.170 2040.110 ;
      LAYER met2 ;
        RECT 1001.060 1714.290 1001.320 1714.610 ;
      LAYER met2 ;
        RECT 1002.860 1704.280 1329.720 2039.830 ;
        RECT 1003.410 1704.000 1016.370 1704.280 ;
        RECT 1017.210 1704.000 1030.170 1704.280 ;
        RECT 1031.010 1704.000 1044.890 1704.280 ;
        RECT 1045.730 1704.000 1058.690 1704.280 ;
        RECT 1059.530 1704.000 1073.410 1704.280 ;
        RECT 1074.250 1704.000 1087.210 1704.280 ;
        RECT 1088.050 1704.000 1101.930 1704.280 ;
        RECT 1102.770 1704.000 1115.730 1704.280 ;
        RECT 1116.570 1704.000 1130.450 1704.280 ;
        RECT 1131.290 1704.000 1144.250 1704.280 ;
        RECT 1145.090 1704.000 1158.970 1704.280 ;
        RECT 1159.810 1704.000 1172.770 1704.280 ;
        RECT 1173.610 1704.000 1187.490 1704.280 ;
        RECT 1188.330 1704.000 1201.290 1704.280 ;
        RECT 1202.130 1704.000 1215.090 1704.280 ;
        RECT 1215.930 1704.000 1229.810 1704.280 ;
        RECT 1230.650 1704.000 1243.610 1704.280 ;
        RECT 1244.450 1704.000 1258.330 1704.280 ;
        RECT 1259.170 1704.000 1272.130 1704.280 ;
        RECT 1272.970 1704.000 1286.850 1704.280 ;
        RECT 1287.690 1704.000 1300.650 1704.280 ;
        RECT 1301.490 1704.000 1315.370 1704.280 ;
        RECT 1316.210 1704.000 1329.170 1704.280 ;
      LAYER met2 ;
        RECT 1002.850 1700.000 1003.130 1704.000 ;
        RECT 1016.650 1700.000 1016.930 1704.000 ;
        RECT 1030.450 1700.000 1030.730 1704.000 ;
        RECT 1045.170 1700.000 1045.450 1704.000 ;
        RECT 1058.970 1700.410 1059.250 1704.000 ;
        RECT 1058.970 1700.270 1062.440 1700.410 ;
        RECT 1058.970 1700.000 1059.250 1700.270 ;
        RECT 1002.960 1689.110 1003.100 1700.000 ;
        RECT 1016.760 1689.450 1016.900 1700.000 ;
        RECT 1016.700 1689.130 1016.960 1689.450 ;
        RECT 1002.900 1688.790 1003.160 1689.110 ;
        RECT 1030.560 1688.430 1030.700 1700.000 ;
        RECT 1045.280 1689.790 1045.420 1700.000 ;
        RECT 1048.900 1694.910 1049.160 1695.230 ;
        RECT 1045.220 1689.470 1045.480 1689.790 ;
        RECT 1030.500 1688.110 1030.760 1688.430 ;
        RECT 1000.140 1013.890 1000.400 1014.210 ;
        RECT 1000.140 1011.510 1000.400 1011.830 ;
        RECT 999.220 1010.150 999.480 1010.470 ;
        RECT 999.680 1010.150 999.940 1010.470 ;
        RECT 998.760 1009.810 999.020 1010.130 ;
        RECT 999.280 1009.530 999.420 1010.150 ;
        RECT 1000.200 1009.530 1000.340 1011.510 ;
        RECT 999.280 1009.390 1000.340 1009.530 ;
        RECT 998.300 1007.770 998.560 1008.090 ;
        RECT 992.780 1007.430 993.040 1007.750 ;
        RECT 1014.400 1007.430 1014.660 1007.750 ;
        RECT 1014.460 1000.010 1014.600 1007.430 ;
        RECT 1048.960 1000.690 1049.100 1694.910 ;
        RECT 1062.300 1051.950 1062.440 1700.270 ;
        RECT 1073.690 1700.000 1073.970 1704.000 ;
        RECT 1087.490 1700.000 1087.770 1704.000 ;
        RECT 1102.210 1700.000 1102.490 1704.000 ;
        RECT 1116.010 1700.000 1116.290 1704.000 ;
        RECT 1130.730 1700.000 1131.010 1704.000 ;
        RECT 1144.530 1700.000 1144.810 1704.000 ;
        RECT 1159.250 1700.000 1159.530 1704.000 ;
        RECT 1173.050 1700.000 1173.330 1704.000 ;
        RECT 1187.770 1700.000 1188.050 1704.000 ;
        RECT 1201.570 1700.410 1201.850 1704.000 ;
        RECT 1200.760 1700.270 1201.850 1700.410 ;
        RECT 1069.600 1694.570 1069.860 1694.890 ;
        RECT 1062.240 1051.630 1062.500 1051.950 ;
        RECT 1058.560 1009.130 1058.820 1009.450 ;
        RECT 1062.690 1009.275 1062.970 1009.645 ;
        RECT 1069.660 1009.450 1069.800 1694.570 ;
        RECT 1073.800 1688.770 1073.940 1700.000 ;
        RECT 1076.500 1694.230 1076.760 1694.550 ;
        RECT 1073.740 1688.450 1074.000 1688.770 ;
        RECT 1075.580 1011.510 1075.840 1011.830 ;
        RECT 1055.790 1007.915 1056.070 1008.285 ;
        RECT 1048.960 1000.550 1050.480 1000.690 ;
        RECT 670.840 1000.000 671.140 1000.010 ;
        RECT 671.760 1000.000 672.980 1000.010 ;
        RECT 673.600 1000.000 675.280 1000.010 ;
        RECT 712.700 1000.000 714.380 1000.010 ;
        RECT 841.960 1000.000 842.720 1000.010 ;
        RECT 843.340 1000.000 845.020 1000.010 ;
        RECT 845.640 1000.000 846.860 1000.010 ;
        RECT 884.740 1000.000 885.960 1000.010 ;
        RECT 890.260 1000.000 890.560 1000.010 ;
        RECT 893.480 1000.000 894.700 1000.010 ;
        RECT 897.620 1000.000 899.300 1000.010 ;
        RECT 901.760 1000.000 903.440 1000.010 ;
        RECT 906.360 1000.000 908.040 1000.010 ;
        RECT 910.960 1000.000 912.180 1000.010 ;
        RECT 1014.300 1000.000 1014.600 1000.010 ;
        RECT 1050.340 1000.010 1050.480 1000.550 ;
        RECT 1055.860 1000.010 1056.000 1007.915 ;
        RECT 1050.340 1000.000 1051.560 1000.010 ;
        RECT 1055.700 1000.000 1056.000 1000.010 ;
        RECT 1058.620 1000.010 1058.760 1009.130 ;
        RECT 1062.760 1000.010 1062.900 1009.275 ;
        RECT 1069.600 1009.130 1069.860 1009.450 ;
        RECT 1071.900 1009.130 1072.160 1009.450 ;
        RECT 1067.290 1008.595 1067.570 1008.965 ;
        RECT 1067.360 1000.010 1067.500 1008.595 ;
        RECT 1071.960 1000.010 1072.100 1009.130 ;
        RECT 1075.640 1007.410 1075.780 1011.510 ;
        RECT 1076.040 1011.170 1076.300 1011.490 ;
        RECT 1075.580 1007.090 1075.840 1007.410 ;
        RECT 1076.100 1007.070 1076.240 1011.170 ;
        RECT 1076.040 1006.750 1076.300 1007.070 ;
        RECT 1076.560 1000.010 1076.700 1694.230 ;
        RECT 1087.600 1689.450 1087.740 1700.000 ;
        RECT 1102.320 1690.130 1102.460 1700.000 ;
        RECT 1104.100 1693.890 1104.360 1694.210 ;
        RECT 1102.260 1689.810 1102.520 1690.130 ;
        RECT 1100.420 1689.470 1100.680 1689.790 ;
        RECT 1079.720 1689.130 1079.980 1689.450 ;
        RECT 1087.540 1689.130 1087.800 1689.450 ;
        RECT 1079.780 1011.830 1079.920 1689.130 ;
        RECT 1098.580 1051.630 1098.840 1051.950 ;
        RECT 1079.720 1011.510 1079.980 1011.830 ;
        RECT 1081.100 1011.510 1081.360 1011.830 ;
        RECT 1076.960 1011.170 1077.220 1011.490 ;
        RECT 1077.020 1007.070 1077.160 1011.170 ;
        RECT 1081.160 1009.790 1081.300 1011.510 ;
        RECT 1090.290 1009.955 1090.570 1010.325 ;
        RECT 1080.180 1009.470 1080.440 1009.790 ;
        RECT 1081.100 1009.470 1081.360 1009.790 ;
        RECT 1077.420 1009.130 1077.680 1009.450 ;
        RECT 1077.480 1007.410 1077.620 1009.130 ;
        RECT 1079.720 1008.790 1079.980 1009.110 ;
        RECT 1079.780 1007.750 1079.920 1008.790 ;
        RECT 1079.720 1007.430 1079.980 1007.750 ;
        RECT 1077.420 1007.090 1077.680 1007.410 ;
        RECT 1076.960 1006.750 1077.220 1007.070 ;
        RECT 1080.240 1000.010 1080.380 1009.470 ;
        RECT 1084.320 1007.770 1084.580 1008.090 ;
        RECT 1084.380 1000.010 1084.520 1007.770 ;
        RECT 1090.360 1000.010 1090.500 1009.955 ;
        RECT 1098.640 1009.110 1098.780 1051.630 ;
        RECT 1100.480 1018.370 1100.620 1689.470 ;
        RECT 1100.480 1018.230 1101.080 1018.370 ;
        RECT 1098.580 1008.790 1098.840 1009.110 ;
        RECT 1100.940 1008.770 1101.080 1018.230 ;
        RECT 1101.790 1014.035 1102.070 1014.405 ;
        RECT 1097.660 1008.450 1097.920 1008.770 ;
        RECT 1100.880 1008.450 1101.140 1008.770 ;
        RECT 1093.060 1008.110 1093.320 1008.430 ;
        RECT 1093.120 1000.010 1093.260 1008.110 ;
        RECT 1097.720 1000.010 1097.860 1008.450 ;
        RECT 1101.860 1000.010 1102.000 1014.035 ;
        RECT 1104.160 1011.830 1104.300 1693.890 ;
        RECT 1111.000 1693.550 1111.260 1693.870 ;
        RECT 1104.100 1011.510 1104.360 1011.830 ;
        RECT 1106.400 1011.510 1106.660 1011.830 ;
        RECT 1106.860 1011.510 1107.120 1011.830 ;
        RECT 1106.460 1000.010 1106.600 1011.510 ;
        RECT 1106.920 1009.450 1107.060 1011.510 ;
        RECT 1106.860 1009.130 1107.120 1009.450 ;
        RECT 1111.060 1000.010 1111.200 1693.550 ;
        RECT 1116.120 1684.350 1116.260 1700.000 ;
        RECT 1130.840 1689.790 1130.980 1700.000 ;
        RECT 1130.780 1689.470 1131.040 1689.790 ;
        RECT 1144.640 1686.390 1144.780 1700.000 ;
        RECT 1159.360 1686.730 1159.500 1700.000 ;
        RECT 1173.160 1689.110 1173.300 1700.000 ;
        RECT 1185.970 1693.355 1186.250 1693.725 ;
        RECT 1186.440 1693.550 1186.700 1693.870 ;
        RECT 1167.580 1688.790 1167.840 1689.110 ;
        RECT 1173.100 1688.790 1173.360 1689.110 ;
        RECT 1159.300 1686.410 1159.560 1686.730 ;
        RECT 1144.580 1686.070 1144.840 1686.390 ;
        RECT 1162.520 1686.070 1162.780 1686.390 ;
        RECT 1116.060 1684.030 1116.320 1684.350 ;
        RECT 1148.720 1684.030 1148.980 1684.350 ;
        RECT 1134.460 1026.470 1134.720 1026.790 ;
        RECT 1119.270 1013.355 1119.550 1013.725 ;
        RECT 1111.460 1008.965 1111.720 1009.110 ;
        RECT 1111.450 1008.595 1111.730 1008.965 ;
        RECT 1115.140 1007.430 1115.400 1007.750 ;
        RECT 1115.200 1000.010 1115.340 1007.430 ;
        RECT 1119.340 1000.010 1119.480 1013.355 ;
        RECT 1125.710 1012.675 1125.990 1013.045 ;
        RECT 1125.780 1000.010 1125.920 1012.675 ;
        RECT 1131.690 1011.995 1131.970 1012.365 ;
        RECT 1131.760 1000.010 1131.900 1011.995 ;
        RECT 1058.620 1000.000 1059.840 1000.010 ;
        RECT 1062.760 1000.000 1064.440 1000.010 ;
        RECT 1067.360 1000.000 1068.580 1000.010 ;
        RECT 1071.960 1000.000 1073.180 1000.010 ;
        RECT 1076.560 1000.000 1077.320 1000.010 ;
        RECT 1080.240 1000.000 1081.920 1000.010 ;
        RECT 1084.380 1000.000 1086.060 1000.010 ;
        RECT 1090.360 1000.000 1090.660 1000.010 ;
        RECT 1093.120 1000.000 1094.800 1000.010 ;
        RECT 1097.720 1000.000 1099.400 1000.010 ;
        RECT 1101.860 1000.000 1103.540 1000.010 ;
        RECT 1106.460 1000.000 1107.680 1000.010 ;
        RECT 1111.060 1000.000 1112.280 1000.010 ;
        RECT 1115.200 1000.000 1116.420 1000.010 ;
        RECT 1119.340 1000.000 1121.020 1000.010 ;
        RECT 1125.780 1000.000 1127.460 1000.010 ;
        RECT 1131.600 1000.000 1131.900 1000.010 ;
        RECT 1134.520 1000.010 1134.660 1026.470 ;
        RECT 1139.520 1026.130 1139.780 1026.450 ;
        RECT 1139.580 1000.010 1139.720 1026.130 ;
        RECT 1143.200 1025.790 1143.460 1026.110 ;
        RECT 1143.260 1000.010 1143.400 1025.790 ;
        RECT 1147.800 1025.450 1148.060 1025.770 ;
        RECT 1145.500 1011.510 1145.760 1011.830 ;
        RECT 1145.560 1007.750 1145.700 1011.510 ;
        RECT 1145.960 1011.170 1146.220 1011.490 ;
        RECT 1146.020 1009.110 1146.160 1011.170 ;
        RECT 1146.420 1010.150 1146.680 1010.470 ;
        RECT 1146.480 1009.645 1146.620 1010.150 ;
        RECT 1146.410 1009.275 1146.690 1009.645 ;
        RECT 1145.960 1008.790 1146.220 1009.110 ;
        RECT 1145.500 1007.430 1145.760 1007.750 ;
        RECT 1147.860 1000.010 1148.000 1025.450 ;
        RECT 1148.780 1008.430 1148.920 1684.030 ;
        RECT 1152.400 1025.110 1152.660 1025.430 ;
        RECT 1151.020 1009.810 1151.280 1010.130 ;
        RECT 1148.720 1008.110 1148.980 1008.430 ;
        RECT 1151.080 1008.090 1151.220 1009.810 ;
        RECT 1151.020 1007.770 1151.280 1008.090 ;
        RECT 1152.460 1000.010 1152.600 1025.110 ;
        RECT 1156.080 1024.770 1156.340 1025.090 ;
        RECT 1156.140 1000.010 1156.280 1024.770 ;
        RECT 1158.370 1011.995 1158.650 1012.365 ;
        RECT 1158.440 1008.965 1158.580 1011.995 ;
        RECT 1160.670 1011.315 1160.950 1011.685 ;
        RECT 1160.210 1009.955 1160.490 1010.325 ;
        RECT 1160.220 1009.810 1160.480 1009.955 ;
        RECT 1158.370 1008.595 1158.650 1008.965 ;
        RECT 1159.290 1008.595 1159.570 1008.965 ;
        RECT 1159.760 1008.790 1160.020 1009.110 ;
        RECT 1159.300 1008.450 1159.560 1008.595 ;
        RECT 1159.820 1008.285 1159.960 1008.790 ;
        RECT 1159.750 1007.915 1160.030 1008.285 ;
        RECT 1160.740 1000.010 1160.880 1011.315 ;
        RECT 1162.580 1009.110 1162.720 1686.070 ;
        RECT 1167.640 1686.050 1167.780 1688.790 ;
        RECT 1167.580 1685.730 1167.840 1686.050 ;
        RECT 1166.200 1024.430 1166.460 1024.750 ;
        RECT 1161.130 1008.595 1161.410 1008.965 ;
        RECT 1162.520 1008.790 1162.780 1009.110 ;
        RECT 1161.140 1008.450 1161.400 1008.595 ;
        RECT 1166.260 1000.010 1166.400 1024.430 ;
        RECT 1169.420 1011.510 1169.680 1011.830 ;
        RECT 1166.660 1011.170 1166.920 1011.490 ;
        RECT 1166.720 1008.285 1166.860 1011.170 ;
        RECT 1167.110 1010.635 1167.390 1011.005 ;
        RECT 1166.650 1007.915 1166.930 1008.285 ;
        RECT 1167.180 1000.010 1167.320 1010.635 ;
        RECT 1169.480 1007.750 1169.620 1011.510 ;
        RECT 1183.220 1009.810 1183.480 1010.130 ;
        RECT 1176.320 1009.645 1176.580 1009.790 ;
        RECT 1176.310 1009.275 1176.590 1009.645 ;
        RECT 1169.420 1007.430 1169.680 1007.750 ;
        RECT 1183.280 1000.010 1183.420 1009.810 ;
        RECT 1183.680 1008.790 1183.940 1009.110 ;
        RECT 1134.520 1000.000 1136.200 1000.010 ;
        RECT 1139.580 1000.000 1140.340 1000.010 ;
        RECT 1143.260 1000.000 1144.940 1000.010 ;
        RECT 1147.860 1000.000 1149.080 1000.010 ;
        RECT 1152.460 1000.000 1153.680 1000.010 ;
        RECT 1156.140 1000.000 1157.820 1000.010 ;
        RECT 1160.740 1000.000 1162.420 1000.010 ;
        RECT 1166.260 1000.000 1166.560 1000.010 ;
        RECT 1167.180 1000.000 1168.860 1000.010 ;
        RECT 1181.740 1000.000 1183.420 1000.010 ;
        RECT 670.840 999.870 671.290 1000.000 ;
        RECT 671.760 999.870 673.130 1000.000 ;
        RECT 673.600 999.870 675.430 1000.000 ;
        RECT 671.010 996.000 671.290 999.870 ;
      LAYER met2 ;
        RECT 671.570 995.720 672.570 998.810 ;
      LAYER met2 ;
        RECT 672.850 996.000 673.130 999.870 ;
      LAYER met2 ;
        RECT 673.410 995.720 674.870 998.810 ;
      LAYER met2 ;
        RECT 675.150 996.000 675.430 999.870 ;
      LAYER met2 ;
        RECT 675.710 995.720 677.170 998.810 ;
      LAYER met2 ;
        RECT 677.450 996.000 677.730 1000.000 ;
      LAYER met2 ;
        RECT 678.010 995.720 679.010 998.810 ;
      LAYER met2 ;
        RECT 679.290 996.000 679.570 1000.000 ;
      LAYER met2 ;
        RECT 679.850 995.720 681.310 998.810 ;
      LAYER met2 ;
        RECT 681.590 996.000 681.870 1000.000 ;
      LAYER met2 ;
        RECT 682.150 995.720 683.610 998.810 ;
      LAYER met2 ;
        RECT 683.890 996.000 684.170 1000.000 ;
      LAYER met2 ;
        RECT 684.450 995.720 685.910 998.810 ;
      LAYER met2 ;
        RECT 686.190 996.000 686.470 1000.000 ;
      LAYER met2 ;
        RECT 686.750 995.720 687.750 998.810 ;
      LAYER met2 ;
        RECT 688.030 996.000 688.310 1000.000 ;
      LAYER met2 ;
        RECT 688.590 995.720 690.050 998.810 ;
      LAYER met2 ;
        RECT 690.330 996.000 690.610 1000.000 ;
      LAYER met2 ;
        RECT 690.890 995.720 692.350 998.810 ;
      LAYER met2 ;
        RECT 692.630 996.000 692.910 1000.000 ;
      LAYER met2 ;
        RECT 693.190 995.720 694.190 998.810 ;
      LAYER met2 ;
        RECT 694.470 996.000 694.750 1000.000 ;
      LAYER met2 ;
        RECT 695.030 995.720 696.490 998.810 ;
      LAYER met2 ;
        RECT 696.770 996.000 697.050 1000.000 ;
      LAYER met2 ;
        RECT 697.330 995.720 698.790 998.810 ;
      LAYER met2 ;
        RECT 699.070 996.000 699.350 1000.000 ;
      LAYER met2 ;
        RECT 699.630 995.720 701.090 998.810 ;
      LAYER met2 ;
        RECT 701.370 996.000 701.650 1000.000 ;
      LAYER met2 ;
        RECT 701.930 995.720 702.930 998.810 ;
      LAYER met2 ;
        RECT 703.210 996.000 703.490 1000.000 ;
      LAYER met2 ;
        RECT 703.770 995.720 705.230 998.810 ;
      LAYER met2 ;
        RECT 705.510 996.000 705.790 1000.000 ;
      LAYER met2 ;
        RECT 706.070 995.720 707.530 998.810 ;
      LAYER met2 ;
        RECT 707.810 996.000 708.090 1000.000 ;
      LAYER met2 ;
        RECT 708.370 995.720 709.830 998.810 ;
      LAYER met2 ;
        RECT 710.110 996.000 710.390 1000.000 ;
      LAYER met2 ;
        RECT 710.670 995.720 711.670 998.810 ;
      LAYER met2 ;
        RECT 711.950 996.000 712.230 1000.000 ;
        RECT 712.700 999.870 714.530 1000.000 ;
      LAYER met2 ;
        RECT 712.510 995.720 713.970 998.810 ;
      LAYER met2 ;
        RECT 714.250 996.000 714.530 999.870 ;
      LAYER met2 ;
        RECT 714.810 995.720 716.270 998.810 ;
      LAYER met2 ;
        RECT 716.550 996.000 716.830 1000.000 ;
      LAYER met2 ;
        RECT 717.110 995.720 718.110 998.810 ;
      LAYER met2 ;
        RECT 718.390 996.000 718.670 1000.000 ;
      LAYER met2 ;
        RECT 718.950 995.720 720.410 998.810 ;
      LAYER met2 ;
        RECT 720.690 996.000 720.970 1000.000 ;
      LAYER met2 ;
        RECT 721.250 995.720 722.710 998.810 ;
      LAYER met2 ;
        RECT 722.990 996.000 723.270 1000.000 ;
      LAYER met2 ;
        RECT 723.550 995.720 725.010 998.810 ;
      LAYER met2 ;
        RECT 725.290 996.000 725.570 1000.000 ;
      LAYER met2 ;
        RECT 725.850 995.720 726.850 998.810 ;
      LAYER met2 ;
        RECT 727.130 996.000 727.410 1000.000 ;
      LAYER met2 ;
        RECT 727.690 995.720 729.150 998.810 ;
      LAYER met2 ;
        RECT 729.430 996.000 729.710 1000.000 ;
      LAYER met2 ;
        RECT 729.990 995.720 731.450 998.810 ;
      LAYER met2 ;
        RECT 731.730 996.000 732.010 1000.000 ;
      LAYER met2 ;
        RECT 732.290 995.720 733.750 998.810 ;
      LAYER met2 ;
        RECT 734.030 996.000 734.310 1000.000 ;
      LAYER met2 ;
        RECT 734.590 995.720 735.590 998.810 ;
      LAYER met2 ;
        RECT 735.870 996.000 736.150 1000.000 ;
      LAYER met2 ;
        RECT 736.430 995.720 737.890 998.810 ;
      LAYER met2 ;
        RECT 738.170 996.000 738.450 1000.000 ;
      LAYER met2 ;
        RECT 738.730 995.720 740.190 998.810 ;
      LAYER met2 ;
        RECT 740.470 996.000 740.750 1000.000 ;
      LAYER met2 ;
        RECT 741.030 995.720 742.030 998.810 ;
      LAYER met2 ;
        RECT 742.310 996.000 742.590 1000.000 ;
      LAYER met2 ;
        RECT 742.870 995.720 744.330 998.810 ;
      LAYER met2 ;
        RECT 744.610 996.000 744.890 1000.000 ;
      LAYER met2 ;
        RECT 745.170 995.720 746.630 998.810 ;
      LAYER met2 ;
        RECT 746.910 996.000 747.190 1000.000 ;
      LAYER met2 ;
        RECT 747.470 995.720 748.930 998.810 ;
      LAYER met2 ;
        RECT 749.210 996.000 749.490 1000.000 ;
      LAYER met2 ;
        RECT 749.770 995.720 750.770 998.810 ;
      LAYER met2 ;
        RECT 751.050 996.000 751.330 1000.000 ;
      LAYER met2 ;
        RECT 751.610 995.720 753.070 998.810 ;
      LAYER met2 ;
        RECT 753.350 996.000 753.630 1000.000 ;
      LAYER met2 ;
        RECT 753.910 995.720 755.370 998.810 ;
      LAYER met2 ;
        RECT 755.650 996.000 755.930 1000.000 ;
      LAYER met2 ;
        RECT 756.210 995.720 757.670 998.810 ;
      LAYER met2 ;
        RECT 757.950 996.000 758.230 1000.000 ;
      LAYER met2 ;
        RECT 758.510 995.720 759.510 998.810 ;
      LAYER met2 ;
        RECT 759.790 996.000 760.070 1000.000 ;
      LAYER met2 ;
        RECT 760.350 995.720 761.810 998.810 ;
      LAYER met2 ;
        RECT 762.090 996.000 762.370 1000.000 ;
      LAYER met2 ;
        RECT 762.650 995.720 764.110 998.810 ;
      LAYER met2 ;
        RECT 764.390 996.000 764.670 1000.000 ;
      LAYER met2 ;
        RECT 764.950 995.720 765.950 998.810 ;
      LAYER met2 ;
        RECT 766.230 996.000 766.510 1000.000 ;
      LAYER met2 ;
        RECT 766.790 995.720 768.250 998.810 ;
      LAYER met2 ;
        RECT 768.530 996.000 768.810 1000.000 ;
      LAYER met2 ;
        RECT 769.090 995.720 770.550 998.810 ;
      LAYER met2 ;
        RECT 770.830 996.000 771.110 1000.000 ;
      LAYER met2 ;
        RECT 771.390 995.720 772.850 998.810 ;
      LAYER met2 ;
        RECT 773.130 996.000 773.410 1000.000 ;
      LAYER met2 ;
        RECT 773.690 995.720 774.690 998.810 ;
      LAYER met2 ;
        RECT 774.970 996.000 775.250 1000.000 ;
      LAYER met2 ;
        RECT 775.530 995.720 776.990 998.810 ;
      LAYER met2 ;
        RECT 777.270 996.000 777.550 1000.000 ;
      LAYER met2 ;
        RECT 777.830 995.720 779.290 998.810 ;
      LAYER met2 ;
        RECT 779.570 996.000 779.850 1000.000 ;
      LAYER met2 ;
        RECT 780.130 995.720 781.590 998.810 ;
      LAYER met2 ;
        RECT 781.870 996.000 782.150 1000.000 ;
      LAYER met2 ;
        RECT 782.430 995.720 783.430 998.810 ;
      LAYER met2 ;
        RECT 783.710 996.000 783.990 1000.000 ;
      LAYER met2 ;
        RECT 784.270 995.720 785.730 998.810 ;
      LAYER met2 ;
        RECT 786.010 996.000 786.290 1000.000 ;
      LAYER met2 ;
        RECT 786.570 995.720 788.030 998.810 ;
      LAYER met2 ;
        RECT 788.310 996.000 788.590 1000.000 ;
      LAYER met2 ;
        RECT 788.870 995.720 789.870 998.810 ;
      LAYER met2 ;
        RECT 790.150 996.000 790.430 1000.000 ;
      LAYER met2 ;
        RECT 790.710 995.720 792.170 998.810 ;
      LAYER met2 ;
        RECT 792.450 996.000 792.730 1000.000 ;
      LAYER met2 ;
        RECT 793.010 995.720 794.470 998.810 ;
      LAYER met2 ;
        RECT 794.750 996.000 795.030 1000.000 ;
      LAYER met2 ;
        RECT 795.310 995.720 796.770 998.810 ;
      LAYER met2 ;
        RECT 797.050 996.000 797.330 1000.000 ;
      LAYER met2 ;
        RECT 797.610 995.720 798.610 998.810 ;
      LAYER met2 ;
        RECT 798.890 996.000 799.170 1000.000 ;
      LAYER met2 ;
        RECT 799.450 995.720 800.910 998.810 ;
      LAYER met2 ;
        RECT 801.190 996.000 801.470 1000.000 ;
      LAYER met2 ;
        RECT 801.750 995.720 803.210 998.810 ;
      LAYER met2 ;
        RECT 803.490 996.000 803.770 1000.000 ;
      LAYER met2 ;
        RECT 804.050 995.720 805.510 998.810 ;
      LAYER met2 ;
        RECT 805.790 996.000 806.070 1000.000 ;
      LAYER met2 ;
        RECT 806.350 995.720 807.350 998.810 ;
      LAYER met2 ;
        RECT 807.630 996.000 807.910 1000.000 ;
      LAYER met2 ;
        RECT 808.190 995.720 809.650 998.810 ;
      LAYER met2 ;
        RECT 809.930 996.000 810.210 1000.000 ;
      LAYER met2 ;
        RECT 810.490 995.720 811.950 998.810 ;
      LAYER met2 ;
        RECT 812.230 996.000 812.510 1000.000 ;
      LAYER met2 ;
        RECT 812.790 995.720 813.790 998.810 ;
      LAYER met2 ;
        RECT 814.070 996.000 814.350 1000.000 ;
      LAYER met2 ;
        RECT 814.630 995.720 816.090 998.810 ;
      LAYER met2 ;
        RECT 816.370 996.000 816.650 1000.000 ;
      LAYER met2 ;
        RECT 816.930 995.720 818.390 998.810 ;
      LAYER met2 ;
        RECT 818.670 996.000 818.950 1000.000 ;
      LAYER met2 ;
        RECT 819.230 995.720 820.690 998.810 ;
      LAYER met2 ;
        RECT 820.970 996.000 821.250 1000.000 ;
      LAYER met2 ;
        RECT 821.530 995.720 822.530 998.810 ;
      LAYER met2 ;
        RECT 822.810 996.000 823.090 1000.000 ;
      LAYER met2 ;
        RECT 823.370 995.720 824.830 998.810 ;
      LAYER met2 ;
        RECT 825.110 996.000 825.390 1000.000 ;
      LAYER met2 ;
        RECT 825.670 995.720 827.130 998.810 ;
      LAYER met2 ;
        RECT 827.410 996.000 827.690 1000.000 ;
      LAYER met2 ;
        RECT 827.970 995.720 829.430 998.810 ;
      LAYER met2 ;
        RECT 829.710 996.000 829.990 1000.000 ;
      LAYER met2 ;
        RECT 830.270 995.720 831.270 998.810 ;
      LAYER met2 ;
        RECT 831.550 996.000 831.830 1000.000 ;
      LAYER met2 ;
        RECT 832.110 995.720 833.570 998.810 ;
      LAYER met2 ;
        RECT 833.850 996.000 834.130 1000.000 ;
      LAYER met2 ;
        RECT 834.410 995.720 835.870 998.810 ;
      LAYER met2 ;
        RECT 836.150 996.000 836.430 1000.000 ;
      LAYER met2 ;
        RECT 836.710 995.720 837.710 998.810 ;
      LAYER met2 ;
        RECT 837.990 996.000 838.270 1000.000 ;
      LAYER met2 ;
        RECT 838.550 995.720 840.010 998.810 ;
      LAYER met2 ;
        RECT 840.290 996.000 840.570 1000.000 ;
        RECT 841.960 999.870 842.870 1000.000 ;
        RECT 843.340 999.870 845.170 1000.000 ;
        RECT 845.640 999.870 847.010 1000.000 ;
      LAYER met2 ;
        RECT 840.850 995.720 842.310 998.810 ;
      LAYER met2 ;
        RECT 842.590 996.000 842.870 999.870 ;
      LAYER met2 ;
        RECT 843.150 995.720 844.610 998.810 ;
      LAYER met2 ;
        RECT 844.890 996.000 845.170 999.870 ;
      LAYER met2 ;
        RECT 845.450 995.720 846.450 998.810 ;
      LAYER met2 ;
        RECT 846.730 996.000 847.010 999.870 ;
      LAYER met2 ;
        RECT 847.290 995.720 848.750 998.810 ;
      LAYER met2 ;
        RECT 849.030 996.000 849.310 1000.000 ;
      LAYER met2 ;
        RECT 849.590 995.720 851.050 998.810 ;
      LAYER met2 ;
        RECT 851.330 996.000 851.610 1000.000 ;
      LAYER met2 ;
        RECT 851.890 995.720 852.890 998.810 ;
      LAYER met2 ;
        RECT 853.170 996.000 853.450 1000.000 ;
      LAYER met2 ;
        RECT 853.730 995.720 855.190 998.810 ;
      LAYER met2 ;
        RECT 855.470 996.000 855.750 1000.000 ;
      LAYER met2 ;
        RECT 856.030 995.720 857.490 998.810 ;
      LAYER met2 ;
        RECT 857.770 996.000 858.050 1000.000 ;
      LAYER met2 ;
        RECT 858.330 995.720 859.790 998.810 ;
      LAYER met2 ;
        RECT 860.070 996.000 860.350 1000.000 ;
      LAYER met2 ;
        RECT 860.630 995.720 861.630 998.810 ;
      LAYER met2 ;
        RECT 861.910 996.000 862.190 1000.000 ;
      LAYER met2 ;
        RECT 862.470 995.720 863.930 998.810 ;
      LAYER met2 ;
        RECT 864.210 996.000 864.490 1000.000 ;
      LAYER met2 ;
        RECT 864.770 995.720 866.230 998.810 ;
      LAYER met2 ;
        RECT 866.510 996.000 866.790 1000.000 ;
      LAYER met2 ;
        RECT 867.070 995.720 868.530 998.810 ;
      LAYER met2 ;
        RECT 868.810 996.000 869.090 1000.000 ;
      LAYER met2 ;
        RECT 869.370 995.720 870.370 998.810 ;
      LAYER met2 ;
        RECT 870.650 996.000 870.930 1000.000 ;
      LAYER met2 ;
        RECT 871.210 995.720 872.670 998.810 ;
      LAYER met2 ;
        RECT 872.950 996.000 873.230 1000.000 ;
      LAYER met2 ;
        RECT 873.510 995.720 874.970 998.810 ;
      LAYER met2 ;
        RECT 875.250 996.000 875.530 1000.000 ;
      LAYER met2 ;
        RECT 875.810 995.720 876.810 998.810 ;
      LAYER met2 ;
        RECT 877.090 996.000 877.370 1000.000 ;
      LAYER met2 ;
        RECT 877.650 995.720 879.110 998.810 ;
      LAYER met2 ;
        RECT 879.390 996.000 879.670 1000.000 ;
      LAYER met2 ;
        RECT 879.950 995.720 881.410 998.810 ;
      LAYER met2 ;
        RECT 881.690 996.000 881.970 1000.000 ;
      LAYER met2 ;
        RECT 882.250 995.720 883.710 998.810 ;
      LAYER met2 ;
        RECT 883.990 996.000 884.270 1000.000 ;
        RECT 884.740 999.870 886.110 1000.000 ;
      LAYER met2 ;
        RECT 884.550 995.720 885.550 998.810 ;
      LAYER met2 ;
        RECT 885.830 996.000 886.110 999.870 ;
      LAYER met2 ;
        RECT 886.390 995.720 887.850 998.810 ;
      LAYER met2 ;
        RECT 888.130 996.000 888.410 1000.000 ;
        RECT 890.260 999.870 890.710 1000.000 ;
      LAYER met2 ;
        RECT 888.690 995.720 890.150 998.810 ;
      LAYER met2 ;
        RECT 890.430 996.000 890.710 999.870 ;
      LAYER met2 ;
        RECT 890.990 995.720 892.450 998.810 ;
      LAYER met2 ;
        RECT 892.730 996.000 893.010 1000.000 ;
        RECT 893.480 999.870 894.850 1000.000 ;
      LAYER met2 ;
        RECT 893.290 995.720 894.290 998.810 ;
      LAYER met2 ;
        RECT 894.570 996.000 894.850 999.870 ;
      LAYER met2 ;
        RECT 895.130 995.720 896.590 998.810 ;
      LAYER met2 ;
        RECT 896.870 996.000 897.150 1000.000 ;
        RECT 897.620 999.870 899.450 1000.000 ;
      LAYER met2 ;
        RECT 897.430 995.720 898.890 998.810 ;
      LAYER met2 ;
        RECT 899.170 996.000 899.450 999.870 ;
      LAYER met2 ;
        RECT 899.730 995.720 900.730 998.810 ;
      LAYER met2 ;
        RECT 901.010 996.000 901.290 1000.000 ;
        RECT 901.760 999.870 903.590 1000.000 ;
      LAYER met2 ;
        RECT 901.570 995.720 903.030 998.810 ;
      LAYER met2 ;
        RECT 903.310 996.000 903.590 999.870 ;
      LAYER met2 ;
        RECT 903.870 995.720 905.330 998.810 ;
      LAYER met2 ;
        RECT 905.610 996.000 905.890 1000.000 ;
        RECT 906.360 999.870 908.190 1000.000 ;
      LAYER met2 ;
        RECT 906.170 995.720 907.630 998.810 ;
      LAYER met2 ;
        RECT 907.910 996.000 908.190 999.870 ;
      LAYER met2 ;
        RECT 908.470 995.720 909.470 998.810 ;
      LAYER met2 ;
        RECT 909.750 996.000 910.030 1000.000 ;
        RECT 910.960 999.870 912.330 1000.000 ;
      LAYER met2 ;
        RECT 910.310 995.720 911.770 998.810 ;
      LAYER met2 ;
        RECT 912.050 996.000 912.330 999.870 ;
      LAYER met2 ;
        RECT 912.610 995.720 914.070 998.810 ;
      LAYER met2 ;
        RECT 914.350 996.000 914.630 1000.000 ;
      LAYER met2 ;
        RECT 914.910 995.720 916.370 998.810 ;
      LAYER met2 ;
        RECT 916.650 996.000 916.930 1000.000 ;
      LAYER met2 ;
        RECT 917.210 995.720 918.210 998.810 ;
      LAYER met2 ;
        RECT 918.490 996.000 918.770 1000.000 ;
      LAYER met2 ;
        RECT 919.050 995.720 920.510 998.810 ;
      LAYER met2 ;
        RECT 920.790 996.000 921.070 1000.000 ;
      LAYER met2 ;
        RECT 921.350 995.720 922.810 998.810 ;
      LAYER met2 ;
        RECT 923.090 996.000 923.370 1000.000 ;
      LAYER met2 ;
        RECT 923.650 995.720 924.650 998.810 ;
      LAYER met2 ;
        RECT 924.930 996.000 925.210 1000.000 ;
      LAYER met2 ;
        RECT 925.490 995.720 926.950 998.810 ;
      LAYER met2 ;
        RECT 927.230 996.000 927.510 1000.000 ;
      LAYER met2 ;
        RECT 927.790 995.720 929.250 998.810 ;
      LAYER met2 ;
        RECT 929.530 996.000 929.810 1000.000 ;
      LAYER met2 ;
        RECT 930.090 995.720 931.550 998.810 ;
      LAYER met2 ;
        RECT 931.830 996.000 932.110 1000.000 ;
      LAYER met2 ;
        RECT 932.390 995.720 933.390 998.810 ;
      LAYER met2 ;
        RECT 933.670 996.000 933.950 1000.000 ;
      LAYER met2 ;
        RECT 934.230 995.720 935.690 998.810 ;
      LAYER met2 ;
        RECT 935.970 996.000 936.250 1000.000 ;
      LAYER met2 ;
        RECT 936.530 995.720 937.990 998.810 ;
      LAYER met2 ;
        RECT 938.270 996.000 938.550 1000.000 ;
      LAYER met2 ;
        RECT 938.830 995.720 940.290 998.810 ;
      LAYER met2 ;
        RECT 940.570 996.000 940.850 1000.000 ;
      LAYER met2 ;
        RECT 941.130 995.720 942.130 998.810 ;
      LAYER met2 ;
        RECT 942.410 996.000 942.690 1000.000 ;
      LAYER met2 ;
        RECT 942.970 995.720 944.430 998.810 ;
      LAYER met2 ;
        RECT 944.710 996.000 944.990 1000.000 ;
      LAYER met2 ;
        RECT 945.270 995.720 946.730 998.810 ;
      LAYER met2 ;
        RECT 947.010 996.000 947.290 1000.000 ;
      LAYER met2 ;
        RECT 947.570 995.720 948.570 998.810 ;
      LAYER met2 ;
        RECT 948.850 996.000 949.130 1000.000 ;
      LAYER met2 ;
        RECT 949.410 995.720 950.870 998.810 ;
      LAYER met2 ;
        RECT 951.150 996.000 951.430 1000.000 ;
      LAYER met2 ;
        RECT 951.710 995.720 953.170 998.810 ;
      LAYER met2 ;
        RECT 953.450 996.000 953.730 1000.000 ;
      LAYER met2 ;
        RECT 954.010 995.720 955.470 998.810 ;
      LAYER met2 ;
        RECT 955.750 996.000 956.030 1000.000 ;
      LAYER met2 ;
        RECT 956.310 995.720 957.310 998.810 ;
      LAYER met2 ;
        RECT 957.590 996.000 957.870 1000.000 ;
      LAYER met2 ;
        RECT 958.150 995.720 959.610 998.810 ;
      LAYER met2 ;
        RECT 959.890 996.000 960.170 1000.000 ;
      LAYER met2 ;
        RECT 960.450 995.720 961.910 998.810 ;
      LAYER met2 ;
        RECT 962.190 996.000 962.470 1000.000 ;
      LAYER met2 ;
        RECT 962.750 995.720 964.210 998.810 ;
      LAYER met2 ;
        RECT 964.490 996.000 964.770 1000.000 ;
      LAYER met2 ;
        RECT 965.050 995.720 966.050 998.810 ;
      LAYER met2 ;
        RECT 966.330 996.000 966.610 1000.000 ;
      LAYER met2 ;
        RECT 966.890 995.720 968.350 998.810 ;
      LAYER met2 ;
        RECT 968.630 996.000 968.910 1000.000 ;
      LAYER met2 ;
        RECT 969.190 995.720 970.650 998.810 ;
      LAYER met2 ;
        RECT 970.930 996.000 971.210 1000.000 ;
      LAYER met2 ;
        RECT 971.490 995.720 972.490 998.810 ;
      LAYER met2 ;
        RECT 972.770 996.000 973.050 1000.000 ;
      LAYER met2 ;
        RECT 973.330 995.720 974.790 998.810 ;
      LAYER met2 ;
        RECT 975.070 996.000 975.350 1000.000 ;
      LAYER met2 ;
        RECT 975.630 995.720 977.090 998.810 ;
      LAYER met2 ;
        RECT 977.370 996.000 977.650 1000.000 ;
      LAYER met2 ;
        RECT 977.930 995.720 979.390 998.810 ;
      LAYER met2 ;
        RECT 979.670 996.000 979.950 1000.000 ;
      LAYER met2 ;
        RECT 980.230 995.720 981.230 998.810 ;
      LAYER met2 ;
        RECT 981.510 996.000 981.790 1000.000 ;
      LAYER met2 ;
        RECT 982.070 995.720 983.530 998.810 ;
      LAYER met2 ;
        RECT 983.810 996.000 984.090 1000.000 ;
      LAYER met2 ;
        RECT 984.370 995.720 985.830 998.810 ;
      LAYER met2 ;
        RECT 986.110 996.000 986.390 1000.000 ;
      LAYER met2 ;
        RECT 986.670 995.720 988.130 998.810 ;
      LAYER met2 ;
        RECT 988.410 996.000 988.690 1000.000 ;
      LAYER met2 ;
        RECT 988.970 995.720 989.970 998.810 ;
      LAYER met2 ;
        RECT 990.250 996.000 990.530 1000.000 ;
      LAYER met2 ;
        RECT 990.810 995.720 992.270 998.810 ;
      LAYER met2 ;
        RECT 992.550 996.000 992.830 1000.000 ;
      LAYER met2 ;
        RECT 993.110 995.720 994.570 998.810 ;
      LAYER met2 ;
        RECT 994.850 996.000 995.130 1000.000 ;
      LAYER met2 ;
        RECT 995.410 995.720 996.410 998.810 ;
      LAYER met2 ;
        RECT 996.690 996.000 996.970 1000.000 ;
      LAYER met2 ;
        RECT 997.250 995.720 998.710 998.810 ;
      LAYER met2 ;
        RECT 998.990 996.000 999.270 1000.000 ;
      LAYER met2 ;
        RECT 999.550 995.720 1001.010 998.810 ;
      LAYER met2 ;
        RECT 1001.290 996.000 1001.570 1000.000 ;
      LAYER met2 ;
        RECT 1001.850 995.720 1003.310 998.810 ;
      LAYER met2 ;
        RECT 1003.590 996.000 1003.870 1000.000 ;
      LAYER met2 ;
        RECT 1004.150 995.720 1005.150 998.810 ;
      LAYER met2 ;
        RECT 1005.430 996.000 1005.710 1000.000 ;
      LAYER met2 ;
        RECT 1005.990 995.720 1007.450 998.810 ;
      LAYER met2 ;
        RECT 1007.730 996.000 1008.010 1000.000 ;
      LAYER met2 ;
        RECT 1008.290 995.720 1009.750 998.810 ;
      LAYER met2 ;
        RECT 1010.030 996.000 1010.310 1000.000 ;
      LAYER met2 ;
        RECT 1010.590 995.720 1011.590 998.810 ;
      LAYER met2 ;
        RECT 1011.870 996.000 1012.150 1000.000 ;
        RECT 1014.170 999.870 1014.600 1000.000 ;
      LAYER met2 ;
        RECT 1012.430 995.720 1013.890 998.810 ;
      LAYER met2 ;
        RECT 1014.170 996.000 1014.450 999.870 ;
      LAYER met2 ;
        RECT 1014.730 995.720 1016.190 998.810 ;
      LAYER met2 ;
        RECT 1016.470 996.000 1016.750 1000.000 ;
      LAYER met2 ;
        RECT 1017.030 995.720 1018.490 998.810 ;
      LAYER met2 ;
        RECT 1018.770 996.000 1019.050 1000.000 ;
      LAYER met2 ;
        RECT 1019.330 995.720 1020.330 998.810 ;
      LAYER met2 ;
        RECT 1020.610 996.000 1020.890 1000.000 ;
      LAYER met2 ;
        RECT 1021.170 995.720 1022.630 998.810 ;
      LAYER met2 ;
        RECT 1022.910 996.000 1023.190 1000.000 ;
      LAYER met2 ;
        RECT 1023.470 995.720 1024.930 998.810 ;
      LAYER met2 ;
        RECT 1025.210 996.000 1025.490 1000.000 ;
      LAYER met2 ;
        RECT 1025.770 995.720 1027.230 998.810 ;
      LAYER met2 ;
        RECT 1027.510 996.000 1027.790 1000.000 ;
      LAYER met2 ;
        RECT 1028.070 995.720 1029.070 998.810 ;
      LAYER met2 ;
        RECT 1029.350 996.000 1029.630 1000.000 ;
      LAYER met2 ;
        RECT 1029.910 995.720 1031.370 998.810 ;
      LAYER met2 ;
        RECT 1031.650 996.000 1031.930 1000.000 ;
      LAYER met2 ;
        RECT 1032.210 995.720 1033.670 998.810 ;
      LAYER met2 ;
        RECT 1033.950 996.000 1034.230 1000.000 ;
      LAYER met2 ;
        RECT 1034.510 995.720 1035.510 998.810 ;
      LAYER met2 ;
        RECT 1035.790 996.000 1036.070 1000.000 ;
      LAYER met2 ;
        RECT 1036.350 995.720 1037.810 998.810 ;
      LAYER met2 ;
        RECT 1038.090 996.000 1038.370 1000.000 ;
      LAYER met2 ;
        RECT 1038.650 995.720 1040.110 998.810 ;
      LAYER met2 ;
        RECT 1040.390 996.000 1040.670 1000.000 ;
      LAYER met2 ;
        RECT 1040.950 995.720 1042.410 998.810 ;
      LAYER met2 ;
        RECT 1042.690 996.000 1042.970 1000.000 ;
      LAYER met2 ;
        RECT 1043.250 995.720 1044.250 998.810 ;
      LAYER met2 ;
        RECT 1044.530 996.000 1044.810 1000.000 ;
      LAYER met2 ;
        RECT 1045.090 995.720 1046.550 998.810 ;
      LAYER met2 ;
        RECT 1046.830 996.000 1047.110 1000.000 ;
      LAYER met2 ;
        RECT 1047.390 995.720 1048.850 998.810 ;
      LAYER met2 ;
        RECT 1049.130 996.000 1049.410 1000.000 ;
        RECT 1050.340 999.870 1051.710 1000.000 ;
      LAYER met2 ;
        RECT 1049.690 995.720 1051.150 998.810 ;
      LAYER met2 ;
        RECT 1051.430 996.000 1051.710 999.870 ;
      LAYER met2 ;
        RECT 1051.990 995.720 1052.990 998.810 ;
      LAYER met2 ;
        RECT 1053.270 996.000 1053.550 1000.000 ;
        RECT 1055.570 999.870 1056.000 1000.000 ;
      LAYER met2 ;
        RECT 1053.830 995.720 1055.290 998.810 ;
      LAYER met2 ;
        RECT 1055.570 996.000 1055.850 999.870 ;
      LAYER met2 ;
        RECT 1056.130 995.720 1057.590 998.810 ;
      LAYER met2 ;
        RECT 1057.870 996.000 1058.150 1000.000 ;
        RECT 1058.620 999.870 1059.990 1000.000 ;
      LAYER met2 ;
        RECT 1058.430 995.720 1059.430 998.810 ;
      LAYER met2 ;
        RECT 1059.710 996.000 1059.990 999.870 ;
      LAYER met2 ;
        RECT 1060.270 995.720 1061.730 998.810 ;
      LAYER met2 ;
        RECT 1062.010 996.000 1062.290 1000.000 ;
        RECT 1062.760 999.870 1064.590 1000.000 ;
      LAYER met2 ;
        RECT 1062.570 995.720 1064.030 998.810 ;
      LAYER met2 ;
        RECT 1064.310 996.000 1064.590 999.870 ;
      LAYER met2 ;
        RECT 1064.870 995.720 1066.330 998.810 ;
      LAYER met2 ;
        RECT 1066.610 996.000 1066.890 1000.000 ;
        RECT 1067.360 999.870 1068.730 1000.000 ;
      LAYER met2 ;
        RECT 1067.170 995.720 1068.170 998.810 ;
      LAYER met2 ;
        RECT 1068.450 996.000 1068.730 999.870 ;
      LAYER met2 ;
        RECT 1069.010 995.720 1070.470 998.810 ;
      LAYER met2 ;
        RECT 1070.750 996.000 1071.030 1000.000 ;
        RECT 1071.960 999.870 1073.330 1000.000 ;
      LAYER met2 ;
        RECT 1071.310 995.720 1072.770 998.810 ;
      LAYER met2 ;
        RECT 1073.050 996.000 1073.330 999.870 ;
      LAYER met2 ;
        RECT 1073.610 995.720 1075.070 998.810 ;
      LAYER met2 ;
        RECT 1075.350 996.000 1075.630 1000.000 ;
        RECT 1076.560 999.870 1077.470 1000.000 ;
      LAYER met2 ;
        RECT 1075.910 995.720 1076.910 998.810 ;
      LAYER met2 ;
        RECT 1077.190 996.000 1077.470 999.870 ;
      LAYER met2 ;
        RECT 1077.750 995.720 1079.210 998.810 ;
      LAYER met2 ;
        RECT 1079.490 996.000 1079.770 1000.000 ;
        RECT 1080.240 999.870 1082.070 1000.000 ;
      LAYER met2 ;
        RECT 1080.050 995.720 1081.510 998.810 ;
      LAYER met2 ;
        RECT 1081.790 996.000 1082.070 999.870 ;
      LAYER met2 ;
        RECT 1082.350 995.720 1083.350 998.810 ;
      LAYER met2 ;
        RECT 1083.630 996.000 1083.910 1000.000 ;
        RECT 1084.380 999.870 1086.210 1000.000 ;
      LAYER met2 ;
        RECT 1084.190 995.720 1085.650 998.810 ;
      LAYER met2 ;
        RECT 1085.930 996.000 1086.210 999.870 ;
      LAYER met2 ;
        RECT 1086.490 995.720 1087.950 998.810 ;
      LAYER met2 ;
        RECT 1088.230 996.000 1088.510 1000.000 ;
        RECT 1090.360 999.870 1090.810 1000.000 ;
      LAYER met2 ;
        RECT 1088.790 995.720 1090.250 998.810 ;
      LAYER met2 ;
        RECT 1090.530 996.000 1090.810 999.870 ;
      LAYER met2 ;
        RECT 1091.090 995.720 1092.090 998.810 ;
      LAYER met2 ;
        RECT 1092.370 996.000 1092.650 1000.000 ;
        RECT 1093.120 999.870 1094.950 1000.000 ;
      LAYER met2 ;
        RECT 1092.930 995.720 1094.390 998.810 ;
      LAYER met2 ;
        RECT 1094.670 996.000 1094.950 999.870 ;
      LAYER met2 ;
        RECT 1095.230 995.720 1096.690 998.810 ;
      LAYER met2 ;
        RECT 1096.970 996.000 1097.250 1000.000 ;
        RECT 1097.720 999.870 1099.550 1000.000 ;
      LAYER met2 ;
        RECT 1097.530 995.720 1098.990 998.810 ;
      LAYER met2 ;
        RECT 1099.270 996.000 1099.550 999.870 ;
      LAYER met2 ;
        RECT 1099.830 995.720 1100.830 998.810 ;
      LAYER met2 ;
        RECT 1101.110 996.000 1101.390 1000.000 ;
        RECT 1101.860 999.870 1103.690 1000.000 ;
      LAYER met2 ;
        RECT 1101.670 995.720 1103.130 998.810 ;
      LAYER met2 ;
        RECT 1103.410 996.000 1103.690 999.870 ;
      LAYER met2 ;
        RECT 1103.970 995.720 1105.430 998.810 ;
      LAYER met2 ;
        RECT 1105.710 996.000 1105.990 1000.000 ;
        RECT 1106.460 999.870 1107.830 1000.000 ;
      LAYER met2 ;
        RECT 1106.270 995.720 1107.270 998.810 ;
      LAYER met2 ;
        RECT 1107.550 996.000 1107.830 999.870 ;
      LAYER met2 ;
        RECT 1108.110 995.720 1109.570 998.810 ;
      LAYER met2 ;
        RECT 1109.850 996.000 1110.130 1000.000 ;
        RECT 1111.060 999.870 1112.430 1000.000 ;
      LAYER met2 ;
        RECT 1110.410 995.720 1111.870 998.810 ;
      LAYER met2 ;
        RECT 1112.150 996.000 1112.430 999.870 ;
      LAYER met2 ;
        RECT 1112.710 995.720 1114.170 998.810 ;
      LAYER met2 ;
        RECT 1114.450 996.000 1114.730 1000.000 ;
        RECT 1115.200 999.870 1116.570 1000.000 ;
      LAYER met2 ;
        RECT 1115.010 995.720 1116.010 998.810 ;
      LAYER met2 ;
        RECT 1116.290 996.000 1116.570 999.870 ;
      LAYER met2 ;
        RECT 1116.850 995.720 1118.310 998.810 ;
      LAYER met2 ;
        RECT 1118.590 996.000 1118.870 1000.000 ;
        RECT 1119.340 999.870 1121.170 1000.000 ;
      LAYER met2 ;
        RECT 1119.150 995.720 1120.610 998.810 ;
      LAYER met2 ;
        RECT 1120.890 996.000 1121.170 999.870 ;
      LAYER met2 ;
        RECT 1121.450 995.720 1122.910 998.810 ;
      LAYER met2 ;
        RECT 1123.190 996.000 1123.470 1000.000 ;
      LAYER met2 ;
        RECT 1123.750 995.720 1124.750 998.810 ;
      LAYER met2 ;
        RECT 1125.030 996.000 1125.310 1000.000 ;
        RECT 1125.780 999.870 1127.610 1000.000 ;
      LAYER met2 ;
        RECT 1125.590 995.720 1127.050 998.810 ;
      LAYER met2 ;
        RECT 1127.330 996.000 1127.610 999.870 ;
      LAYER met2 ;
        RECT 1127.890 995.720 1129.350 998.810 ;
      LAYER met2 ;
        RECT 1129.630 996.000 1129.910 1000.000 ;
        RECT 1131.470 999.870 1131.900 1000.000 ;
      LAYER met2 ;
        RECT 1130.190 995.720 1131.190 998.810 ;
      LAYER met2 ;
        RECT 1131.470 996.000 1131.750 999.870 ;
      LAYER met2 ;
        RECT 1132.030 995.720 1133.490 998.810 ;
      LAYER met2 ;
        RECT 1133.770 996.000 1134.050 1000.000 ;
        RECT 1134.520 999.870 1136.350 1000.000 ;
      LAYER met2 ;
        RECT 1134.330 995.720 1135.790 998.810 ;
      LAYER met2 ;
        RECT 1136.070 996.000 1136.350 999.870 ;
      LAYER met2 ;
        RECT 1136.630 995.720 1138.090 998.810 ;
      LAYER met2 ;
        RECT 1138.370 996.000 1138.650 1000.000 ;
        RECT 1139.580 999.870 1140.490 1000.000 ;
      LAYER met2 ;
        RECT 1138.930 995.720 1139.930 998.810 ;
      LAYER met2 ;
        RECT 1140.210 996.000 1140.490 999.870 ;
      LAYER met2 ;
        RECT 1140.770 995.720 1142.230 998.810 ;
      LAYER met2 ;
        RECT 1142.510 996.000 1142.790 1000.000 ;
        RECT 1143.260 999.870 1145.090 1000.000 ;
      LAYER met2 ;
        RECT 1143.070 995.720 1144.530 998.810 ;
      LAYER met2 ;
        RECT 1144.810 996.000 1145.090 999.870 ;
      LAYER met2 ;
        RECT 1145.370 995.720 1146.830 998.810 ;
      LAYER met2 ;
        RECT 1147.110 996.000 1147.390 1000.000 ;
        RECT 1147.860 999.870 1149.230 1000.000 ;
      LAYER met2 ;
        RECT 1147.670 995.720 1148.670 998.810 ;
      LAYER met2 ;
        RECT 1148.950 996.000 1149.230 999.870 ;
      LAYER met2 ;
        RECT 1149.510 995.720 1150.970 998.810 ;
      LAYER met2 ;
        RECT 1151.250 996.000 1151.530 1000.000 ;
        RECT 1152.460 999.870 1153.830 1000.000 ;
      LAYER met2 ;
        RECT 1151.810 995.720 1153.270 998.810 ;
      LAYER met2 ;
        RECT 1153.550 996.000 1153.830 999.870 ;
      LAYER met2 ;
        RECT 1154.110 995.720 1155.110 998.810 ;
      LAYER met2 ;
        RECT 1155.390 996.000 1155.670 1000.000 ;
        RECT 1156.140 999.870 1157.970 1000.000 ;
      LAYER met2 ;
        RECT 1155.950 995.720 1157.410 998.810 ;
      LAYER met2 ;
        RECT 1157.690 996.000 1157.970 999.870 ;
      LAYER met2 ;
        RECT 1158.250 995.720 1159.710 998.810 ;
      LAYER met2 ;
        RECT 1159.990 996.000 1160.270 1000.000 ;
        RECT 1160.740 999.870 1162.570 1000.000 ;
      LAYER met2 ;
        RECT 1160.550 995.720 1162.010 998.810 ;
      LAYER met2 ;
        RECT 1162.290 996.000 1162.570 999.870 ;
      LAYER met2 ;
        RECT 1162.850 995.720 1163.850 998.810 ;
      LAYER met2 ;
        RECT 1164.130 996.000 1164.410 1000.000 ;
        RECT 1166.260 999.870 1166.710 1000.000 ;
        RECT 1167.180 999.870 1169.010 1000.000 ;
      LAYER met2 ;
        RECT 1164.690 995.720 1166.150 998.810 ;
      LAYER met2 ;
        RECT 1166.430 996.000 1166.710 999.870 ;
      LAYER met2 ;
        RECT 1166.990 995.720 1168.450 998.810 ;
      LAYER met2 ;
        RECT 1168.730 996.000 1169.010 999.870 ;
      LAYER met2 ;
        RECT 1169.290 995.720 1170.750 998.810 ;
      LAYER met2 ;
        RECT 1171.030 996.000 1171.310 1000.000 ;
      LAYER met2 ;
        RECT 1171.590 995.720 1172.590 998.810 ;
      LAYER met2 ;
        RECT 1172.870 996.000 1173.150 1000.000 ;
      LAYER met2 ;
        RECT 1173.430 995.720 1174.890 998.810 ;
      LAYER met2 ;
        RECT 1175.170 996.000 1175.450 1000.000 ;
      LAYER met2 ;
        RECT 1175.730 995.720 1177.190 998.810 ;
      LAYER met2 ;
        RECT 1177.470 996.000 1177.750 1000.000 ;
      LAYER met2 ;
        RECT 1178.030 995.720 1179.030 998.810 ;
      LAYER met2 ;
        RECT 1179.310 996.000 1179.590 1000.000 ;
        RECT 1181.610 999.870 1183.420 1000.000 ;
        RECT 1183.740 1000.010 1183.880 1008.790 ;
        RECT 1186.040 1000.010 1186.180 1693.355 ;
        RECT 1186.500 1010.130 1186.640 1693.550 ;
        RECT 1187.880 1686.390 1188.020 1700.000 ;
        RECT 1190.580 1689.810 1190.840 1690.130 ;
        RECT 1188.740 1688.790 1189.000 1689.110 ;
        RECT 1187.820 1686.070 1188.080 1686.390 ;
        RECT 1186.440 1009.810 1186.700 1010.130 ;
        RECT 1186.900 1008.110 1187.160 1008.430 ;
        RECT 1186.960 1000.010 1187.100 1008.110 ;
        RECT 1188.800 1000.010 1188.940 1688.790 ;
        RECT 1190.120 1685.730 1190.380 1686.050 ;
        RECT 1190.180 1008.430 1190.320 1685.730 ;
        RECT 1190.640 1009.110 1190.780 1689.810 ;
        RECT 1195.180 1689.130 1195.440 1689.450 ;
        RECT 1195.240 1686.050 1195.380 1689.130 ;
        RECT 1200.240 1688.790 1200.500 1689.110 ;
        RECT 1195.180 1685.730 1195.440 1686.050 ;
        RECT 1200.300 1025.430 1200.440 1688.790 ;
        RECT 1196.100 1025.110 1196.360 1025.430 ;
        RECT 1200.240 1025.110 1200.500 1025.430 ;
        RECT 1193.800 1019.670 1194.060 1019.990 ;
        RECT 1191.490 1009.955 1191.770 1010.325 ;
        RECT 1190.580 1008.790 1190.840 1009.110 ;
        RECT 1190.120 1008.110 1190.380 1008.430 ;
        RECT 1191.560 1008.090 1191.700 1009.955 ;
        RECT 1191.040 1007.770 1191.300 1008.090 ;
        RECT 1191.500 1007.770 1191.760 1008.090 ;
        RECT 1191.100 1000.010 1191.240 1007.770 ;
        RECT 1183.740 1000.000 1184.040 1000.010 ;
        RECT 1186.040 1000.000 1186.340 1000.010 ;
        RECT 1186.960 1000.000 1188.180 1000.010 ;
        RECT 1188.800 1000.000 1190.480 1000.010 ;
        RECT 1191.100 1000.000 1192.780 1000.010 ;
        RECT 1183.740 999.870 1184.190 1000.000 ;
        RECT 1186.040 999.870 1186.490 1000.000 ;
        RECT 1186.960 999.870 1188.330 1000.000 ;
        RECT 1188.800 999.870 1190.630 1000.000 ;
        RECT 1191.100 999.870 1192.930 1000.000 ;
      LAYER met2 ;
        RECT 1179.870 995.720 1181.330 998.810 ;
      LAYER met2 ;
        RECT 1181.610 996.000 1181.890 999.870 ;
      LAYER met2 ;
        RECT 1182.170 995.720 1183.630 998.810 ;
      LAYER met2 ;
        RECT 1183.910 996.000 1184.190 999.870 ;
      LAYER met2 ;
        RECT 1184.470 995.720 1185.930 998.810 ;
      LAYER met2 ;
        RECT 1186.210 996.000 1186.490 999.870 ;
      LAYER met2 ;
        RECT 1186.770 995.720 1187.770 998.810 ;
      LAYER met2 ;
        RECT 1188.050 996.000 1188.330 999.870 ;
      LAYER met2 ;
        RECT 1188.610 995.720 1190.070 998.810 ;
      LAYER met2 ;
        RECT 1190.350 996.000 1190.630 999.870 ;
      LAYER met2 ;
        RECT 1190.910 995.720 1192.370 998.810 ;
      LAYER met2 ;
        RECT 1192.650 996.000 1192.930 999.870 ;
        RECT 1193.860 999.590 1194.000 1019.670 ;
        RECT 1196.160 1000.010 1196.300 1025.110 ;
        RECT 1200.760 1014.210 1200.900 1700.270 ;
        RECT 1201.570 1700.000 1201.850 1700.270 ;
        RECT 1215.370 1700.000 1215.650 1704.000 ;
        RECT 1230.090 1700.000 1230.370 1704.000 ;
        RECT 1243.890 1700.410 1244.170 1704.000 ;
        RECT 1243.080 1700.270 1244.170 1700.410 ;
        RECT 1207.140 1689.130 1207.400 1689.450 ;
        RECT 1207.200 1014.210 1207.340 1689.130 ;
        RECT 1215.480 1689.110 1215.620 1700.000 ;
        RECT 1220.940 1693.890 1221.200 1694.210 ;
        RECT 1215.420 1688.790 1215.680 1689.110 ;
        RECT 1215.420 1686.070 1215.680 1686.390 ;
        RECT 1197.940 1013.890 1198.200 1014.210 ;
        RECT 1198.400 1013.890 1198.660 1014.210 ;
        RECT 1200.700 1013.890 1200.960 1014.210 ;
        RECT 1202.540 1013.890 1202.800 1014.210 ;
        RECT 1207.140 1013.890 1207.400 1014.210 ;
        RECT 1214.960 1013.890 1215.220 1014.210 ;
        RECT 1198.000 1013.530 1198.140 1013.890 ;
        RECT 1197.480 1013.210 1197.740 1013.530 ;
        RECT 1197.940 1013.210 1198.200 1013.530 ;
        RECT 1197.540 1007.750 1197.680 1013.210 ;
        RECT 1197.480 1007.430 1197.740 1007.750 ;
        RECT 1198.460 1000.010 1198.600 1013.890 ;
        RECT 1200.230 1011.995 1200.510 1012.365 ;
        RECT 1200.300 1009.450 1200.440 1011.995 ;
        RECT 1200.240 1009.130 1200.500 1009.450 ;
        RECT 1202.600 1000.010 1202.740 1013.890 ;
        RECT 1208.980 1013.550 1209.240 1013.870 ;
        RECT 1204.840 1010.150 1205.100 1010.470 ;
        RECT 1204.900 1000.010 1205.040 1010.150 ;
        RECT 1205.300 1009.470 1205.560 1009.790 ;
        RECT 1194.620 1000.000 1196.300 1000.010 ;
        RECT 1196.920 1000.000 1198.600 1000.010 ;
        RECT 1201.520 1000.000 1202.740 1000.010 ;
        RECT 1203.360 1000.000 1205.040 1000.010 ;
        RECT 1194.490 999.870 1196.300 1000.000 ;
        RECT 1196.790 999.870 1198.600 1000.000 ;
        RECT 1193.800 999.270 1194.060 999.590 ;
      LAYER met2 ;
        RECT 1193.210 995.720 1194.210 998.810 ;
      LAYER met2 ;
        RECT 1194.490 996.000 1194.770 999.870 ;
      LAYER met2 ;
        RECT 1195.050 995.720 1196.510 998.810 ;
      LAYER met2 ;
        RECT 1196.790 996.000 1197.070 999.870 ;
        RECT 1197.480 999.330 1197.740 999.590 ;
        RECT 1199.090 999.330 1199.370 1000.000 ;
        RECT 1197.480 999.270 1199.370 999.330 ;
        RECT 1197.540 999.190 1199.370 999.270 ;
      LAYER met2 ;
        RECT 1197.350 995.720 1198.810 998.810 ;
      LAYER met2 ;
        RECT 1199.090 996.000 1199.370 999.190 ;
        RECT 1201.390 999.870 1202.740 1000.000 ;
        RECT 1203.230 999.870 1205.040 1000.000 ;
        RECT 1205.360 1000.010 1205.500 1009.470 ;
        RECT 1207.600 1008.965 1207.860 1009.110 ;
        RECT 1207.590 1008.595 1207.870 1008.965 ;
        RECT 1207.600 1008.285 1207.860 1008.430 ;
        RECT 1207.590 1007.915 1207.870 1008.285 ;
        RECT 1208.060 1008.110 1208.320 1008.430 ;
        RECT 1208.120 1001.290 1208.260 1008.110 ;
        RECT 1208.060 1000.970 1208.320 1001.290 ;
        RECT 1209.040 1000.010 1209.180 1013.550 ;
        RECT 1210.360 1009.470 1210.620 1009.790 ;
        RECT 1209.440 1008.965 1209.700 1009.110 ;
        RECT 1209.430 1008.595 1209.710 1008.965 ;
        RECT 1209.440 1008.285 1209.700 1008.430 ;
        RECT 1209.430 1007.915 1209.710 1008.285 ;
        RECT 1210.420 1000.010 1210.560 1009.470 ;
        RECT 1210.820 1009.130 1211.080 1009.450 ;
        RECT 1205.360 1000.000 1205.660 1000.010 ;
        RECT 1207.960 1000.000 1209.180 1000.010 ;
        RECT 1210.260 1000.000 1210.560 1000.010 ;
        RECT 1205.360 999.870 1205.810 1000.000 ;
      LAYER met2 ;
        RECT 1199.650 995.720 1201.110 998.810 ;
      LAYER met2 ;
        RECT 1201.390 996.000 1201.670 999.870 ;
      LAYER met2 ;
        RECT 1201.950 995.720 1202.950 998.810 ;
      LAYER met2 ;
        RECT 1203.230 996.000 1203.510 999.870 ;
      LAYER met2 ;
        RECT 1203.790 995.720 1205.250 998.810 ;
      LAYER met2 ;
        RECT 1205.530 996.000 1205.810 999.870 ;
        RECT 1207.830 999.870 1209.180 1000.000 ;
        RECT 1210.130 999.870 1210.560 1000.000 ;
        RECT 1210.880 1000.010 1211.020 1009.130 ;
        RECT 1215.020 1000.010 1215.160 1013.890 ;
        RECT 1210.880 1000.000 1212.100 1000.010 ;
        RECT 1214.400 1000.000 1215.160 1000.010 ;
        RECT 1210.880 999.870 1212.250 1000.000 ;
      LAYER met2 ;
        RECT 1206.090 995.720 1207.550 998.810 ;
      LAYER met2 ;
        RECT 1207.830 996.000 1208.110 999.870 ;
      LAYER met2 ;
        RECT 1208.390 995.720 1209.850 998.810 ;
      LAYER met2 ;
        RECT 1210.130 996.000 1210.410 999.870 ;
      LAYER met2 ;
        RECT 1210.690 995.720 1211.690 998.810 ;
      LAYER met2 ;
        RECT 1211.970 996.000 1212.250 999.870 ;
        RECT 1214.270 999.870 1215.160 1000.000 ;
      LAYER met2 ;
        RECT 1212.530 995.720 1213.990 998.810 ;
      LAYER met2 ;
        RECT 1214.270 996.000 1214.550 999.870 ;
        RECT 1215.480 999.590 1215.620 1686.070 ;
        RECT 1220.480 1684.030 1220.740 1684.350 ;
        RECT 1220.020 1048.570 1220.280 1048.890 ;
        RECT 1216.570 1000.970 1216.830 1001.290 ;
        RECT 1216.630 1000.000 1216.770 1000.970 ;
        RECT 1220.080 1000.010 1220.220 1048.570 ;
        RECT 1220.540 1014.210 1220.680 1684.030 ;
        RECT 1221.000 1048.890 1221.140 1693.890 ;
        RECT 1230.200 1689.450 1230.340 1700.000 ;
        RECT 1230.140 1689.130 1230.400 1689.450 ;
        RECT 1238.420 1688.790 1238.680 1689.110 ;
        RECT 1224.620 1685.730 1224.880 1686.050 ;
        RECT 1220.940 1048.570 1221.200 1048.890 ;
        RECT 1220.480 1013.890 1220.740 1014.210 ;
        RECT 1223.700 1012.870 1223.960 1013.190 ;
        RECT 1224.160 1012.870 1224.420 1013.190 ;
        RECT 1223.240 1009.810 1223.500 1010.130 ;
        RECT 1223.300 1000.010 1223.440 1009.810 ;
        RECT 1218.540 1000.000 1220.220 1000.010 ;
        RECT 1223.140 1000.000 1223.440 1000.010 ;
        RECT 1215.420 999.270 1215.680 999.590 ;
      LAYER met2 ;
        RECT 1214.830 995.720 1216.290 998.810 ;
      LAYER met2 ;
        RECT 1216.570 996.000 1216.850 1000.000 ;
        RECT 1218.410 999.870 1220.220 1000.000 ;
      LAYER met2 ;
        RECT 1217.130 995.720 1218.130 998.810 ;
      LAYER met2 ;
        RECT 1218.410 996.000 1218.690 999.870 ;
        RECT 1219.100 999.330 1219.360 999.590 ;
        RECT 1220.710 999.330 1220.990 1000.000 ;
        RECT 1219.100 999.270 1220.990 999.330 ;
        RECT 1219.160 999.190 1220.990 999.270 ;
      LAYER met2 ;
        RECT 1218.970 995.720 1220.430 998.810 ;
      LAYER met2 ;
        RECT 1220.710 996.000 1220.990 999.190 ;
        RECT 1223.010 999.870 1223.440 1000.000 ;
        RECT 1223.760 1000.010 1223.900 1012.870 ;
        RECT 1224.220 1012.510 1224.360 1012.870 ;
        RECT 1224.680 1012.510 1224.820 1685.730 ;
        RECT 1237.960 1019.670 1238.220 1019.990 ;
        RECT 1226.000 1013.210 1226.260 1013.530 ;
        RECT 1224.160 1012.190 1224.420 1012.510 ;
        RECT 1224.620 1012.190 1224.880 1012.510 ;
        RECT 1226.060 1000.010 1226.200 1013.210 ;
        RECT 1228.300 1012.530 1228.560 1012.850 ;
        RECT 1237.500 1012.530 1237.760 1012.850 ;
        RECT 1228.360 1000.010 1228.500 1012.530 ;
        RECT 1230.140 1012.190 1230.400 1012.510 ;
        RECT 1230.200 1000.010 1230.340 1012.190 ;
        RECT 1232.440 1007.430 1232.700 1007.750 ;
        RECT 1232.500 1000.010 1232.640 1007.430 ;
        RECT 1237.560 1000.010 1237.700 1012.530 ;
        RECT 1223.760 1000.000 1225.440 1000.010 ;
        RECT 1226.060 1000.000 1227.280 1000.010 ;
        RECT 1228.360 1000.000 1229.580 1000.010 ;
        RECT 1230.200 1000.000 1231.880 1000.010 ;
        RECT 1232.500 1000.000 1234.180 1000.010 ;
        RECT 1236.020 1000.000 1237.700 1000.010 ;
        RECT 1223.760 999.870 1225.590 1000.000 ;
        RECT 1226.060 999.870 1227.430 1000.000 ;
        RECT 1228.360 999.870 1229.730 1000.000 ;
        RECT 1230.200 999.870 1232.030 1000.000 ;
        RECT 1232.500 999.870 1234.330 1000.000 ;
      LAYER met2 ;
        RECT 1221.270 995.720 1222.730 998.810 ;
      LAYER met2 ;
        RECT 1223.010 996.000 1223.290 999.870 ;
      LAYER met2 ;
        RECT 1223.570 995.720 1225.030 998.810 ;
      LAYER met2 ;
        RECT 1225.310 996.000 1225.590 999.870 ;
      LAYER met2 ;
        RECT 1225.870 995.720 1226.870 998.810 ;
      LAYER met2 ;
        RECT 1227.150 996.000 1227.430 999.870 ;
      LAYER met2 ;
        RECT 1227.710 995.720 1229.170 998.810 ;
      LAYER met2 ;
        RECT 1229.450 996.000 1229.730 999.870 ;
      LAYER met2 ;
        RECT 1230.010 995.720 1231.470 998.810 ;
      LAYER met2 ;
        RECT 1231.750 996.000 1232.030 999.870 ;
      LAYER met2 ;
        RECT 1232.310 995.720 1233.770 998.810 ;
      LAYER met2 ;
        RECT 1234.050 996.000 1234.330 999.870 ;
        RECT 1235.890 999.870 1237.700 1000.000 ;
        RECT 1238.020 1000.010 1238.160 1019.670 ;
        RECT 1238.480 1009.790 1238.620 1688.790 ;
        RECT 1243.080 1684.350 1243.220 1700.270 ;
        RECT 1243.890 1700.000 1244.170 1700.270 ;
        RECT 1258.610 1700.000 1258.890 1704.000 ;
        RECT 1272.410 1700.000 1272.690 1704.000 ;
        RECT 1287.130 1700.000 1287.410 1704.000 ;
        RECT 1300.930 1700.000 1301.210 1704.000 ;
        RECT 1315.650 1700.000 1315.930 1704.000 ;
        RECT 1329.450 1700.410 1329.730 1704.000 ;
        RECT 1329.450 1700.270 1331.540 1700.410 ;
        RECT 1329.450 1700.000 1329.730 1700.270 ;
        RECT 1243.480 1689.470 1243.740 1689.790 ;
        RECT 1254.980 1689.470 1255.240 1689.790 ;
        RECT 1243.020 1684.030 1243.280 1684.350 ;
        RECT 1238.420 1009.470 1238.680 1009.790 ;
        RECT 1238.880 1007.770 1239.140 1008.090 ;
        RECT 1238.940 1000.010 1239.080 1007.770 ;
        RECT 1243.540 1000.010 1243.680 1689.470 ;
        RECT 1243.940 1686.410 1244.200 1686.730 ;
        RECT 1244.000 1014.120 1244.140 1686.410 ;
        RECT 1252.680 1020.010 1252.940 1020.330 ;
        RECT 1244.000 1013.980 1246.440 1014.120 ;
        RECT 1244.860 1013.210 1245.120 1013.530 ;
        RECT 1243.940 1012.190 1244.200 1012.510 ;
        RECT 1244.000 1011.490 1244.140 1012.190 ;
        RECT 1243.940 1011.170 1244.200 1011.490 ;
        RECT 1244.920 1000.010 1245.060 1013.210 ;
        RECT 1238.020 1000.000 1238.320 1000.010 ;
        RECT 1238.940 1000.000 1240.620 1000.010 ;
        RECT 1242.460 1000.000 1243.680 1000.010 ;
        RECT 1244.760 1000.000 1245.060 1000.010 ;
        RECT 1238.020 999.870 1238.470 1000.000 ;
        RECT 1238.940 999.870 1240.770 1000.000 ;
      LAYER met2 ;
        RECT 1234.610 995.720 1235.610 998.810 ;
      LAYER met2 ;
        RECT 1235.890 996.000 1236.170 999.870 ;
      LAYER met2 ;
        RECT 1236.450 995.720 1237.910 998.810 ;
      LAYER met2 ;
        RECT 1238.190 996.000 1238.470 999.870 ;
      LAYER met2 ;
        RECT 1238.750 995.720 1240.210 998.810 ;
      LAYER met2 ;
        RECT 1240.490 996.000 1240.770 999.870 ;
        RECT 1242.330 999.870 1243.680 1000.000 ;
        RECT 1244.630 999.870 1245.060 1000.000 ;
        RECT 1246.300 1000.010 1246.440 1013.980 ;
        RECT 1250.380 1007.770 1250.640 1008.090 ;
        RECT 1250.440 1000.010 1250.580 1007.770 ;
        RECT 1252.740 1000.010 1252.880 1020.010 ;
        RECT 1255.040 1008.090 1255.180 1689.470 ;
        RECT 1258.720 1688.430 1258.860 1700.000 ;
        RECT 1268.320 1694.230 1268.580 1694.550 ;
        RECT 1258.200 1688.110 1258.460 1688.430 ;
        RECT 1258.660 1688.110 1258.920 1688.430 ;
        RECT 1262.340 1688.110 1262.600 1688.430 ;
        RECT 1258.260 1686.730 1258.400 1688.110 ;
        RECT 1258.200 1686.410 1258.460 1686.730 ;
        RECT 1259.120 1013.890 1259.380 1014.210 ;
        RECT 1254.980 1007.770 1255.240 1008.090 ;
        RECT 1254.520 1007.430 1254.780 1007.750 ;
        RECT 1257.280 1007.430 1257.540 1007.750 ;
        RECT 1254.580 1000.010 1254.720 1007.430 ;
        RECT 1257.340 1000.010 1257.480 1007.430 ;
        RECT 1259.180 1000.010 1259.320 1013.890 ;
        RECT 1262.400 1013.870 1262.540 1688.110 ;
        RECT 1267.860 1020.350 1268.120 1020.670 ;
        RECT 1262.340 1013.550 1262.600 1013.870 ;
        RECT 1259.580 1012.870 1259.840 1013.190 ;
        RECT 1265.560 1012.870 1265.820 1013.190 ;
        RECT 1246.300 1000.000 1247.060 1000.010 ;
        RECT 1249.360 1000.000 1250.580 1000.010 ;
        RECT 1251.200 1000.000 1252.880 1000.010 ;
        RECT 1253.500 1000.000 1254.720 1000.010 ;
        RECT 1255.800 1000.000 1257.480 1000.010 ;
        RECT 1258.100 1000.000 1259.320 1000.010 ;
        RECT 1246.300 999.870 1247.210 1000.000 ;
      LAYER met2 ;
        RECT 1241.050 995.720 1242.050 998.810 ;
      LAYER met2 ;
        RECT 1242.330 996.000 1242.610 999.870 ;
      LAYER met2 ;
        RECT 1242.890 995.720 1244.350 998.810 ;
      LAYER met2 ;
        RECT 1244.630 996.000 1244.910 999.870 ;
      LAYER met2 ;
        RECT 1245.190 995.720 1246.650 998.810 ;
      LAYER met2 ;
        RECT 1246.930 996.000 1247.210 999.870 ;
        RECT 1249.230 999.870 1250.580 1000.000 ;
        RECT 1251.070 999.870 1252.880 1000.000 ;
        RECT 1253.370 999.870 1254.720 1000.000 ;
        RECT 1255.670 999.870 1257.480 1000.000 ;
        RECT 1257.970 999.870 1259.320 1000.000 ;
        RECT 1259.640 1000.010 1259.780 1012.870 ;
        RECT 1262.340 1011.510 1262.600 1011.830 ;
        RECT 1262.400 1000.010 1262.540 1011.510 ;
        RECT 1265.620 1000.010 1265.760 1012.870 ;
        RECT 1267.920 1000.010 1268.060 1020.350 ;
        RECT 1259.640 1000.000 1259.940 1000.010 ;
        RECT 1262.240 1000.000 1262.540 1000.010 ;
        RECT 1264.540 1000.000 1265.760 1000.010 ;
        RECT 1266.380 1000.000 1268.060 1000.010 ;
        RECT 1259.640 999.870 1260.090 1000.000 ;
      LAYER met2 ;
        RECT 1247.490 995.720 1248.950 998.810 ;
      LAYER met2 ;
        RECT 1249.230 996.000 1249.510 999.870 ;
      LAYER met2 ;
        RECT 1249.790 995.720 1250.790 998.810 ;
      LAYER met2 ;
        RECT 1251.070 996.000 1251.350 999.870 ;
      LAYER met2 ;
        RECT 1251.630 995.720 1253.090 998.810 ;
      LAYER met2 ;
        RECT 1253.370 996.000 1253.650 999.870 ;
      LAYER met2 ;
        RECT 1253.930 995.720 1255.390 998.810 ;
      LAYER met2 ;
        RECT 1255.670 996.000 1255.950 999.870 ;
      LAYER met2 ;
        RECT 1256.230 995.720 1257.690 998.810 ;
      LAYER met2 ;
        RECT 1257.970 996.000 1258.250 999.870 ;
      LAYER met2 ;
        RECT 1258.530 995.720 1259.530 998.810 ;
      LAYER met2 ;
        RECT 1259.810 996.000 1260.090 999.870 ;
        RECT 1262.110 999.870 1262.540 1000.000 ;
        RECT 1264.410 999.870 1265.760 1000.000 ;
        RECT 1266.250 999.870 1268.060 1000.000 ;
        RECT 1268.380 1000.010 1268.520 1694.230 ;
        RECT 1268.780 1689.130 1269.040 1689.450 ;
        RECT 1268.840 1013.190 1268.980 1689.130 ;
        RECT 1272.520 1684.350 1272.660 1700.000 ;
        RECT 1287.240 1689.110 1287.380 1700.000 ;
        RECT 1288.560 1694.570 1288.820 1694.890 ;
        RECT 1287.180 1688.790 1287.440 1689.110 ;
        RECT 1276.600 1686.410 1276.860 1686.730 ;
        RECT 1272.460 1684.030 1272.720 1684.350 ;
        RECT 1276.660 1021.770 1276.800 1686.410 ;
        RECT 1288.620 1656.470 1288.760 1694.570 ;
        RECT 1301.040 1689.790 1301.180 1700.000 ;
        RECT 1310.640 1695.590 1310.900 1695.910 ;
        RECT 1300.980 1689.470 1301.240 1689.790 ;
        RECT 1293.620 1688.450 1293.880 1688.770 ;
        RECT 1291.320 1684.030 1291.580 1684.350 ;
        RECT 1288.560 1656.150 1288.820 1656.470 ;
        RECT 1289.020 1655.470 1289.280 1655.790 ;
        RECT 1289.080 1595.270 1289.220 1655.470 ;
        RECT 1289.020 1594.950 1289.280 1595.270 ;
        RECT 1289.020 1593.590 1289.280 1593.910 ;
        RECT 1289.080 1587.110 1289.220 1593.590 ;
        RECT 1289.020 1586.790 1289.280 1587.110 ;
        RECT 1290.400 1586.790 1290.660 1587.110 ;
        RECT 1290.460 1558.890 1290.600 1586.790 ;
        RECT 1289.020 1558.570 1289.280 1558.890 ;
        RECT 1290.400 1558.570 1290.660 1558.890 ;
        RECT 1289.080 1538.830 1289.220 1558.570 ;
        RECT 1288.560 1538.510 1288.820 1538.830 ;
        RECT 1289.020 1538.510 1289.280 1538.830 ;
        RECT 1288.620 1490.890 1288.760 1538.510 ;
        RECT 1288.560 1490.570 1288.820 1490.890 ;
        RECT 1289.480 1490.570 1289.740 1490.890 ;
        RECT 1289.540 1442.270 1289.680 1490.570 ;
        RECT 1289.020 1441.950 1289.280 1442.270 ;
        RECT 1289.480 1441.950 1289.740 1442.270 ;
        RECT 1289.080 1414.730 1289.220 1441.950 ;
        RECT 1289.020 1414.410 1289.280 1414.730 ;
        RECT 1289.940 1414.410 1290.200 1414.730 ;
        RECT 1290.000 1414.130 1290.140 1414.410 ;
        RECT 1289.540 1413.990 1290.140 1414.130 ;
        RECT 1289.540 1366.530 1289.680 1413.990 ;
        RECT 1289.080 1366.390 1289.680 1366.530 ;
        RECT 1289.080 1352.510 1289.220 1366.390 ;
        RECT 1289.020 1352.190 1289.280 1352.510 ;
        RECT 1289.940 1352.190 1290.200 1352.510 ;
        RECT 1290.000 1317.830 1290.140 1352.190 ;
        RECT 1289.020 1317.510 1289.280 1317.830 ;
        RECT 1289.940 1317.510 1290.200 1317.830 ;
        RECT 1289.080 1304.230 1289.220 1317.510 ;
        RECT 1289.020 1303.910 1289.280 1304.230 ;
        RECT 1290.400 1303.910 1290.660 1304.230 ;
        RECT 1290.460 1269.210 1290.600 1303.910 ;
        RECT 1289.020 1268.890 1289.280 1269.210 ;
        RECT 1290.400 1268.890 1290.660 1269.210 ;
        RECT 1289.080 1255.950 1289.220 1268.890 ;
        RECT 1287.640 1255.630 1287.900 1255.950 ;
        RECT 1289.020 1255.630 1289.280 1255.950 ;
        RECT 1287.700 1207.670 1287.840 1255.630 ;
        RECT 1287.640 1207.350 1287.900 1207.670 ;
        RECT 1288.560 1207.350 1288.820 1207.670 ;
        RECT 1288.620 1173.330 1288.760 1207.350 ;
        RECT 1288.560 1173.010 1288.820 1173.330 ;
        RECT 1289.020 1172.330 1289.280 1172.650 ;
        RECT 1289.080 1159.130 1289.220 1172.330 ;
        RECT 1288.620 1158.990 1289.220 1159.130 ;
        RECT 1288.620 1125.050 1288.760 1158.990 ;
        RECT 1288.560 1124.730 1288.820 1125.050 ;
        RECT 1289.020 1124.390 1289.280 1124.710 ;
        RECT 1289.080 1111.110 1289.220 1124.390 ;
        RECT 1288.560 1110.790 1288.820 1111.110 ;
        RECT 1289.020 1110.790 1289.280 1111.110 ;
        RECT 1288.620 1076.770 1288.760 1110.790 ;
        RECT 1288.560 1076.450 1288.820 1076.770 ;
        RECT 1289.020 1075.770 1289.280 1076.090 ;
        RECT 1289.080 1062.570 1289.220 1075.770 ;
        RECT 1288.620 1062.430 1289.220 1062.570 ;
        RECT 1288.620 1028.490 1288.760 1062.430 ;
        RECT 1288.560 1028.170 1288.820 1028.490 ;
        RECT 1289.020 1027.830 1289.280 1028.150 ;
        RECT 1276.660 1021.630 1280.940 1021.770 ;
        RECT 1278.900 1020.690 1279.160 1021.010 ;
        RECT 1269.240 1013.550 1269.500 1013.870 ;
        RECT 1268.780 1012.870 1269.040 1013.190 ;
        RECT 1269.300 1008.770 1269.440 1013.550 ;
        RECT 1270.160 1011.850 1270.420 1012.170 ;
        RECT 1276.140 1011.850 1276.400 1012.170 ;
        RECT 1269.240 1008.450 1269.500 1008.770 ;
        RECT 1270.220 1000.010 1270.360 1011.850 ;
        RECT 1274.300 1009.470 1274.560 1009.790 ;
        RECT 1274.360 1000.010 1274.500 1009.470 ;
        RECT 1276.200 1000.010 1276.340 1011.850 ;
        RECT 1278.960 1000.010 1279.100 1020.690 ;
        RECT 1279.820 1009.130 1280.080 1009.450 ;
        RECT 1279.880 1000.010 1280.020 1009.130 ;
        RECT 1268.380 1000.000 1268.680 1000.010 ;
        RECT 1270.220 1000.000 1270.980 1000.010 ;
        RECT 1273.280 1000.000 1274.500 1000.010 ;
        RECT 1275.120 1000.000 1276.340 1000.010 ;
        RECT 1277.420 1000.000 1279.100 1000.010 ;
        RECT 1279.720 1000.000 1280.020 1000.010 ;
        RECT 1268.380 999.870 1268.830 1000.000 ;
        RECT 1270.220 999.870 1271.130 1000.000 ;
      LAYER met2 ;
        RECT 1260.370 995.720 1261.830 998.810 ;
      LAYER met2 ;
        RECT 1262.110 996.000 1262.390 999.870 ;
      LAYER met2 ;
        RECT 1262.670 995.720 1264.130 998.810 ;
      LAYER met2 ;
        RECT 1264.410 996.000 1264.690 999.870 ;
      LAYER met2 ;
        RECT 1264.970 995.720 1265.970 998.810 ;
      LAYER met2 ;
        RECT 1266.250 996.000 1266.530 999.870 ;
      LAYER met2 ;
        RECT 1266.810 995.720 1268.270 998.810 ;
      LAYER met2 ;
        RECT 1268.550 996.000 1268.830 999.870 ;
      LAYER met2 ;
        RECT 1269.110 995.720 1270.570 998.810 ;
      LAYER met2 ;
        RECT 1270.850 996.000 1271.130 999.870 ;
        RECT 1273.150 999.870 1274.500 1000.000 ;
        RECT 1274.990 999.870 1276.340 1000.000 ;
        RECT 1277.290 999.870 1279.100 1000.000 ;
        RECT 1279.590 999.870 1280.020 1000.000 ;
        RECT 1280.800 1000.010 1280.940 1021.630 ;
        RECT 1285.800 1019.330 1286.060 1019.650 ;
        RECT 1284.880 1013.890 1285.140 1014.210 ;
        RECT 1284.940 1012.510 1285.080 1013.890 ;
        RECT 1284.880 1012.190 1285.140 1012.510 ;
        RECT 1285.330 1010.635 1285.610 1011.005 ;
        RECT 1285.400 1000.010 1285.540 1010.635 ;
        RECT 1280.800 1000.000 1282.020 1000.010 ;
        RECT 1283.860 1000.000 1285.540 1000.010 ;
        RECT 1280.800 999.870 1282.170 1000.000 ;
      LAYER met2 ;
        RECT 1271.410 995.720 1272.870 998.810 ;
      LAYER met2 ;
        RECT 1273.150 996.000 1273.430 999.870 ;
      LAYER met2 ;
        RECT 1273.710 995.720 1274.710 998.810 ;
      LAYER met2 ;
        RECT 1274.990 996.000 1275.270 999.870 ;
      LAYER met2 ;
        RECT 1275.550 995.720 1277.010 998.810 ;
      LAYER met2 ;
        RECT 1277.290 996.000 1277.570 999.870 ;
      LAYER met2 ;
        RECT 1277.850 995.720 1279.310 998.810 ;
      LAYER met2 ;
        RECT 1279.590 996.000 1279.870 999.870 ;
      LAYER met2 ;
        RECT 1280.150 995.720 1281.610 998.810 ;
      LAYER met2 ;
        RECT 1281.890 996.000 1282.170 999.870 ;
        RECT 1283.730 999.870 1285.540 1000.000 ;
        RECT 1285.860 1000.010 1286.000 1019.330 ;
        RECT 1289.080 1014.550 1289.220 1027.830 ;
        RECT 1288.560 1014.230 1288.820 1014.550 ;
        RECT 1289.020 1014.230 1289.280 1014.550 ;
        RECT 1288.620 1001.370 1288.760 1014.230 ;
        RECT 1289.540 1011.490 1291.060 1011.570 ;
        RECT 1289.480 1011.430 1291.060 1011.490 ;
        RECT 1289.480 1011.170 1289.740 1011.430 ;
        RECT 1290.400 1010.830 1290.660 1011.150 ;
        RECT 1288.390 1001.230 1288.760 1001.370 ;
        RECT 1285.860 1000.000 1286.160 1000.010 ;
        RECT 1288.390 1000.000 1288.530 1001.230 ;
        RECT 1290.460 1000.010 1290.600 1010.830 ;
        RECT 1290.300 1000.000 1290.600 1000.010 ;
        RECT 1285.860 999.870 1286.310 1000.000 ;
      LAYER met2 ;
        RECT 1282.450 995.720 1283.450 998.810 ;
      LAYER met2 ;
        RECT 1283.730 996.000 1284.010 999.870 ;
      LAYER met2 ;
        RECT 1284.290 995.720 1285.750 998.810 ;
      LAYER met2 ;
        RECT 1286.030 996.000 1286.310 999.870 ;
      LAYER met2 ;
        RECT 1286.590 995.720 1288.050 998.810 ;
      LAYER met2 ;
        RECT 1288.330 996.000 1288.610 1000.000 ;
        RECT 1290.170 999.870 1290.600 1000.000 ;
        RECT 1290.920 1000.010 1291.060 1011.430 ;
        RECT 1291.380 1000.690 1291.520 1684.030 ;
        RECT 1292.700 1013.210 1292.960 1013.530 ;
        RECT 1292.760 1008.090 1292.900 1013.210 ;
        RECT 1293.680 1008.090 1293.820 1688.450 ;
        RECT 1301.900 1018.990 1302.160 1019.310 ;
        RECT 1300.980 1014.230 1301.240 1014.550 ;
        RECT 1294.080 1013.890 1294.340 1014.210 ;
        RECT 1292.700 1007.770 1292.960 1008.090 ;
        RECT 1293.620 1007.770 1293.880 1008.090 ;
        RECT 1294.140 1007.750 1294.280 1013.890 ;
        RECT 1294.540 1012.250 1294.800 1012.510 ;
        RECT 1294.540 1012.190 1296.120 1012.250 ;
        RECT 1294.600 1012.170 1296.120 1012.190 ;
        RECT 1294.600 1012.110 1296.180 1012.170 ;
        RECT 1295.920 1011.850 1296.180 1012.110 ;
        RECT 1297.300 1008.110 1297.560 1008.430 ;
        RECT 1300.520 1008.110 1300.780 1008.430 ;
        RECT 1294.080 1007.430 1294.340 1007.750 ;
        RECT 1291.380 1000.550 1293.820 1000.690 ;
        RECT 1293.680 1000.010 1293.820 1000.550 ;
        RECT 1297.360 1000.010 1297.500 1008.110 ;
        RECT 1300.580 1000.010 1300.720 1008.110 ;
        RECT 1290.920 1000.000 1292.600 1000.010 ;
        RECT 1293.680 1000.000 1294.900 1000.010 ;
        RECT 1297.200 1000.000 1297.500 1000.010 ;
        RECT 1299.040 1000.000 1300.720 1000.010 ;
        RECT 1290.920 999.870 1292.750 1000.000 ;
        RECT 1293.680 999.870 1295.050 1000.000 ;
      LAYER met2 ;
        RECT 1288.890 995.720 1289.890 998.810 ;
      LAYER met2 ;
        RECT 1290.170 996.000 1290.450 999.870 ;
      LAYER met2 ;
        RECT 1290.730 995.720 1292.190 998.810 ;
      LAYER met2 ;
        RECT 1292.470 996.000 1292.750 999.870 ;
      LAYER met2 ;
        RECT 1293.030 995.720 1294.490 998.810 ;
      LAYER met2 ;
        RECT 1294.770 996.000 1295.050 999.870 ;
        RECT 1297.070 999.870 1297.500 1000.000 ;
        RECT 1298.910 999.870 1300.720 1000.000 ;
        RECT 1301.040 1000.010 1301.180 1014.230 ;
        RECT 1301.960 1000.010 1302.100 1018.990 ;
        RECT 1310.700 1012.250 1310.840 1695.590 ;
        RECT 1315.760 1689.450 1315.900 1700.000 ;
        RECT 1315.700 1689.130 1315.960 1689.450 ;
        RECT 1313.860 1018.650 1314.120 1018.970 ;
        RECT 1308.860 1012.110 1310.840 1012.250 ;
        RECT 1304.200 1008.790 1304.460 1009.110 ;
        RECT 1304.260 1000.010 1304.400 1008.790 ;
        RECT 1308.860 1000.010 1309.000 1012.110 ;
        RECT 1309.720 1011.170 1309.980 1011.490 ;
        RECT 1301.040 1000.000 1301.340 1000.010 ;
        RECT 1301.960 1000.000 1303.640 1000.010 ;
        RECT 1304.260 1000.000 1305.940 1000.010 ;
        RECT 1307.780 1000.000 1309.000 1000.010 ;
        RECT 1301.040 999.870 1301.490 1000.000 ;
        RECT 1301.960 999.870 1303.790 1000.000 ;
        RECT 1304.260 999.870 1306.090 1000.000 ;
      LAYER met2 ;
        RECT 1295.330 995.720 1296.790 998.810 ;
      LAYER met2 ;
        RECT 1297.070 996.000 1297.350 999.870 ;
      LAYER met2 ;
        RECT 1297.630 995.720 1298.630 998.810 ;
      LAYER met2 ;
        RECT 1298.910 996.000 1299.190 999.870 ;
      LAYER met2 ;
        RECT 1299.470 995.720 1300.930 998.810 ;
      LAYER met2 ;
        RECT 1301.210 996.000 1301.490 999.870 ;
      LAYER met2 ;
        RECT 1301.770 995.720 1303.230 998.810 ;
      LAYER met2 ;
        RECT 1303.510 996.000 1303.790 999.870 ;
      LAYER met2 ;
        RECT 1304.070 995.720 1305.530 998.810 ;
      LAYER met2 ;
        RECT 1305.810 996.000 1306.090 999.870 ;
        RECT 1307.650 999.870 1309.000 1000.000 ;
        RECT 1309.780 1000.010 1309.920 1011.170 ;
        RECT 1313.390 1007.915 1313.670 1008.285 ;
        RECT 1313.460 1000.010 1313.600 1007.915 ;
        RECT 1309.780 1000.000 1310.080 1000.010 ;
        RECT 1312.380 1000.000 1313.600 1000.010 ;
        RECT 1309.780 999.870 1310.230 1000.000 ;
      LAYER met2 ;
        RECT 1306.370 995.720 1307.370 998.810 ;
      LAYER met2 ;
        RECT 1307.650 996.000 1307.930 999.870 ;
      LAYER met2 ;
        RECT 1308.210 995.720 1309.670 998.810 ;
      LAYER met2 ;
        RECT 1309.950 996.000 1310.230 999.870 ;
        RECT 1312.250 999.870 1313.600 1000.000 ;
        RECT 1313.920 1000.010 1314.060 1018.650 ;
        RECT 1314.780 1018.310 1315.040 1018.630 ;
        RECT 1314.840 1000.010 1314.980 1018.310 ;
        RECT 1326.280 1017.970 1326.540 1018.290 ;
        RECT 1320.300 1010.830 1320.560 1011.150 ;
        RECT 1320.360 1009.450 1320.500 1010.830 ;
        RECT 1320.300 1009.130 1320.560 1009.450 ;
        RECT 1318.000 1008.450 1318.260 1008.770 ;
        RECT 1325.820 1008.450 1326.080 1008.770 ;
        RECT 1318.060 1000.010 1318.200 1008.450 ;
        RECT 1319.380 1007.770 1319.640 1008.090 ;
        RECT 1319.440 1000.010 1319.580 1007.770 ;
        RECT 1324.440 1007.430 1324.700 1007.750 ;
        RECT 1324.500 1000.010 1324.640 1007.430 ;
        RECT 1325.880 1000.010 1326.020 1008.450 ;
        RECT 1313.920 1000.000 1314.220 1000.010 ;
        RECT 1314.840 1000.000 1316.520 1000.010 ;
        RECT 1318.060 1000.000 1318.820 1000.010 ;
        RECT 1319.440 1000.000 1321.120 1000.010 ;
        RECT 1322.960 1000.000 1324.640 1000.010 ;
        RECT 1325.260 1000.000 1326.020 1000.010 ;
        RECT 1313.920 999.870 1314.370 1000.000 ;
        RECT 1314.840 999.870 1316.670 1000.000 ;
        RECT 1318.060 999.870 1318.970 1000.000 ;
        RECT 1319.440 999.870 1321.270 1000.000 ;
      LAYER met2 ;
        RECT 1310.510 995.720 1311.970 998.810 ;
      LAYER met2 ;
        RECT 1312.250 996.000 1312.530 999.870 ;
      LAYER met2 ;
        RECT 1312.810 995.720 1313.810 998.810 ;
      LAYER met2 ;
        RECT 1314.090 996.000 1314.370 999.870 ;
      LAYER met2 ;
        RECT 1314.650 995.720 1316.110 998.810 ;
      LAYER met2 ;
        RECT 1316.390 996.000 1316.670 999.870 ;
      LAYER met2 ;
        RECT 1316.950 995.720 1318.410 998.810 ;
      LAYER met2 ;
        RECT 1318.690 996.000 1318.970 999.870 ;
      LAYER met2 ;
        RECT 1319.250 995.720 1320.710 998.810 ;
      LAYER met2 ;
        RECT 1320.990 996.000 1321.270 999.870 ;
        RECT 1322.830 999.870 1324.640 1000.000 ;
        RECT 1325.130 999.870 1326.020 1000.000 ;
        RECT 1326.340 1000.010 1326.480 1017.970 ;
        RECT 1331.400 1009.110 1331.540 1700.270 ;
        RECT 1331.340 1008.790 1331.600 1009.110 ;
        RECT 1330.870 1007.235 1331.150 1007.605 ;
        RECT 1330.940 1000.010 1331.080 1007.235 ;
        RECT 1331.860 1000.690 1332.000 2051.910 ;
        RECT 1332.260 2049.870 1332.520 2050.190 ;
        RECT 1332.320 1006.050 1332.460 2049.870 ;
        RECT 1332.780 1007.750 1332.920 2053.950 ;
        RECT 1338.700 2053.610 1338.960 2053.930 ;
        RECT 1333.180 2053.270 1333.440 2053.590 ;
        RECT 1333.240 1013.530 1333.380 2053.270 ;
        RECT 1335.020 2052.930 1335.280 2053.250 ;
        RECT 1334.560 2052.590 1334.820 2052.910 ;
        RECT 1334.100 2051.570 1334.360 2051.890 ;
        RECT 1333.640 2051.230 1333.900 2051.550 ;
        RECT 1333.700 1014.210 1333.840 2051.230 ;
        RECT 1333.640 1013.890 1333.900 1014.210 ;
        RECT 1333.180 1013.210 1333.440 1013.530 ;
        RECT 1334.160 1011.830 1334.300 2051.570 ;
        RECT 1334.100 1011.510 1334.360 1011.830 ;
        RECT 1334.620 1009.790 1334.760 2052.590 ;
        RECT 1334.560 1009.470 1334.820 1009.790 ;
        RECT 1335.080 1008.090 1335.220 2052.930 ;
        RECT 1335.480 2052.250 1335.740 2052.570 ;
        RECT 1335.540 1008.430 1335.680 2052.250 ;
        RECT 1338.240 2050.890 1338.500 2051.210 ;
        RECT 1337.780 2049.530 1338.040 2049.850 ;
        RECT 1335.930 1997.995 1336.210 1998.365 ;
        RECT 1336.000 1008.770 1336.140 1997.995 ;
        RECT 1336.390 1787.195 1336.670 1787.565 ;
        RECT 1335.940 1008.450 1336.200 1008.770 ;
        RECT 1335.480 1008.110 1335.740 1008.430 ;
        RECT 1335.020 1007.770 1335.280 1008.090 ;
        RECT 1336.460 1007.750 1336.600 1787.195 ;
        RECT 1336.850 1766.795 1337.130 1767.165 ;
        RECT 1336.920 1010.470 1337.060 1766.795 ;
        RECT 1337.310 1745.035 1337.590 1745.405 ;
        RECT 1336.860 1010.150 1337.120 1010.470 ;
        RECT 1337.380 1009.450 1337.520 1745.035 ;
        RECT 1337.840 1694.890 1337.980 2049.530 ;
        RECT 1337.780 1694.570 1338.040 1694.890 ;
        RECT 1338.300 1693.870 1338.440 2050.890 ;
        RECT 1338.240 1693.550 1338.500 1693.870 ;
        RECT 1337.780 1017.630 1338.040 1017.950 ;
        RECT 1337.320 1009.130 1337.580 1009.450 ;
        RECT 1332.720 1007.430 1332.980 1007.750 ;
        RECT 1333.180 1007.430 1333.440 1007.750 ;
        RECT 1336.400 1007.430 1336.660 1007.750 ;
        RECT 1332.260 1005.730 1332.520 1006.050 ;
        RECT 1331.860 1000.610 1332.460 1000.690 ;
        RECT 1331.860 1000.550 1332.520 1000.610 ;
        RECT 1332.260 1000.290 1332.520 1000.550 ;
        RECT 1332.320 1000.135 1332.460 1000.290 ;
        RECT 1326.340 1000.000 1327.560 1000.010 ;
        RECT 1329.860 1000.000 1331.080 1000.010 ;
        RECT 1326.340 999.870 1327.710 1000.000 ;
      LAYER met2 ;
        RECT 1321.550 995.720 1322.550 998.810 ;
      LAYER met2 ;
        RECT 1322.830 996.000 1323.110 999.870 ;
      LAYER met2 ;
        RECT 1323.390 995.720 1324.850 998.810 ;
      LAYER met2 ;
        RECT 1325.130 996.000 1325.410 999.870 ;
      LAYER met2 ;
        RECT 1325.690 995.720 1327.150 998.810 ;
      LAYER met2 ;
        RECT 1327.430 996.000 1327.710 999.870 ;
        RECT 1329.730 999.870 1331.080 1000.000 ;
      LAYER met2 ;
        RECT 1327.990 995.720 1329.450 998.810 ;
      LAYER met2 ;
        RECT 1329.730 996.000 1330.010 999.870 ;
        RECT 1331.570 999.330 1331.850 1000.000 ;
        RECT 1333.240 999.330 1333.380 1007.430 ;
        RECT 1337.840 1000.690 1337.980 1017.630 ;
        RECT 1338.760 1012.850 1338.900 2053.610 ;
        RECT 1343.760 2050.550 1344.020 2050.870 ;
        RECT 1339.150 2018.395 1339.430 2018.765 ;
        RECT 1339.220 1013.870 1339.360 2018.395 ;
        RECT 1339.610 1976.235 1339.890 1976.605 ;
        RECT 1339.680 1020.330 1339.820 1976.235 ;
        RECT 1340.070 1955.835 1340.350 1956.205 ;
        RECT 1339.620 1020.010 1339.880 1020.330 ;
        RECT 1339.160 1013.550 1339.420 1013.870 ;
        RECT 1338.700 1012.530 1338.960 1012.850 ;
        RECT 1340.140 1010.130 1340.280 1955.835 ;
        RECT 1340.530 1934.075 1340.810 1934.445 ;
        RECT 1340.600 1019.990 1340.740 1934.075 ;
        RECT 1340.990 1913.675 1341.270 1914.045 ;
        RECT 1341.060 1021.010 1341.200 1913.675 ;
        RECT 1341.450 1891.915 1341.730 1892.285 ;
        RECT 1341.000 1020.690 1341.260 1021.010 ;
        RECT 1340.540 1019.670 1340.800 1019.990 ;
        RECT 1341.520 1013.190 1341.660 1891.915 ;
        RECT 1341.910 1871.515 1342.190 1871.885 ;
        RECT 1341.460 1012.870 1341.720 1013.190 ;
        RECT 1341.980 1012.510 1342.120 1871.515 ;
        RECT 1342.370 1849.755 1342.650 1850.125 ;
        RECT 1341.920 1012.190 1342.180 1012.510 ;
        RECT 1342.440 1012.170 1342.580 1849.755 ;
        RECT 1342.830 1829.355 1343.110 1829.725 ;
        RECT 1342.380 1011.850 1342.640 1012.170 ;
        RECT 1342.900 1011.150 1343.040 1829.355 ;
        RECT 1343.290 1807.595 1343.570 1807.965 ;
        RECT 1342.840 1010.830 1343.100 1011.150 ;
        RECT 1340.080 1009.810 1340.340 1010.130 ;
        RECT 1341.000 1008.110 1341.260 1008.430 ;
        RECT 1338.700 1007.770 1338.960 1008.090 ;
        RECT 1338.240 1005.730 1338.500 1006.050 ;
        RECT 1333.640 1000.290 1333.900 1000.610 ;
        RECT 1337.380 1000.550 1337.980 1000.690 ;
        RECT 1333.700 1000.010 1333.840 1000.290 ;
        RECT 1337.380 1000.010 1337.520 1000.550 ;
        RECT 1338.300 1000.010 1338.440 1005.730 ;
        RECT 1333.700 1000.000 1334.000 1000.010 ;
        RECT 1336.300 1000.000 1337.520 1000.010 ;
        RECT 1338.140 1000.000 1338.440 1000.010 ;
        RECT 1333.700 999.870 1334.150 1000.000 ;
        RECT 1331.570 999.190 1333.380 999.330 ;
      LAYER met2 ;
        RECT 1330.290 995.720 1331.290 998.810 ;
      LAYER met2 ;
        RECT 1331.570 996.000 1331.850 999.190 ;
      LAYER met2 ;
        RECT 1332.130 995.720 1333.590 998.810 ;
      LAYER met2 ;
        RECT 1333.870 996.000 1334.150 999.870 ;
        RECT 1336.170 999.870 1337.520 1000.000 ;
        RECT 1338.010 999.870 1338.440 1000.000 ;
        RECT 1338.760 1000.010 1338.900 1007.770 ;
        RECT 1341.060 1000.010 1341.200 1008.110 ;
        RECT 1343.360 1000.010 1343.500 1807.595 ;
        RECT 1343.820 1694.210 1343.960 2050.550 ;
        RECT 1344.220 2050.210 1344.480 2050.530 ;
        RECT 1344.280 1694.550 1344.420 2050.210 ;
        RECT 1344.680 2049.190 1344.940 2049.510 ;
        RECT 1344.740 1695.910 1344.880 2049.190 ;
        RECT 1345.130 1724.635 1345.410 1725.005 ;
        RECT 1344.680 1695.590 1344.940 1695.910 ;
        RECT 1344.220 1694.230 1344.480 1694.550 ;
        RECT 1343.760 1693.890 1344.020 1694.210 ;
        RECT 1345.200 1020.670 1345.340 1724.635 ;
        RECT 1345.140 1020.350 1345.400 1020.670 ;
        RECT 1347.440 1010.490 1347.700 1010.810 ;
        RECT 1345.600 1008.790 1345.860 1009.110 ;
        RECT 1345.660 1000.010 1345.800 1008.790 ;
        RECT 1347.500 1000.010 1347.640 1010.490 ;
        RECT 1352.100 1000.010 1352.240 2917.890 ;
        RECT 1431.620 2917.550 1431.880 2917.870 ;
        RECT 1406.780 2914.830 1407.040 2915.150 ;
        RECT 1372.730 2912.595 1373.010 2912.965 ;
        RECT 1362.620 2849.550 1362.880 2849.870 ;
        RECT 1358.940 1017.970 1359.200 1018.290 ;
        RECT 1357.100 1012.530 1357.360 1012.850 ;
        RECT 1354.800 1010.830 1355.060 1011.150 ;
        RECT 1354.860 1000.010 1355.000 1010.830 ;
        RECT 1357.160 1000.010 1357.300 1012.530 ;
        RECT 1359.000 1000.010 1359.140 1017.970 ;
        RECT 1361.240 1013.890 1361.500 1014.210 ;
        RECT 1361.300 1000.010 1361.440 1013.890 ;
        RECT 1362.680 1012.850 1362.820 2849.550 ;
        RECT 1365.840 2780.870 1366.100 2781.190 ;
        RECT 1365.900 1014.210 1366.040 2780.870 ;
        RECT 1365.840 1013.890 1366.100 1014.210 ;
        RECT 1362.620 1012.530 1362.880 1012.850 ;
        RECT 1372.800 1012.510 1372.940 2912.595 ;
        RECT 1400.340 2608.150 1400.600 2608.470 ;
        RECT 1397.120 2594.550 1397.380 2594.870 ;
        RECT 1386.540 2486.090 1386.800 2486.410 ;
        RECT 1383.320 2485.750 1383.580 2486.070 ;
        RECT 1369.980 1012.190 1370.240 1012.510 ;
        RECT 1372.740 1012.190 1373.000 1012.510 ;
        RECT 1368.140 1008.110 1368.400 1008.430 ;
        RECT 1368.200 1000.010 1368.340 1008.110 ;
        RECT 1370.040 1000.010 1370.180 1012.190 ;
        RECT 1376.420 1011.850 1376.680 1012.170 ;
        RECT 1376.480 1000.010 1376.620 1011.850 ;
        RECT 1378.720 1011.510 1378.980 1011.830 ;
        RECT 1378.780 1000.010 1378.920 1011.510 ;
        RECT 1383.380 1008.430 1383.520 2485.750 ;
        RECT 1386.600 1012.510 1386.740 2486.090 ;
        RECT 1397.180 1012.510 1397.320 2594.550 ;
        RECT 1384.700 1012.190 1384.960 1012.510 ;
        RECT 1386.540 1012.190 1386.800 1012.510 ;
        RECT 1393.440 1012.190 1393.700 1012.510 ;
        RECT 1397.120 1012.190 1397.380 1012.510 ;
        RECT 1383.320 1008.110 1383.580 1008.430 ;
        RECT 1384.760 1000.010 1384.900 1012.190 ;
        RECT 1386.540 1011.170 1386.800 1011.490 ;
        RECT 1386.600 1000.010 1386.740 1011.170 ;
        RECT 1393.500 1000.010 1393.640 1012.190 ;
        RECT 1400.400 1008.090 1400.540 2608.150 ;
        RECT 1402.640 1017.630 1402.900 1017.950 ;
        RECT 1396.200 1007.770 1396.460 1008.090 ;
        RECT 1400.340 1007.770 1400.600 1008.090 ;
        RECT 1396.260 1000.010 1396.400 1007.770 ;
        RECT 1402.700 1000.010 1402.840 1017.630 ;
        RECT 1406.840 1012.510 1406.980 2914.830 ;
        RECT 1424.720 2580.610 1424.980 2580.930 ;
        RECT 1420.580 2488.810 1420.840 2489.130 ;
        RECT 1404.940 1012.190 1405.200 1012.510 ;
        RECT 1406.780 1012.190 1407.040 1012.510 ;
        RECT 1405.000 1000.010 1405.140 1012.190 ;
        RECT 1417.820 1010.490 1418.080 1010.810 ;
        RECT 1413.220 1007.770 1413.480 1008.090 ;
        RECT 1411.380 1007.430 1411.640 1007.750 ;
        RECT 1411.440 1000.010 1411.580 1007.430 ;
        RECT 1413.280 1000.010 1413.420 1007.770 ;
        RECT 1417.880 1000.010 1418.020 1010.490 ;
        RECT 1420.640 1000.690 1420.780 2488.810 ;
        RECT 1421.040 2488.130 1421.300 2488.450 ;
        RECT 1420.180 1000.550 1420.780 1000.690 ;
        RECT 1420.180 1000.010 1420.320 1000.550 ;
        RECT 1421.100 1000.010 1421.240 2488.130 ;
        RECT 1424.780 1007.750 1424.920 2580.610 ;
        RECT 1427.940 2486.770 1428.200 2487.090 ;
        RECT 1424.720 1007.430 1424.980 1007.750 ;
        RECT 1428.000 1000.010 1428.140 2486.770 ;
        RECT 1431.680 1011.830 1431.820 2917.550 ;
        RECT 1459.220 2915.850 1459.480 2916.170 ;
        RECT 1455.540 2913.810 1455.800 2914.130 ;
        RECT 1438.520 2912.110 1438.780 2912.430 ;
        RECT 1434.380 2691.110 1434.640 2691.430 ;
        RECT 1432.080 2484.730 1432.340 2485.050 ;
        RECT 1432.140 1012.170 1432.280 2484.730 ;
        RECT 1432.080 1011.850 1432.340 1012.170 ;
        RECT 1431.620 1011.510 1431.880 1011.830 ;
        RECT 1431.160 1007.430 1431.420 1007.750 ;
        RECT 1431.220 1000.010 1431.360 1007.430 ;
        RECT 1434.440 1000.010 1434.580 2691.110 ;
        RECT 1434.840 1018.650 1435.100 1018.970 ;
        RECT 1434.900 1007.750 1435.040 1018.650 ;
        RECT 1437.600 1018.310 1437.860 1018.630 ;
        RECT 1434.840 1007.430 1435.100 1007.750 ;
        RECT 1437.660 1000.010 1437.800 1018.310 ;
        RECT 1438.580 1008.090 1438.720 2912.110 ;
        RECT 1455.080 2488.470 1455.340 2488.790 ;
        RECT 1442.660 2485.410 1442.920 2485.730 ;
        RECT 1442.720 2463.485 1442.860 2485.410 ;
        RECT 1441.730 2463.115 1442.010 2463.485 ;
        RECT 1442.650 2463.115 1442.930 2463.485 ;
        RECT 1441.800 2429.630 1441.940 2463.115 ;
        RECT 1441.740 2429.310 1442.000 2429.630 ;
        RECT 1441.280 2428.290 1441.540 2428.610 ;
        RECT 1441.340 2415.010 1441.480 2428.290 ;
        RECT 1441.280 2414.690 1441.540 2415.010 ;
        RECT 1441.740 2414.690 1442.000 2415.010 ;
        RECT 1441.800 2380.670 1441.940 2414.690 ;
        RECT 1441.740 2380.350 1442.000 2380.670 ;
        RECT 1441.280 2380.010 1441.540 2380.330 ;
        RECT 1441.340 2366.810 1441.480 2380.010 ;
        RECT 1441.340 2366.670 1441.940 2366.810 ;
        RECT 1441.800 2342.590 1441.940 2366.670 ;
        RECT 1440.360 2342.270 1440.620 2342.590 ;
        RECT 1441.740 2342.270 1442.000 2342.590 ;
        RECT 1440.420 2319.130 1440.560 2342.270 ;
        RECT 1440.360 2318.810 1440.620 2319.130 ;
        RECT 1441.280 2318.810 1441.540 2319.130 ;
        RECT 1441.340 2318.450 1441.480 2318.810 ;
        RECT 1441.280 2318.130 1441.540 2318.450 ;
        RECT 1441.740 2318.130 1442.000 2318.450 ;
        RECT 1441.800 2284.110 1441.940 2318.130 ;
        RECT 1441.740 2283.790 1442.000 2284.110 ;
        RECT 1441.280 2283.450 1441.540 2283.770 ;
        RECT 1441.340 2270.250 1441.480 2283.450 ;
        RECT 1441.340 2270.110 1441.940 2270.250 ;
        RECT 1441.800 2246.030 1441.940 2270.110 ;
        RECT 1440.360 2245.710 1440.620 2246.030 ;
        RECT 1441.740 2245.710 1442.000 2246.030 ;
        RECT 1440.420 2222.570 1440.560 2245.710 ;
        RECT 1440.360 2222.250 1440.620 2222.570 ;
        RECT 1441.280 2222.250 1441.540 2222.570 ;
        RECT 1441.340 2221.890 1441.480 2222.250 ;
        RECT 1441.280 2221.570 1441.540 2221.890 ;
        RECT 1441.740 2221.570 1442.000 2221.890 ;
        RECT 1441.800 2187.550 1441.940 2221.570 ;
        RECT 1441.740 2187.230 1442.000 2187.550 ;
        RECT 1441.280 2186.890 1441.540 2187.210 ;
        RECT 1441.340 2173.690 1441.480 2186.890 ;
        RECT 1441.340 2173.550 1441.940 2173.690 ;
        RECT 1441.800 2149.470 1441.940 2173.550 ;
        RECT 1440.360 2149.150 1440.620 2149.470 ;
        RECT 1441.740 2149.150 1442.000 2149.470 ;
        RECT 1440.420 2126.010 1440.560 2149.150 ;
        RECT 1440.360 2125.690 1440.620 2126.010 ;
        RECT 1441.280 2125.690 1441.540 2126.010 ;
        RECT 1441.340 2125.330 1441.480 2125.690 ;
        RECT 1440.360 2125.010 1440.620 2125.330 ;
        RECT 1441.280 2125.010 1441.540 2125.330 ;
        RECT 1440.420 2090.845 1440.560 2125.010 ;
        RECT 1439.430 2090.475 1439.710 2090.845 ;
        RECT 1440.350 2090.475 1440.630 2090.845 ;
        RECT 1439.500 2042.710 1439.640 2090.475 ;
        RECT 1439.440 2042.390 1439.700 2042.710 ;
        RECT 1439.900 2042.565 1440.160 2042.710 ;
        RECT 1439.890 2042.195 1440.170 2042.565 ;
        RECT 1441.730 2042.195 1442.010 2042.565 ;
        RECT 1441.800 1994.090 1441.940 2042.195 ;
        RECT 1441.740 1993.770 1442.000 1994.090 ;
        RECT 1442.660 1993.770 1442.920 1994.090 ;
        RECT 1442.720 1946.005 1442.860 1993.770 ;
        RECT 1441.730 1945.635 1442.010 1946.005 ;
        RECT 1442.650 1945.635 1442.930 1946.005 ;
        RECT 1441.800 1897.530 1441.940 1945.635 ;
        RECT 1441.740 1897.210 1442.000 1897.530 ;
        RECT 1442.660 1897.210 1442.920 1897.530 ;
        RECT 1442.720 1849.445 1442.860 1897.210 ;
        RECT 1441.730 1849.075 1442.010 1849.445 ;
        RECT 1442.650 1849.075 1442.930 1849.445 ;
        RECT 1441.800 1663.125 1441.940 1849.075 ;
        RECT 1441.730 1662.755 1442.010 1663.125 ;
        RECT 1443.110 1662.755 1443.390 1663.125 ;
        RECT 1443.180 1642.530 1443.320 1662.755 ;
        RECT 1441.740 1642.210 1442.000 1642.530 ;
        RECT 1443.120 1642.210 1443.380 1642.530 ;
        RECT 1441.800 1618.050 1441.940 1642.210 ;
        RECT 1441.740 1617.730 1442.000 1618.050 ;
        RECT 1442.660 1617.730 1442.920 1618.050 ;
        RECT 1442.720 1594.250 1442.860 1617.730 ;
        RECT 1441.740 1593.930 1442.000 1594.250 ;
        RECT 1442.660 1593.930 1442.920 1594.250 ;
        RECT 1441.800 1569.770 1441.940 1593.930 ;
        RECT 1440.360 1569.450 1440.620 1569.770 ;
        RECT 1441.740 1569.450 1442.000 1569.770 ;
        RECT 1440.420 1545.970 1440.560 1569.450 ;
        RECT 1440.360 1545.650 1440.620 1545.970 ;
        RECT 1440.820 1545.650 1441.080 1545.970 ;
        RECT 1440.880 1545.290 1441.020 1545.650 ;
        RECT 1440.360 1544.970 1440.620 1545.290 ;
        RECT 1440.820 1544.970 1441.080 1545.290 ;
        RECT 1440.420 1497.690 1440.560 1544.970 ;
        RECT 1440.360 1497.370 1440.620 1497.690 ;
        RECT 1441.740 1497.370 1442.000 1497.690 ;
        RECT 1441.800 1473.210 1441.940 1497.370 ;
        RECT 1440.360 1472.890 1440.620 1473.210 ;
        RECT 1441.740 1472.890 1442.000 1473.210 ;
        RECT 1440.420 1449.410 1440.560 1472.890 ;
        RECT 1440.360 1449.090 1440.620 1449.410 ;
        RECT 1440.820 1449.090 1441.080 1449.410 ;
        RECT 1440.880 1448.730 1441.020 1449.090 ;
        RECT 1440.820 1448.410 1441.080 1448.730 ;
        RECT 1442.660 1448.410 1442.920 1448.730 ;
        RECT 1442.720 1387.190 1442.860 1448.410 ;
        RECT 1441.740 1386.870 1442.000 1387.190 ;
        RECT 1442.660 1386.870 1442.920 1387.190 ;
        RECT 1441.800 1338.765 1441.940 1386.870 ;
        RECT 1441.730 1338.395 1442.010 1338.765 ;
        RECT 1442.650 1338.395 1442.930 1338.765 ;
        RECT 1442.720 1290.485 1442.860 1338.395 ;
        RECT 1440.820 1289.970 1441.080 1290.290 ;
        RECT 1441.730 1290.115 1442.010 1290.485 ;
        RECT 1442.650 1290.115 1442.930 1290.485 ;
        RECT 1441.740 1289.970 1442.000 1290.115 ;
        RECT 1440.880 1242.350 1441.020 1289.970 ;
        RECT 1440.360 1242.030 1440.620 1242.350 ;
        RECT 1440.820 1242.030 1441.080 1242.350 ;
        RECT 1440.420 1220.930 1440.560 1242.030 ;
        RECT 1440.360 1220.610 1440.620 1220.930 ;
        RECT 1441.740 1220.610 1442.000 1220.930 ;
        RECT 1441.800 1159.245 1441.940 1220.610 ;
        RECT 1441.730 1158.875 1442.010 1159.245 ;
        RECT 1442.650 1158.875 1442.930 1159.245 ;
        RECT 1442.720 1111.110 1442.860 1158.875 ;
        RECT 1441.740 1110.790 1442.000 1111.110 ;
        RECT 1442.660 1110.790 1442.920 1111.110 ;
        RECT 1441.800 1076.850 1441.940 1110.790 ;
        RECT 1440.880 1076.710 1441.940 1076.850 ;
        RECT 1440.880 1062.830 1441.020 1076.710 ;
        RECT 1440.360 1062.510 1440.620 1062.830 ;
        RECT 1440.820 1062.510 1441.080 1062.830 ;
        RECT 1440.420 1028.570 1440.560 1062.510 ;
        RECT 1454.620 1051.970 1454.880 1052.290 ;
        RECT 1439.960 1028.430 1440.560 1028.570 ;
        RECT 1438.520 1007.770 1438.780 1008.090 ;
        RECT 1439.960 1000.010 1440.100 1028.430 ;
        RECT 1452.780 1013.890 1453.040 1014.210 ;
        RECT 1446.340 1013.550 1446.600 1013.870 ;
        RECT 1444.040 1012.870 1444.300 1013.190 ;
        RECT 1444.100 1000.010 1444.240 1012.870 ;
        RECT 1446.400 1000.010 1446.540 1013.550 ;
        RECT 1447.720 1010.150 1447.980 1010.470 ;
        RECT 1447.780 1000.010 1447.920 1010.150 ;
        RECT 1452.840 1000.010 1452.980 1013.890 ;
        RECT 1454.680 1000.690 1454.820 1051.970 ;
        RECT 1455.140 1014.210 1455.280 2488.470 ;
        RECT 1455.600 1052.290 1455.740 2913.810 ;
        RECT 1455.540 1051.970 1455.800 1052.290 ;
        RECT 1455.080 1013.890 1455.340 1014.210 ;
        RECT 1456.920 1013.890 1457.180 1014.210 ;
        RECT 1454.680 1000.550 1455.280 1000.690 ;
        RECT 1455.140 1000.010 1455.280 1000.550 ;
        RECT 1456.980 1000.010 1457.120 1013.890 ;
        RECT 1459.280 1013.870 1459.420 2915.850 ;
        RECT 1494.640 2915.510 1494.900 2915.830 ;
        RECT 1473.020 2915.170 1473.280 2915.490 ;
        RECT 1469.340 2546.270 1469.600 2546.590 ;
        RECT 1461.520 2486.430 1461.780 2486.750 ;
        RECT 1461.060 1019.330 1461.320 1019.650 ;
        RECT 1459.220 1013.550 1459.480 1013.870 ;
        RECT 1461.120 1000.690 1461.260 1019.330 ;
        RECT 1461.580 1014.210 1461.720 2486.430 ;
        RECT 1462.440 1018.990 1462.700 1019.310 ;
        RECT 1461.520 1013.890 1461.780 1014.210 ;
        RECT 1461.120 1000.550 1461.720 1000.690 ;
        RECT 1461.580 1000.010 1461.720 1000.550 ;
        RECT 1462.500 1000.010 1462.640 1018.990 ;
        RECT 1465.660 1013.890 1465.920 1014.210 ;
        RECT 1465.720 1000.010 1465.860 1013.890 ;
        RECT 1469.400 1000.010 1469.540 2546.270 ;
        RECT 1472.100 1021.030 1472.360 1021.350 ;
        RECT 1472.160 1000.010 1472.300 1021.030 ;
        RECT 1473.080 1014.210 1473.220 2915.170 ;
        RECT 1493.260 2914.150 1493.520 2914.470 ;
        RECT 1492.340 2912.450 1492.600 2912.770 ;
        RECT 1483.590 2850.035 1483.870 2850.405 ;
        RECT 1483.660 2849.870 1483.800 2850.035 ;
        RECT 1483.600 2849.550 1483.860 2849.870 ;
        RECT 1482.210 2830.315 1482.490 2830.685 ;
        RECT 1474.400 1019.670 1474.660 1019.990 ;
        RECT 1473.020 1013.890 1473.280 1014.210 ;
        RECT 1474.460 1000.010 1474.600 1019.670 ;
        RECT 1480.840 1016.950 1481.100 1017.270 ;
        RECT 1479.000 1013.890 1479.260 1014.210 ;
        RECT 1479.060 1000.010 1479.200 1013.890 ;
        RECT 1480.900 1000.010 1481.040 1016.950 ;
        RECT 1482.280 1014.210 1482.420 2830.315 ;
        RECT 1490.030 2801.755 1490.310 2802.125 ;
        RECT 1485.430 2784.075 1485.710 2784.445 ;
        RECT 1485.500 2781.190 1485.640 2784.075 ;
        RECT 1485.440 2780.870 1485.700 2781.190 ;
        RECT 1489.570 2767.755 1489.850 2768.125 ;
        RECT 1489.110 2720.835 1489.390 2721.205 ;
        RECT 1488.650 2691.595 1488.930 2691.965 ;
        RECT 1488.720 2691.430 1488.860 2691.595 ;
        RECT 1488.660 2691.110 1488.920 2691.430 ;
        RECT 1482.670 2657.595 1482.950 2657.965 ;
        RECT 1482.220 1013.890 1482.480 1014.210 ;
        RECT 1482.740 1000.010 1482.880 2657.595 ;
        RECT 1485.430 2610.675 1485.710 2611.045 ;
        RECT 1485.500 2608.470 1485.640 2610.675 ;
        RECT 1485.440 2608.150 1485.700 2608.470 ;
        RECT 1488.650 2595.715 1488.930 2596.085 ;
        RECT 1488.720 2594.870 1488.860 2595.715 ;
        RECT 1488.660 2594.550 1488.920 2594.870 ;
        RECT 1488.650 2580.755 1488.930 2581.125 ;
        RECT 1488.660 2580.610 1488.920 2580.755 ;
        RECT 1488.650 2567.155 1488.930 2567.525 ;
        RECT 1483.590 2547.435 1483.870 2547.805 ;
        RECT 1483.660 2546.590 1483.800 2547.435 ;
        RECT 1483.600 2546.270 1483.860 2546.590 ;
        RECT 1488.720 1012.510 1488.860 2567.155 ;
        RECT 1488.660 1012.190 1488.920 1012.510 ;
        RECT 1489.180 1009.790 1489.320 2720.835 ;
        RECT 1489.640 1021.010 1489.780 2767.755 ;
        RECT 1489.580 1020.690 1489.840 1021.010 ;
        RECT 1490.100 1016.250 1490.240 2801.755 ;
        RECT 1492.400 2494.230 1492.540 2912.450 ;
        RECT 1492.800 2911.770 1493.060 2912.090 ;
        RECT 1492.340 2493.910 1492.600 2494.230 ;
        RECT 1492.860 2491.510 1493.000 2911.770 ;
        RECT 1493.320 2494.910 1493.460 2914.150 ;
        RECT 1493.720 2913.470 1493.980 2913.790 ;
        RECT 1493.260 2494.590 1493.520 2494.910 ;
        RECT 1492.800 2491.190 1493.060 2491.510 ;
        RECT 1490.040 1015.930 1490.300 1016.250 ;
        RECT 1493.780 1014.210 1493.920 2913.470 ;
        RECT 1494.180 2912.790 1494.440 2913.110 ;
        RECT 1494.240 2494.570 1494.380 2912.790 ;
        RECT 1494.700 2495.590 1494.840 2915.510 ;
        RECT 1495.100 2914.490 1495.360 2914.810 ;
        RECT 1494.640 2495.270 1494.900 2495.590 ;
        RECT 1495.160 2495.250 1495.300 2914.490 ;
        RECT 1500.620 2913.130 1500.880 2913.450 ;
        RECT 1496.940 2898.170 1497.200 2898.490 ;
        RECT 1496.470 2753.475 1496.750 2753.845 ;
        RECT 1496.010 2739.195 1496.290 2739.565 ;
        RECT 1495.550 2629.035 1495.830 2629.405 ;
        RECT 1495.100 2494.930 1495.360 2495.250 ;
        RECT 1494.180 2494.250 1494.440 2494.570 ;
        RECT 1495.100 1020.010 1495.360 1020.330 ;
        RECT 1489.580 1013.890 1489.840 1014.210 ;
        RECT 1493.720 1013.890 1493.980 1014.210 ;
        RECT 1494.640 1013.890 1494.900 1014.210 ;
        RECT 1489.120 1009.470 1489.380 1009.790 ;
        RECT 1487.740 1009.130 1488.000 1009.450 ;
        RECT 1487.800 1000.010 1487.940 1009.130 ;
        RECT 1489.640 1000.010 1489.780 1013.890 ;
        RECT 1491.880 1008.450 1492.140 1008.770 ;
        RECT 1491.940 1000.010 1492.080 1008.450 ;
        RECT 1338.760 1000.000 1340.440 1000.010 ;
        RECT 1341.060 1000.000 1342.740 1000.010 ;
        RECT 1343.360 1000.000 1345.040 1000.010 ;
        RECT 1345.660 1000.000 1346.880 1000.010 ;
        RECT 1347.500 1000.000 1349.180 1000.010 ;
        RECT 1351.480 1000.000 1352.240 1000.010 ;
        RECT 1353.320 1000.000 1355.000 1000.010 ;
        RECT 1355.620 1000.000 1357.300 1000.010 ;
        RECT 1357.920 1000.000 1359.140 1000.010 ;
        RECT 1360.220 1000.000 1361.440 1000.010 ;
        RECT 1366.660 1000.000 1368.340 1000.010 ;
        RECT 1368.960 1000.000 1370.180 1000.010 ;
        RECT 1375.400 1000.000 1376.620 1000.010 ;
        RECT 1377.240 1000.000 1378.920 1000.010 ;
        RECT 1384.140 1000.000 1384.900 1000.010 ;
        RECT 1385.980 1000.000 1386.740 1000.010 ;
        RECT 1392.880 1000.000 1393.640 1000.010 ;
        RECT 1394.720 1000.000 1396.400 1000.010 ;
        RECT 1401.160 1000.000 1402.840 1000.010 ;
        RECT 1403.460 1000.000 1405.140 1000.010 ;
        RECT 1409.900 1000.000 1411.580 1000.010 ;
        RECT 1412.200 1000.000 1413.420 1000.010 ;
        RECT 1416.800 1000.000 1418.020 1000.010 ;
        RECT 1418.640 1000.000 1420.320 1000.010 ;
        RECT 1420.940 1000.000 1421.240 1000.010 ;
        RECT 1427.380 1000.000 1428.140 1000.010 ;
        RECT 1429.680 1000.000 1431.360 1000.010 ;
        RECT 1433.820 1000.000 1434.580 1000.010 ;
        RECT 1436.120 1000.000 1437.800 1000.010 ;
        RECT 1438.420 1000.000 1440.100 1000.010 ;
        RECT 1442.560 1000.000 1444.240 1000.010 ;
        RECT 1444.860 1000.000 1446.540 1000.010 ;
        RECT 1447.160 1000.000 1447.920 1000.010 ;
        RECT 1451.300 1000.000 1452.980 1000.010 ;
        RECT 1453.600 1000.000 1455.280 1000.010 ;
        RECT 1455.900 1000.000 1457.120 1000.010 ;
        RECT 1460.040 1000.000 1461.720 1000.010 ;
        RECT 1462.340 1000.000 1462.640 1000.010 ;
        RECT 1464.640 1000.000 1465.860 1000.010 ;
        RECT 1468.780 1000.000 1469.540 1000.010 ;
        RECT 1471.080 1000.000 1472.300 1000.010 ;
        RECT 1472.920 1000.000 1474.600 1000.010 ;
        RECT 1477.520 1000.000 1479.200 1000.010 ;
        RECT 1479.820 1000.000 1481.040 1000.010 ;
        RECT 1481.660 1000.000 1482.880 1000.010 ;
        RECT 1486.260 1000.000 1487.940 1000.010 ;
        RECT 1488.560 1000.000 1489.780 1000.010 ;
        RECT 1490.400 1000.000 1492.080 1000.010 ;
        RECT 1494.700 1000.010 1494.840 1013.890 ;
        RECT 1495.160 1010.210 1495.300 1020.010 ;
        RECT 1495.620 1013.870 1495.760 2629.035 ;
        RECT 1495.560 1013.550 1495.820 1013.870 ;
        RECT 1496.080 1013.530 1496.220 2739.195 ;
        RECT 1496.020 1013.210 1496.280 1013.530 ;
        RECT 1495.160 1010.070 1495.760 1010.210 ;
        RECT 1495.620 1000.010 1495.760 1010.070 ;
        RECT 1496.540 1008.090 1496.680 2753.475 ;
        RECT 1497.000 1012.850 1497.140 2898.170 ;
        RECT 1497.400 2896.470 1497.660 2896.790 ;
        RECT 1496.940 1012.530 1497.200 1012.850 ;
        RECT 1497.460 1008.430 1497.600 2896.470 ;
        RECT 1500.680 2884.405 1500.820 2913.130 ;
        RECT 1535.180 2900.055 1535.320 2917.890 ;
        RECT 1598.600 2917.550 1598.860 2917.870 ;
        RECT 1567.320 2912.110 1567.580 2912.430 ;
        RECT 1546.160 2911.770 1546.420 2912.090 ;
        RECT 1546.220 2900.055 1546.360 2911.770 ;
        RECT 1567.380 2900.055 1567.520 2912.110 ;
        RECT 1598.660 2900.055 1598.800 2917.550 ;
        RECT 1641.840 2915.850 1642.100 2916.170 ;
        RECT 1630.800 2914.830 1631.060 2915.150 ;
        RECT 1609.640 2912.450 1609.900 2912.770 ;
        RECT 1609.700 2900.055 1609.840 2912.450 ;
        RECT 1630.860 2900.055 1631.000 2914.830 ;
        RECT 1641.900 2900.055 1642.040 2915.850 ;
        RECT 1705.320 2915.510 1705.580 2915.830 ;
        RECT 1694.280 2915.170 1694.540 2915.490 ;
        RECT 1663.000 2912.790 1663.260 2913.110 ;
        RECT 1663.060 2900.055 1663.200 2912.790 ;
        RECT 1694.340 2900.055 1694.480 2915.170 ;
        RECT 1705.380 2900.055 1705.520 2915.510 ;
        RECT 1768.800 2914.490 1769.060 2914.810 ;
        RECT 1758.680 2913.810 1758.940 2914.130 ;
        RECT 1758.740 2900.055 1758.880 2913.810 ;
        RECT 1768.860 2900.055 1769.000 2914.490 ;
        RECT 1779.840 2914.150 1780.100 2914.470 ;
        RECT 1779.900 2900.055 1780.040 2914.150 ;
        RECT 1801.000 2913.470 1801.260 2913.790 ;
        RECT 1789.960 2912.790 1790.220 2913.110 ;
        RECT 1790.020 2900.055 1790.160 2912.790 ;
        RECT 1801.060 2900.055 1801.200 2913.470 ;
        RECT 1812.040 2913.130 1812.300 2913.450 ;
        RECT 1833.200 2913.130 1833.460 2913.450 ;
        RECT 1894.380 2913.130 1894.640 2913.450 ;
        RECT 1812.100 2900.055 1812.240 2913.130 ;
        RECT 1833.260 2900.055 1833.400 2913.130 ;
        RECT 1843.310 2912.595 1843.590 2912.965 ;
        RECT 1892.080 2912.790 1892.340 2913.110 ;
        RECT 1843.380 2900.055 1843.520 2912.595 ;
        RECT 1854.360 2912.450 1854.620 2912.770 ;
        RECT 1854.420 2900.055 1854.560 2912.450 ;
        RECT 1864.480 2911.770 1864.740 2912.090 ;
        RECT 1864.540 2900.055 1864.680 2911.770 ;
        RECT 1502.850 2896.530 1503.130 2900.055 ;
        RECT 1524.930 2898.570 1525.210 2900.055 ;
        RECT 1524.140 2898.490 1525.210 2898.570 ;
        RECT 1524.080 2898.430 1525.210 2898.490 ;
        RECT 1524.080 2898.170 1524.340 2898.430 ;
        RECT 1503.380 2896.530 1503.640 2896.790 ;
        RECT 1502.850 2896.470 1503.640 2896.530 ;
        RECT 1502.850 2896.390 1503.580 2896.470 ;
        RECT 1502.850 2896.055 1503.130 2896.390 ;
        RECT 1524.930 2896.055 1525.210 2898.430 ;
        RECT 1535.050 2896.055 1535.330 2900.055 ;
        RECT 1546.090 2896.055 1546.370 2900.055 ;
        RECT 1567.250 2896.055 1567.530 2900.055 ;
        RECT 1598.530 2896.055 1598.810 2900.055 ;
        RECT 1609.570 2896.055 1609.850 2900.055 ;
        RECT 1630.730 2896.055 1631.010 2900.055 ;
        RECT 1641.770 2896.055 1642.050 2900.055 ;
        RECT 1662.930 2896.055 1663.210 2900.055 ;
        RECT 1694.210 2896.055 1694.490 2900.055 ;
        RECT 1705.250 2896.055 1705.530 2900.055 ;
        RECT 1758.610 2896.055 1758.890 2900.055 ;
        RECT 1768.730 2896.055 1769.010 2900.055 ;
        RECT 1779.770 2896.055 1780.050 2900.055 ;
        RECT 1789.890 2896.055 1790.170 2900.055 ;
        RECT 1800.930 2896.055 1801.210 2900.055 ;
        RECT 1811.970 2896.055 1812.250 2900.055 ;
        RECT 1833.130 2896.055 1833.410 2900.055 ;
        RECT 1843.250 2896.055 1843.530 2900.055 ;
        RECT 1854.290 2896.055 1854.570 2900.055 ;
        RECT 1864.410 2896.055 1864.690 2900.055 ;
        RECT 1875.450 2896.530 1875.730 2900.055 ;
        RECT 1876.900 2896.530 1877.160 2896.790 ;
        RECT 1875.450 2896.470 1877.160 2896.530 ;
        RECT 1885.570 2896.530 1885.850 2900.055 ;
        RECT 1875.450 2896.390 1877.100 2896.470 ;
        RECT 1885.570 2896.390 1886.300 2896.530 ;
        RECT 1875.450 2896.055 1875.730 2896.390 ;
        RECT 1885.570 2896.055 1885.850 2896.390 ;
      LAYER met2 ;
        RECT 1503.410 2895.775 1513.610 2896.055 ;
        RECT 1514.450 2895.775 1524.650 2896.055 ;
        RECT 1525.490 2895.775 1534.770 2896.055 ;
        RECT 1535.610 2895.775 1545.810 2896.055 ;
        RECT 1546.650 2895.775 1555.930 2896.055 ;
        RECT 1556.770 2895.775 1566.970 2896.055 ;
        RECT 1567.810 2895.775 1577.090 2896.055 ;
        RECT 1577.930 2895.775 1588.130 2896.055 ;
        RECT 1588.970 2895.775 1598.250 2896.055 ;
        RECT 1599.090 2895.775 1609.290 2896.055 ;
        RECT 1610.130 2895.775 1620.330 2896.055 ;
        RECT 1621.170 2895.775 1630.450 2896.055 ;
        RECT 1631.290 2895.775 1641.490 2896.055 ;
        RECT 1642.330 2895.775 1651.610 2896.055 ;
        RECT 1652.450 2895.775 1662.650 2896.055 ;
        RECT 1663.490 2895.775 1672.770 2896.055 ;
        RECT 1673.610 2895.775 1683.810 2896.055 ;
        RECT 1684.650 2895.775 1693.930 2896.055 ;
        RECT 1694.770 2895.775 1704.970 2896.055 ;
        RECT 1705.810 2895.775 1716.010 2896.055 ;
        RECT 1716.850 2895.775 1726.130 2896.055 ;
        RECT 1726.970 2895.775 1737.170 2896.055 ;
        RECT 1738.010 2895.775 1747.290 2896.055 ;
        RECT 1748.130 2895.775 1758.330 2896.055 ;
        RECT 1759.170 2895.775 1768.450 2896.055 ;
        RECT 1769.290 2895.775 1779.490 2896.055 ;
        RECT 1780.330 2895.775 1789.610 2896.055 ;
        RECT 1790.450 2895.775 1800.650 2896.055 ;
        RECT 1801.490 2895.775 1811.690 2896.055 ;
        RECT 1812.530 2895.775 1821.810 2896.055 ;
        RECT 1822.650 2895.775 1832.850 2896.055 ;
        RECT 1833.690 2895.775 1842.970 2896.055 ;
        RECT 1843.810 2895.775 1854.010 2896.055 ;
        RECT 1854.850 2895.775 1864.130 2896.055 ;
        RECT 1864.970 2895.775 1875.170 2896.055 ;
        RECT 1876.010 2895.775 1885.290 2896.055 ;
      LAYER met2 ;
        RECT 1500.610 2884.035 1500.890 2884.405 ;
        RECT 1501.990 2884.035 1502.270 2884.405 ;
        RECT 1502.060 2843.070 1502.200 2884.035 ;
        RECT 1501.540 2842.750 1501.800 2843.070 ;
        RECT 1502.000 2842.750 1502.260 2843.070 ;
        RECT 1501.600 2816.210 1501.740 2842.750 ;
        RECT 1501.540 2815.890 1501.800 2816.210 ;
        RECT 1501.540 2815.210 1501.800 2815.530 ;
        RECT 1501.600 2794.790 1501.740 2815.210 ;
        RECT 1501.540 2794.470 1501.800 2794.790 ;
        RECT 1502.000 2794.470 1502.260 2794.790 ;
        RECT 1502.060 2767.250 1502.200 2794.470 ;
        RECT 1502.000 2766.930 1502.260 2767.250 ;
        RECT 1502.000 2766.250 1502.260 2766.570 ;
        RECT 1502.060 2753.310 1502.200 2766.250 ;
        RECT 1501.540 2752.990 1501.800 2753.310 ;
        RECT 1502.000 2752.990 1502.260 2753.310 ;
        RECT 1501.600 2719.310 1501.740 2752.990 ;
        RECT 1501.540 2718.990 1501.800 2719.310 ;
        RECT 1501.540 2718.310 1501.800 2718.630 ;
        RECT 1497.850 2676.975 1498.130 2677.345 ;
        RECT 1497.920 1009.110 1498.060 2676.975 ;
        RECT 1501.600 2670.690 1501.740 2718.310 ;
        RECT 1501.540 2670.370 1501.800 2670.690 ;
        RECT 1502.000 2670.030 1502.260 2670.350 ;
        RECT 1502.060 2656.750 1502.200 2670.030 ;
        RECT 1501.540 2656.430 1501.800 2656.750 ;
        RECT 1502.000 2656.430 1502.260 2656.750 ;
        RECT 1501.600 2622.750 1501.740 2656.430 ;
        RECT 1501.540 2622.430 1501.800 2622.750 ;
        RECT 1501.540 2621.750 1501.800 2622.070 ;
        RECT 1501.600 2608.210 1501.740 2621.750 ;
        RECT 1501.600 2608.070 1502.200 2608.210 ;
        RECT 1502.060 2560.045 1502.200 2608.070 ;
        RECT 1501.990 2559.675 1502.270 2560.045 ;
        RECT 1500.150 2558.995 1500.430 2559.365 ;
        RECT 1498.310 2519.215 1498.590 2519.585 ;
        RECT 1498.380 1013.190 1498.520 2519.215 ;
        RECT 1500.220 2512.250 1500.360 2558.995 ;
        RECT 1500.160 2511.930 1500.420 2512.250 ;
        RECT 1502.000 2511.930 1502.260 2512.250 ;
        RECT 1502.060 2495.930 1502.200 2511.930 ;
      LAYER met2 ;
        RECT 1502.860 2504.280 1885.840 2895.775 ;
        RECT 1503.410 2504.000 1512.690 2504.280 ;
        RECT 1513.530 2504.000 1523.730 2504.280 ;
        RECT 1524.570 2504.000 1533.850 2504.280 ;
        RECT 1534.690 2504.000 1544.890 2504.280 ;
        RECT 1545.730 2504.000 1555.010 2504.280 ;
        RECT 1555.850 2504.000 1566.050 2504.280 ;
        RECT 1566.890 2504.000 1576.170 2504.280 ;
        RECT 1577.010 2504.000 1587.210 2504.280 ;
        RECT 1588.050 2504.000 1598.250 2504.280 ;
        RECT 1599.090 2504.000 1608.370 2504.280 ;
        RECT 1609.210 2504.000 1619.410 2504.280 ;
        RECT 1620.250 2504.000 1629.530 2504.280 ;
        RECT 1630.370 2504.000 1640.570 2504.280 ;
        RECT 1641.410 2504.000 1650.690 2504.280 ;
        RECT 1651.530 2504.000 1661.730 2504.280 ;
        RECT 1662.570 2504.000 1671.850 2504.280 ;
        RECT 1672.690 2504.000 1682.890 2504.280 ;
        RECT 1683.730 2504.000 1693.930 2504.280 ;
        RECT 1694.770 2504.000 1704.050 2504.280 ;
        RECT 1704.890 2504.000 1715.090 2504.280 ;
        RECT 1715.930 2504.000 1725.210 2504.280 ;
        RECT 1726.050 2504.000 1736.250 2504.280 ;
        RECT 1737.090 2504.000 1746.370 2504.280 ;
        RECT 1747.210 2504.000 1757.410 2504.280 ;
        RECT 1758.250 2504.000 1767.530 2504.280 ;
        RECT 1768.370 2504.000 1778.570 2504.280 ;
        RECT 1779.410 2504.000 1789.610 2504.280 ;
        RECT 1790.450 2504.000 1799.730 2504.280 ;
        RECT 1800.570 2504.000 1810.770 2504.280 ;
        RECT 1811.610 2504.000 1820.890 2504.280 ;
        RECT 1821.730 2504.000 1831.930 2504.280 ;
        RECT 1832.770 2504.000 1842.050 2504.280 ;
        RECT 1842.890 2504.000 1853.090 2504.280 ;
        RECT 1853.930 2504.000 1863.210 2504.280 ;
        RECT 1864.050 2504.000 1874.250 2504.280 ;
        RECT 1875.090 2504.000 1885.290 2504.280 ;
      LAYER met2 ;
        RECT 1524.010 2500.770 1524.290 2504.000 ;
        RECT 1524.010 2500.630 1524.740 2500.770 ;
        RECT 1524.010 2500.000 1524.290 2500.630 ;
        RECT 1502.000 2495.610 1502.260 2495.930 ;
        RECT 1512.120 2491.190 1512.380 2491.510 ;
        RECT 1507.520 2485.070 1507.780 2485.390 ;
        RECT 1507.060 1020.350 1507.320 1020.670 ;
        RECT 1498.320 1012.870 1498.580 1013.190 ;
        RECT 1500.620 1011.510 1500.880 1011.830 ;
        RECT 1497.860 1008.790 1498.120 1009.110 ;
        RECT 1497.400 1008.110 1497.660 1008.430 ;
        RECT 1496.480 1007.770 1496.740 1008.090 ;
        RECT 1500.680 1000.010 1500.820 1011.510 ;
        RECT 1503.840 1009.810 1504.100 1010.130 ;
        RECT 1503.900 1000.010 1504.040 1009.810 ;
        RECT 1507.120 1000.010 1507.260 1020.350 ;
        RECT 1507.580 1014.210 1507.720 2485.070 ;
        RECT 1507.520 1013.890 1507.780 1014.210 ;
        RECT 1511.660 1013.550 1511.920 1013.870 ;
        RECT 1509.360 1011.850 1509.620 1012.170 ;
        RECT 1509.420 1000.010 1509.560 1011.850 ;
        RECT 1511.720 1007.750 1511.860 1013.550 ;
        RECT 1511.660 1007.430 1511.920 1007.750 ;
        RECT 1512.180 1000.010 1512.320 2491.190 ;
        RECT 1520.850 2463.115 1521.130 2463.485 ;
        RECT 1520.920 2429.290 1521.060 2463.115 ;
        RECT 1520.860 2428.970 1521.120 2429.290 ;
        RECT 1521.320 2428.290 1521.580 2428.610 ;
        RECT 1521.380 2415.010 1521.520 2428.290 ;
        RECT 1519.940 2414.690 1520.200 2415.010 ;
        RECT 1521.320 2414.690 1521.580 2415.010 ;
        RECT 1520.000 2366.925 1520.140 2414.690 ;
        RECT 1519.930 2366.555 1520.210 2366.925 ;
        RECT 1520.850 2366.555 1521.130 2366.925 ;
        RECT 1520.920 2332.390 1521.060 2366.555 ;
        RECT 1520.860 2332.070 1521.120 2332.390 ;
        RECT 1521.320 2331.730 1521.580 2332.050 ;
        RECT 1521.380 2284.450 1521.520 2331.730 ;
        RECT 1521.320 2284.130 1521.580 2284.450 ;
        RECT 1521.320 2283.450 1521.580 2283.770 ;
        RECT 1521.380 2270.170 1521.520 2283.450 ;
        RECT 1521.320 2269.850 1521.580 2270.170 ;
        RECT 1521.780 2269.850 1522.040 2270.170 ;
        RECT 1521.840 2263.030 1521.980 2269.850 ;
        RECT 1520.860 2262.710 1521.120 2263.030 ;
        RECT 1521.780 2262.710 1522.040 2263.030 ;
        RECT 1520.920 2215.090 1521.060 2262.710 ;
        RECT 1520.400 2214.770 1520.660 2215.090 ;
        RECT 1520.860 2214.770 1521.120 2215.090 ;
        RECT 1520.460 2173.950 1520.600 2214.770 ;
        RECT 1520.400 2173.630 1520.660 2173.950 ;
        RECT 1520.860 2173.630 1521.120 2173.950 ;
        RECT 1520.920 2163.070 1521.060 2173.630 ;
        RECT 1520.860 2162.750 1521.120 2163.070 ;
        RECT 1521.780 2162.750 1522.040 2163.070 ;
        RECT 1521.840 2100.930 1521.980 2162.750 ;
        RECT 1520.460 2100.790 1521.980 2100.930 ;
        RECT 1520.460 2077.050 1520.600 2100.790 ;
        RECT 1519.940 2076.730 1520.200 2077.050 ;
        RECT 1520.400 2076.730 1520.660 2077.050 ;
        RECT 1520.000 2069.910 1520.140 2076.730 ;
        RECT 1519.020 2069.590 1519.280 2069.910 ;
        RECT 1519.940 2069.590 1520.200 2069.910 ;
        RECT 1519.080 2025.450 1519.220 2069.590 ;
        RECT 1519.080 2025.310 1520.140 2025.450 ;
        RECT 1520.000 1994.090 1520.140 2025.310 ;
        RECT 1519.940 1993.770 1520.200 1994.090 ;
        RECT 1521.320 1993.770 1521.580 1994.090 ;
        RECT 1521.380 1946.150 1521.520 1993.770 ;
        RECT 1521.320 1945.830 1521.580 1946.150 ;
        RECT 1520.860 1945.490 1521.120 1945.810 ;
        RECT 1520.920 1932.290 1521.060 1945.490 ;
        RECT 1520.920 1932.150 1521.520 1932.290 ;
        RECT 1521.380 1931.870 1521.520 1932.150 ;
        RECT 1521.320 1931.550 1521.580 1931.870 ;
        RECT 1522.240 1931.550 1522.500 1931.870 ;
        RECT 1522.300 1896.250 1522.440 1931.550 ;
        RECT 1521.380 1896.110 1522.440 1896.250 ;
        RECT 1521.380 1859.790 1521.520 1896.110 ;
        RECT 1521.320 1859.470 1521.580 1859.790 ;
        RECT 1522.240 1859.470 1522.500 1859.790 ;
        RECT 1522.300 1800.370 1522.440 1859.470 ;
        RECT 1521.380 1800.230 1522.440 1800.370 ;
        RECT 1521.380 1763.230 1521.520 1800.230 ;
        RECT 1521.320 1762.910 1521.580 1763.230 ;
        RECT 1522.240 1762.910 1522.500 1763.230 ;
        RECT 1522.300 1690.810 1522.440 1762.910 ;
        RECT 1520.860 1690.490 1521.120 1690.810 ;
        RECT 1522.240 1690.490 1522.500 1690.810 ;
        RECT 1520.920 1690.210 1521.060 1690.490 ;
        RECT 1520.920 1690.070 1521.520 1690.210 ;
        RECT 1521.380 1656.470 1521.520 1690.070 ;
        RECT 1521.320 1656.150 1521.580 1656.470 ;
        RECT 1520.860 1655.810 1521.120 1656.130 ;
        RECT 1520.920 1607.850 1521.060 1655.810 ;
        RECT 1520.860 1607.530 1521.120 1607.850 ;
        RECT 1521.320 1607.530 1521.580 1607.850 ;
        RECT 1521.380 1593.910 1521.520 1607.530 ;
        RECT 1521.320 1593.590 1521.580 1593.910 ;
        RECT 1522.700 1593.590 1522.960 1593.910 ;
        RECT 1522.760 1546.310 1522.900 1593.590 ;
        RECT 1521.320 1545.990 1521.580 1546.310 ;
        RECT 1522.700 1545.990 1522.960 1546.310 ;
        RECT 1521.380 1545.630 1521.520 1545.990 ;
        RECT 1521.320 1545.310 1521.580 1545.630 ;
        RECT 1522.240 1545.310 1522.500 1545.630 ;
        RECT 1522.300 1507.970 1522.440 1545.310 ;
        RECT 1521.380 1507.830 1522.440 1507.970 ;
        RECT 1521.380 1497.350 1521.520 1507.830 ;
        RECT 1521.320 1497.030 1521.580 1497.350 ;
        RECT 1522.700 1497.030 1522.960 1497.350 ;
        RECT 1522.760 1449.750 1522.900 1497.030 ;
        RECT 1521.320 1449.430 1521.580 1449.750 ;
        RECT 1522.700 1449.430 1522.960 1449.750 ;
        RECT 1521.380 1449.070 1521.520 1449.430 ;
        RECT 1521.320 1448.750 1521.580 1449.070 ;
        RECT 1522.240 1448.750 1522.500 1449.070 ;
        RECT 1522.300 1413.450 1522.440 1448.750 ;
        RECT 1521.380 1413.310 1522.440 1413.450 ;
        RECT 1521.380 1400.790 1521.520 1413.310 ;
        RECT 1521.320 1400.470 1521.580 1400.790 ;
        RECT 1522.700 1400.470 1522.960 1400.790 ;
        RECT 1522.760 1353.190 1522.900 1400.470 ;
        RECT 1521.320 1352.870 1521.580 1353.190 ;
        RECT 1522.700 1352.870 1522.960 1353.190 ;
        RECT 1521.380 1352.510 1521.520 1352.870 ;
        RECT 1521.320 1352.190 1521.580 1352.510 ;
        RECT 1522.700 1352.190 1522.960 1352.510 ;
        RECT 1522.760 1317.490 1522.900 1352.190 ;
        RECT 1521.320 1317.170 1521.580 1317.490 ;
        RECT 1522.700 1317.170 1522.960 1317.490 ;
        RECT 1521.380 1304.230 1521.520 1317.170 ;
        RECT 1521.320 1303.910 1521.580 1304.230 ;
        RECT 1522.700 1303.910 1522.960 1304.230 ;
        RECT 1522.760 1257.165 1522.900 1303.910 ;
        RECT 1522.690 1256.795 1522.970 1257.165 ;
        RECT 1521.770 1255.435 1522.050 1255.805 ;
        RECT 1521.840 1207.670 1521.980 1255.435 ;
        RECT 1520.860 1207.350 1521.120 1207.670 ;
        RECT 1521.780 1207.350 1522.040 1207.670 ;
        RECT 1520.920 1206.990 1521.060 1207.350 ;
        RECT 1519.480 1206.670 1519.740 1206.990 ;
        RECT 1520.860 1206.670 1521.120 1206.990 ;
        RECT 1519.540 1159.390 1519.680 1206.670 ;
        RECT 1519.480 1159.070 1519.740 1159.390 ;
        RECT 1520.860 1159.130 1521.120 1159.390 ;
        RECT 1520.860 1159.070 1521.520 1159.130 ;
        RECT 1520.920 1158.990 1521.520 1159.070 ;
        RECT 1521.380 1125.050 1521.520 1158.990 ;
        RECT 1521.320 1124.730 1521.580 1125.050 ;
        RECT 1521.780 1124.050 1522.040 1124.370 ;
        RECT 1521.840 1104.050 1521.980 1124.050 ;
        RECT 1521.380 1103.910 1521.980 1104.050 ;
        RECT 1521.380 1080.170 1521.520 1103.910 ;
        RECT 1520.400 1079.850 1520.660 1080.170 ;
        RECT 1521.320 1079.850 1521.580 1080.170 ;
        RECT 1520.460 1055.885 1520.600 1079.850 ;
        RECT 1520.390 1055.515 1520.670 1055.885 ;
        RECT 1521.310 1055.515 1521.590 1055.885 ;
        RECT 1521.380 1038.770 1521.520 1055.515 ;
        RECT 1520.920 1038.630 1521.520 1038.770 ;
        RECT 1514.420 1016.270 1514.680 1016.590 ;
        RECT 1514.480 1000.010 1514.620 1016.270 ;
        RECT 1517.180 1013.550 1517.440 1013.870 ;
        RECT 1517.240 1012.850 1517.380 1013.550 ;
        RECT 1518.560 1013.210 1518.820 1013.530 ;
        RECT 1517.180 1012.530 1517.440 1012.850 ;
        RECT 1516.720 1012.190 1516.980 1012.510 ;
        RECT 1516.780 1011.570 1516.920 1012.190 ;
        RECT 1518.620 1012.170 1518.760 1013.210 ;
        RECT 1518.560 1011.850 1518.820 1012.170 ;
        RECT 1516.780 1011.430 1518.300 1011.570 ;
        RECT 1518.160 1010.890 1518.300 1011.430 ;
        RECT 1518.160 1010.750 1519.680 1010.890 ;
        RECT 1514.880 1007.430 1515.140 1007.750 ;
        RECT 1494.700 1000.000 1495.000 1000.010 ;
        RECT 1495.620 1000.000 1496.840 1000.010 ;
        RECT 1499.140 1000.000 1500.820 1000.010 ;
        RECT 1503.740 1000.000 1504.040 1000.010 ;
        RECT 1505.580 1000.000 1507.260 1000.010 ;
        RECT 1507.880 1000.000 1509.560 1000.010 ;
        RECT 1512.020 1000.000 1512.320 1000.010 ;
        RECT 1514.320 1000.000 1514.620 1000.010 ;
        RECT 1338.760 999.870 1340.590 1000.000 ;
        RECT 1341.060 999.870 1342.890 1000.000 ;
        RECT 1343.360 999.870 1345.190 1000.000 ;
        RECT 1345.660 999.870 1347.030 1000.000 ;
        RECT 1347.500 999.870 1349.330 1000.000 ;
      LAYER met2 ;
        RECT 1334.430 995.720 1335.890 998.810 ;
      LAYER met2 ;
        RECT 1336.170 996.000 1336.450 999.870 ;
      LAYER met2 ;
        RECT 1336.730 995.720 1337.730 998.810 ;
      LAYER met2 ;
        RECT 1338.010 996.000 1338.290 999.870 ;
      LAYER met2 ;
        RECT 1338.570 995.720 1340.030 998.810 ;
      LAYER met2 ;
        RECT 1340.310 996.000 1340.590 999.870 ;
      LAYER met2 ;
        RECT 1340.870 995.720 1342.330 998.810 ;
      LAYER met2 ;
        RECT 1342.610 996.000 1342.890 999.870 ;
      LAYER met2 ;
        RECT 1343.170 995.720 1344.630 998.810 ;
      LAYER met2 ;
        RECT 1344.910 996.000 1345.190 999.870 ;
      LAYER met2 ;
        RECT 1345.470 995.720 1346.470 998.810 ;
      LAYER met2 ;
        RECT 1346.750 996.000 1347.030 999.870 ;
      LAYER met2 ;
        RECT 1347.310 995.720 1348.770 998.810 ;
      LAYER met2 ;
        RECT 1349.050 996.000 1349.330 999.870 ;
        RECT 1351.350 999.870 1352.240 1000.000 ;
        RECT 1353.190 999.870 1355.000 1000.000 ;
        RECT 1355.490 999.870 1357.300 1000.000 ;
        RECT 1357.790 999.870 1359.140 1000.000 ;
        RECT 1360.090 999.870 1361.440 1000.000 ;
      LAYER met2 ;
        RECT 1349.610 995.720 1351.070 998.810 ;
      LAYER met2 ;
        RECT 1351.350 996.000 1351.630 999.870 ;
      LAYER met2 ;
        RECT 1351.910 995.720 1352.910 998.810 ;
      LAYER met2 ;
        RECT 1353.190 996.000 1353.470 999.870 ;
      LAYER met2 ;
        RECT 1353.750 995.720 1355.210 998.810 ;
      LAYER met2 ;
        RECT 1355.490 996.000 1355.770 999.870 ;
      LAYER met2 ;
        RECT 1356.050 995.720 1357.510 998.810 ;
      LAYER met2 ;
        RECT 1357.790 996.000 1358.070 999.870 ;
      LAYER met2 ;
        RECT 1358.350 995.720 1359.810 998.810 ;
      LAYER met2 ;
        RECT 1360.090 996.000 1360.370 999.870 ;
      LAYER met2 ;
        RECT 1360.650 995.720 1361.650 998.810 ;
      LAYER met2 ;
        RECT 1361.930 996.000 1362.210 1000.000 ;
      LAYER met2 ;
        RECT 1362.490 995.720 1363.950 998.810 ;
      LAYER met2 ;
        RECT 1364.230 996.000 1364.510 1000.000 ;
        RECT 1366.530 999.870 1368.340 1000.000 ;
        RECT 1368.830 999.870 1370.180 1000.000 ;
      LAYER met2 ;
        RECT 1364.790 995.720 1366.250 998.810 ;
      LAYER met2 ;
        RECT 1366.530 996.000 1366.810 999.870 ;
      LAYER met2 ;
        RECT 1367.090 995.720 1368.550 998.810 ;
      LAYER met2 ;
        RECT 1368.830 996.000 1369.110 999.870 ;
      LAYER met2 ;
        RECT 1369.390 995.720 1370.390 998.810 ;
      LAYER met2 ;
        RECT 1370.670 996.000 1370.950 1000.000 ;
      LAYER met2 ;
        RECT 1371.230 995.720 1372.690 998.810 ;
      LAYER met2 ;
        RECT 1372.970 996.000 1373.250 1000.000 ;
        RECT 1375.270 999.870 1376.620 1000.000 ;
        RECT 1377.110 999.870 1378.920 1000.000 ;
      LAYER met2 ;
        RECT 1373.530 995.720 1374.990 998.810 ;
      LAYER met2 ;
        RECT 1375.270 996.000 1375.550 999.870 ;
      LAYER met2 ;
        RECT 1375.830 995.720 1376.830 998.810 ;
      LAYER met2 ;
        RECT 1377.110 996.000 1377.390 999.870 ;
      LAYER met2 ;
        RECT 1377.670 995.720 1379.130 998.810 ;
      LAYER met2 ;
        RECT 1379.410 996.000 1379.690 1000.000 ;
      LAYER met2 ;
        RECT 1379.970 995.720 1381.430 998.810 ;
      LAYER met2 ;
        RECT 1381.710 996.000 1381.990 1000.000 ;
        RECT 1384.010 999.870 1384.900 1000.000 ;
        RECT 1385.850 999.870 1386.740 1000.000 ;
      LAYER met2 ;
        RECT 1382.270 995.720 1383.730 998.810 ;
      LAYER met2 ;
        RECT 1384.010 996.000 1384.290 999.870 ;
      LAYER met2 ;
        RECT 1384.570 995.720 1385.570 998.810 ;
      LAYER met2 ;
        RECT 1385.850 996.000 1386.130 999.870 ;
      LAYER met2 ;
        RECT 1386.410 995.720 1387.870 998.810 ;
      LAYER met2 ;
        RECT 1388.150 996.000 1388.430 1000.000 ;
      LAYER met2 ;
        RECT 1388.710 995.720 1390.170 998.810 ;
      LAYER met2 ;
        RECT 1390.450 996.000 1390.730 1000.000 ;
        RECT 1392.750 999.870 1393.640 1000.000 ;
        RECT 1394.590 999.870 1396.400 1000.000 ;
      LAYER met2 ;
        RECT 1391.010 995.720 1392.470 998.810 ;
      LAYER met2 ;
        RECT 1392.750 996.000 1393.030 999.870 ;
      LAYER met2 ;
        RECT 1393.310 995.720 1394.310 998.810 ;
      LAYER met2 ;
        RECT 1394.590 996.000 1394.870 999.870 ;
      LAYER met2 ;
        RECT 1395.150 995.720 1396.610 998.810 ;
      LAYER met2 ;
        RECT 1396.890 996.000 1397.170 1000.000 ;
      LAYER met2 ;
        RECT 1397.450 995.720 1398.910 998.810 ;
      LAYER met2 ;
        RECT 1399.190 996.000 1399.470 1000.000 ;
        RECT 1401.030 999.870 1402.840 1000.000 ;
        RECT 1403.330 999.870 1405.140 1000.000 ;
      LAYER met2 ;
        RECT 1399.750 995.720 1400.750 998.810 ;
      LAYER met2 ;
        RECT 1401.030 996.000 1401.310 999.870 ;
      LAYER met2 ;
        RECT 1401.590 995.720 1403.050 998.810 ;
      LAYER met2 ;
        RECT 1403.330 996.000 1403.610 999.870 ;
      LAYER met2 ;
        RECT 1403.890 995.720 1405.350 998.810 ;
      LAYER met2 ;
        RECT 1405.630 996.000 1405.910 1000.000 ;
      LAYER met2 ;
        RECT 1406.190 995.720 1407.650 998.810 ;
      LAYER met2 ;
        RECT 1407.930 996.000 1408.210 1000.000 ;
        RECT 1409.770 999.870 1411.580 1000.000 ;
        RECT 1412.070 999.870 1413.420 1000.000 ;
      LAYER met2 ;
        RECT 1408.490 995.720 1409.490 998.810 ;
      LAYER met2 ;
        RECT 1409.770 996.000 1410.050 999.870 ;
      LAYER met2 ;
        RECT 1410.330 995.720 1411.790 998.810 ;
      LAYER met2 ;
        RECT 1412.070 996.000 1412.350 999.870 ;
      LAYER met2 ;
        RECT 1412.630 995.720 1414.090 998.810 ;
      LAYER met2 ;
        RECT 1414.370 996.000 1414.650 1000.000 ;
        RECT 1416.670 999.870 1418.020 1000.000 ;
        RECT 1418.510 999.870 1420.320 1000.000 ;
        RECT 1420.810 999.870 1421.240 1000.000 ;
      LAYER met2 ;
        RECT 1414.930 995.720 1416.390 998.810 ;
      LAYER met2 ;
        RECT 1416.670 996.000 1416.950 999.870 ;
      LAYER met2 ;
        RECT 1417.230 995.720 1418.230 998.810 ;
      LAYER met2 ;
        RECT 1418.510 996.000 1418.790 999.870 ;
      LAYER met2 ;
        RECT 1419.070 995.720 1420.530 998.810 ;
      LAYER met2 ;
        RECT 1420.810 996.000 1421.090 999.870 ;
      LAYER met2 ;
        RECT 1421.370 995.720 1422.830 998.810 ;
      LAYER met2 ;
        RECT 1423.110 996.000 1423.390 1000.000 ;
      LAYER met2 ;
        RECT 1423.670 995.720 1424.670 998.810 ;
      LAYER met2 ;
        RECT 1424.950 996.000 1425.230 1000.000 ;
        RECT 1427.250 999.870 1428.140 1000.000 ;
        RECT 1429.550 999.870 1431.360 1000.000 ;
      LAYER met2 ;
        RECT 1425.510 995.720 1426.970 998.810 ;
      LAYER met2 ;
        RECT 1427.250 996.000 1427.530 999.870 ;
      LAYER met2 ;
        RECT 1427.810 995.720 1429.270 998.810 ;
      LAYER met2 ;
        RECT 1429.550 996.000 1429.830 999.870 ;
      LAYER met2 ;
        RECT 1430.110 995.720 1431.570 998.810 ;
      LAYER met2 ;
        RECT 1431.850 996.000 1432.130 1000.000 ;
        RECT 1433.690 999.870 1434.580 1000.000 ;
        RECT 1435.990 999.870 1437.800 1000.000 ;
        RECT 1438.290 999.870 1440.100 1000.000 ;
      LAYER met2 ;
        RECT 1432.410 995.720 1433.410 998.810 ;
      LAYER met2 ;
        RECT 1433.690 996.000 1433.970 999.870 ;
      LAYER met2 ;
        RECT 1434.250 995.720 1435.710 998.810 ;
      LAYER met2 ;
        RECT 1435.990 996.000 1436.270 999.870 ;
      LAYER met2 ;
        RECT 1436.550 995.720 1438.010 998.810 ;
      LAYER met2 ;
        RECT 1438.290 996.000 1438.570 999.870 ;
      LAYER met2 ;
        RECT 1438.850 995.720 1440.310 998.810 ;
      LAYER met2 ;
        RECT 1440.590 996.000 1440.870 1000.000 ;
        RECT 1442.430 999.870 1444.240 1000.000 ;
        RECT 1444.730 999.870 1446.540 1000.000 ;
        RECT 1447.030 999.870 1447.920 1000.000 ;
      LAYER met2 ;
        RECT 1441.150 995.720 1442.150 998.810 ;
      LAYER met2 ;
        RECT 1442.430 996.000 1442.710 999.870 ;
      LAYER met2 ;
        RECT 1442.990 995.720 1444.450 998.810 ;
      LAYER met2 ;
        RECT 1444.730 996.000 1445.010 999.870 ;
      LAYER met2 ;
        RECT 1445.290 995.720 1446.750 998.810 ;
      LAYER met2 ;
        RECT 1447.030 996.000 1447.310 999.870 ;
      LAYER met2 ;
        RECT 1447.590 995.720 1448.590 998.810 ;
      LAYER met2 ;
        RECT 1448.870 996.000 1449.150 1000.000 ;
        RECT 1451.170 999.870 1452.980 1000.000 ;
        RECT 1453.470 999.870 1455.280 1000.000 ;
        RECT 1455.770 999.870 1457.120 1000.000 ;
      LAYER met2 ;
        RECT 1449.430 995.720 1450.890 998.810 ;
      LAYER met2 ;
        RECT 1451.170 996.000 1451.450 999.870 ;
      LAYER met2 ;
        RECT 1451.730 995.720 1453.190 998.810 ;
      LAYER met2 ;
        RECT 1453.470 996.000 1453.750 999.870 ;
      LAYER met2 ;
        RECT 1454.030 995.720 1455.490 998.810 ;
      LAYER met2 ;
        RECT 1455.770 996.000 1456.050 999.870 ;
      LAYER met2 ;
        RECT 1456.330 995.720 1457.330 998.810 ;
      LAYER met2 ;
        RECT 1457.610 996.000 1457.890 1000.000 ;
        RECT 1459.910 999.870 1461.720 1000.000 ;
        RECT 1462.210 999.870 1462.640 1000.000 ;
        RECT 1464.510 999.870 1465.860 1000.000 ;
      LAYER met2 ;
        RECT 1458.170 995.720 1459.630 998.810 ;
      LAYER met2 ;
        RECT 1459.910 996.000 1460.190 999.870 ;
      LAYER met2 ;
        RECT 1460.470 995.720 1461.930 998.810 ;
      LAYER met2 ;
        RECT 1462.210 996.000 1462.490 999.870 ;
      LAYER met2 ;
        RECT 1462.770 995.720 1464.230 998.810 ;
      LAYER met2 ;
        RECT 1464.510 996.000 1464.790 999.870 ;
      LAYER met2 ;
        RECT 1465.070 995.720 1466.070 998.810 ;
      LAYER met2 ;
        RECT 1466.350 996.000 1466.630 1000.000 ;
        RECT 1468.650 999.870 1469.540 1000.000 ;
        RECT 1470.950 999.870 1472.300 1000.000 ;
        RECT 1472.790 999.870 1474.600 1000.000 ;
      LAYER met2 ;
        RECT 1466.910 995.720 1468.370 998.810 ;
      LAYER met2 ;
        RECT 1468.650 996.000 1468.930 999.870 ;
      LAYER met2 ;
        RECT 1469.210 995.720 1470.670 998.810 ;
      LAYER met2 ;
        RECT 1470.950 996.000 1471.230 999.870 ;
      LAYER met2 ;
        RECT 1471.510 995.720 1472.510 998.810 ;
      LAYER met2 ;
        RECT 1472.790 996.000 1473.070 999.870 ;
      LAYER met2 ;
        RECT 1473.350 995.720 1474.810 998.810 ;
      LAYER met2 ;
        RECT 1475.090 996.000 1475.370 1000.000 ;
        RECT 1477.390 999.870 1479.200 1000.000 ;
        RECT 1479.690 999.870 1481.040 1000.000 ;
        RECT 1481.530 999.870 1482.880 1000.000 ;
      LAYER met2 ;
        RECT 1475.650 995.720 1477.110 998.810 ;
      LAYER met2 ;
        RECT 1477.390 996.000 1477.670 999.870 ;
      LAYER met2 ;
        RECT 1477.950 995.720 1479.410 998.810 ;
      LAYER met2 ;
        RECT 1479.690 996.000 1479.970 999.870 ;
      LAYER met2 ;
        RECT 1480.250 995.720 1481.250 998.810 ;
      LAYER met2 ;
        RECT 1481.530 996.000 1481.810 999.870 ;
      LAYER met2 ;
        RECT 1482.090 995.720 1483.550 998.810 ;
      LAYER met2 ;
        RECT 1483.830 996.000 1484.110 1000.000 ;
        RECT 1486.130 999.870 1487.940 1000.000 ;
        RECT 1488.430 999.870 1489.780 1000.000 ;
        RECT 1490.270 999.870 1492.080 1000.000 ;
      LAYER met2 ;
        RECT 1484.390 995.720 1485.850 998.810 ;
      LAYER met2 ;
        RECT 1486.130 996.000 1486.410 999.870 ;
      LAYER met2 ;
        RECT 1486.690 995.720 1488.150 998.810 ;
      LAYER met2 ;
        RECT 1488.430 996.000 1488.710 999.870 ;
      LAYER met2 ;
        RECT 1488.990 995.720 1489.990 998.810 ;
      LAYER met2 ;
        RECT 1490.270 996.000 1490.550 999.870 ;
      LAYER met2 ;
        RECT 1490.830 995.720 1492.290 998.810 ;
      LAYER met2 ;
        RECT 1492.570 996.000 1492.850 1000.000 ;
        RECT 1494.700 999.870 1495.150 1000.000 ;
        RECT 1495.620 999.870 1496.990 1000.000 ;
      LAYER met2 ;
        RECT 1493.130 995.720 1494.590 998.810 ;
      LAYER met2 ;
        RECT 1494.870 996.000 1495.150 999.870 ;
      LAYER met2 ;
        RECT 1495.430 995.720 1496.430 998.810 ;
      LAYER met2 ;
        RECT 1496.710 996.000 1496.990 999.870 ;
        RECT 1499.010 999.870 1500.820 1000.000 ;
      LAYER met2 ;
        RECT 1497.270 995.720 1498.730 998.810 ;
      LAYER met2 ;
        RECT 1499.010 996.000 1499.290 999.870 ;
      LAYER met2 ;
        RECT 1499.570 995.720 1501.030 998.810 ;
      LAYER met2 ;
        RECT 1501.310 996.000 1501.590 1000.000 ;
        RECT 1503.610 999.870 1504.040 1000.000 ;
        RECT 1505.450 999.870 1507.260 1000.000 ;
        RECT 1507.750 999.870 1509.560 1000.000 ;
      LAYER met2 ;
        RECT 1501.870 995.720 1503.330 998.810 ;
      LAYER met2 ;
        RECT 1503.610 996.000 1503.890 999.870 ;
      LAYER met2 ;
        RECT 1504.170 995.720 1505.170 998.810 ;
      LAYER met2 ;
        RECT 1505.450 996.000 1505.730 999.870 ;
      LAYER met2 ;
        RECT 1506.010 995.720 1507.470 998.810 ;
      LAYER met2 ;
        RECT 1507.750 996.000 1508.030 999.870 ;
      LAYER met2 ;
        RECT 1508.310 995.720 1509.770 998.810 ;
      LAYER met2 ;
        RECT 1510.050 996.000 1510.330 1000.000 ;
        RECT 1511.890 999.870 1512.320 1000.000 ;
        RECT 1514.190 999.870 1514.620 1000.000 ;
        RECT 1514.940 1000.010 1515.080 1007.430 ;
        RECT 1519.540 1000.010 1519.680 1010.750 ;
        RECT 1520.920 1010.470 1521.060 1038.630 ;
        RECT 1521.320 1020.690 1521.580 1021.010 ;
        RECT 1520.860 1010.150 1521.120 1010.470 ;
        RECT 1521.380 1000.010 1521.520 1020.690 ;
        RECT 1524.080 1012.870 1524.340 1013.190 ;
        RECT 1524.140 1008.770 1524.280 1012.870 ;
        RECT 1524.600 1012.510 1524.740 2500.630 ;
        RECT 1534.130 2500.000 1534.410 2504.000 ;
        RECT 1545.170 2500.090 1545.450 2504.000 ;
        RECT 1544.840 2500.000 1545.450 2500.090 ;
        RECT 1555.290 2500.000 1555.570 2504.000 ;
        RECT 1576.450 2500.000 1576.730 2504.000 ;
        RECT 1587.490 2500.000 1587.770 2504.000 ;
        RECT 1608.650 2500.000 1608.930 2504.000 ;
        RECT 1619.690 2500.000 1619.970 2504.000 ;
        RECT 1629.810 2500.000 1630.090 2504.000 ;
        RECT 1640.850 2500.090 1641.130 2504.000 ;
        RECT 1662.010 2500.090 1662.290 2504.000 ;
        RECT 1635.460 2500.000 1641.130 2500.090 ;
        RECT 1656.160 2500.000 1662.290 2500.090 ;
        RECT 1683.170 2500.000 1683.450 2504.000 ;
        RECT 1704.330 2500.000 1704.610 2504.000 ;
        RECT 1715.370 2500.000 1715.650 2504.000 ;
        RECT 1725.490 2500.000 1725.770 2504.000 ;
        RECT 1746.650 2500.000 1746.930 2504.000 ;
        RECT 1757.690 2500.000 1757.970 2504.000 ;
        RECT 1767.810 2500.090 1768.090 2504.000 ;
        RECT 1766.560 2500.000 1768.090 2500.090 ;
        RECT 1778.850 2500.000 1779.130 2504.000 ;
        RECT 1789.890 2500.000 1790.170 2504.000 ;
        RECT 1811.050 2500.000 1811.330 2504.000 ;
        RECT 1832.210 2500.000 1832.490 2504.000 ;
        RECT 1842.330 2500.000 1842.610 2504.000 ;
        RECT 1853.370 2500.090 1853.650 2504.000 ;
        RECT 1849.360 2500.000 1853.650 2500.090 ;
        RECT 1874.530 2500.000 1874.810 2504.000 ;
        RECT 1885.570 2500.000 1885.850 2504.000 ;
        RECT 1532.360 2493.910 1532.620 2494.230 ;
        RECT 1530.060 2487.790 1530.320 2488.110 ;
        RECT 1528.220 2484.390 1528.480 2484.710 ;
        RECT 1528.280 1014.210 1528.420 2484.390 ;
        RECT 1530.120 2463.485 1530.260 2487.790 ;
        RECT 1530.050 2463.115 1530.330 2463.485 ;
        RECT 1528.220 1013.890 1528.480 1014.210 ;
        RECT 1524.540 1012.190 1524.800 1012.510 ;
        RECT 1525.460 1011.850 1525.720 1012.170 ;
        RECT 1524.540 1009.530 1524.800 1009.790 ;
        RECT 1524.540 1009.470 1525.200 1009.530 ;
        RECT 1524.600 1009.390 1525.200 1009.470 ;
        RECT 1525.060 1008.770 1525.200 1009.390 ;
        RECT 1524.080 1008.450 1524.340 1008.770 ;
        RECT 1525.000 1008.450 1525.260 1008.770 ;
        RECT 1525.520 1000.010 1525.660 1011.850 ;
        RECT 1531.900 1009.530 1532.160 1009.790 ;
        RECT 1531.040 1009.470 1532.160 1009.530 ;
        RECT 1531.040 1009.450 1532.100 1009.470 ;
        RECT 1530.980 1009.390 1532.100 1009.450 ;
        RECT 1530.980 1009.130 1531.240 1009.390 ;
        RECT 1532.420 1008.770 1532.560 2493.910 ;
        RECT 1534.260 2485.050 1534.400 2500.000 ;
        RECT 1544.840 2499.950 1545.370 2500.000 ;
        RECT 1544.840 2485.050 1544.980 2499.950 ;
        RECT 1553.060 2495.270 1553.320 2495.590 ;
        RECT 1545.700 2494.250 1545.960 2494.570 ;
        RECT 1552.140 2494.250 1552.400 2494.570 ;
        RECT 1545.240 2493.910 1545.500 2494.230 ;
        RECT 1534.200 2484.730 1534.460 2485.050 ;
        RECT 1544.780 2484.730 1545.040 2485.050 ;
        RECT 1542.020 2484.050 1542.280 2484.370 ;
        RECT 1533.280 1020.690 1533.540 1021.010 ;
        RECT 1528.220 1008.450 1528.480 1008.770 ;
        RECT 1532.360 1008.450 1532.620 1008.770 ;
        RECT 1514.940 1000.000 1516.620 1000.010 ;
        RECT 1519.540 1000.000 1520.760 1000.010 ;
        RECT 1521.380 1000.000 1523.060 1000.010 ;
        RECT 1525.360 1000.000 1525.660 1000.010 ;
        RECT 1528.280 1000.010 1528.420 1008.450 ;
        RECT 1533.340 1000.010 1533.480 1020.690 ;
        RECT 1542.080 1012.170 1542.220 2484.050 ;
        RECT 1545.300 1076.170 1545.440 2493.910 ;
        RECT 1544.380 1076.030 1545.440 1076.170 ;
        RECT 1544.380 1028.570 1544.520 1076.030 ;
        RECT 1543.920 1028.430 1544.520 1028.570 ;
        RECT 1535.120 1011.850 1535.380 1012.170 ;
        RECT 1542.020 1011.850 1542.280 1012.170 ;
        RECT 1542.480 1011.850 1542.740 1012.170 ;
        RECT 1535.180 1000.010 1535.320 1011.850 ;
        RECT 1542.540 1009.790 1542.680 1011.850 ;
        RECT 1542.480 1009.470 1542.740 1009.790 ;
        RECT 1536.500 1008.450 1536.760 1008.770 ;
        RECT 1542.020 1008.450 1542.280 1008.770 ;
        RECT 1528.280 1000.000 1529.500 1000.010 ;
        RECT 1531.800 1000.000 1533.480 1000.010 ;
        RECT 1534.100 1000.000 1535.320 1000.010 ;
        RECT 1536.560 1000.010 1536.700 1008.450 ;
        RECT 1542.080 1000.010 1542.220 1008.450 ;
        RECT 1543.920 1000.010 1544.060 1028.430 ;
        RECT 1545.760 1014.210 1545.900 2494.250 ;
        RECT 1545.700 1013.890 1545.960 1014.210 ;
        RECT 1548.000 1013.890 1548.260 1014.210 ;
        RECT 1545.700 1012.190 1545.960 1012.510 ;
        RECT 1536.560 1000.000 1538.240 1000.010 ;
        RECT 1540.540 1000.000 1542.220 1000.010 ;
        RECT 1542.840 1000.000 1544.060 1000.010 ;
        RECT 1545.760 1000.010 1545.900 1012.190 ;
        RECT 1548.060 1000.010 1548.200 1013.890 ;
        RECT 1552.200 1000.010 1552.340 2494.250 ;
        RECT 1553.120 1012.510 1553.260 2495.270 ;
        RECT 1555.420 2486.070 1555.560 2500.000 ;
        RECT 1559.500 2495.610 1559.760 2495.930 ;
        RECT 1555.360 2485.750 1555.620 2486.070 ;
        RECT 1559.560 1014.210 1559.700 2495.610 ;
        RECT 1574.220 2494.930 1574.480 2495.250 ;
        RECT 1567.780 1017.290 1568.040 1017.610 ;
        RECT 1559.500 1013.890 1559.760 1014.210 ;
        RECT 1562.720 1013.890 1562.980 1014.210 ;
        RECT 1553.060 1012.190 1553.320 1012.510 ;
        RECT 1556.280 1012.190 1556.540 1012.510 ;
        RECT 1556.740 1012.190 1557.000 1012.510 ;
        RECT 1555.820 1009.470 1556.080 1009.790 ;
        RECT 1555.880 1000.010 1556.020 1009.470 ;
        RECT 1545.760 1000.000 1546.980 1000.010 ;
        RECT 1548.060 1000.000 1549.280 1000.010 ;
        RECT 1551.580 1000.000 1552.340 1000.010 ;
        RECT 1555.720 1000.000 1556.020 1000.010 ;
        RECT 1514.940 999.870 1516.770 1000.000 ;
      LAYER met2 ;
        RECT 1510.610 995.720 1511.610 998.810 ;
      LAYER met2 ;
        RECT 1511.890 996.000 1512.170 999.870 ;
      LAYER met2 ;
        RECT 1512.450 995.720 1513.910 998.810 ;
      LAYER met2 ;
        RECT 1514.190 996.000 1514.470 999.870 ;
      LAYER met2 ;
        RECT 1514.750 995.720 1516.210 998.810 ;
      LAYER met2 ;
        RECT 1516.490 996.000 1516.770 999.870 ;
      LAYER met2 ;
        RECT 1517.050 995.720 1518.510 998.810 ;
      LAYER met2 ;
        RECT 1518.790 996.000 1519.070 1000.000 ;
        RECT 1519.540 999.870 1520.910 1000.000 ;
        RECT 1521.380 999.870 1523.210 1000.000 ;
      LAYER met2 ;
        RECT 1519.350 995.720 1520.350 998.810 ;
      LAYER met2 ;
        RECT 1520.630 996.000 1520.910 999.870 ;
      LAYER met2 ;
        RECT 1521.190 995.720 1522.650 998.810 ;
      LAYER met2 ;
        RECT 1522.930 996.000 1523.210 999.870 ;
        RECT 1525.230 999.870 1525.660 1000.000 ;
      LAYER met2 ;
        RECT 1523.490 995.720 1524.950 998.810 ;
      LAYER met2 ;
        RECT 1525.230 996.000 1525.510 999.870 ;
      LAYER met2 ;
        RECT 1525.790 995.720 1527.250 998.810 ;
      LAYER met2 ;
        RECT 1527.530 996.000 1527.810 1000.000 ;
        RECT 1528.280 999.870 1529.650 1000.000 ;
      LAYER met2 ;
        RECT 1528.090 995.720 1529.090 998.810 ;
      LAYER met2 ;
        RECT 1529.370 996.000 1529.650 999.870 ;
        RECT 1531.670 999.870 1533.480 1000.000 ;
        RECT 1533.970 999.870 1535.320 1000.000 ;
      LAYER met2 ;
        RECT 1529.930 995.720 1531.390 998.810 ;
      LAYER met2 ;
        RECT 1531.670 996.000 1531.950 999.870 ;
      LAYER met2 ;
        RECT 1532.230 995.720 1533.690 998.810 ;
      LAYER met2 ;
        RECT 1533.970 996.000 1534.250 999.870 ;
      LAYER met2 ;
        RECT 1534.530 995.720 1535.530 998.810 ;
      LAYER met2 ;
        RECT 1535.810 996.000 1536.090 1000.000 ;
        RECT 1536.560 999.870 1538.390 1000.000 ;
      LAYER met2 ;
        RECT 1536.370 995.720 1537.830 998.810 ;
      LAYER met2 ;
        RECT 1538.110 996.000 1538.390 999.870 ;
        RECT 1540.410 999.870 1542.220 1000.000 ;
        RECT 1542.710 999.870 1544.060 1000.000 ;
      LAYER met2 ;
        RECT 1538.670 995.720 1540.130 998.810 ;
      LAYER met2 ;
        RECT 1540.410 996.000 1540.690 999.870 ;
      LAYER met2 ;
        RECT 1540.970 995.720 1542.430 998.810 ;
      LAYER met2 ;
        RECT 1542.710 996.000 1542.990 999.870 ;
      LAYER met2 ;
        RECT 1543.270 995.720 1544.270 998.810 ;
      LAYER met2 ;
        RECT 1544.550 996.000 1544.830 1000.000 ;
        RECT 1545.760 999.870 1547.130 1000.000 ;
        RECT 1548.060 999.870 1549.430 1000.000 ;
      LAYER met2 ;
        RECT 1545.110 995.720 1546.570 998.810 ;
      LAYER met2 ;
        RECT 1546.850 996.000 1547.130 999.870 ;
      LAYER met2 ;
        RECT 1547.410 995.720 1548.870 998.810 ;
      LAYER met2 ;
        RECT 1549.150 996.000 1549.430 999.870 ;
        RECT 1551.450 999.870 1552.340 1000.000 ;
      LAYER met2 ;
        RECT 1549.710 995.720 1551.170 998.810 ;
      LAYER met2 ;
        RECT 1551.450 996.000 1551.730 999.870 ;
      LAYER met2 ;
        RECT 1552.010 995.720 1553.010 998.810 ;
      LAYER met2 ;
        RECT 1553.290 996.000 1553.570 1000.000 ;
        RECT 1555.590 999.870 1556.020 1000.000 ;
        RECT 1556.340 1000.010 1556.480 1012.190 ;
        RECT 1556.800 1010.470 1556.940 1012.190 ;
        RECT 1556.740 1010.150 1557.000 1010.470 ;
        RECT 1559.960 1008.790 1560.220 1009.110 ;
        RECT 1560.020 1000.010 1560.160 1008.790 ;
        RECT 1556.340 1000.000 1558.020 1000.010 ;
        RECT 1559.860 1000.000 1560.160 1000.010 ;
        RECT 1562.780 1000.010 1562.920 1013.890 ;
        RECT 1567.840 1000.010 1567.980 1017.290 ;
        RECT 1574.280 1014.210 1574.420 2494.930 ;
        RECT 1576.580 2484.370 1576.720 2500.000 ;
        RECT 1580.200 2494.590 1580.460 2494.910 ;
        RECT 1586.640 2494.590 1586.900 2494.910 ;
        RECT 1579.740 2485.750 1580.000 2486.070 ;
        RECT 1576.520 2484.050 1576.780 2484.370 ;
        RECT 1574.220 1013.890 1574.480 1014.210 ;
        RECT 1577.900 1013.890 1578.160 1014.210 ;
        RECT 1578.360 1013.890 1578.620 1014.210 ;
        RECT 1576.520 1010.150 1576.780 1010.470 ;
        RECT 1568.240 1009.130 1568.500 1009.450 ;
        RECT 1562.780 1000.000 1564.460 1000.010 ;
        RECT 1566.760 1000.000 1567.980 1000.010 ;
        RECT 1556.340 999.870 1558.170 1000.000 ;
      LAYER met2 ;
        RECT 1553.850 995.720 1555.310 998.810 ;
      LAYER met2 ;
        RECT 1555.590 996.000 1555.870 999.870 ;
      LAYER met2 ;
        RECT 1556.150 995.720 1557.610 998.810 ;
      LAYER met2 ;
        RECT 1557.890 996.000 1558.170 999.870 ;
        RECT 1559.730 999.870 1560.160 1000.000 ;
      LAYER met2 ;
        RECT 1558.450 995.720 1559.450 998.810 ;
      LAYER met2 ;
        RECT 1559.730 996.000 1560.010 999.870 ;
      LAYER met2 ;
        RECT 1560.290 995.720 1561.750 998.810 ;
      LAYER met2 ;
        RECT 1562.030 996.000 1562.310 1000.000 ;
        RECT 1562.780 999.870 1564.610 1000.000 ;
      LAYER met2 ;
        RECT 1562.590 995.720 1564.050 998.810 ;
      LAYER met2 ;
        RECT 1564.330 996.000 1564.610 999.870 ;
        RECT 1566.630 999.870 1567.980 1000.000 ;
        RECT 1568.300 1000.010 1568.440 1009.130 ;
        RECT 1574.680 1007.770 1574.940 1008.090 ;
        RECT 1574.740 1000.010 1574.880 1007.770 ;
        RECT 1576.580 1000.010 1576.720 1010.150 ;
        RECT 1576.980 1009.810 1577.240 1010.130 ;
        RECT 1568.300 1000.000 1568.600 1000.010 ;
        RECT 1573.200 1000.000 1574.880 1000.010 ;
        RECT 1575.500 1000.000 1576.720 1000.010 ;
        RECT 1568.300 999.870 1568.750 1000.000 ;
      LAYER met2 ;
        RECT 1564.890 995.720 1566.350 998.810 ;
      LAYER met2 ;
        RECT 1566.630 996.000 1566.910 999.870 ;
      LAYER met2 ;
        RECT 1567.190 995.720 1568.190 998.810 ;
      LAYER met2 ;
        RECT 1568.470 996.000 1568.750 999.870 ;
      LAYER met2 ;
        RECT 1569.030 995.720 1570.490 998.810 ;
      LAYER met2 ;
        RECT 1570.770 996.000 1571.050 1000.000 ;
        RECT 1573.070 999.870 1574.880 1000.000 ;
        RECT 1575.370 999.870 1576.720 1000.000 ;
        RECT 1577.040 1000.010 1577.180 1009.810 ;
        RECT 1577.960 1000.010 1578.100 1013.890 ;
        RECT 1578.420 1008.770 1578.560 1013.890 ;
        RECT 1579.800 1010.470 1579.940 2485.750 ;
        RECT 1580.260 1010.470 1580.400 2494.590 ;
        RECT 1586.700 1023.810 1586.840 2494.590 ;
        RECT 1587.620 2486.410 1587.760 2500.000 ;
        RECT 1607.340 2494.930 1607.600 2495.250 ;
        RECT 1600.440 2489.490 1600.700 2489.810 ;
        RECT 1587.560 2486.090 1587.820 2486.410 ;
        RECT 1585.320 1023.670 1586.840 1023.810 ;
        RECT 1579.740 1010.150 1580.000 1010.470 ;
        RECT 1580.200 1010.150 1580.460 1010.470 ;
        RECT 1578.360 1008.450 1578.620 1008.770 ;
        RECT 1585.320 1000.010 1585.460 1023.670 ;
        RECT 1600.500 1013.870 1600.640 2489.490 ;
        RECT 1591.700 1013.550 1591.960 1013.870 ;
        RECT 1596.300 1013.550 1596.560 1013.870 ;
        RECT 1600.440 1013.550 1600.700 1013.870 ;
        RECT 1585.720 1010.150 1585.980 1010.470 ;
        RECT 1577.040 1000.000 1577.340 1000.010 ;
        RECT 1577.960 1000.000 1579.640 1000.010 ;
        RECT 1583.780 1000.000 1585.460 1000.010 ;
        RECT 1577.040 999.870 1577.490 1000.000 ;
        RECT 1577.960 999.870 1579.790 1000.000 ;
      LAYER met2 ;
        RECT 1571.330 995.720 1572.790 998.810 ;
      LAYER met2 ;
        RECT 1573.070 996.000 1573.350 999.870 ;
      LAYER met2 ;
        RECT 1573.630 995.720 1575.090 998.810 ;
      LAYER met2 ;
        RECT 1575.370 996.000 1575.650 999.870 ;
      LAYER met2 ;
        RECT 1575.930 995.720 1576.930 998.810 ;
      LAYER met2 ;
        RECT 1577.210 996.000 1577.490 999.870 ;
      LAYER met2 ;
        RECT 1577.770 995.720 1579.230 998.810 ;
      LAYER met2 ;
        RECT 1579.510 996.000 1579.790 999.870 ;
      LAYER met2 ;
        RECT 1580.070 995.720 1581.530 998.810 ;
      LAYER met2 ;
        RECT 1581.810 996.000 1582.090 1000.000 ;
        RECT 1583.650 999.870 1585.460 1000.000 ;
        RECT 1585.780 1000.010 1585.920 1010.150 ;
        RECT 1591.760 1010.130 1591.900 1013.550 ;
        RECT 1593.080 1010.150 1593.340 1010.470 ;
        RECT 1591.700 1009.810 1591.960 1010.130 ;
        RECT 1593.140 1000.010 1593.280 1010.150 ;
        RECT 1596.360 1000.010 1596.500 1013.550 ;
        RECT 1603.200 1009.810 1603.460 1010.130 ;
        RECT 1602.740 1009.130 1603.000 1009.450 ;
        RECT 1602.800 1000.010 1602.940 1009.130 ;
        RECT 1585.780 1000.000 1586.080 1000.010 ;
        RECT 1592.520 1000.000 1593.280 1000.010 ;
        RECT 1594.820 1000.000 1596.500 1000.010 ;
        RECT 1601.260 1000.000 1602.940 1000.010 ;
        RECT 1585.780 999.870 1586.230 1000.000 ;
      LAYER met2 ;
        RECT 1582.370 995.720 1583.370 998.810 ;
      LAYER met2 ;
        RECT 1583.650 996.000 1583.930 999.870 ;
      LAYER met2 ;
        RECT 1584.210 995.720 1585.670 998.810 ;
      LAYER met2 ;
        RECT 1585.950 996.000 1586.230 999.870 ;
      LAYER met2 ;
        RECT 1586.510 995.720 1587.970 998.810 ;
      LAYER met2 ;
        RECT 1588.250 996.000 1588.530 1000.000 ;
      LAYER met2 ;
        RECT 1588.810 995.720 1590.270 998.810 ;
      LAYER met2 ;
        RECT 1590.550 996.000 1590.830 1000.000 ;
        RECT 1592.390 999.870 1593.280 1000.000 ;
        RECT 1594.690 999.870 1596.500 1000.000 ;
      LAYER met2 ;
        RECT 1591.110 995.720 1592.110 998.810 ;
      LAYER met2 ;
        RECT 1592.390 996.000 1592.670 999.870 ;
      LAYER met2 ;
        RECT 1592.950 995.720 1594.410 998.810 ;
      LAYER met2 ;
        RECT 1594.690 996.000 1594.970 999.870 ;
      LAYER met2 ;
        RECT 1595.250 995.720 1596.710 998.810 ;
      LAYER met2 ;
        RECT 1596.990 996.000 1597.270 1000.000 ;
      LAYER met2 ;
        RECT 1597.550 995.720 1599.010 998.810 ;
      LAYER met2 ;
        RECT 1599.290 996.000 1599.570 1000.000 ;
        RECT 1601.130 999.870 1602.940 1000.000 ;
        RECT 1603.260 1000.010 1603.400 1009.810 ;
        RECT 1607.400 1009.450 1607.540 2494.930 ;
        RECT 1608.780 2485.730 1608.920 2500.000 ;
        RECT 1608.720 2485.410 1608.980 2485.730 ;
        RECT 1608.720 2484.730 1608.980 2485.050 ;
        RECT 1607.340 1009.130 1607.600 1009.450 ;
        RECT 1608.780 1000.010 1608.920 2484.730 ;
        RECT 1619.820 2484.710 1619.960 2500.000 ;
        RECT 1621.140 2495.270 1621.400 2495.590 ;
        RECT 1619.760 2484.390 1620.020 2484.710 ;
        RECT 1614.700 1016.610 1614.960 1016.930 ;
        RECT 1614.760 1012.170 1614.900 1016.610 ;
        RECT 1614.700 1011.850 1614.960 1012.170 ;
        RECT 1613.780 1009.130 1614.040 1009.450 ;
        RECT 1613.840 1000.010 1613.980 1009.130 ;
        RECT 1620.220 1007.430 1620.480 1007.750 ;
        RECT 1620.280 1000.010 1620.420 1007.430 ;
        RECT 1621.200 1000.010 1621.340 2495.270 ;
        RECT 1629.940 2485.390 1630.080 2500.000 ;
        RECT 1635.460 2499.950 1641.050 2500.000 ;
        RECT 1656.160 2499.950 1662.210 2500.000 ;
        RECT 1629.880 2485.070 1630.140 2485.390 ;
        RECT 1625.740 1015.930 1626.000 1016.250 ;
        RECT 1603.260 1000.000 1603.560 1000.010 ;
        RECT 1608.780 1000.000 1610.000 1000.010 ;
        RECT 1612.300 1000.000 1613.980 1000.010 ;
        RECT 1618.740 1000.000 1620.420 1000.010 ;
        RECT 1621.040 1000.000 1621.340 1000.010 ;
        RECT 1625.800 1000.010 1625.940 1015.930 ;
        RECT 1628.500 1013.210 1628.760 1013.530 ;
        RECT 1628.560 1000.010 1628.700 1013.210 ;
        RECT 1635.460 1007.750 1635.600 2499.950 ;
        RECT 1652.420 2484.050 1652.680 2484.370 ;
        RECT 1652.480 1009.790 1652.620 2484.050 ;
        RECT 1656.160 1016.590 1656.300 2499.950 ;
        RECT 1683.300 2484.370 1683.440 2500.000 ;
        RECT 1693.820 2489.150 1694.080 2489.470 ;
        RECT 1686.920 2486.090 1687.180 2486.410 ;
        RECT 1683.240 2484.050 1683.500 2484.370 ;
        RECT 1669.440 1814.590 1669.700 1814.910 ;
        RECT 1668.980 1735.030 1669.240 1735.350 ;
        RECT 1656.100 1016.270 1656.360 1016.590 ;
        RECT 1665.760 1013.550 1666.020 1013.870 ;
        RECT 1662.540 1011.850 1662.800 1012.170 ;
        RECT 1652.420 1009.470 1652.680 1009.790 ;
        RECT 1635.400 1007.430 1635.660 1007.750 ;
        RECT 1662.600 1000.010 1662.740 1011.850 ;
        RECT 1665.820 1000.010 1665.960 1013.550 ;
        RECT 1669.040 1001.370 1669.180 1735.030 ;
        RECT 1669.500 1013.870 1669.640 1814.590 ;
        RECT 1669.440 1013.550 1669.700 1013.870 ;
        RECT 1686.980 1010.470 1687.120 2486.090 ;
        RECT 1693.880 1013.190 1694.020 2489.150 ;
        RECT 1700.720 2484.050 1700.980 2484.370 ;
        RECT 1693.820 1012.870 1694.080 1013.190 ;
        RECT 1700.780 1010.810 1700.920 2484.050 ;
        RECT 1704.460 1021.350 1704.600 2500.000 ;
        RECT 1715.500 2484.370 1715.640 2500.000 ;
        RECT 1725.620 2487.090 1725.760 2500.000 ;
        RECT 1725.560 2486.770 1725.820 2487.090 ;
        RECT 1746.780 2486.070 1746.920 2500.000 ;
        RECT 1757.820 2486.750 1757.960 2500.000 ;
        RECT 1766.560 2499.950 1768.010 2500.000 ;
        RECT 1757.760 2486.430 1758.020 2486.750 ;
        RECT 1746.720 2485.750 1746.980 2486.070 ;
        RECT 1715.440 2484.050 1715.700 2484.370 ;
        RECT 1724.640 1928.830 1724.900 1929.150 ;
        RECT 1717.740 1925.770 1718.000 1926.090 ;
        RECT 1710.840 1736.390 1711.100 1736.710 ;
        RECT 1704.400 1021.030 1704.660 1021.350 ;
        RECT 1710.900 1013.190 1711.040 1736.390 ;
        RECT 1717.800 1013.190 1717.940 1925.770 ;
        RECT 1720.040 1013.210 1720.300 1013.530 ;
        RECT 1707.160 1012.870 1707.420 1013.190 ;
        RECT 1710.840 1012.870 1711.100 1013.190 ;
        RECT 1715.440 1012.870 1715.700 1013.190 ;
        RECT 1717.740 1012.870 1718.000 1013.190 ;
        RECT 1700.720 1010.490 1700.980 1010.810 ;
        RECT 1686.920 1010.150 1687.180 1010.470 ;
        RECT 1668.580 1001.230 1669.180 1001.370 ;
        RECT 1668.580 1000.690 1668.720 1001.230 ;
        RECT 1668.120 1000.550 1668.720 1000.690 ;
        RECT 1668.120 1000.010 1668.260 1000.550 ;
        RECT 1707.220 1000.010 1707.360 1012.870 ;
        RECT 1710.840 1010.490 1711.100 1010.810 ;
        RECT 1710.900 1000.010 1711.040 1010.490 ;
        RECT 1715.500 1000.010 1715.640 1012.870 ;
        RECT 1720.100 1000.010 1720.240 1013.210 ;
        RECT 1724.700 1000.010 1724.840 1928.830 ;
        RECT 1745.340 1927.470 1745.600 1927.790 ;
        RECT 1738.440 1926.110 1738.700 1926.430 ;
        RECT 1737.980 1849.270 1738.240 1849.590 ;
        RECT 1728.780 1021.030 1729.040 1021.350 ;
        RECT 1728.840 1000.010 1728.980 1021.030 ;
        RECT 1738.040 1013.190 1738.180 1849.270 ;
        RECT 1733.380 1012.870 1733.640 1013.190 ;
        RECT 1737.980 1012.870 1738.240 1013.190 ;
        RECT 1733.440 1000.010 1733.580 1012.870 ;
        RECT 1738.500 1000.690 1738.640 1926.110 ;
        RECT 1738.900 1012.870 1739.160 1013.190 ;
        RECT 1738.960 1010.810 1739.100 1012.870 ;
        RECT 1738.900 1010.490 1739.160 1010.810 ;
        RECT 1741.660 1010.490 1741.920 1010.810 ;
        RECT 1737.580 1000.550 1738.640 1000.690 ;
        RECT 1737.580 1000.010 1737.720 1000.550 ;
        RECT 1741.720 1000.010 1741.860 1010.490 ;
        RECT 1745.400 1000.010 1745.540 1927.470 ;
        RECT 1766.040 1926.450 1766.300 1926.770 ;
        RECT 1759.140 1883.610 1759.400 1883.930 ;
        RECT 1752.240 1736.730 1752.500 1737.050 ;
        RECT 1752.300 1010.470 1752.440 1736.730 ;
        RECT 1759.200 1013.870 1759.340 1883.610 ;
        RECT 1755.000 1013.550 1755.260 1013.870 ;
        RECT 1759.140 1013.550 1759.400 1013.870 ;
        RECT 1759.600 1013.550 1759.860 1013.870 ;
        RECT 1749.940 1010.150 1750.200 1010.470 ;
        RECT 1752.240 1010.150 1752.500 1010.470 ;
        RECT 1750.000 1000.010 1750.140 1010.150 ;
        RECT 1755.060 1000.010 1755.200 1013.550 ;
        RECT 1759.660 1010.810 1759.800 1013.550 ;
        RECT 1759.600 1010.490 1759.860 1010.810 ;
        RECT 1766.100 1010.470 1766.240 1926.450 ;
        RECT 1766.560 1017.270 1766.700 2499.950 ;
        RECT 1778.980 2486.410 1779.120 2500.000 ;
        RECT 1790.020 2489.810 1790.160 2500.000 ;
        RECT 1789.960 2489.490 1790.220 2489.810 ;
        RECT 1811.180 2489.470 1811.320 2500.000 ;
        RECT 1811.120 2489.150 1811.380 2489.470 ;
        RECT 1832.340 2488.110 1832.480 2500.000 ;
        RECT 1842.460 2489.130 1842.600 2500.000 ;
        RECT 1849.360 2499.950 1853.570 2500.000 ;
        RECT 1842.400 2488.810 1842.660 2489.130 ;
        RECT 1832.280 2487.790 1832.540 2488.110 ;
        RECT 1778.920 2486.090 1779.180 2486.410 ;
        RECT 1845.620 1927.810 1845.880 1928.130 ;
        RECT 1779.380 1927.130 1779.640 1927.450 ;
        RECT 1772.940 1766.310 1773.200 1766.630 ;
        RECT 1772.480 1735.710 1772.740 1736.030 ;
        RECT 1766.500 1016.950 1766.760 1017.270 ;
        RECT 1767.880 1010.490 1768.140 1010.810 ;
        RECT 1763.740 1010.150 1764.000 1010.470 ;
        RECT 1766.040 1010.150 1766.300 1010.470 ;
        RECT 1758.680 1009.810 1758.940 1010.130 ;
        RECT 1758.740 1000.010 1758.880 1009.810 ;
        RECT 1763.800 1000.010 1763.940 1010.150 ;
        RECT 1767.940 1000.010 1768.080 1010.490 ;
        RECT 1772.540 1000.010 1772.680 1735.710 ;
        RECT 1773.000 1010.810 1773.140 1766.310 ;
        RECT 1772.940 1010.490 1773.200 1010.810 ;
        RECT 1776.620 1007.430 1776.880 1007.750 ;
        RECT 1776.680 1000.010 1776.820 1007.430 ;
        RECT 1625.800 1000.000 1627.480 1000.010 ;
        RECT 1628.560 1000.000 1629.780 1000.010 ;
        RECT 1662.440 1000.000 1662.740 1000.010 ;
        RECT 1664.280 1000.000 1665.960 1000.010 ;
        RECT 1666.580 1000.000 1668.260 1000.010 ;
        RECT 1705.680 1000.000 1707.360 1000.010 ;
        RECT 1710.280 1000.000 1711.040 1000.010 ;
        RECT 1714.420 1000.000 1715.640 1000.010 ;
        RECT 1718.560 1000.000 1720.240 1000.010 ;
        RECT 1723.160 1000.000 1724.840 1000.010 ;
        RECT 1727.300 1000.000 1728.980 1000.010 ;
        RECT 1731.900 1000.000 1733.580 1000.010 ;
        RECT 1736.040 1000.000 1737.720 1000.010 ;
        RECT 1740.640 1000.000 1741.860 1000.010 ;
        RECT 1744.780 1000.000 1745.540 1000.010 ;
        RECT 1749.380 1000.000 1750.140 1000.010 ;
        RECT 1753.520 1000.000 1755.200 1000.010 ;
        RECT 1758.120 1000.000 1758.880 1000.010 ;
        RECT 1762.260 1000.000 1763.940 1000.010 ;
        RECT 1766.400 1000.000 1768.080 1000.010 ;
        RECT 1771.000 1000.000 1772.680 1000.010 ;
        RECT 1775.140 1000.000 1776.820 1000.010 ;
        RECT 1779.440 1000.010 1779.580 1927.130 ;
        RECT 1786.740 1926.790 1787.000 1927.110 ;
        RECT 1779.840 1925.430 1780.100 1925.750 ;
        RECT 1779.900 1007.750 1780.040 1925.430 ;
        RECT 1779.840 1007.430 1780.100 1007.750 ;
        RECT 1786.800 1000.690 1786.940 1926.790 ;
        RECT 1835.040 1925.090 1835.300 1925.410 ;
        RECT 1821.240 1870.010 1821.500 1870.330 ;
        RECT 1800.540 1738.090 1800.800 1738.410 ;
        RECT 1793.640 1737.410 1793.900 1737.730 ;
        RECT 1789.500 1009.470 1789.760 1009.790 ;
        RECT 1785.420 1000.550 1786.940 1000.690 ;
        RECT 1785.420 1000.010 1785.560 1000.550 ;
        RECT 1789.560 1000.010 1789.700 1009.470 ;
        RECT 1793.700 1000.010 1793.840 1737.410 ;
        RECT 1800.600 1007.750 1800.740 1738.090 ;
        RECT 1814.340 1737.750 1814.600 1738.070 ;
        RECT 1813.880 1737.070 1814.140 1737.390 ;
        RECT 1807.440 1736.050 1807.700 1736.370 ;
        RECT 1806.980 1735.370 1807.240 1735.690 ;
        RECT 1807.040 1007.750 1807.180 1735.370 ;
        RECT 1798.240 1007.430 1798.500 1007.750 ;
        RECT 1800.540 1007.430 1800.800 1007.750 ;
        RECT 1802.840 1007.430 1803.100 1007.750 ;
        RECT 1806.980 1007.430 1807.240 1007.750 ;
        RECT 1798.300 1000.010 1798.440 1007.430 ;
        RECT 1802.900 1000.010 1803.040 1007.430 ;
        RECT 1807.500 1000.690 1807.640 1736.050 ;
        RECT 1813.940 1007.750 1814.080 1737.070 ;
        RECT 1811.580 1007.430 1811.840 1007.750 ;
        RECT 1813.880 1007.430 1814.140 1007.750 ;
        RECT 1807.040 1000.550 1807.640 1000.690 ;
        RECT 1807.040 1000.010 1807.180 1000.550 ;
        RECT 1811.640 1000.010 1811.780 1007.430 ;
        RECT 1814.400 1000.010 1814.540 1737.750 ;
        RECT 1821.300 1000.690 1821.440 1870.010 ;
        RECT 1835.100 1010.810 1835.240 1925.090 ;
        RECT 1830.900 1010.490 1831.160 1010.810 ;
        RECT 1835.040 1010.490 1835.300 1010.810 ;
        RECT 1826.760 1009.810 1827.020 1010.130 ;
        RECT 1824.460 1008.450 1824.720 1008.770 ;
        RECT 1820.380 1000.550 1821.440 1000.690 ;
        RECT 1820.380 1000.010 1820.520 1000.550 ;
        RECT 1824.520 1000.010 1824.660 1008.450 ;
        RECT 1826.820 1000.010 1826.960 1009.810 ;
        RECT 1830.960 1000.010 1831.100 1010.490 ;
        RECT 1845.680 1010.130 1845.820 1927.810 ;
        RECT 1849.360 1018.290 1849.500 2499.950 ;
        RECT 1874.660 2488.450 1874.800 2500.000 ;
        RECT 1885.700 2488.790 1885.840 2500.000 ;
        RECT 1885.640 2488.470 1885.900 2488.790 ;
        RECT 1874.600 2488.130 1874.860 2488.450 ;
        RECT 1876.440 1935.290 1876.700 1935.610 ;
        RECT 1849.300 1017.970 1849.560 1018.290 ;
        RECT 1866.320 1012.530 1866.580 1012.850 ;
        RECT 1866.380 1011.830 1866.520 1012.530 ;
        RECT 1876.500 1012.510 1876.640 1935.290 ;
        RECT 1886.160 1014.210 1886.300 2896.390 ;
        RECT 1886.550 2828.955 1886.830 2829.325 ;
        RECT 1886.620 1018.970 1886.760 2828.955 ;
        RECT 1887.010 2815.355 1887.290 2815.725 ;
        RECT 1887.080 1019.990 1887.220 2815.355 ;
        RECT 1890.690 2800.735 1890.970 2801.105 ;
        RECT 1887.470 2782.715 1887.750 2783.085 ;
        RECT 1887.020 1019.670 1887.280 1019.990 ;
        RECT 1886.560 1018.650 1886.820 1018.970 ;
        RECT 1886.100 1013.890 1886.360 1014.210 ;
        RECT 1887.540 1012.850 1887.680 2782.715 ;
        RECT 1887.480 1012.530 1887.740 1012.850 ;
        RECT 1872.300 1012.190 1872.560 1012.510 ;
        RECT 1876.440 1012.190 1876.700 1012.510 ;
        RECT 1865.860 1011.510 1866.120 1011.830 ;
        RECT 1866.320 1011.510 1866.580 1011.830 ;
        RECT 1865.920 1010.810 1866.060 1011.510 ;
        RECT 1865.860 1010.490 1866.120 1010.810 ;
        RECT 1845.620 1009.810 1845.880 1010.130 ;
        RECT 1834.580 1008.790 1834.840 1009.110 ;
        RECT 1834.640 1000.010 1834.780 1008.790 ;
        RECT 1872.360 1000.010 1872.500 1012.190 ;
        RECT 1890.760 1011.490 1890.900 2800.735 ;
        RECT 1891.150 2753.135 1891.430 2753.505 ;
        RECT 1890.700 1011.170 1890.960 1011.490 ;
        RECT 1873.220 1010.830 1873.480 1011.150 ;
        RECT 1873.280 1008.430 1873.420 1010.830 ;
        RECT 1883.340 1010.490 1883.600 1010.810 ;
        RECT 1878.740 1009.810 1879.000 1010.130 ;
        RECT 1873.220 1008.110 1873.480 1008.430 ;
        RECT 1878.800 1000.010 1878.940 1009.810 ;
        RECT 1883.400 1000.010 1883.540 1010.490 ;
        RECT 1891.220 1009.450 1891.360 2753.135 ;
        RECT 1891.610 2738.175 1891.890 2738.545 ;
        RECT 1891.680 1011.150 1891.820 2738.175 ;
        RECT 1892.140 2495.590 1892.280 2912.790 ;
        RECT 1893.460 2912.450 1893.720 2912.770 ;
        RECT 1893.000 2911.770 1893.260 2912.090 ;
        RECT 1892.540 2896.470 1892.800 2896.790 ;
        RECT 1892.080 2495.270 1892.340 2495.590 ;
        RECT 1892.600 2495.250 1892.740 2896.470 ;
        RECT 1892.540 2494.930 1892.800 2495.250 ;
        RECT 1893.060 2494.230 1893.200 2911.770 ;
        RECT 1893.520 2494.570 1893.660 2912.450 ;
        RECT 1893.920 2780.870 1894.180 2781.190 ;
        RECT 1893.460 2494.250 1893.720 2494.570 ;
        RECT 1893.000 2493.910 1893.260 2494.230 ;
        RECT 1891.620 1010.830 1891.880 1011.150 ;
        RECT 1893.980 1010.130 1894.120 2780.870 ;
        RECT 1894.440 2494.910 1894.580 2913.130 ;
        RECT 1897.590 2845.275 1897.870 2845.645 ;
        RECT 1894.830 2577.355 1895.110 2577.725 ;
        RECT 1894.380 2494.590 1894.640 2494.910 ;
        RECT 1894.900 1011.830 1895.040 2577.355 ;
        RECT 1897.660 1017.610 1897.800 2845.275 ;
        RECT 2100.920 2781.210 2101.180 2781.530 ;
        RECT 2556.320 2781.210 2556.580 2781.530 ;
        RECT 1898.050 2767.075 1898.330 2767.445 ;
        RECT 1898.120 1020.670 1898.260 2767.075 ;
        RECT 1898.510 2718.795 1898.790 2719.165 ;
        RECT 1898.060 1020.350 1898.320 1020.670 ;
        RECT 1898.580 1018.630 1898.720 2718.795 ;
        RECT 1898.970 2687.515 1899.250 2687.885 ;
        RECT 1899.040 1019.650 1899.180 2687.515 ;
        RECT 1899.430 2672.555 1899.710 2672.925 ;
        RECT 1898.980 1019.330 1899.240 1019.650 ;
        RECT 1899.500 1019.310 1899.640 2672.555 ;
        RECT 1899.890 2656.915 1900.170 2657.285 ;
        RECT 1899.440 1018.990 1899.700 1019.310 ;
        RECT 1898.520 1018.310 1898.780 1018.630 ;
        RECT 1899.960 1017.950 1900.100 2656.915 ;
        RECT 1900.350 2624.955 1900.630 2625.325 ;
        RECT 1899.900 1017.630 1900.160 1017.950 ;
        RECT 1897.600 1017.290 1897.860 1017.610 ;
        RECT 1894.840 1011.510 1895.100 1011.830 ;
        RECT 1893.920 1009.810 1894.180 1010.130 ;
        RECT 1891.160 1009.130 1891.420 1009.450 ;
        RECT 1900.420 1008.430 1900.560 2624.955 ;
        RECT 1900.810 2608.635 1901.090 2609.005 ;
        RECT 1900.880 1016.930 1901.020 2608.635 ;
        RECT 1901.270 2562.395 1901.550 2562.765 ;
        RECT 1900.820 1016.610 1901.080 1016.930 ;
        RECT 1900.360 1008.110 1900.620 1008.430 ;
        RECT 1901.340 1008.090 1901.480 2562.395 ;
        RECT 1901.730 2546.755 1902.010 2547.125 ;
        RECT 1901.800 1020.330 1901.940 2546.755 ;
        RECT 1903.570 2514.795 1903.850 2515.165 ;
        RECT 1903.640 2504.090 1903.780 2514.795 ;
        RECT 1902.200 2503.770 1902.460 2504.090 ;
        RECT 1903.580 2503.770 1903.840 2504.090 ;
        RECT 1902.260 1021.010 1902.400 2503.770 ;
        RECT 2082.980 1946.850 2083.240 1947.170 ;
        RECT 2073.320 1946.510 2073.580 1946.830 ;
        RECT 2044.340 1928.830 2044.600 1929.150 ;
        RECT 1964.300 1927.810 1964.560 1928.130 ;
        RECT 1929.340 1927.470 1929.600 1927.790 ;
        RECT 1929.400 1917.095 1929.540 1927.470 ;
        RECT 1952.340 1925.090 1952.600 1925.410 ;
        RECT 1952.400 1917.095 1952.540 1925.090 ;
        RECT 1964.360 1917.095 1964.500 1927.810 ;
        RECT 1998.340 1927.130 1998.600 1927.450 ;
        RECT 1987.300 1926.110 1987.560 1926.430 ;
        RECT 1975.340 1925.770 1975.600 1926.090 ;
        RECT 1975.400 1917.095 1975.540 1925.770 ;
        RECT 1987.360 1917.095 1987.500 1926.110 ;
        RECT 1998.400 1917.095 1998.540 1927.130 ;
        RECT 2033.300 1926.790 2033.560 1927.110 ;
        RECT 2010.300 1926.450 2010.560 1926.770 ;
        RECT 2010.360 1917.095 2010.500 1926.450 ;
        RECT 2033.360 1917.095 2033.500 1926.790 ;
        RECT 2044.400 1917.095 2044.540 1928.830 ;
        RECT 2067.340 1925.430 2067.600 1925.750 ;
        RECT 2067.400 1917.095 2067.540 1925.430 ;
        RECT 1929.290 1913.095 1929.570 1917.095 ;
        RECT 1952.290 1913.095 1952.570 1917.095 ;
        RECT 1964.250 1913.095 1964.530 1917.095 ;
        RECT 1975.290 1913.095 1975.570 1917.095 ;
        RECT 1987.250 1913.095 1987.530 1917.095 ;
        RECT 1998.290 1913.095 1998.570 1917.095 ;
        RECT 2010.250 1913.095 2010.530 1917.095 ;
        RECT 2033.250 1913.095 2033.530 1917.095 ;
        RECT 2044.290 1913.095 2044.570 1917.095 ;
        RECT 2067.290 1913.095 2067.570 1917.095 ;
      LAYER met2 ;
        RECT 1922.860 1912.815 1929.010 1913.095 ;
        RECT 1929.850 1912.815 1940.970 1913.095 ;
        RECT 1941.810 1912.815 1952.010 1913.095 ;
        RECT 1952.850 1912.815 1963.970 1913.095 ;
        RECT 1964.810 1912.815 1975.010 1913.095 ;
        RECT 1975.850 1912.815 1986.970 1913.095 ;
        RECT 1987.810 1912.815 1998.010 1913.095 ;
        RECT 1998.850 1912.815 2009.970 1913.095 ;
        RECT 2010.810 1912.815 2021.010 1913.095 ;
        RECT 2021.850 1912.815 2032.970 1913.095 ;
        RECT 2033.810 1912.815 2044.010 1913.095 ;
        RECT 2044.850 1912.815 2055.970 1913.095 ;
        RECT 2056.810 1912.815 2067.010 1913.095 ;
        RECT 2067.850 1912.815 2072.160 1913.095 ;
      LAYER met2 ;
        RECT 1904.490 1885.795 1904.770 1886.165 ;
        RECT 1904.560 1883.930 1904.700 1885.795 ;
        RECT 1904.500 1883.610 1904.760 1883.930 ;
        RECT 1904.490 1870.155 1904.770 1870.525 ;
        RECT 1904.500 1870.010 1904.760 1870.155 ;
        RECT 1904.490 1851.795 1904.770 1852.165 ;
        RECT 1904.560 1849.590 1904.700 1851.795 ;
        RECT 1904.500 1849.270 1904.760 1849.590 ;
        RECT 1904.490 1817.795 1904.770 1818.165 ;
        RECT 1904.560 1814.910 1904.700 1817.795 ;
        RECT 1904.500 1814.590 1904.760 1814.910 ;
        RECT 1904.490 1767.475 1904.770 1767.845 ;
        RECT 1904.560 1766.630 1904.700 1767.475 ;
        RECT 1904.500 1766.310 1904.760 1766.630 ;
      LAYER met2 ;
        RECT 1922.860 1754.280 2072.160 1912.815 ;
        RECT 1923.410 1754.000 1933.610 1754.280 ;
        RECT 1934.450 1754.000 1944.650 1754.280 ;
        RECT 1945.490 1754.000 1956.610 1754.280 ;
        RECT 1957.450 1754.000 1967.650 1754.280 ;
        RECT 1968.490 1754.000 1979.610 1754.280 ;
        RECT 1980.450 1754.000 1990.650 1754.280 ;
        RECT 1991.490 1754.000 2002.610 1754.280 ;
        RECT 2003.450 1754.000 2013.650 1754.280 ;
        RECT 2014.490 1754.000 2025.610 1754.280 ;
        RECT 2026.450 1754.000 2036.650 1754.280 ;
        RECT 2037.490 1754.000 2048.610 1754.280 ;
        RECT 2049.450 1754.000 2059.650 1754.280 ;
        RECT 2060.490 1754.000 2071.610 1754.280 ;
      LAYER met2 ;
        RECT 1933.890 1750.000 1934.170 1754.000 ;
        RECT 1944.930 1750.000 1945.210 1754.000 ;
        RECT 1956.890 1750.000 1957.170 1754.000 ;
        RECT 1967.930 1750.000 1968.210 1754.000 ;
        RECT 1979.890 1750.000 1980.170 1754.000 ;
        RECT 1990.930 1750.000 1991.210 1754.000 ;
        RECT 2002.890 1750.000 2003.170 1754.000 ;
        RECT 2013.930 1750.000 2014.210 1754.000 ;
        RECT 2036.930 1750.000 2037.210 1754.000 ;
        RECT 2059.930 1750.000 2060.210 1754.000 ;
        RECT 2071.890 1750.000 2072.170 1754.000 ;
        RECT 1934.000 1738.750 1934.140 1750.000 ;
        RECT 1907.720 1738.430 1907.980 1738.750 ;
        RECT 1933.940 1738.430 1934.200 1738.750 ;
        RECT 1902.200 1020.690 1902.460 1021.010 ;
        RECT 1901.740 1020.010 1902.000 1020.330 ;
        RECT 1907.780 1008.770 1907.920 1738.430 ;
        RECT 1945.040 1736.710 1945.180 1750.000 ;
        RECT 1957.000 1738.410 1957.140 1750.000 ;
        RECT 1956.940 1738.090 1957.200 1738.410 ;
        RECT 1968.040 1737.730 1968.180 1750.000 ;
        RECT 1967.980 1737.410 1968.240 1737.730 ;
        RECT 1980.000 1737.050 1980.140 1750.000 ;
        RECT 1991.040 1738.070 1991.180 1750.000 ;
        RECT 1990.980 1737.750 1991.240 1738.070 ;
        RECT 1979.940 1736.730 1980.200 1737.050 ;
        RECT 1944.980 1736.390 1945.240 1736.710 ;
        RECT 2003.000 1736.030 2003.140 1750.000 ;
        RECT 2014.040 1737.390 2014.180 1750.000 ;
        RECT 2013.980 1737.070 2014.240 1737.390 ;
        RECT 2037.040 1736.370 2037.180 1750.000 ;
        RECT 2036.980 1736.050 2037.240 1736.370 ;
        RECT 2002.940 1735.710 2003.200 1736.030 ;
        RECT 2060.040 1735.350 2060.180 1750.000 ;
        RECT 2072.000 1735.690 2072.140 1750.000 ;
        RECT 2071.940 1735.370 2072.200 1735.690 ;
        RECT 2059.980 1735.030 2060.240 1735.350 ;
        RECT 2007.540 1687.770 2007.800 1688.090 ;
        RECT 2007.600 1014.210 2007.740 1687.770 ;
        RECT 2055.840 1687.430 2056.100 1687.750 ;
        RECT 2042.040 1687.090 2042.300 1687.410 ;
        RECT 2002.940 1013.890 2003.200 1014.210 ;
        RECT 2007.540 1013.890 2007.800 1014.210 ;
        RECT 1907.720 1008.450 1907.980 1008.770 ;
        RECT 1901.280 1007.770 1901.540 1008.090 ;
        RECT 2003.000 1000.010 2003.140 1013.890 ;
        RECT 2004.780 1012.530 2005.040 1012.850 ;
        RECT 2004.840 1000.010 2004.980 1012.530 ;
        RECT 2042.100 1000.010 2042.240 1687.090 ;
        RECT 2055.380 1010.830 2055.640 1011.150 ;
        RECT 2046.180 1009.130 2046.440 1009.450 ;
        RECT 2046.240 1000.010 2046.380 1009.130 ;
        RECT 2050.780 1008.450 2051.040 1008.770 ;
        RECT 2050.840 1000.010 2050.980 1008.450 ;
        RECT 1779.440 1000.000 1779.740 1000.010 ;
        RECT 1783.880 1000.000 1785.560 1000.010 ;
        RECT 1788.480 1000.000 1789.700 1000.010 ;
        RECT 1792.620 1000.000 1793.840 1000.010 ;
        RECT 1797.220 1000.000 1798.440 1000.010 ;
        RECT 1801.360 1000.000 1803.040 1000.010 ;
        RECT 1805.960 1000.000 1807.180 1000.010 ;
        RECT 1810.100 1000.000 1811.780 1000.010 ;
        RECT 1814.240 1000.000 1814.540 1000.010 ;
        RECT 1818.840 1000.000 1820.520 1000.010 ;
        RECT 1822.980 1000.000 1824.660 1000.010 ;
        RECT 1825.280 1000.000 1826.960 1000.010 ;
        RECT 1829.880 1000.000 1831.100 1000.010 ;
        RECT 1834.020 1000.000 1834.780 1000.010 ;
        RECT 1870.820 1000.000 1872.500 1000.010 ;
        RECT 1877.260 1000.000 1878.940 1000.010 ;
        RECT 1881.860 1000.000 1883.540 1000.010 ;
        RECT 2001.460 1000.000 2003.140 1000.010 ;
        RECT 2003.760 1000.000 2004.980 1000.010 ;
        RECT 2040.560 1000.000 2042.240 1000.010 ;
        RECT 2044.700 1000.000 2046.380 1000.010 ;
        RECT 2049.300 1000.000 2050.980 1000.010 ;
        RECT 2055.440 1000.010 2055.580 1010.830 ;
        RECT 2055.900 1008.770 2056.040 1687.430 ;
        RECT 2069.640 1686.750 2069.900 1687.070 ;
        RECT 2061.360 1011.850 2061.620 1012.170 ;
        RECT 2055.840 1008.450 2056.100 1008.770 ;
        RECT 2061.420 1000.010 2061.560 1011.850 ;
        RECT 2065.960 1008.450 2066.220 1008.770 ;
        RECT 2066.020 1000.010 2066.160 1008.450 ;
        RECT 2069.700 1000.010 2069.840 1686.750 ;
        RECT 2073.380 1012.850 2073.520 1946.510 ;
        RECT 2080.220 1870.010 2080.480 1870.330 ;
        RECT 2076.990 1819.495 2077.270 1819.865 ;
        RECT 2077.060 1013.190 2077.200 1819.495 ;
        RECT 2077.000 1012.870 2077.260 1013.190 ;
        RECT 2073.320 1012.530 2073.580 1012.850 ;
        RECT 2078.840 1011.850 2079.100 1012.170 ;
        RECT 2074.700 1011.170 2074.960 1011.490 ;
        RECT 2074.760 1000.010 2074.900 1011.170 ;
        RECT 2078.900 1000.010 2079.040 1011.850 ;
        RECT 2080.280 1008.770 2080.420 1870.010 ;
        RECT 2082.060 1062.510 2082.320 1062.830 ;
        RECT 2080.220 1008.450 2080.480 1008.770 ;
        RECT 2082.120 1000.010 2082.260 1062.510 ;
        RECT 2083.040 1012.170 2083.180 1946.850 ;
        RECT 2090.340 1946.170 2090.600 1946.490 ;
        RECT 2083.440 1945.830 2083.700 1946.150 ;
        RECT 2083.500 1062.830 2083.640 1945.830 ;
        RECT 2083.890 1884.435 2084.170 1884.805 ;
        RECT 2083.440 1062.510 2083.700 1062.830 ;
        RECT 2082.980 1011.850 2083.240 1012.170 ;
        RECT 2083.960 1011.830 2084.100 1884.435 ;
        RECT 2084.350 1850.435 2084.630 1850.805 ;
        RECT 2084.420 1013.530 2084.560 1850.435 ;
        RECT 2084.810 1835.475 2085.090 1835.845 ;
        RECT 2084.360 1013.210 2084.620 1013.530 ;
        RECT 2083.900 1011.510 2084.160 1011.830 ;
        RECT 2084.880 1009.790 2085.020 1835.475 ;
        RECT 2085.270 1800.795 2085.550 1801.165 ;
        RECT 2085.340 1021.350 2085.480 1800.795 ;
        RECT 2085.730 1782.435 2086.010 1782.805 ;
        RECT 2085.280 1021.030 2085.540 1021.350 ;
        RECT 2085.800 1013.870 2085.940 1782.435 ;
        RECT 2086.190 1766.795 2086.470 1767.165 ;
        RECT 2085.740 1013.550 2086.000 1013.870 ;
        RECT 2085.280 1010.830 2085.540 1011.150 ;
        RECT 2084.820 1009.470 2085.080 1009.790 ;
        RECT 2085.340 1009.450 2085.480 1010.830 ;
        RECT 2086.260 1010.470 2086.400 1766.795 ;
        RECT 2090.400 1012.170 2090.540 1946.170 ;
        RECT 2087.580 1011.850 2087.840 1012.170 ;
        RECT 2090.340 1011.850 2090.600 1012.170 ;
        RECT 2086.200 1010.150 2086.460 1010.470 ;
        RECT 2085.280 1009.130 2085.540 1009.450 ;
        RECT 2087.640 1000.010 2087.780 1011.850 ;
        RECT 2100.980 1009.110 2101.120 2781.210 ;
        RECT 2422.000 2780.870 2422.260 2781.190 ;
        RECT 2422.060 2773.820 2422.200 2780.870 ;
        RECT 2556.380 2773.820 2556.520 2781.210 ;
        RECT 2422.060 2773.380 2422.380 2773.820 ;
        RECT 2556.380 2773.380 2556.700 2773.820 ;
        RECT 2422.100 2769.820 2422.380 2773.380 ;
        RECT 2556.420 2769.820 2556.700 2773.380 ;
      LAYER met2 ;
        RECT 2400.030 2769.540 2421.820 2769.820 ;
        RECT 2422.660 2769.540 2556.140 2769.820 ;
        RECT 2400.030 2604.280 2556.690 2769.540 ;
        RECT 2400.580 2604.000 2534.060 2604.280 ;
        RECT 2534.900 2604.000 2556.690 2604.280 ;
      LAYER met2 ;
        RECT 2400.020 2600.730 2400.300 2604.000 ;
        RECT 2534.340 2600.730 2534.620 2604.000 ;
        RECT 2394.460 2600.590 2400.300 2600.730 ;
        RECT 2321.260 1946.850 2321.520 1947.170 ;
        RECT 2321.320 1937.745 2321.460 1946.850 ;
        RECT 2379.220 1946.510 2379.480 1946.830 ;
        RECT 2379.280 1937.745 2379.420 1946.510 ;
        RECT 2321.250 1933.745 2321.530 1937.745 ;
        RECT 2379.210 1933.745 2379.490 1937.745 ;
        RECT 2394.460 1935.610 2394.600 2600.590 ;
        RECT 2400.020 2600.000 2400.300 2600.590 ;
        RECT 2532.460 2600.590 2534.620 2600.730 ;
        RECT 2437.180 1946.170 2437.440 1946.490 ;
        RECT 2437.240 1937.745 2437.380 1946.170 ;
        RECT 2495.140 1945.830 2495.400 1946.150 ;
        RECT 2495.200 1937.745 2495.340 1945.830 ;
        RECT 2394.400 1935.290 2394.660 1935.610 ;
        RECT 2437.170 1933.745 2437.450 1937.745 ;
        RECT 2495.130 1933.745 2495.410 1937.745 ;
      LAYER met2 ;
        RECT 2302.860 1933.465 2320.970 1933.745 ;
        RECT 2321.810 1933.465 2378.930 1933.745 ;
        RECT 2379.770 1933.465 2436.890 1933.745 ;
        RECT 2437.730 1933.465 2494.850 1933.745 ;
        RECT 2495.690 1933.465 2514.720 1933.745 ;
      LAYER met2 ;
        RECT 2283.990 1875.595 2284.270 1875.965 ;
        RECT 2284.060 1870.330 2284.200 1875.595 ;
        RECT 2284.000 1870.010 2284.260 1870.330 ;
        RECT 2287.210 1789.915 2287.490 1790.285 ;
        RECT 2287.280 1012.510 2287.420 1789.915 ;
      LAYER met2 ;
        RECT 2302.860 1704.280 2514.720 1933.465 ;
      LAYER met2 ;
        RECT 2523.650 1892.170 2523.930 1892.285 ;
        RECT 2518.660 1892.030 2523.930 1892.170 ;
        RECT 2518.660 1807.170 2518.800 1892.030 ;
        RECT 2523.650 1891.915 2523.930 1892.030 ;
        RECT 2518.200 1807.030 2518.800 1807.170 ;
        RECT 2518.200 1800.370 2518.340 1807.030 ;
        RECT 2523.650 1802.410 2523.930 1802.525 ;
        RECT 2521.880 1802.270 2523.930 1802.410 ;
        RECT 2518.200 1800.230 2518.800 1800.370 ;
        RECT 2518.660 1799.690 2518.800 1800.230 ;
        RECT 2518.660 1799.550 2519.260 1799.690 ;
        RECT 2519.120 1752.770 2519.260 1799.550 ;
        RECT 2521.880 1759.570 2522.020 1802.270 ;
        RECT 2523.650 1802.155 2523.930 1802.270 ;
        RECT 2520.500 1759.430 2522.020 1759.570 ;
        RECT 2520.500 1752.770 2520.640 1759.430 ;
        RECT 2519.120 1752.630 2520.180 1752.770 ;
        RECT 2520.500 1752.630 2521.100 1752.770 ;
        RECT 2520.040 1724.890 2520.180 1752.630 ;
        RECT 2519.580 1724.750 2520.180 1724.890 ;
        RECT 2519.060 1709.870 2519.320 1710.190 ;
      LAYER met2 ;
        RECT 2303.410 1704.000 2360.530 1704.280 ;
        RECT 2361.370 1704.000 2418.490 1704.280 ;
        RECT 2419.330 1704.000 2476.450 1704.280 ;
        RECT 2477.290 1704.000 2514.720 1704.280 ;
      LAYER met2 ;
        RECT 2518.590 1704.235 2518.870 1704.605 ;
        RECT 2302.850 1700.000 2303.130 1704.000 ;
        RECT 2360.810 1700.000 2361.090 1704.000 ;
        RECT 2418.770 1700.000 2419.050 1704.000 ;
        RECT 2476.730 1700.000 2477.010 1704.000 ;
        RECT 2302.920 1688.090 2303.060 1700.000 ;
        RECT 2302.860 1687.770 2303.120 1688.090 ;
        RECT 2360.880 1687.750 2361.020 1700.000 ;
        RECT 2360.820 1687.430 2361.080 1687.750 ;
        RECT 2418.840 1687.410 2418.980 1700.000 ;
        RECT 2418.780 1687.090 2419.040 1687.410 ;
        RECT 2476.800 1687.070 2476.940 1700.000 ;
        RECT 2476.740 1686.750 2477.000 1687.070 ;
        RECT 2518.660 1656.890 2518.800 1704.235 ;
        RECT 2518.200 1656.750 2518.800 1656.890 ;
        RECT 2518.200 1656.130 2518.340 1656.750 ;
        RECT 2518.140 1655.810 2518.400 1656.130 ;
        RECT 2519.120 1655.530 2519.260 1709.870 ;
        RECT 2519.580 1704.605 2519.720 1724.750 ;
        RECT 2520.960 1710.190 2521.100 1752.630 ;
        RECT 2523.650 1717.835 2523.930 1718.205 ;
        RECT 2520.900 1709.870 2521.160 1710.190 ;
        RECT 2519.510 1704.235 2519.790 1704.605 ;
        RECT 2523.720 1704.410 2523.860 1717.835 ;
        RECT 2523.660 1704.090 2523.920 1704.410 ;
        RECT 2519.520 1703.750 2519.780 1704.070 ;
        RECT 2518.660 1655.390 2519.260 1655.530 ;
        RECT 2518.660 1642.190 2518.800 1655.390 ;
        RECT 2517.680 1641.870 2517.940 1642.190 ;
        RECT 2518.600 1641.870 2518.860 1642.190 ;
        RECT 2517.740 1594.250 2517.880 1641.870 ;
        RECT 2519.580 1608.725 2519.720 1703.750 ;
        RECT 2519.980 1655.810 2520.240 1656.130 ;
        RECT 2520.040 1618.050 2520.180 1655.810 ;
        RECT 2519.980 1617.730 2520.240 1618.050 ;
        RECT 2520.900 1617.730 2521.160 1618.050 ;
        RECT 2519.510 1608.355 2519.790 1608.725 ;
        RECT 2519.510 1606.995 2519.790 1607.365 ;
        RECT 2517.680 1593.930 2517.940 1594.250 ;
        RECT 2518.600 1593.930 2518.860 1594.250 ;
        RECT 2518.660 1569.770 2518.800 1593.930 ;
        RECT 2517.220 1569.450 2517.480 1569.770 ;
        RECT 2518.600 1569.450 2518.860 1569.770 ;
        RECT 2517.280 1545.970 2517.420 1569.450 ;
        RECT 2518.140 1559.250 2518.400 1559.570 ;
        RECT 2518.200 1558.890 2518.340 1559.250 ;
        RECT 2518.140 1558.570 2518.400 1558.890 ;
        RECT 2517.220 1545.650 2517.480 1545.970 ;
        RECT 2519.060 1545.650 2519.320 1545.970 ;
        RECT 2519.120 1462.410 2519.260 1545.650 ;
        RECT 2518.660 1462.270 2519.260 1462.410 ;
        RECT 2518.660 1415.410 2518.800 1462.270 ;
        RECT 2518.600 1415.090 2518.860 1415.410 ;
        RECT 2519.060 1414.750 2519.320 1415.070 ;
        RECT 2518.140 1366.470 2518.400 1366.790 ;
        RECT 2518.200 1366.110 2518.340 1366.470 ;
        RECT 2518.140 1365.790 2518.400 1366.110 ;
        RECT 2518.600 1318.190 2518.860 1318.510 ;
        RECT 2518.660 1317.830 2518.800 1318.190 ;
        RECT 2518.600 1317.510 2518.860 1317.830 ;
        RECT 2518.140 1269.910 2518.400 1270.230 ;
        RECT 2518.200 1269.550 2518.340 1269.910 ;
        RECT 2518.140 1269.230 2518.400 1269.550 ;
        RECT 2519.120 1269.290 2519.260 1414.750 ;
        RECT 2518.660 1269.150 2519.260 1269.290 ;
        RECT 2518.660 1222.290 2518.800 1269.150 ;
        RECT 2518.600 1221.970 2518.860 1222.290 ;
        RECT 2519.060 1221.630 2519.320 1221.950 ;
        RECT 2518.140 1173.350 2518.400 1173.670 ;
        RECT 2518.200 1172.990 2518.340 1173.350 ;
        RECT 2518.140 1172.670 2518.400 1172.990 ;
        RECT 2519.120 1172.730 2519.260 1221.630 ;
        RECT 2518.660 1172.590 2519.260 1172.730 ;
        RECT 2518.660 1125.730 2518.800 1172.590 ;
        RECT 2518.600 1125.410 2518.860 1125.730 ;
        RECT 2519.060 1125.070 2519.320 1125.390 ;
        RECT 2518.140 1076.790 2518.400 1077.110 ;
        RECT 2518.200 1076.430 2518.340 1076.790 ;
        RECT 2518.140 1076.110 2518.400 1076.430 ;
        RECT 2519.120 1076.170 2519.260 1125.070 ;
        RECT 2518.660 1076.030 2519.260 1076.170 ;
        RECT 2518.660 1029.170 2518.800 1076.030 ;
        RECT 2518.600 1028.850 2518.860 1029.170 ;
        RECT 2519.060 1028.510 2519.320 1028.830 ;
        RECT 2518.600 1028.170 2518.860 1028.490 ;
        RECT 2287.220 1012.190 2287.480 1012.510 ;
        RECT 2518.660 1011.150 2518.800 1028.170 ;
        RECT 2519.120 1011.490 2519.260 1028.510 ;
        RECT 2519.580 1011.830 2519.720 1606.995 ;
        RECT 2520.960 1594.250 2521.100 1617.730 ;
        RECT 2519.980 1593.930 2520.240 1594.250 ;
        RECT 2520.900 1593.930 2521.160 1594.250 ;
        RECT 2520.040 1559.570 2520.180 1593.930 ;
        RECT 2519.980 1559.250 2520.240 1559.570 ;
        RECT 2519.980 1558.570 2520.240 1558.890 ;
        RECT 2520.040 1366.790 2520.180 1558.570 ;
        RECT 2519.980 1366.470 2520.240 1366.790 ;
        RECT 2519.980 1365.790 2520.240 1366.110 ;
        RECT 2520.040 1318.510 2520.180 1365.790 ;
        RECT 2519.980 1318.190 2520.240 1318.510 ;
        RECT 2519.980 1317.510 2520.240 1317.830 ;
        RECT 2520.040 1270.230 2520.180 1317.510 ;
        RECT 2519.980 1269.910 2520.240 1270.230 ;
        RECT 2519.980 1269.230 2520.240 1269.550 ;
        RECT 2520.040 1173.670 2520.180 1269.230 ;
        RECT 2519.980 1173.350 2520.240 1173.670 ;
        RECT 2519.980 1172.670 2520.240 1172.990 ;
        RECT 2520.040 1077.110 2520.180 1172.670 ;
        RECT 2519.980 1076.790 2520.240 1077.110 ;
        RECT 2519.980 1076.110 2520.240 1076.430 ;
        RECT 2520.040 1028.490 2520.180 1076.110 ;
        RECT 2519.980 1028.170 2520.240 1028.490 ;
        RECT 2519.520 1011.510 2519.780 1011.830 ;
        RECT 2519.060 1011.170 2519.320 1011.490 ;
        RECT 2518.600 1010.830 2518.860 1011.150 ;
        RECT 2532.460 1010.810 2532.600 2600.590 ;
        RECT 2534.340 2600.000 2534.620 2600.590 ;
        RECT 2532.400 1010.490 2532.660 1010.810 ;
        RECT 2100.920 1008.790 2101.180 1009.110 ;
        RECT 2055.440 1000.000 2055.740 1000.010 ;
        RECT 2059.880 1000.000 2061.560 1000.010 ;
        RECT 2064.480 1000.000 2066.160 1000.010 ;
        RECT 2068.620 1000.000 2069.840 1000.010 ;
        RECT 2073.220 1000.000 2074.900 1000.010 ;
        RECT 2077.360 1000.000 2079.040 1000.010 ;
        RECT 2081.960 1000.000 2082.260 1000.010 ;
        RECT 2086.100 1000.000 2087.780 1000.010 ;
        RECT 1603.260 999.870 1603.710 1000.000 ;
      LAYER met2 ;
        RECT 1599.850 995.720 1600.850 998.810 ;
      LAYER met2 ;
        RECT 1601.130 996.000 1601.410 999.870 ;
      LAYER met2 ;
        RECT 1601.690 995.720 1603.150 998.810 ;
      LAYER met2 ;
        RECT 1603.430 996.000 1603.710 999.870 ;
      LAYER met2 ;
        RECT 1603.990 995.720 1605.450 998.810 ;
      LAYER met2 ;
        RECT 1605.730 996.000 1606.010 1000.000 ;
      LAYER met2 ;
        RECT 1606.290 995.720 1607.290 998.810 ;
      LAYER met2 ;
        RECT 1607.570 996.000 1607.850 1000.000 ;
        RECT 1608.780 999.870 1610.150 1000.000 ;
      LAYER met2 ;
        RECT 1608.130 995.720 1609.590 998.810 ;
      LAYER met2 ;
        RECT 1609.870 996.000 1610.150 999.870 ;
        RECT 1612.170 999.870 1613.980 1000.000 ;
      LAYER met2 ;
        RECT 1610.430 995.720 1611.890 998.810 ;
      LAYER met2 ;
        RECT 1612.170 996.000 1612.450 999.870 ;
      LAYER met2 ;
        RECT 1612.730 995.720 1614.190 998.810 ;
      LAYER met2 ;
        RECT 1614.470 996.000 1614.750 1000.000 ;
      LAYER met2 ;
        RECT 1615.030 995.720 1616.030 998.810 ;
      LAYER met2 ;
        RECT 1616.310 996.000 1616.590 1000.000 ;
        RECT 1618.610 999.870 1620.420 1000.000 ;
        RECT 1620.910 999.870 1621.340 1000.000 ;
      LAYER met2 ;
        RECT 1616.870 995.720 1618.330 998.810 ;
      LAYER met2 ;
        RECT 1618.610 996.000 1618.890 999.870 ;
      LAYER met2 ;
        RECT 1619.170 995.720 1620.630 998.810 ;
      LAYER met2 ;
        RECT 1620.910 996.000 1621.190 999.870 ;
      LAYER met2 ;
        RECT 1621.470 995.720 1622.930 998.810 ;
      LAYER met2 ;
        RECT 1623.210 996.000 1623.490 1000.000 ;
      LAYER met2 ;
        RECT 1623.770 995.720 1624.770 998.810 ;
      LAYER met2 ;
        RECT 1625.050 996.000 1625.330 1000.000 ;
        RECT 1625.800 999.870 1627.630 1000.000 ;
        RECT 1628.560 999.870 1629.930 1000.000 ;
      LAYER met2 ;
        RECT 1625.610 995.720 1627.070 998.810 ;
      LAYER met2 ;
        RECT 1627.350 996.000 1627.630 999.870 ;
      LAYER met2 ;
        RECT 1627.910 995.720 1629.370 998.810 ;
      LAYER met2 ;
        RECT 1629.650 996.000 1629.930 999.870 ;
      LAYER met2 ;
        RECT 1630.210 995.720 1631.210 998.810 ;
      LAYER met2 ;
        RECT 1631.490 996.000 1631.770 1000.000 ;
      LAYER met2 ;
        RECT 1632.050 995.720 1633.510 998.810 ;
      LAYER met2 ;
        RECT 1633.790 996.000 1634.070 1000.000 ;
      LAYER met2 ;
        RECT 1634.350 995.720 1635.810 998.810 ;
      LAYER met2 ;
        RECT 1636.090 996.000 1636.370 1000.000 ;
      LAYER met2 ;
        RECT 1636.650 995.720 1638.110 998.810 ;
      LAYER met2 ;
        RECT 1638.390 996.000 1638.670 1000.000 ;
      LAYER met2 ;
        RECT 1638.950 995.720 1639.950 998.810 ;
      LAYER met2 ;
        RECT 1640.230 996.000 1640.510 1000.000 ;
      LAYER met2 ;
        RECT 1640.790 995.720 1642.250 998.810 ;
      LAYER met2 ;
        RECT 1642.530 996.000 1642.810 1000.000 ;
      LAYER met2 ;
        RECT 1643.090 995.720 1644.550 998.810 ;
      LAYER met2 ;
        RECT 1644.830 996.000 1645.110 1000.000 ;
      LAYER met2 ;
        RECT 1645.390 995.720 1646.850 998.810 ;
      LAYER met2 ;
        RECT 1647.130 996.000 1647.410 1000.000 ;
      LAYER met2 ;
        RECT 1647.690 995.720 1648.690 998.810 ;
      LAYER met2 ;
        RECT 1648.970 996.000 1649.250 1000.000 ;
      LAYER met2 ;
        RECT 1649.530 995.720 1650.990 998.810 ;
      LAYER met2 ;
        RECT 1651.270 996.000 1651.550 1000.000 ;
      LAYER met2 ;
        RECT 1651.830 995.720 1653.290 998.810 ;
      LAYER met2 ;
        RECT 1653.570 996.000 1653.850 1000.000 ;
      LAYER met2 ;
        RECT 1654.130 995.720 1655.130 998.810 ;
      LAYER met2 ;
        RECT 1655.410 996.000 1655.690 1000.000 ;
      LAYER met2 ;
        RECT 1655.970 995.720 1657.430 998.810 ;
      LAYER met2 ;
        RECT 1657.710 996.000 1657.990 1000.000 ;
      LAYER met2 ;
        RECT 1658.270 995.720 1659.730 998.810 ;
      LAYER met2 ;
        RECT 1660.010 996.000 1660.290 1000.000 ;
        RECT 1662.310 999.870 1662.740 1000.000 ;
        RECT 1664.150 999.870 1665.960 1000.000 ;
        RECT 1666.450 999.870 1668.260 1000.000 ;
      LAYER met2 ;
        RECT 1660.570 995.720 1662.030 998.810 ;
      LAYER met2 ;
        RECT 1662.310 996.000 1662.590 999.870 ;
      LAYER met2 ;
        RECT 1662.870 995.720 1663.870 998.810 ;
      LAYER met2 ;
        RECT 1664.150 996.000 1664.430 999.870 ;
      LAYER met2 ;
        RECT 1664.710 995.720 1666.170 998.810 ;
      LAYER met2 ;
        RECT 1666.450 996.000 1666.730 999.870 ;
      LAYER met2 ;
        RECT 1667.010 995.720 1668.470 998.810 ;
      LAYER met2 ;
        RECT 1668.750 996.000 1669.030 1000.000 ;
      LAYER met2 ;
        RECT 1669.310 995.720 1670.770 998.810 ;
      LAYER met2 ;
        RECT 1671.050 996.000 1671.330 1000.000 ;
      LAYER met2 ;
        RECT 1671.610 995.720 1672.610 998.810 ;
      LAYER met2 ;
        RECT 1672.890 996.000 1673.170 1000.000 ;
      LAYER met2 ;
        RECT 1673.450 995.720 1674.910 998.810 ;
      LAYER met2 ;
        RECT 1675.190 996.000 1675.470 1000.000 ;
      LAYER met2 ;
        RECT 1675.750 995.720 1677.210 998.810 ;
      LAYER met2 ;
        RECT 1677.490 996.000 1677.770 1000.000 ;
      LAYER met2 ;
        RECT 1678.050 995.720 1679.050 998.810 ;
      LAYER met2 ;
        RECT 1679.330 996.000 1679.610 1000.000 ;
      LAYER met2 ;
        RECT 1679.890 995.720 1681.350 998.810 ;
      LAYER met2 ;
        RECT 1681.630 996.000 1681.910 1000.000 ;
      LAYER met2 ;
        RECT 1682.190 995.720 1683.650 998.810 ;
      LAYER met2 ;
        RECT 1683.930 996.000 1684.210 1000.000 ;
      LAYER met2 ;
        RECT 1684.490 995.720 1685.950 998.810 ;
      LAYER met2 ;
        RECT 1686.230 996.000 1686.510 1000.000 ;
      LAYER met2 ;
        RECT 1686.790 995.720 1687.790 998.810 ;
      LAYER met2 ;
        RECT 1688.070 996.000 1688.350 1000.000 ;
      LAYER met2 ;
        RECT 1688.630 995.720 1690.090 998.810 ;
      LAYER met2 ;
        RECT 1690.370 996.000 1690.650 1000.000 ;
      LAYER met2 ;
        RECT 1690.930 995.720 1692.390 998.810 ;
      LAYER met2 ;
        RECT 1692.670 996.000 1692.950 1000.000 ;
      LAYER met2 ;
        RECT 1693.230 995.720 1694.230 998.810 ;
      LAYER met2 ;
        RECT 1694.510 996.000 1694.790 1000.000 ;
      LAYER met2 ;
        RECT 1695.070 995.720 1696.530 998.810 ;
      LAYER met2 ;
        RECT 1696.810 996.000 1697.090 1000.000 ;
      LAYER met2 ;
        RECT 1697.370 995.720 1698.830 998.810 ;
      LAYER met2 ;
        RECT 1699.110 996.000 1699.390 1000.000 ;
      LAYER met2 ;
        RECT 1699.670 995.720 1701.130 998.810 ;
      LAYER met2 ;
        RECT 1701.410 996.000 1701.690 1000.000 ;
      LAYER met2 ;
        RECT 1701.970 995.720 1702.970 998.810 ;
      LAYER met2 ;
        RECT 1703.250 996.000 1703.530 1000.000 ;
        RECT 1705.550 999.870 1707.360 1000.000 ;
      LAYER met2 ;
        RECT 1703.810 995.720 1705.270 998.810 ;
      LAYER met2 ;
        RECT 1705.550 996.000 1705.830 999.870 ;
      LAYER met2 ;
        RECT 1706.110 995.720 1707.570 998.810 ;
      LAYER met2 ;
        RECT 1707.850 996.000 1708.130 1000.000 ;
        RECT 1710.150 999.870 1711.040 1000.000 ;
      LAYER met2 ;
        RECT 1708.410 995.720 1709.870 998.810 ;
      LAYER met2 ;
        RECT 1710.150 996.000 1710.430 999.870 ;
      LAYER met2 ;
        RECT 1710.710 995.720 1711.710 998.810 ;
      LAYER met2 ;
        RECT 1711.990 996.000 1712.270 1000.000 ;
        RECT 1714.290 999.870 1715.640 1000.000 ;
      LAYER met2 ;
        RECT 1712.550 995.720 1714.010 998.810 ;
      LAYER met2 ;
        RECT 1714.290 996.000 1714.570 999.870 ;
      LAYER met2 ;
        RECT 1714.850 995.720 1716.310 998.810 ;
      LAYER met2 ;
        RECT 1716.590 996.000 1716.870 1000.000 ;
        RECT 1718.430 999.870 1720.240 1000.000 ;
      LAYER met2 ;
        RECT 1717.150 995.720 1718.150 998.810 ;
      LAYER met2 ;
        RECT 1718.430 996.000 1718.710 999.870 ;
      LAYER met2 ;
        RECT 1718.990 995.720 1720.450 998.810 ;
      LAYER met2 ;
        RECT 1720.730 996.000 1721.010 1000.000 ;
        RECT 1723.030 999.870 1724.840 1000.000 ;
      LAYER met2 ;
        RECT 1721.290 995.720 1722.750 998.810 ;
      LAYER met2 ;
        RECT 1723.030 996.000 1723.310 999.870 ;
      LAYER met2 ;
        RECT 1723.590 995.720 1725.050 998.810 ;
      LAYER met2 ;
        RECT 1725.330 996.000 1725.610 1000.000 ;
        RECT 1727.170 999.870 1728.980 1000.000 ;
      LAYER met2 ;
        RECT 1725.890 995.720 1726.890 998.810 ;
      LAYER met2 ;
        RECT 1727.170 996.000 1727.450 999.870 ;
      LAYER met2 ;
        RECT 1727.730 995.720 1729.190 998.810 ;
      LAYER met2 ;
        RECT 1729.470 996.000 1729.750 1000.000 ;
        RECT 1731.770 999.870 1733.580 1000.000 ;
      LAYER met2 ;
        RECT 1730.030 995.720 1731.490 998.810 ;
      LAYER met2 ;
        RECT 1731.770 996.000 1732.050 999.870 ;
      LAYER met2 ;
        RECT 1732.330 995.720 1733.790 998.810 ;
      LAYER met2 ;
        RECT 1734.070 996.000 1734.350 1000.000 ;
        RECT 1735.910 999.870 1737.720 1000.000 ;
      LAYER met2 ;
        RECT 1734.630 995.720 1735.630 998.810 ;
      LAYER met2 ;
        RECT 1735.910 996.000 1736.190 999.870 ;
      LAYER met2 ;
        RECT 1736.470 995.720 1737.930 998.810 ;
      LAYER met2 ;
        RECT 1738.210 996.000 1738.490 1000.000 ;
        RECT 1740.510 999.870 1741.860 1000.000 ;
      LAYER met2 ;
        RECT 1738.770 995.720 1740.230 998.810 ;
      LAYER met2 ;
        RECT 1740.510 996.000 1740.790 999.870 ;
      LAYER met2 ;
        RECT 1741.070 995.720 1742.070 998.810 ;
      LAYER met2 ;
        RECT 1742.350 996.000 1742.630 1000.000 ;
        RECT 1744.650 999.870 1745.540 1000.000 ;
      LAYER met2 ;
        RECT 1742.910 995.720 1744.370 998.810 ;
      LAYER met2 ;
        RECT 1744.650 996.000 1744.930 999.870 ;
      LAYER met2 ;
        RECT 1745.210 995.720 1746.670 998.810 ;
      LAYER met2 ;
        RECT 1746.950 996.000 1747.230 1000.000 ;
        RECT 1749.250 999.870 1750.140 1000.000 ;
      LAYER met2 ;
        RECT 1747.510 995.720 1748.970 998.810 ;
      LAYER met2 ;
        RECT 1749.250 996.000 1749.530 999.870 ;
      LAYER met2 ;
        RECT 1749.810 995.720 1750.810 998.810 ;
      LAYER met2 ;
        RECT 1751.090 996.000 1751.370 1000.000 ;
        RECT 1753.390 999.870 1755.200 1000.000 ;
      LAYER met2 ;
        RECT 1751.650 995.720 1753.110 998.810 ;
      LAYER met2 ;
        RECT 1753.390 996.000 1753.670 999.870 ;
      LAYER met2 ;
        RECT 1753.950 995.720 1755.410 998.810 ;
      LAYER met2 ;
        RECT 1755.690 996.000 1755.970 1000.000 ;
        RECT 1757.990 999.870 1758.880 1000.000 ;
      LAYER met2 ;
        RECT 1756.250 995.720 1757.710 998.810 ;
      LAYER met2 ;
        RECT 1757.990 996.000 1758.270 999.870 ;
      LAYER met2 ;
        RECT 1758.550 995.720 1759.550 998.810 ;
      LAYER met2 ;
        RECT 1759.830 996.000 1760.110 1000.000 ;
        RECT 1762.130 999.870 1763.940 1000.000 ;
      LAYER met2 ;
        RECT 1760.390 995.720 1761.850 998.810 ;
      LAYER met2 ;
        RECT 1762.130 996.000 1762.410 999.870 ;
      LAYER met2 ;
        RECT 1762.690 995.720 1764.150 998.810 ;
      LAYER met2 ;
        RECT 1764.430 996.000 1764.710 1000.000 ;
        RECT 1766.270 999.870 1768.080 1000.000 ;
      LAYER met2 ;
        RECT 1764.990 995.720 1765.990 998.810 ;
      LAYER met2 ;
        RECT 1766.270 996.000 1766.550 999.870 ;
      LAYER met2 ;
        RECT 1766.830 995.720 1768.290 998.810 ;
      LAYER met2 ;
        RECT 1768.570 996.000 1768.850 1000.000 ;
        RECT 1770.870 999.870 1772.680 1000.000 ;
      LAYER met2 ;
        RECT 1769.130 995.720 1770.590 998.810 ;
      LAYER met2 ;
        RECT 1770.870 996.000 1771.150 999.870 ;
      LAYER met2 ;
        RECT 1771.430 995.720 1772.890 998.810 ;
      LAYER met2 ;
        RECT 1773.170 996.000 1773.450 1000.000 ;
        RECT 1775.010 999.870 1776.820 1000.000 ;
      LAYER met2 ;
        RECT 1773.730 995.720 1774.730 998.810 ;
      LAYER met2 ;
        RECT 1775.010 996.000 1775.290 999.870 ;
      LAYER met2 ;
        RECT 1775.570 995.720 1777.030 998.810 ;
      LAYER met2 ;
        RECT 1777.310 996.000 1777.590 1000.000 ;
        RECT 1779.440 999.870 1779.890 1000.000 ;
      LAYER met2 ;
        RECT 1777.870 995.720 1779.330 998.810 ;
      LAYER met2 ;
        RECT 1779.610 996.000 1779.890 999.870 ;
      LAYER met2 ;
        RECT 1780.170 995.720 1781.630 998.810 ;
      LAYER met2 ;
        RECT 1781.910 996.000 1782.190 1000.000 ;
        RECT 1783.750 999.870 1785.560 1000.000 ;
      LAYER met2 ;
        RECT 1782.470 995.720 1783.470 998.810 ;
      LAYER met2 ;
        RECT 1783.750 996.000 1784.030 999.870 ;
      LAYER met2 ;
        RECT 1784.310 995.720 1785.770 998.810 ;
      LAYER met2 ;
        RECT 1786.050 996.000 1786.330 1000.000 ;
        RECT 1788.350 999.870 1789.700 1000.000 ;
      LAYER met2 ;
        RECT 1786.610 995.720 1788.070 998.810 ;
      LAYER met2 ;
        RECT 1788.350 996.000 1788.630 999.870 ;
      LAYER met2 ;
        RECT 1788.910 995.720 1789.910 998.810 ;
      LAYER met2 ;
        RECT 1790.190 996.000 1790.470 1000.000 ;
        RECT 1792.490 999.870 1793.840 1000.000 ;
      LAYER met2 ;
        RECT 1790.750 995.720 1792.210 998.810 ;
      LAYER met2 ;
        RECT 1792.490 996.000 1792.770 999.870 ;
      LAYER met2 ;
        RECT 1793.050 995.720 1794.510 998.810 ;
      LAYER met2 ;
        RECT 1794.790 996.000 1795.070 1000.000 ;
        RECT 1797.090 999.870 1798.440 1000.000 ;
      LAYER met2 ;
        RECT 1795.350 995.720 1796.810 998.810 ;
      LAYER met2 ;
        RECT 1797.090 996.000 1797.370 999.870 ;
      LAYER met2 ;
        RECT 1797.650 995.720 1798.650 998.810 ;
      LAYER met2 ;
        RECT 1798.930 996.000 1799.210 1000.000 ;
        RECT 1801.230 999.870 1803.040 1000.000 ;
      LAYER met2 ;
        RECT 1799.490 995.720 1800.950 998.810 ;
      LAYER met2 ;
        RECT 1801.230 996.000 1801.510 999.870 ;
      LAYER met2 ;
        RECT 1801.790 995.720 1803.250 998.810 ;
      LAYER met2 ;
        RECT 1803.530 996.000 1803.810 1000.000 ;
        RECT 1805.830 999.870 1807.180 1000.000 ;
      LAYER met2 ;
        RECT 1804.090 995.720 1805.550 998.810 ;
      LAYER met2 ;
        RECT 1805.830 996.000 1806.110 999.870 ;
      LAYER met2 ;
        RECT 1806.390 995.720 1807.390 998.810 ;
      LAYER met2 ;
        RECT 1807.670 996.000 1807.950 1000.000 ;
        RECT 1809.970 999.870 1811.780 1000.000 ;
      LAYER met2 ;
        RECT 1808.230 995.720 1809.690 998.810 ;
      LAYER met2 ;
        RECT 1809.970 996.000 1810.250 999.870 ;
      LAYER met2 ;
        RECT 1810.530 995.720 1811.990 998.810 ;
      LAYER met2 ;
        RECT 1812.270 996.000 1812.550 1000.000 ;
        RECT 1814.110 999.870 1814.540 1000.000 ;
      LAYER met2 ;
        RECT 1812.830 995.720 1813.830 998.810 ;
      LAYER met2 ;
        RECT 1814.110 996.000 1814.390 999.870 ;
      LAYER met2 ;
        RECT 1814.670 995.720 1816.130 998.810 ;
      LAYER met2 ;
        RECT 1816.410 996.000 1816.690 1000.000 ;
        RECT 1818.710 999.870 1820.520 1000.000 ;
      LAYER met2 ;
        RECT 1816.970 995.720 1818.430 998.810 ;
      LAYER met2 ;
        RECT 1818.710 996.000 1818.990 999.870 ;
      LAYER met2 ;
        RECT 1819.270 995.720 1820.730 998.810 ;
      LAYER met2 ;
        RECT 1821.010 996.000 1821.290 1000.000 ;
        RECT 1822.850 999.870 1824.660 1000.000 ;
        RECT 1825.150 999.870 1826.960 1000.000 ;
      LAYER met2 ;
        RECT 1821.570 995.720 1822.570 998.810 ;
      LAYER met2 ;
        RECT 1822.850 996.000 1823.130 999.870 ;
      LAYER met2 ;
        RECT 1823.410 995.720 1824.870 998.810 ;
      LAYER met2 ;
        RECT 1825.150 996.000 1825.430 999.870 ;
      LAYER met2 ;
        RECT 1825.710 995.720 1827.170 998.810 ;
      LAYER met2 ;
        RECT 1827.450 996.000 1827.730 1000.000 ;
        RECT 1829.750 999.870 1831.100 1000.000 ;
      LAYER met2 ;
        RECT 1828.010 995.720 1829.470 998.810 ;
      LAYER met2 ;
        RECT 1829.750 996.000 1830.030 999.870 ;
      LAYER met2 ;
        RECT 1830.310 995.720 1831.310 998.810 ;
      LAYER met2 ;
        RECT 1831.590 996.000 1831.870 1000.000 ;
        RECT 1833.890 999.870 1834.780 1000.000 ;
      LAYER met2 ;
        RECT 1832.150 995.720 1833.610 998.810 ;
      LAYER met2 ;
        RECT 1833.890 996.000 1834.170 999.870 ;
      LAYER met2 ;
        RECT 1834.450 995.720 1835.910 998.810 ;
      LAYER met2 ;
        RECT 1836.190 996.000 1836.470 1000.000 ;
      LAYER met2 ;
        RECT 1836.750 995.720 1837.750 998.810 ;
      LAYER met2 ;
        RECT 1838.030 996.000 1838.310 1000.000 ;
      LAYER met2 ;
        RECT 1838.590 995.720 1840.050 998.810 ;
      LAYER met2 ;
        RECT 1840.330 996.000 1840.610 1000.000 ;
      LAYER met2 ;
        RECT 1840.890 995.720 1842.350 998.810 ;
      LAYER met2 ;
        RECT 1842.630 996.000 1842.910 1000.000 ;
      LAYER met2 ;
        RECT 1843.190 995.720 1844.650 998.810 ;
      LAYER met2 ;
        RECT 1844.930 996.000 1845.210 1000.000 ;
      LAYER met2 ;
        RECT 1845.490 995.720 1846.490 998.810 ;
      LAYER met2 ;
        RECT 1846.770 996.000 1847.050 1000.000 ;
      LAYER met2 ;
        RECT 1847.330 995.720 1848.790 998.810 ;
      LAYER met2 ;
        RECT 1849.070 996.000 1849.350 1000.000 ;
      LAYER met2 ;
        RECT 1849.630 995.720 1851.090 998.810 ;
      LAYER met2 ;
        RECT 1851.370 996.000 1851.650 1000.000 ;
      LAYER met2 ;
        RECT 1851.930 995.720 1852.930 998.810 ;
      LAYER met2 ;
        RECT 1853.210 996.000 1853.490 1000.000 ;
      LAYER met2 ;
        RECT 1853.770 995.720 1855.230 998.810 ;
      LAYER met2 ;
        RECT 1855.510 996.000 1855.790 1000.000 ;
      LAYER met2 ;
        RECT 1856.070 995.720 1857.530 998.810 ;
      LAYER met2 ;
        RECT 1857.810 996.000 1858.090 1000.000 ;
      LAYER met2 ;
        RECT 1858.370 995.720 1859.830 998.810 ;
      LAYER met2 ;
        RECT 1860.110 996.000 1860.390 1000.000 ;
      LAYER met2 ;
        RECT 1860.670 995.720 1861.670 998.810 ;
      LAYER met2 ;
        RECT 1861.950 996.000 1862.230 1000.000 ;
      LAYER met2 ;
        RECT 1862.510 995.720 1863.970 998.810 ;
      LAYER met2 ;
        RECT 1864.250 996.000 1864.530 1000.000 ;
      LAYER met2 ;
        RECT 1864.810 995.720 1866.270 998.810 ;
      LAYER met2 ;
        RECT 1866.550 996.000 1866.830 1000.000 ;
      LAYER met2 ;
        RECT 1867.110 995.720 1868.570 998.810 ;
      LAYER met2 ;
        RECT 1868.850 996.000 1869.130 1000.000 ;
        RECT 1870.690 999.870 1872.500 1000.000 ;
      LAYER met2 ;
        RECT 1869.410 995.720 1870.410 998.810 ;
      LAYER met2 ;
        RECT 1870.690 996.000 1870.970 999.870 ;
      LAYER met2 ;
        RECT 1871.250 995.720 1872.710 998.810 ;
      LAYER met2 ;
        RECT 1872.990 996.000 1873.270 1000.000 ;
      LAYER met2 ;
        RECT 1873.550 995.720 1875.010 998.810 ;
      LAYER met2 ;
        RECT 1875.290 996.000 1875.570 1000.000 ;
        RECT 1877.130 999.870 1878.940 1000.000 ;
      LAYER met2 ;
        RECT 1875.850 995.720 1876.850 998.810 ;
      LAYER met2 ;
        RECT 1877.130 996.000 1877.410 999.870 ;
      LAYER met2 ;
        RECT 1877.690 995.720 1879.150 998.810 ;
      LAYER met2 ;
        RECT 1879.430 996.000 1879.710 1000.000 ;
        RECT 1881.730 999.870 1883.540 1000.000 ;
      LAYER met2 ;
        RECT 1879.990 995.720 1881.450 998.810 ;
      LAYER met2 ;
        RECT 1881.730 996.000 1882.010 999.870 ;
      LAYER met2 ;
        RECT 1882.290 995.720 1883.750 998.810 ;
      LAYER met2 ;
        RECT 1884.030 996.000 1884.310 1000.000 ;
      LAYER met2 ;
        RECT 1884.590 995.720 1885.590 998.810 ;
      LAYER met2 ;
        RECT 1885.870 996.000 1886.150 1000.000 ;
      LAYER met2 ;
        RECT 1886.430 995.720 1887.890 998.810 ;
      LAYER met2 ;
        RECT 1888.170 996.000 1888.450 1000.000 ;
      LAYER met2 ;
        RECT 1888.730 995.720 1890.190 998.810 ;
      LAYER met2 ;
        RECT 1890.470 996.000 1890.750 1000.000 ;
      LAYER met2 ;
        RECT 1891.030 995.720 1892.490 998.810 ;
      LAYER met2 ;
        RECT 1892.770 996.000 1893.050 1000.000 ;
      LAYER met2 ;
        RECT 1893.330 995.720 1894.330 998.810 ;
      LAYER met2 ;
        RECT 1894.610 996.000 1894.890 1000.000 ;
      LAYER met2 ;
        RECT 1895.170 995.720 1896.630 998.810 ;
      LAYER met2 ;
        RECT 1896.910 996.000 1897.190 1000.000 ;
      LAYER met2 ;
        RECT 1897.470 995.720 1898.930 998.810 ;
      LAYER met2 ;
        RECT 1899.210 996.000 1899.490 1000.000 ;
      LAYER met2 ;
        RECT 1899.770 995.720 1900.770 998.810 ;
      LAYER met2 ;
        RECT 1901.050 996.000 1901.330 1000.000 ;
      LAYER met2 ;
        RECT 1901.610 995.720 1903.070 998.810 ;
      LAYER met2 ;
        RECT 1903.350 996.000 1903.630 1000.000 ;
      LAYER met2 ;
        RECT 1903.910 995.720 1905.370 998.810 ;
      LAYER met2 ;
        RECT 1905.650 996.000 1905.930 1000.000 ;
      LAYER met2 ;
        RECT 1906.210 995.720 1907.670 998.810 ;
      LAYER met2 ;
        RECT 1907.950 996.000 1908.230 1000.000 ;
      LAYER met2 ;
        RECT 1908.510 995.720 1909.510 998.810 ;
      LAYER met2 ;
        RECT 1909.790 996.000 1910.070 1000.000 ;
      LAYER met2 ;
        RECT 1910.350 995.720 1911.810 998.810 ;
      LAYER met2 ;
        RECT 1912.090 996.000 1912.370 1000.000 ;
      LAYER met2 ;
        RECT 1912.650 995.720 1914.110 998.810 ;
      LAYER met2 ;
        RECT 1914.390 996.000 1914.670 1000.000 ;
      LAYER met2 ;
        RECT 1914.950 995.720 1916.410 998.810 ;
      LAYER met2 ;
        RECT 1916.690 996.000 1916.970 1000.000 ;
      LAYER met2 ;
        RECT 1917.250 995.720 1918.250 998.810 ;
      LAYER met2 ;
        RECT 1918.530 996.000 1918.810 1000.000 ;
      LAYER met2 ;
        RECT 1919.090 995.720 1920.550 998.810 ;
      LAYER met2 ;
        RECT 1920.830 996.000 1921.110 1000.000 ;
      LAYER met2 ;
        RECT 1921.390 995.720 1922.850 998.810 ;
      LAYER met2 ;
        RECT 1923.130 996.000 1923.410 1000.000 ;
      LAYER met2 ;
        RECT 1923.690 995.720 1924.690 998.810 ;
      LAYER met2 ;
        RECT 1924.970 996.000 1925.250 1000.000 ;
      LAYER met2 ;
        RECT 1925.530 995.720 1926.990 998.810 ;
      LAYER met2 ;
        RECT 1927.270 996.000 1927.550 1000.000 ;
      LAYER met2 ;
        RECT 1927.830 995.720 1929.290 998.810 ;
      LAYER met2 ;
        RECT 1929.570 996.000 1929.850 1000.000 ;
      LAYER met2 ;
        RECT 1930.130 995.720 1931.590 998.810 ;
      LAYER met2 ;
        RECT 1931.870 996.000 1932.150 1000.000 ;
      LAYER met2 ;
        RECT 1932.430 995.720 1933.430 998.810 ;
      LAYER met2 ;
        RECT 1933.710 996.000 1933.990 1000.000 ;
      LAYER met2 ;
        RECT 1934.270 995.720 1935.730 998.810 ;
      LAYER met2 ;
        RECT 1936.010 996.000 1936.290 1000.000 ;
      LAYER met2 ;
        RECT 1936.570 995.720 1938.030 998.810 ;
      LAYER met2 ;
        RECT 1938.310 996.000 1938.590 1000.000 ;
      LAYER met2 ;
        RECT 1938.870 995.720 1940.330 998.810 ;
      LAYER met2 ;
        RECT 1940.610 996.000 1940.890 1000.000 ;
      LAYER met2 ;
        RECT 1941.170 995.720 1942.170 998.810 ;
      LAYER met2 ;
        RECT 1942.450 996.000 1942.730 1000.000 ;
      LAYER met2 ;
        RECT 1943.010 995.720 1944.470 998.810 ;
      LAYER met2 ;
        RECT 1944.750 996.000 1945.030 1000.000 ;
      LAYER met2 ;
        RECT 1945.310 995.720 1946.770 998.810 ;
      LAYER met2 ;
        RECT 1947.050 996.000 1947.330 1000.000 ;
      LAYER met2 ;
        RECT 1947.610 995.720 1948.610 998.810 ;
      LAYER met2 ;
        RECT 1948.890 996.000 1949.170 1000.000 ;
      LAYER met2 ;
        RECT 1949.450 995.720 1950.910 998.810 ;
      LAYER met2 ;
        RECT 1951.190 996.000 1951.470 1000.000 ;
      LAYER met2 ;
        RECT 1951.750 995.720 1953.210 998.810 ;
      LAYER met2 ;
        RECT 1953.490 996.000 1953.770 1000.000 ;
      LAYER met2 ;
        RECT 1954.050 995.720 1955.510 998.810 ;
      LAYER met2 ;
        RECT 1955.790 996.000 1956.070 1000.000 ;
      LAYER met2 ;
        RECT 1956.350 995.720 1957.350 998.810 ;
      LAYER met2 ;
        RECT 1957.630 996.000 1957.910 1000.000 ;
      LAYER met2 ;
        RECT 1958.190 995.720 1959.650 998.810 ;
      LAYER met2 ;
        RECT 1959.930 996.000 1960.210 1000.000 ;
      LAYER met2 ;
        RECT 1960.490 995.720 1961.950 998.810 ;
      LAYER met2 ;
        RECT 1962.230 996.000 1962.510 1000.000 ;
      LAYER met2 ;
        RECT 1962.790 995.720 1964.250 998.810 ;
      LAYER met2 ;
        RECT 1964.530 996.000 1964.810 1000.000 ;
      LAYER met2 ;
        RECT 1965.090 995.720 1966.090 998.810 ;
      LAYER met2 ;
        RECT 1966.370 996.000 1966.650 1000.000 ;
      LAYER met2 ;
        RECT 1966.930 995.720 1968.390 998.810 ;
      LAYER met2 ;
        RECT 1968.670 996.000 1968.950 1000.000 ;
      LAYER met2 ;
        RECT 1969.230 995.720 1970.690 998.810 ;
      LAYER met2 ;
        RECT 1970.970 996.000 1971.250 1000.000 ;
      LAYER met2 ;
        RECT 1971.530 995.720 1972.530 998.810 ;
      LAYER met2 ;
        RECT 1972.810 996.000 1973.090 1000.000 ;
      LAYER met2 ;
        RECT 1973.370 995.720 1974.830 998.810 ;
      LAYER met2 ;
        RECT 1975.110 996.000 1975.390 1000.000 ;
      LAYER met2 ;
        RECT 1975.670 995.720 1977.130 998.810 ;
      LAYER met2 ;
        RECT 1977.410 996.000 1977.690 1000.000 ;
      LAYER met2 ;
        RECT 1977.970 995.720 1979.430 998.810 ;
      LAYER met2 ;
        RECT 1979.710 996.000 1979.990 1000.000 ;
      LAYER met2 ;
        RECT 1980.270 995.720 1981.270 998.810 ;
      LAYER met2 ;
        RECT 1981.550 996.000 1981.830 1000.000 ;
      LAYER met2 ;
        RECT 1982.110 995.720 1983.570 998.810 ;
      LAYER met2 ;
        RECT 1983.850 996.000 1984.130 1000.000 ;
      LAYER met2 ;
        RECT 1984.410 995.720 1985.870 998.810 ;
      LAYER met2 ;
        RECT 1986.150 996.000 1986.430 1000.000 ;
      LAYER met2 ;
        RECT 1986.710 995.720 1988.170 998.810 ;
      LAYER met2 ;
        RECT 1988.450 996.000 1988.730 1000.000 ;
      LAYER met2 ;
        RECT 1989.010 995.720 1990.010 998.810 ;
      LAYER met2 ;
        RECT 1990.290 996.000 1990.570 1000.000 ;
      LAYER met2 ;
        RECT 1990.850 995.720 1992.310 998.810 ;
      LAYER met2 ;
        RECT 1992.590 996.000 1992.870 1000.000 ;
      LAYER met2 ;
        RECT 1993.150 995.720 1994.610 998.810 ;
      LAYER met2 ;
        RECT 1994.890 996.000 1995.170 1000.000 ;
      LAYER met2 ;
        RECT 1995.450 995.720 1996.450 998.810 ;
      LAYER met2 ;
        RECT 1996.730 996.000 1997.010 1000.000 ;
      LAYER met2 ;
        RECT 1997.290 995.720 1998.750 998.810 ;
      LAYER met2 ;
        RECT 1999.030 996.000 1999.310 1000.000 ;
        RECT 2001.330 999.870 2003.140 1000.000 ;
        RECT 2003.630 999.870 2004.980 1000.000 ;
      LAYER met2 ;
        RECT 1999.590 995.720 2001.050 998.810 ;
      LAYER met2 ;
        RECT 2001.330 996.000 2001.610 999.870 ;
      LAYER met2 ;
        RECT 2001.890 995.720 2003.350 998.810 ;
      LAYER met2 ;
        RECT 2003.630 996.000 2003.910 999.870 ;
      LAYER met2 ;
        RECT 2004.190 995.720 2005.190 998.810 ;
      LAYER met2 ;
        RECT 2005.470 996.000 2005.750 1000.000 ;
      LAYER met2 ;
        RECT 2006.030 995.720 2007.490 998.810 ;
      LAYER met2 ;
        RECT 2007.770 996.000 2008.050 1000.000 ;
      LAYER met2 ;
        RECT 2008.330 995.720 2009.790 998.810 ;
      LAYER met2 ;
        RECT 2010.070 996.000 2010.350 1000.000 ;
      LAYER met2 ;
        RECT 2010.630 995.720 2011.630 998.810 ;
      LAYER met2 ;
        RECT 2011.910 996.000 2012.190 1000.000 ;
      LAYER met2 ;
        RECT 2012.470 995.720 2013.930 998.810 ;
      LAYER met2 ;
        RECT 2014.210 996.000 2014.490 1000.000 ;
      LAYER met2 ;
        RECT 2014.770 995.720 2016.230 998.810 ;
      LAYER met2 ;
        RECT 2016.510 996.000 2016.790 1000.000 ;
      LAYER met2 ;
        RECT 2017.070 995.720 2018.530 998.810 ;
      LAYER met2 ;
        RECT 2018.810 996.000 2019.090 1000.000 ;
      LAYER met2 ;
        RECT 2019.370 995.720 2020.370 998.810 ;
      LAYER met2 ;
        RECT 2020.650 996.000 2020.930 1000.000 ;
      LAYER met2 ;
        RECT 2021.210 995.720 2022.670 998.810 ;
      LAYER met2 ;
        RECT 2022.950 996.000 2023.230 1000.000 ;
      LAYER met2 ;
        RECT 2023.510 995.720 2024.970 998.810 ;
      LAYER met2 ;
        RECT 2025.250 996.000 2025.530 1000.000 ;
      LAYER met2 ;
        RECT 2025.810 995.720 2027.270 998.810 ;
      LAYER met2 ;
        RECT 2027.550 996.000 2027.830 1000.000 ;
      LAYER met2 ;
        RECT 2028.110 995.720 2029.110 998.810 ;
      LAYER met2 ;
        RECT 2029.390 996.000 2029.670 1000.000 ;
      LAYER met2 ;
        RECT 2029.950 995.720 2031.410 998.810 ;
      LAYER met2 ;
        RECT 2031.690 996.000 2031.970 1000.000 ;
      LAYER met2 ;
        RECT 2032.250 995.720 2033.710 998.810 ;
      LAYER met2 ;
        RECT 2033.990 996.000 2034.270 1000.000 ;
      LAYER met2 ;
        RECT 2034.550 995.720 2035.550 998.810 ;
      LAYER met2 ;
        RECT 2035.830 996.000 2036.110 1000.000 ;
      LAYER met2 ;
        RECT 2036.390 995.720 2037.850 998.810 ;
      LAYER met2 ;
        RECT 2038.130 996.000 2038.410 1000.000 ;
        RECT 2040.430 999.870 2042.240 1000.000 ;
      LAYER met2 ;
        RECT 2038.690 995.720 2040.150 998.810 ;
      LAYER met2 ;
        RECT 2040.430 996.000 2040.710 999.870 ;
      LAYER met2 ;
        RECT 2040.990 995.720 2042.450 998.810 ;
      LAYER met2 ;
        RECT 2042.730 996.000 2043.010 1000.000 ;
        RECT 2044.570 999.870 2046.380 1000.000 ;
      LAYER met2 ;
        RECT 2043.290 995.720 2044.290 998.810 ;
      LAYER met2 ;
        RECT 2044.570 996.000 2044.850 999.870 ;
      LAYER met2 ;
        RECT 2045.130 995.720 2046.590 998.810 ;
      LAYER met2 ;
        RECT 2046.870 996.000 2047.150 1000.000 ;
        RECT 2049.170 999.870 2050.980 1000.000 ;
      LAYER met2 ;
        RECT 2047.430 995.720 2048.890 998.810 ;
      LAYER met2 ;
        RECT 2049.170 996.000 2049.450 999.870 ;
      LAYER met2 ;
        RECT 2049.730 995.720 2051.190 998.810 ;
      LAYER met2 ;
        RECT 2051.470 996.000 2051.750 1000.000 ;
      LAYER met2 ;
        RECT 2052.030 995.720 2053.030 998.810 ;
      LAYER met2 ;
        RECT 2053.310 996.000 2053.590 1000.000 ;
        RECT 2055.440 999.870 2055.890 1000.000 ;
      LAYER met2 ;
        RECT 2053.870 995.720 2055.330 998.810 ;
      LAYER met2 ;
        RECT 2055.610 996.000 2055.890 999.870 ;
      LAYER met2 ;
        RECT 2056.170 995.720 2057.630 998.810 ;
      LAYER met2 ;
        RECT 2057.910 996.000 2058.190 1000.000 ;
        RECT 2059.750 999.870 2061.560 1000.000 ;
      LAYER met2 ;
        RECT 2058.470 995.720 2059.470 998.810 ;
      LAYER met2 ;
        RECT 2059.750 996.000 2060.030 999.870 ;
      LAYER met2 ;
        RECT 2060.310 995.720 2061.770 998.810 ;
      LAYER met2 ;
        RECT 2062.050 996.000 2062.330 1000.000 ;
        RECT 2064.350 999.870 2066.160 1000.000 ;
      LAYER met2 ;
        RECT 2062.610 995.720 2064.070 998.810 ;
      LAYER met2 ;
        RECT 2064.350 996.000 2064.630 999.870 ;
      LAYER met2 ;
        RECT 2064.910 995.720 2066.370 998.810 ;
      LAYER met2 ;
        RECT 2066.650 996.000 2066.930 1000.000 ;
        RECT 2068.490 999.870 2069.840 1000.000 ;
      LAYER met2 ;
        RECT 2067.210 995.720 2068.210 998.810 ;
      LAYER met2 ;
        RECT 2068.490 996.000 2068.770 999.870 ;
      LAYER met2 ;
        RECT 2069.050 995.720 2070.510 998.810 ;
      LAYER met2 ;
        RECT 2070.790 996.000 2071.070 1000.000 ;
        RECT 2073.090 999.870 2074.900 1000.000 ;
      LAYER met2 ;
        RECT 2071.350 995.720 2072.810 998.810 ;
      LAYER met2 ;
        RECT 2073.090 996.000 2073.370 999.870 ;
      LAYER met2 ;
        RECT 2073.650 995.720 2075.110 998.810 ;
      LAYER met2 ;
        RECT 2075.390 996.000 2075.670 1000.000 ;
        RECT 2077.230 999.870 2079.040 1000.000 ;
      LAYER met2 ;
        RECT 2075.950 995.720 2076.950 998.810 ;
      LAYER met2 ;
        RECT 2077.230 996.000 2077.510 999.870 ;
      LAYER met2 ;
        RECT 2077.790 995.720 2079.250 998.810 ;
      LAYER met2 ;
        RECT 2079.530 996.000 2079.810 1000.000 ;
        RECT 2081.830 999.870 2082.260 1000.000 ;
      LAYER met2 ;
        RECT 2080.090 995.720 2081.550 998.810 ;
      LAYER met2 ;
        RECT 2081.830 996.000 2082.110 999.870 ;
      LAYER met2 ;
        RECT 2082.390 995.720 2083.390 998.810 ;
      LAYER met2 ;
        RECT 2083.670 996.000 2083.950 1000.000 ;
        RECT 2085.970 999.870 2087.780 1000.000 ;
      LAYER met2 ;
        RECT 2084.230 995.720 2085.690 998.810 ;
      LAYER met2 ;
        RECT 2085.970 996.000 2086.250 999.870 ;
      LAYER met2 ;
        RECT 2086.530 995.720 2087.990 998.810 ;
      LAYER met2 ;
        RECT 2088.270 996.000 2088.550 1000.000 ;
      LAYER met2 ;
        RECT 2088.830 995.720 2090.290 998.810 ;
      LAYER met2 ;
        RECT 2090.570 996.000 2090.850 1000.000 ;
      LAYER met2 ;
        RECT 2091.130 995.720 2092.130 998.810 ;
      LAYER met2 ;
        RECT 2092.410 996.000 2092.690 1000.000 ;
      LAYER met2 ;
        RECT 2092.970 995.720 2094.430 998.810 ;
      LAYER met2 ;
        RECT 2094.710 996.000 2094.990 1000.000 ;
      LAYER met2 ;
        RECT 2095.270 995.720 2096.730 998.810 ;
      LAYER met2 ;
        RECT 2097.010 996.000 2097.290 1000.000 ;
      LAYER met2 ;
        RECT 2097.570 995.720 2099.030 998.810 ;
      LAYER met2 ;
        RECT 2099.310 996.000 2099.590 1000.000 ;
      LAYER met2 ;
        RECT 2099.870 995.720 2100.870 998.810 ;
      LAYER met2 ;
        RECT 2101.150 996.000 2101.430 1000.000 ;
      LAYER met2 ;
        RECT 2101.710 995.720 2103.170 998.810 ;
      LAYER met2 ;
        RECT 2103.450 996.000 2103.730 1000.000 ;
      LAYER met2 ;
        RECT 2104.010 995.720 2105.470 998.810 ;
      LAYER met2 ;
        RECT 2105.750 996.000 2106.030 1000.000 ;
      LAYER met2 ;
        RECT 2106.310 995.720 2107.310 998.810 ;
      LAYER met2 ;
        RECT 2107.590 996.000 2107.870 1000.000 ;
      LAYER met2 ;
        RECT 2108.150 995.720 2109.610 998.810 ;
      LAYER met2 ;
        RECT 2109.890 996.000 2110.170 1000.000 ;
      LAYER met2 ;
        RECT 2110.450 995.720 2111.910 998.810 ;
      LAYER met2 ;
        RECT 2112.190 996.000 2112.470 1000.000 ;
      LAYER met2 ;
        RECT 2112.750 995.720 2114.210 998.810 ;
      LAYER met2 ;
        RECT 2114.490 996.000 2114.770 1000.000 ;
      LAYER met2 ;
        RECT 2115.050 995.720 2116.050 998.810 ;
      LAYER met2 ;
        RECT 2116.330 996.000 2116.610 1000.000 ;
      LAYER met2 ;
        RECT 2116.890 995.720 2118.350 998.810 ;
      LAYER met2 ;
        RECT 2118.630 996.000 2118.910 1000.000 ;
      LAYER met2 ;
        RECT 2119.190 995.720 2120.650 998.810 ;
      LAYER met2 ;
        RECT 2120.930 996.000 2121.210 1000.000 ;
      LAYER met2 ;
        RECT 2121.490 995.720 2122.950 998.810 ;
      LAYER met2 ;
        RECT 2123.230 996.000 2123.510 1000.000 ;
      LAYER met2 ;
        RECT 2123.790 995.720 2124.790 998.810 ;
      LAYER met2 ;
        RECT 2125.070 996.000 2125.350 1000.000 ;
      LAYER met2 ;
        RECT 2125.630 995.720 2127.090 998.810 ;
      LAYER met2 ;
        RECT 2127.370 996.000 2127.650 1000.000 ;
      LAYER met2 ;
        RECT 2127.930 995.720 2129.390 998.810 ;
      LAYER met2 ;
        RECT 2129.670 996.000 2129.950 1000.000 ;
      LAYER met2 ;
        RECT 2130.230 995.720 2131.230 998.810 ;
      LAYER met2 ;
        RECT 2131.510 996.000 2131.790 1000.000 ;
      LAYER met2 ;
        RECT 2132.070 995.720 2133.530 998.810 ;
      LAYER met2 ;
        RECT 2133.810 996.000 2134.090 1000.000 ;
      LAYER met2 ;
        RECT 2134.370 995.720 2135.830 998.810 ;
      LAYER met2 ;
        RECT 2136.110 996.000 2136.390 1000.000 ;
      LAYER met2 ;
        RECT 2136.670 995.720 2138.130 998.810 ;
      LAYER met2 ;
        RECT 2138.410 996.000 2138.690 1000.000 ;
      LAYER met2 ;
        RECT 2138.970 995.720 2139.970 998.810 ;
      LAYER met2 ;
        RECT 2140.250 996.000 2140.530 1000.000 ;
      LAYER met2 ;
        RECT 2140.810 995.720 2142.270 998.810 ;
      LAYER met2 ;
        RECT 2142.550 996.000 2142.830 1000.000 ;
      LAYER met2 ;
        RECT 2143.110 995.720 2144.570 998.810 ;
      LAYER met2 ;
        RECT 2144.850 996.000 2145.130 1000.000 ;
      LAYER met2 ;
        RECT 2145.410 995.720 2146.870 998.810 ;
      LAYER met2 ;
        RECT 2147.150 996.000 2147.430 1000.000 ;
      LAYER met2 ;
        RECT 2147.710 995.720 2148.710 998.810 ;
      LAYER met2 ;
        RECT 2148.990 996.000 2149.270 1000.000 ;
      LAYER met2 ;
        RECT 2149.550 995.720 2151.010 998.810 ;
      LAYER met2 ;
        RECT 2151.290 996.000 2151.570 1000.000 ;
      LAYER met2 ;
        RECT 2151.850 995.720 2153.310 998.810 ;
      LAYER met2 ;
        RECT 2153.590 996.000 2153.870 1000.000 ;
      LAYER met2 ;
        RECT 2154.150 995.720 2155.150 998.810 ;
      LAYER met2 ;
        RECT 2155.430 996.000 2155.710 1000.000 ;
      LAYER met2 ;
        RECT 2155.990 995.720 2157.450 998.810 ;
      LAYER met2 ;
        RECT 2157.730 996.000 2158.010 1000.000 ;
      LAYER met2 ;
        RECT 2158.290 995.720 2159.750 998.810 ;
      LAYER met2 ;
        RECT 2160.030 996.000 2160.310 1000.000 ;
      LAYER met2 ;
        RECT 2160.590 995.720 2162.050 998.810 ;
      LAYER met2 ;
        RECT 2162.330 996.000 2162.610 1000.000 ;
      LAYER met2 ;
        RECT 2162.890 995.720 2163.890 998.810 ;
      LAYER met2 ;
        RECT 2164.170 996.000 2164.450 1000.000 ;
      LAYER met2 ;
        RECT 2164.730 995.720 2166.190 998.810 ;
      LAYER met2 ;
        RECT 2166.470 996.000 2166.750 1000.000 ;
      LAYER met2 ;
        RECT 2167.030 995.720 2168.490 998.810 ;
      LAYER met2 ;
        RECT 2168.770 996.000 2169.050 1000.000 ;
      LAYER met2 ;
        RECT 671.020 604.280 2169.040 995.720 ;
        RECT 671.020 602.195 671.190 604.280 ;
        RECT 672.030 602.195 673.950 604.280 ;
        RECT 674.790 602.195 677.170 604.280 ;
        RECT 678.010 602.195 679.930 604.280 ;
        RECT 680.770 602.195 683.150 604.280 ;
        RECT 683.990 602.195 686.370 604.280 ;
        RECT 687.210 602.195 689.130 604.280 ;
        RECT 689.970 602.195 692.350 604.280 ;
        RECT 693.190 602.195 695.570 604.280 ;
        RECT 696.410 602.195 698.330 604.280 ;
        RECT 699.170 602.195 701.550 604.280 ;
        RECT 702.390 602.195 704.770 604.280 ;
        RECT 705.610 602.195 707.530 604.280 ;
        RECT 708.370 602.195 710.750 604.280 ;
        RECT 711.590 602.195 713.970 604.280 ;
        RECT 714.810 602.195 716.730 604.280 ;
        RECT 717.570 602.195 719.950 604.280 ;
        RECT 720.790 602.195 723.170 604.280 ;
        RECT 724.010 602.195 725.930 604.280 ;
        RECT 726.770 602.195 729.150 604.280 ;
        RECT 729.990 602.195 732.370 604.280 ;
        RECT 733.210 602.195 735.130 604.280 ;
        RECT 735.970 602.195 738.350 604.280 ;
        RECT 739.190 602.195 741.570 604.280 ;
        RECT 742.410 602.195 744.330 604.280 ;
        RECT 745.170 602.195 747.550 604.280 ;
        RECT 748.390 602.195 750.770 604.280 ;
        RECT 751.610 602.195 753.530 604.280 ;
        RECT 754.370 602.195 756.750 604.280 ;
        RECT 757.590 602.195 759.510 604.280 ;
        RECT 760.350 602.195 762.730 604.280 ;
        RECT 763.570 602.195 765.950 604.280 ;
        RECT 766.790 602.195 768.710 604.280 ;
        RECT 769.550 602.195 771.930 604.280 ;
        RECT 772.770 602.195 775.150 604.280 ;
        RECT 775.990 602.195 777.910 604.280 ;
        RECT 778.750 602.195 781.130 604.280 ;
        RECT 781.970 602.195 784.350 604.280 ;
        RECT 785.190 602.195 787.110 604.280 ;
        RECT 787.950 602.195 790.330 604.280 ;
        RECT 791.170 602.195 793.550 604.280 ;
        RECT 794.390 602.195 796.310 604.280 ;
        RECT 797.150 602.195 799.530 604.280 ;
        RECT 800.370 602.195 802.750 604.280 ;
        RECT 803.590 602.195 805.510 604.280 ;
        RECT 806.350 602.195 808.730 604.280 ;
        RECT 809.570 602.195 811.950 604.280 ;
        RECT 812.790 602.195 814.710 604.280 ;
        RECT 815.550 602.195 817.930 604.280 ;
        RECT 818.770 602.195 821.150 604.280 ;
        RECT 821.990 602.195 823.910 604.280 ;
        RECT 824.750 602.195 827.130 604.280 ;
        RECT 827.970 602.195 830.350 604.280 ;
        RECT 831.190 602.195 833.110 604.280 ;
        RECT 833.950 602.195 836.330 604.280 ;
        RECT 837.170 602.195 839.550 604.280 ;
        RECT 840.390 602.195 842.310 604.280 ;
        RECT 843.150 602.195 845.530 604.280 ;
        RECT 846.370 602.195 848.290 604.280 ;
        RECT 849.130 602.195 851.510 604.280 ;
        RECT 852.350 602.195 854.730 604.280 ;
        RECT 855.570 602.195 857.490 604.280 ;
        RECT 858.330 602.195 860.710 604.280 ;
        RECT 861.550 602.195 863.930 604.280 ;
        RECT 864.770 602.195 866.690 604.280 ;
        RECT 867.530 602.195 869.910 604.280 ;
        RECT 870.750 602.195 873.130 604.280 ;
        RECT 873.970 602.195 875.890 604.280 ;
        RECT 876.730 602.195 879.110 604.280 ;
        RECT 879.950 602.195 882.330 604.280 ;
        RECT 883.170 602.195 885.090 604.280 ;
        RECT 885.930 602.195 888.310 604.280 ;
        RECT 889.150 602.195 891.530 604.280 ;
        RECT 892.370 602.195 894.290 604.280 ;
        RECT 895.130 602.195 897.510 604.280 ;
        RECT 898.350 602.195 900.730 604.280 ;
        RECT 901.570 602.195 903.490 604.280 ;
        RECT 904.330 602.195 906.710 604.280 ;
        RECT 907.550 602.195 909.930 604.280 ;
        RECT 910.770 602.195 912.690 604.280 ;
        RECT 913.530 602.195 915.910 604.280 ;
        RECT 916.750 602.195 919.130 604.280 ;
        RECT 919.970 602.195 921.890 604.280 ;
        RECT 922.730 602.195 925.110 604.280 ;
        RECT 925.950 602.195 928.330 604.280 ;
        RECT 929.170 602.195 931.090 604.280 ;
        RECT 931.930 602.195 934.310 604.280 ;
        RECT 935.150 602.195 937.070 604.280 ;
        RECT 937.910 602.195 940.290 604.280 ;
        RECT 941.130 602.195 943.510 604.280 ;
        RECT 944.350 602.195 946.270 604.280 ;
        RECT 947.110 602.195 949.490 604.280 ;
        RECT 950.330 602.195 952.710 604.280 ;
        RECT 953.550 602.195 955.470 604.280 ;
        RECT 956.310 602.195 958.690 604.280 ;
        RECT 959.530 602.195 961.910 604.280 ;
        RECT 962.750 602.195 964.670 604.280 ;
        RECT 965.510 602.195 967.890 604.280 ;
        RECT 968.730 602.195 971.110 604.280 ;
        RECT 971.950 602.195 973.870 604.280 ;
        RECT 974.710 602.195 977.090 604.280 ;
        RECT 977.930 602.195 980.310 604.280 ;
        RECT 981.150 602.195 983.070 604.280 ;
        RECT 983.910 602.195 986.290 604.280 ;
        RECT 987.130 602.195 989.510 604.280 ;
        RECT 990.350 602.195 992.270 604.280 ;
        RECT 993.110 602.195 995.490 604.280 ;
        RECT 996.330 602.195 998.710 604.280 ;
        RECT 999.550 602.195 1001.470 604.280 ;
        RECT 1002.310 602.195 1004.690 604.280 ;
        RECT 1005.530 602.195 1007.910 604.280 ;
        RECT 1008.750 602.195 1010.670 604.280 ;
        RECT 1011.510 602.195 1013.890 604.280 ;
        RECT 1014.730 602.195 1017.110 604.280 ;
        RECT 1017.950 602.195 1019.870 604.280 ;
        RECT 1020.710 602.195 1023.090 604.280 ;
        RECT 1023.930 602.195 1025.850 604.280 ;
        RECT 1026.690 602.195 1029.070 604.280 ;
        RECT 1029.910 602.195 1032.290 604.280 ;
        RECT 1033.130 602.195 1035.050 604.280 ;
        RECT 1035.890 602.195 1038.270 604.280 ;
        RECT 1039.110 602.195 1041.490 604.280 ;
        RECT 1042.330 602.195 1044.250 604.280 ;
        RECT 1045.090 602.195 1047.470 604.280 ;
        RECT 1048.310 602.195 1050.690 604.280 ;
        RECT 1051.530 602.195 1053.450 604.280 ;
        RECT 1054.290 602.195 1056.670 604.280 ;
        RECT 1057.510 602.195 1059.890 604.280 ;
        RECT 1060.730 602.195 1062.650 604.280 ;
        RECT 1063.490 602.195 1065.870 604.280 ;
        RECT 1066.710 602.195 1069.090 604.280 ;
        RECT 1069.930 602.195 1071.850 604.280 ;
        RECT 1072.690 602.195 1075.070 604.280 ;
        RECT 1075.910 602.195 1078.290 604.280 ;
        RECT 1079.130 602.195 1081.050 604.280 ;
        RECT 1081.890 602.195 1084.270 604.280 ;
        RECT 1085.110 602.195 1087.490 604.280 ;
        RECT 1088.330 602.195 1090.250 604.280 ;
        RECT 1091.090 602.195 1093.470 604.280 ;
        RECT 1094.310 602.195 1096.690 604.280 ;
        RECT 1097.530 602.195 1099.450 604.280 ;
        RECT 1100.290 602.195 1102.670 604.280 ;
        RECT 1103.510 602.195 1105.890 604.280 ;
        RECT 1106.730 602.195 1108.650 604.280 ;
        RECT 1109.490 602.195 1111.870 604.280 ;
        RECT 1112.710 602.195 1114.630 604.280 ;
        RECT 1115.470 602.195 1117.850 604.280 ;
        RECT 1118.690 602.195 1121.070 604.280 ;
        RECT 1121.910 602.195 1123.830 604.280 ;
        RECT 1124.670 602.195 1127.050 604.280 ;
        RECT 1127.890 602.195 1130.270 604.280 ;
        RECT 1131.110 602.195 1133.030 604.280 ;
        RECT 1133.870 602.195 1136.250 604.280 ;
        RECT 1137.090 602.195 1139.470 604.280 ;
        RECT 1140.310 602.195 1142.230 604.280 ;
        RECT 1143.070 602.195 1145.450 604.280 ;
        RECT 1146.290 602.195 1148.670 604.280 ;
        RECT 1149.510 602.195 1151.430 604.280 ;
        RECT 1152.270 602.195 1154.650 604.280 ;
        RECT 1155.490 602.195 1157.870 604.280 ;
        RECT 1158.710 602.195 1160.630 604.280 ;
        RECT 1161.470 602.195 1163.850 604.280 ;
        RECT 1164.690 602.195 1167.070 604.280 ;
        RECT 1167.910 602.195 1169.830 604.280 ;
        RECT 1170.670 602.195 1173.050 604.280 ;
        RECT 1173.890 602.195 1176.270 604.280 ;
        RECT 1177.110 602.195 1179.030 604.280 ;
        RECT 1179.870 602.195 1182.250 604.280 ;
        RECT 1183.090 602.195 1185.470 604.280 ;
        RECT 1186.310 602.195 1188.230 604.280 ;
        RECT 1189.070 602.195 1191.450 604.280 ;
        RECT 1192.290 602.195 1194.670 604.280 ;
        RECT 1195.510 602.195 1197.430 604.280 ;
        RECT 1198.270 602.195 1200.650 604.280 ;
        RECT 1201.490 602.195 1203.410 604.280 ;
        RECT 1204.250 602.195 1206.630 604.280 ;
        RECT 1207.470 602.195 1209.850 604.280 ;
        RECT 1210.690 602.195 1212.610 604.280 ;
        RECT 1213.450 602.195 1215.830 604.280 ;
        RECT 1216.670 602.195 1219.050 604.280 ;
        RECT 1219.890 602.195 1221.810 604.280 ;
        RECT 1222.650 602.195 1225.030 604.280 ;
        RECT 1225.870 602.195 1228.250 604.280 ;
        RECT 1229.090 602.195 1231.010 604.280 ;
        RECT 1231.850 602.195 1234.230 604.280 ;
        RECT 1235.070 602.195 1237.450 604.280 ;
        RECT 1238.290 602.195 1240.210 604.280 ;
        RECT 1241.050 602.195 1243.430 604.280 ;
        RECT 1244.270 602.195 1246.650 604.280 ;
        RECT 1247.490 602.195 1249.410 604.280 ;
        RECT 1250.250 602.195 1252.630 604.280 ;
        RECT 1253.470 602.195 1255.850 604.280 ;
        RECT 1256.690 602.195 1258.610 604.280 ;
        RECT 1259.450 602.195 1261.830 604.280 ;
        RECT 1262.670 602.195 1265.050 604.280 ;
        RECT 1265.890 602.195 1267.810 604.280 ;
        RECT 1268.650 602.195 1271.030 604.280 ;
        RECT 1271.870 602.195 1274.250 604.280 ;
        RECT 1275.090 602.195 1277.010 604.280 ;
        RECT 1277.850 602.195 1280.230 604.280 ;
        RECT 1281.070 602.195 1283.450 604.280 ;
        RECT 1284.290 602.195 1286.210 604.280 ;
        RECT 1287.050 602.195 1289.430 604.280 ;
        RECT 1290.270 602.195 1292.190 604.280 ;
        RECT 1293.030 602.195 1295.410 604.280 ;
        RECT 1296.250 602.195 1298.630 604.280 ;
        RECT 1299.470 602.195 1301.390 604.280 ;
        RECT 1302.230 602.195 1304.610 604.280 ;
        RECT 1305.450 602.195 1307.830 604.280 ;
        RECT 1308.670 602.195 1310.590 604.280 ;
        RECT 1311.430 602.195 1313.810 604.280 ;
        RECT 1314.650 602.195 1317.030 604.280 ;
        RECT 1317.870 602.195 1319.790 604.280 ;
        RECT 1320.630 602.195 1323.010 604.280 ;
        RECT 1323.850 602.195 1326.230 604.280 ;
        RECT 1327.070 602.195 1328.990 604.280 ;
        RECT 1329.830 602.195 1332.210 604.280 ;
        RECT 1333.050 602.195 1335.430 604.280 ;
        RECT 1336.270 602.195 1338.190 604.280 ;
        RECT 1339.030 602.195 1341.410 604.280 ;
        RECT 1342.250 602.195 1344.630 604.280 ;
        RECT 1345.470 602.195 1347.390 604.280 ;
        RECT 1348.230 602.195 1350.610 604.280 ;
        RECT 1351.450 602.195 1353.830 604.280 ;
        RECT 1354.670 602.195 1356.590 604.280 ;
        RECT 1357.430 602.195 1359.810 604.280 ;
        RECT 1360.650 602.195 1363.030 604.280 ;
        RECT 1363.870 602.195 1365.790 604.280 ;
        RECT 1366.630 602.195 1369.010 604.280 ;
        RECT 1369.850 602.195 1372.230 604.280 ;
        RECT 1373.070 602.195 1374.990 604.280 ;
        RECT 1375.830 602.195 1378.210 604.280 ;
        RECT 1379.050 602.195 1380.970 604.280 ;
        RECT 1381.810 602.195 1384.190 604.280 ;
        RECT 1385.030 602.195 1387.410 604.280 ;
        RECT 1388.250 602.195 1390.170 604.280 ;
        RECT 1391.010 602.195 1393.390 604.280 ;
        RECT 1394.230 602.195 1396.610 604.280 ;
        RECT 1397.450 602.195 1399.370 604.280 ;
        RECT 1400.210 602.195 1402.590 604.280 ;
        RECT 1403.430 602.195 1405.810 604.280 ;
        RECT 1406.650 602.195 1408.570 604.280 ;
        RECT 1409.410 602.195 1411.790 604.280 ;
        RECT 1412.630 602.195 1415.010 604.280 ;
        RECT 1415.850 602.195 1417.770 604.280 ;
        RECT 1418.610 602.195 1420.990 604.280 ;
        RECT 1421.830 602.195 1424.210 604.280 ;
        RECT 1425.050 602.195 1426.970 604.280 ;
        RECT 1427.810 602.195 1430.190 604.280 ;
        RECT 1431.030 602.195 1433.410 604.280 ;
        RECT 1434.250 602.195 1436.170 604.280 ;
        RECT 1437.010 602.195 1439.390 604.280 ;
        RECT 1440.230 602.195 1442.610 604.280 ;
        RECT 1443.450 602.195 1445.370 604.280 ;
        RECT 1446.210 602.195 1448.590 604.280 ;
        RECT 1449.430 602.195 1451.810 604.280 ;
        RECT 1452.650 602.195 1454.570 604.280 ;
        RECT 1455.410 602.195 1457.790 604.280 ;
        RECT 1458.630 602.195 1461.010 604.280 ;
        RECT 1461.850 602.195 1463.770 604.280 ;
        RECT 1464.610 602.195 1466.990 604.280 ;
        RECT 1467.830 602.195 1469.750 604.280 ;
        RECT 1470.590 602.195 1472.970 604.280 ;
        RECT 1473.810 602.195 1476.190 604.280 ;
        RECT 1477.030 602.195 1478.950 604.280 ;
        RECT 1479.790 602.195 1482.170 604.280 ;
        RECT 1483.010 602.195 1485.390 604.280 ;
        RECT 1486.230 602.195 1488.150 604.280 ;
        RECT 1488.990 602.195 1491.370 604.280 ;
        RECT 1492.210 602.195 1494.590 604.280 ;
        RECT 1495.430 602.195 1497.350 604.280 ;
        RECT 1498.190 602.195 1500.570 604.280 ;
        RECT 1501.410 602.195 1503.790 604.280 ;
        RECT 1504.630 602.195 1506.550 604.280 ;
        RECT 1507.390 602.195 1509.770 604.280 ;
        RECT 1510.610 602.195 1512.990 604.280 ;
        RECT 1513.830 602.195 1515.750 604.280 ;
        RECT 1516.590 602.195 1518.970 604.280 ;
        RECT 1519.810 602.195 1522.190 604.280 ;
        RECT 1523.030 602.195 1524.950 604.280 ;
        RECT 1525.790 602.195 1528.170 604.280 ;
        RECT 1529.010 602.195 1531.390 604.280 ;
        RECT 1532.230 602.195 1534.150 604.280 ;
        RECT 1534.990 602.195 1537.370 604.280 ;
        RECT 1538.210 602.195 1540.590 604.280 ;
        RECT 1541.430 602.195 1543.350 604.280 ;
        RECT 1544.190 602.195 1546.570 604.280 ;
        RECT 1547.410 602.195 1549.790 604.280 ;
        RECT 1550.630 602.195 1552.550 604.280 ;
        RECT 1553.390 602.195 1555.770 604.280 ;
        RECT 1556.610 602.195 1558.530 604.280 ;
        RECT 1559.370 602.195 1561.750 604.280 ;
        RECT 1562.590 602.195 1564.970 604.280 ;
        RECT 1565.810 602.195 1567.730 604.280 ;
        RECT 1568.570 602.195 1570.950 604.280 ;
        RECT 1571.790 602.195 1574.170 604.280 ;
        RECT 1575.010 602.195 1576.930 604.280 ;
        RECT 1577.770 602.195 1580.150 604.280 ;
        RECT 1580.990 602.195 1583.370 604.280 ;
        RECT 1584.210 602.195 1586.130 604.280 ;
        RECT 1586.970 602.195 1589.350 604.280 ;
        RECT 1590.190 602.195 1592.570 604.280 ;
        RECT 1593.410 602.195 1595.330 604.280 ;
        RECT 1596.170 602.195 1598.550 604.280 ;
        RECT 1599.390 602.195 1601.770 604.280 ;
        RECT 1602.610 602.195 1604.530 604.280 ;
        RECT 1605.370 602.195 1607.750 604.280 ;
        RECT 1608.590 602.195 1610.970 604.280 ;
        RECT 1611.810 602.195 1613.730 604.280 ;
        RECT 1614.570 602.195 1616.950 604.280 ;
        RECT 1617.790 602.195 1620.170 604.280 ;
        RECT 1621.010 602.195 1622.930 604.280 ;
        RECT 1623.770 602.195 1626.150 604.280 ;
        RECT 1626.990 602.195 1629.370 604.280 ;
        RECT 1630.210 602.195 1632.130 604.280 ;
        RECT 1632.970 602.195 1635.350 604.280 ;
        RECT 1636.190 602.195 1638.570 604.280 ;
        RECT 1639.410 602.195 1641.330 604.280 ;
        RECT 1642.170 602.195 1644.550 604.280 ;
        RECT 1645.390 602.195 1647.310 604.280 ;
        RECT 1648.150 602.195 1650.530 604.280 ;
        RECT 1651.370 602.195 1653.750 604.280 ;
        RECT 1654.590 602.195 1656.510 604.280 ;
        RECT 1657.350 602.195 1659.730 604.280 ;
        RECT 1660.570 602.195 1662.950 604.280 ;
        RECT 1663.790 602.195 1665.710 604.280 ;
        RECT 1666.550 602.195 1668.930 604.280 ;
        RECT 1669.770 602.195 1672.150 604.280 ;
        RECT 1672.990 602.195 1674.910 604.280 ;
        RECT 1675.750 602.195 1678.130 604.280 ;
        RECT 1678.970 602.195 1681.350 604.280 ;
        RECT 1682.190 602.195 1684.110 604.280 ;
        RECT 1684.950 602.195 1687.330 604.280 ;
        RECT 1688.170 602.195 1690.550 604.280 ;
        RECT 1691.390 602.195 1693.310 604.280 ;
        RECT 1694.150 602.195 1696.530 604.280 ;
        RECT 1697.370 602.195 1699.750 604.280 ;
        RECT 1700.590 602.195 1702.510 604.280 ;
        RECT 1703.350 602.195 1705.730 604.280 ;
        RECT 1706.570 602.195 1708.950 604.280 ;
        RECT 1709.790 602.195 1711.710 604.280 ;
        RECT 1712.550 602.195 1714.930 604.280 ;
        RECT 1715.770 602.195 1718.150 604.280 ;
        RECT 1718.990 602.195 1720.910 604.280 ;
        RECT 1721.750 602.195 1724.130 604.280 ;
        RECT 1724.970 602.195 1727.350 604.280 ;
        RECT 1728.190 602.195 1730.110 604.280 ;
        RECT 1730.950 602.195 1733.330 604.280 ;
        RECT 1734.170 602.195 1736.090 604.280 ;
        RECT 1736.930 602.195 1739.310 604.280 ;
        RECT 1740.150 602.195 1742.530 604.280 ;
        RECT 1743.370 602.195 1745.290 604.280 ;
        RECT 1746.130 602.195 1748.510 604.280 ;
        RECT 1749.350 602.195 1751.730 604.280 ;
        RECT 1752.570 602.195 1754.490 604.280 ;
        RECT 1755.330 602.195 1757.710 604.280 ;
        RECT 1758.550 602.195 1760.930 604.280 ;
        RECT 1761.770 602.195 1763.690 604.280 ;
        RECT 1764.530 602.195 1766.910 604.280 ;
        RECT 1767.750 602.195 1770.130 604.280 ;
        RECT 1770.970 602.195 1772.890 604.280 ;
        RECT 1773.730 602.195 1776.110 604.280 ;
        RECT 1776.950 602.195 1779.330 604.280 ;
        RECT 1780.170 602.195 1782.090 604.280 ;
        RECT 1782.930 602.195 1785.310 604.280 ;
        RECT 1786.150 602.195 1788.530 604.280 ;
        RECT 1789.370 602.195 1791.290 604.280 ;
        RECT 1792.130 602.195 1794.510 604.280 ;
        RECT 1795.350 602.195 1797.730 604.280 ;
        RECT 1798.570 602.195 1800.490 604.280 ;
        RECT 1801.330 602.195 1803.710 604.280 ;
        RECT 1804.550 602.195 1806.930 604.280 ;
        RECT 1807.770 602.195 1809.690 604.280 ;
        RECT 1810.530 602.195 1812.910 604.280 ;
        RECT 1813.750 602.195 1816.130 604.280 ;
        RECT 1816.970 602.195 1818.890 604.280 ;
        RECT 1819.730 602.195 1822.110 604.280 ;
        RECT 1822.950 602.195 1824.870 604.280 ;
        RECT 1825.710 602.195 1828.090 604.280 ;
        RECT 1828.930 602.195 1831.310 604.280 ;
        RECT 1832.150 602.195 1834.070 604.280 ;
        RECT 1834.910 602.195 1837.290 604.280 ;
        RECT 1838.130 602.195 1840.510 604.280 ;
        RECT 1841.350 602.195 1843.270 604.280 ;
        RECT 1844.110 602.195 1846.490 604.280 ;
        RECT 1847.330 602.195 1849.710 604.280 ;
        RECT 1850.550 602.195 1852.470 604.280 ;
        RECT 1853.310 602.195 1855.690 604.280 ;
        RECT 1856.530 602.195 1858.910 604.280 ;
        RECT 1859.750 602.195 1861.670 604.280 ;
        RECT 1862.510 602.195 1864.890 604.280 ;
        RECT 1865.730 602.195 1868.110 604.280 ;
        RECT 1868.950 602.195 1870.870 604.280 ;
        RECT 1871.710 602.195 1874.090 604.280 ;
        RECT 1874.930 602.195 1877.310 604.280 ;
        RECT 1878.150 602.195 1880.070 604.280 ;
        RECT 1880.910 602.195 1883.290 604.280 ;
        RECT 1884.130 602.195 1886.510 604.280 ;
        RECT 1887.350 602.195 1889.270 604.280 ;
        RECT 1890.110 602.195 1892.490 604.280 ;
        RECT 1893.330 602.195 1895.710 604.280 ;
        RECT 1896.550 602.195 1898.470 604.280 ;
        RECT 1899.310 602.195 1901.690 604.280 ;
        RECT 1902.530 602.195 1904.910 604.280 ;
        RECT 1905.750 602.195 1907.670 604.280 ;
        RECT 1908.510 602.195 1910.890 604.280 ;
        RECT 1911.730 602.195 1913.650 604.280 ;
        RECT 1914.490 602.195 1916.870 604.280 ;
        RECT 1917.710 602.195 1920.090 604.280 ;
        RECT 1920.930 602.195 1922.850 604.280 ;
        RECT 1923.690 602.195 1926.070 604.280 ;
        RECT 1926.910 602.195 1929.290 604.280 ;
        RECT 1930.130 602.195 1932.050 604.280 ;
        RECT 1932.890 602.195 1935.270 604.280 ;
        RECT 1936.110 602.195 1938.490 604.280 ;
        RECT 1939.330 602.195 1941.250 604.280 ;
        RECT 1942.090 602.195 1944.470 604.280 ;
        RECT 1945.310 602.195 1947.690 604.280 ;
        RECT 1948.530 602.195 1950.450 604.280 ;
        RECT 1951.290 602.195 1953.670 604.280 ;
        RECT 1954.510 602.195 1956.890 604.280 ;
        RECT 1957.730 602.195 1959.650 604.280 ;
        RECT 1960.490 602.195 1962.870 604.280 ;
        RECT 1963.710 602.195 1966.090 604.280 ;
        RECT 1966.930 602.195 1968.850 604.280 ;
        RECT 1969.690 602.195 1972.070 604.280 ;
        RECT 1972.910 602.195 1975.290 604.280 ;
        RECT 1976.130 602.195 1978.050 604.280 ;
        RECT 1978.890 602.195 1981.270 604.280 ;
        RECT 1982.110 602.195 1984.490 604.280 ;
        RECT 1985.330 602.195 1987.250 604.280 ;
        RECT 1988.090 602.195 1990.470 604.280 ;
        RECT 1991.310 602.195 1993.690 604.280 ;
        RECT 1994.530 602.195 1996.450 604.280 ;
        RECT 1997.290 602.195 1999.670 604.280 ;
        RECT 2000.510 602.195 2002.430 604.280 ;
        RECT 2003.270 602.195 2005.650 604.280 ;
        RECT 2006.490 602.195 2008.870 604.280 ;
        RECT 2009.710 602.195 2011.630 604.280 ;
        RECT 2012.470 602.195 2014.850 604.280 ;
        RECT 2015.690 602.195 2018.070 604.280 ;
        RECT 2018.910 602.195 2020.830 604.280 ;
        RECT 2021.670 602.195 2024.050 604.280 ;
        RECT 2024.890 602.195 2027.270 604.280 ;
        RECT 2028.110 602.195 2030.030 604.280 ;
        RECT 2030.870 602.195 2033.250 604.280 ;
        RECT 2034.090 602.195 2036.470 604.280 ;
        RECT 2037.310 602.195 2039.230 604.280 ;
        RECT 2040.070 602.195 2042.450 604.280 ;
        RECT 2043.290 602.195 2045.670 604.280 ;
        RECT 2046.510 602.195 2048.430 604.280 ;
        RECT 2049.270 602.195 2051.650 604.280 ;
        RECT 2052.490 602.195 2054.870 604.280 ;
        RECT 2055.710 602.195 2057.630 604.280 ;
        RECT 2058.470 602.195 2060.850 604.280 ;
        RECT 2061.690 602.195 2064.070 604.280 ;
        RECT 2064.910 602.195 2066.830 604.280 ;
        RECT 2067.670 602.195 2070.050 604.280 ;
        RECT 2070.890 602.195 2073.270 604.280 ;
        RECT 2074.110 602.195 2076.030 604.280 ;
        RECT 2076.870 602.195 2079.250 604.280 ;
        RECT 2080.090 602.195 2082.470 604.280 ;
        RECT 2083.310 602.195 2085.230 604.280 ;
        RECT 2086.070 602.195 2088.450 604.280 ;
        RECT 2089.290 602.195 2091.210 604.280 ;
        RECT 2092.050 602.195 2094.430 604.280 ;
        RECT 2095.270 602.195 2097.650 604.280 ;
        RECT 2098.490 602.195 2100.410 604.280 ;
        RECT 2101.250 602.195 2103.630 604.280 ;
        RECT 2104.470 602.195 2106.850 604.280 ;
        RECT 2107.690 602.195 2109.610 604.280 ;
        RECT 2110.450 602.195 2112.830 604.280 ;
        RECT 2113.670 602.195 2116.050 604.280 ;
        RECT 2116.890 602.195 2118.810 604.280 ;
        RECT 2119.650 602.195 2122.030 604.280 ;
        RECT 2122.870 602.195 2125.250 604.280 ;
        RECT 2126.090 602.195 2128.010 604.280 ;
        RECT 2128.850 602.195 2131.230 604.280 ;
        RECT 2132.070 602.195 2134.450 604.280 ;
        RECT 2135.290 602.195 2137.210 604.280 ;
        RECT 2138.050 602.195 2140.430 604.280 ;
        RECT 2141.270 602.195 2143.650 604.280 ;
        RECT 2144.490 602.195 2146.410 604.280 ;
        RECT 2147.250 602.195 2149.630 604.280 ;
        RECT 2150.470 602.195 2152.850 604.280 ;
        RECT 2153.690 602.195 2155.610 604.280 ;
        RECT 2156.450 602.195 2158.830 604.280 ;
        RECT 2159.670 602.195 2162.050 604.280 ;
        RECT 2162.890 602.195 2164.810 604.280 ;
        RECT 2165.650 602.195 2168.030 604.280 ;
        RECT 2168.870 602.195 2169.040 604.280 ;
      LAYER via2 ;
        RECT 420.530 2729.040 420.810 2729.320 ;
        RECT 420.070 2707.280 420.350 2707.560 ;
        RECT 586.590 2686.880 586.870 2687.160 ;
        RECT 586.590 2666.480 586.870 2666.760 ;
        RECT 985.410 1014.080 985.690 1014.360 ;
        RECT 984.950 1013.400 985.230 1013.680 ;
        RECT 1058.090 2808.600 1058.370 2808.880 ;
        RECT 993.230 2670.560 993.510 2670.840 ;
        RECT 992.770 2622.960 993.050 2623.240 ;
        RECT 990.010 1893.320 990.290 1893.600 ;
        RECT 989.550 1871.560 989.830 1871.840 ;
        RECT 989.090 1851.160 989.370 1851.440 ;
        RECT 988.630 1809.000 988.910 1809.280 ;
        RECT 987.710 1787.240 987.990 1787.520 ;
        RECT 987.250 1766.840 987.530 1767.120 ;
        RECT 986.790 1745.080 987.070 1745.360 ;
        RECT 988.170 1724.680 988.450 1724.960 ;
        RECT 986.330 1012.040 986.610 1012.320 ;
        RECT 985.870 1010.680 986.150 1010.960 ;
        RECT 992.310 1998.040 992.590 1998.320 ;
        RECT 991.850 1935.480 992.130 1935.760 ;
        RECT 993.690 2646.080 993.970 2646.360 ;
        RECT 994.150 2018.440 994.430 2018.720 ;
        RECT 994.610 1976.280 994.890 1976.560 ;
        RECT 995.070 1955.880 995.350 1956.160 ;
        RECT 995.530 1913.720 995.810 1914.000 ;
        RECT 995.990 1829.400 996.270 1829.680 ;
        RECT 1110.990 2780.720 1111.270 2781.000 ;
        RECT 1016.690 2051.760 1016.970 2052.040 ;
        RECT 1111.450 2760.320 1111.730 2760.600 ;
        RECT 1112.830 2734.480 1113.110 2734.760 ;
        RECT 1112.370 2712.720 1112.650 2713.000 ;
        RECT 1111.910 2691.640 1112.190 2691.920 ;
        RECT 1113.290 2666.480 1113.570 2666.760 ;
        RECT 1113.750 2644.720 1114.030 2645.000 ;
        RECT 1114.210 2622.280 1114.490 2622.560 ;
        RECT 1130.770 2050.400 1131.050 2050.680 ;
        RECT 1159.290 2051.080 1159.570 2051.360 ;
        RECT 1315.690 2049.720 1315.970 2050.000 ;
        RECT 1062.690 1009.320 1062.970 1009.600 ;
        RECT 1055.790 1007.960 1056.070 1008.240 ;
        RECT 1067.290 1008.640 1067.570 1008.920 ;
        RECT 1090.290 1010.000 1090.570 1010.280 ;
        RECT 1101.790 1014.080 1102.070 1014.360 ;
        RECT 1185.970 1693.400 1186.250 1693.680 ;
        RECT 1119.270 1013.400 1119.550 1013.680 ;
        RECT 1111.450 1008.640 1111.730 1008.920 ;
        RECT 1125.710 1012.720 1125.990 1013.000 ;
        RECT 1131.690 1012.040 1131.970 1012.320 ;
        RECT 1146.410 1009.320 1146.690 1009.600 ;
        RECT 1158.370 1012.040 1158.650 1012.320 ;
        RECT 1160.670 1011.360 1160.950 1011.640 ;
        RECT 1160.210 1010.000 1160.490 1010.280 ;
        RECT 1158.370 1008.640 1158.650 1008.920 ;
        RECT 1159.290 1008.640 1159.570 1008.920 ;
        RECT 1159.750 1007.960 1160.030 1008.240 ;
        RECT 1161.130 1008.640 1161.410 1008.920 ;
        RECT 1167.110 1010.680 1167.390 1010.960 ;
        RECT 1166.650 1007.960 1166.930 1008.240 ;
        RECT 1176.310 1009.320 1176.590 1009.600 ;
        RECT 1191.490 1010.000 1191.770 1010.280 ;
        RECT 1200.230 1012.040 1200.510 1012.320 ;
        RECT 1207.590 1008.640 1207.870 1008.920 ;
        RECT 1207.590 1007.960 1207.870 1008.240 ;
        RECT 1209.430 1008.640 1209.710 1008.920 ;
        RECT 1209.430 1007.960 1209.710 1008.240 ;
        RECT 1285.330 1010.680 1285.610 1010.960 ;
        RECT 1313.390 1007.960 1313.670 1008.240 ;
        RECT 1330.870 1007.280 1331.150 1007.560 ;
        RECT 1335.930 1998.040 1336.210 1998.320 ;
        RECT 1336.390 1787.240 1336.670 1787.520 ;
        RECT 1336.850 1766.840 1337.130 1767.120 ;
        RECT 1337.310 1745.080 1337.590 1745.360 ;
        RECT 1339.150 2018.440 1339.430 2018.720 ;
        RECT 1339.610 1976.280 1339.890 1976.560 ;
        RECT 1340.070 1955.880 1340.350 1956.160 ;
        RECT 1340.530 1934.120 1340.810 1934.400 ;
        RECT 1340.990 1913.720 1341.270 1914.000 ;
        RECT 1341.450 1891.960 1341.730 1892.240 ;
        RECT 1341.910 1871.560 1342.190 1871.840 ;
        RECT 1342.370 1849.800 1342.650 1850.080 ;
        RECT 1342.830 1829.400 1343.110 1829.680 ;
        RECT 1343.290 1807.640 1343.570 1807.920 ;
        RECT 1345.130 1724.680 1345.410 1724.960 ;
        RECT 1372.730 2912.640 1373.010 2912.920 ;
        RECT 1441.730 2463.160 1442.010 2463.440 ;
        RECT 1442.650 2463.160 1442.930 2463.440 ;
        RECT 1439.430 2090.520 1439.710 2090.800 ;
        RECT 1440.350 2090.520 1440.630 2090.800 ;
        RECT 1439.890 2042.240 1440.170 2042.520 ;
        RECT 1441.730 2042.240 1442.010 2042.520 ;
        RECT 1441.730 1945.680 1442.010 1945.960 ;
        RECT 1442.650 1945.680 1442.930 1945.960 ;
        RECT 1441.730 1849.120 1442.010 1849.400 ;
        RECT 1442.650 1849.120 1442.930 1849.400 ;
        RECT 1441.730 1662.800 1442.010 1663.080 ;
        RECT 1443.110 1662.800 1443.390 1663.080 ;
        RECT 1441.730 1338.440 1442.010 1338.720 ;
        RECT 1442.650 1338.440 1442.930 1338.720 ;
        RECT 1441.730 1290.160 1442.010 1290.440 ;
        RECT 1442.650 1290.160 1442.930 1290.440 ;
        RECT 1441.730 1158.920 1442.010 1159.200 ;
        RECT 1442.650 1158.920 1442.930 1159.200 ;
        RECT 1483.590 2850.080 1483.870 2850.360 ;
        RECT 1482.210 2830.360 1482.490 2830.640 ;
        RECT 1490.030 2801.800 1490.310 2802.080 ;
        RECT 1485.430 2784.120 1485.710 2784.400 ;
        RECT 1489.570 2767.800 1489.850 2768.080 ;
        RECT 1489.110 2720.880 1489.390 2721.160 ;
        RECT 1488.650 2691.640 1488.930 2691.920 ;
        RECT 1482.670 2657.640 1482.950 2657.920 ;
        RECT 1485.430 2610.720 1485.710 2611.000 ;
        RECT 1488.650 2595.760 1488.930 2596.040 ;
        RECT 1488.650 2580.800 1488.930 2581.080 ;
        RECT 1488.650 2567.200 1488.930 2567.480 ;
        RECT 1483.590 2547.480 1483.870 2547.760 ;
        RECT 1496.470 2753.520 1496.750 2753.800 ;
        RECT 1496.010 2739.240 1496.290 2739.520 ;
        RECT 1495.550 2629.080 1495.830 2629.360 ;
        RECT 1843.310 2912.640 1843.590 2912.920 ;
        RECT 1500.610 2884.080 1500.890 2884.360 ;
        RECT 1501.990 2884.080 1502.270 2884.360 ;
        RECT 1497.850 2677.020 1498.130 2677.300 ;
        RECT 1501.990 2559.720 1502.270 2560.000 ;
        RECT 1500.150 2559.040 1500.430 2559.320 ;
        RECT 1498.310 2519.260 1498.590 2519.540 ;
        RECT 1520.850 2463.160 1521.130 2463.440 ;
        RECT 1519.930 2366.600 1520.210 2366.880 ;
        RECT 1520.850 2366.600 1521.130 2366.880 ;
        RECT 1522.690 1256.840 1522.970 1257.120 ;
        RECT 1521.770 1255.480 1522.050 1255.760 ;
        RECT 1520.390 1055.560 1520.670 1055.840 ;
        RECT 1521.310 1055.560 1521.590 1055.840 ;
        RECT 1530.050 2463.160 1530.330 2463.440 ;
        RECT 1886.550 2829.000 1886.830 2829.280 ;
        RECT 1887.010 2815.400 1887.290 2815.680 ;
        RECT 1890.690 2800.780 1890.970 2801.060 ;
        RECT 1887.470 2782.760 1887.750 2783.040 ;
        RECT 1891.150 2753.180 1891.430 2753.460 ;
        RECT 1891.610 2738.220 1891.890 2738.500 ;
        RECT 1897.590 2845.320 1897.870 2845.600 ;
        RECT 1894.830 2577.400 1895.110 2577.680 ;
        RECT 1898.050 2767.120 1898.330 2767.400 ;
        RECT 1898.510 2718.840 1898.790 2719.120 ;
        RECT 1898.970 2687.560 1899.250 2687.840 ;
        RECT 1899.430 2672.600 1899.710 2672.880 ;
        RECT 1899.890 2656.960 1900.170 2657.240 ;
        RECT 1900.350 2625.000 1900.630 2625.280 ;
        RECT 1900.810 2608.680 1901.090 2608.960 ;
        RECT 1901.270 2562.440 1901.550 2562.720 ;
        RECT 1901.730 2546.800 1902.010 2547.080 ;
        RECT 1903.570 2514.840 1903.850 2515.120 ;
        RECT 1904.490 1885.840 1904.770 1886.120 ;
        RECT 1904.490 1870.200 1904.770 1870.480 ;
        RECT 1904.490 1851.840 1904.770 1852.120 ;
        RECT 1904.490 1817.840 1904.770 1818.120 ;
        RECT 1904.490 1767.520 1904.770 1767.800 ;
        RECT 2076.990 1819.540 2077.270 1819.820 ;
        RECT 2083.890 1884.480 2084.170 1884.760 ;
        RECT 2084.350 1850.480 2084.630 1850.760 ;
        RECT 2084.810 1835.520 2085.090 1835.800 ;
        RECT 2085.270 1800.840 2085.550 1801.120 ;
        RECT 2085.730 1782.480 2086.010 1782.760 ;
        RECT 2086.190 1766.840 2086.470 1767.120 ;
        RECT 2283.990 1875.640 2284.270 1875.920 ;
        RECT 2287.210 1789.960 2287.490 1790.240 ;
        RECT 2523.650 1891.960 2523.930 1892.240 ;
        RECT 2523.650 1802.200 2523.930 1802.480 ;
        RECT 2518.590 1704.280 2518.870 1704.560 ;
        RECT 2523.650 1717.880 2523.930 1718.160 ;
        RECT 2519.510 1704.280 2519.790 1704.560 ;
        RECT 2519.510 1608.400 2519.790 1608.680 ;
        RECT 2519.510 1607.040 2519.790 1607.320 ;
      LAYER met3 ;
        RECT 1372.705 2912.930 1373.035 2912.945 ;
        RECT 1843.285 2912.930 1843.615 2912.945 ;
        RECT 1372.705 2912.630 1843.615 2912.930 ;
        RECT 1372.705 2912.615 1373.035 2912.630 ;
        RECT 1843.285 2912.615 1843.615 2912.630 ;
        RECT 1500.585 2884.370 1500.915 2884.385 ;
        RECT 1501.965 2884.370 1502.295 2884.385 ;
        RECT 1500.585 2884.070 1502.295 2884.370 ;
        RECT 1500.585 2884.055 1500.915 2884.070 ;
        RECT 1501.965 2884.055 1502.295 2884.070 ;
      LAYER met3 ;
        RECT 1504.000 2881.840 1885.335 2889.125 ;
        RECT 1504.400 2880.480 1885.335 2881.840 ;
        RECT 1504.400 2880.440 1884.935 2880.480 ;
        RECT 1504.000 2879.080 1884.935 2880.440 ;
        RECT 1504.000 2865.520 1885.335 2879.080 ;
        RECT 1504.400 2864.160 1885.335 2865.520 ;
        RECT 1504.400 2864.120 1884.935 2864.160 ;
        RECT 1504.000 2862.760 1884.935 2864.120 ;
        RECT 1504.000 2850.560 1885.335 2862.760 ;
      LAYER met3 ;
        RECT 1483.565 2850.370 1483.895 2850.385 ;
        RECT 1483.565 2850.160 1500.210 2850.370 ;
        RECT 1483.565 2850.070 1504.000 2850.160 ;
        RECT 1483.565 2850.055 1483.895 2850.070 ;
        RECT 1499.910 2849.880 1504.000 2850.070 ;
        RECT 1500.000 2849.560 1504.000 2849.880 ;
      LAYER met3 ;
        RECT 1504.400 2849.200 1885.335 2850.560 ;
        RECT 1504.400 2849.160 1884.935 2849.200 ;
        RECT 1504.000 2847.800 1884.935 2849.160 ;
      LAYER met3 ;
        RECT 1885.335 2848.520 1889.335 2848.800 ;
        RECT 1885.335 2848.200 1889.370 2848.520 ;
      LAYER met3 ;
        RECT 1504.000 2834.240 1885.335 2847.800 ;
      LAYER met3 ;
        RECT 1889.070 2845.610 1889.370 2848.200 ;
        RECT 1897.565 2845.610 1897.895 2845.625 ;
        RECT 1889.070 2845.310 1897.895 2845.610 ;
        RECT 1897.565 2845.295 1897.895 2845.310 ;
        RECT 1500.000 2833.560 1504.000 2833.840 ;
        RECT 1499.910 2833.240 1504.000 2833.560 ;
        RECT 1482.185 2830.650 1482.515 2830.665 ;
        RECT 1499.910 2830.650 1500.210 2833.240 ;
      LAYER met3 ;
        RECT 1504.400 2832.880 1885.335 2834.240 ;
        RECT 1504.400 2832.840 1884.935 2832.880 ;
      LAYER met3 ;
        RECT 1482.185 2830.350 1500.210 2830.650 ;
      LAYER met3 ;
        RECT 1504.000 2831.480 1884.935 2832.840 ;
      LAYER met3 ;
        RECT 1885.335 2831.880 1889.335 2832.480 ;
        RECT 1482.185 2830.335 1482.515 2830.350 ;
      LAYER met3 ;
        RECT 1504.000 2819.280 1885.335 2831.480 ;
      LAYER met3 ;
        RECT 1886.310 2829.305 1886.610 2831.880 ;
        RECT 1886.310 2828.990 1886.855 2829.305 ;
        RECT 1886.525 2828.975 1886.855 2828.990 ;
      LAYER met3 ;
        RECT 1504.400 2817.920 1885.335 2819.280 ;
        RECT 1504.400 2817.880 1884.935 2817.920 ;
        RECT 1504.000 2816.520 1884.935 2817.880 ;
      LAYER met3 ;
        RECT 1885.335 2816.920 1889.335 2817.520 ;
        RECT 998.470 2808.890 998.850 2808.900 ;
        RECT 1058.065 2808.890 1058.395 2808.905 ;
        RECT 998.470 2808.590 1058.395 2808.890 ;
        RECT 998.470 2808.580 998.850 2808.590 ;
        RECT 1058.065 2808.575 1058.395 2808.590 ;
      LAYER met3 ;
        RECT 1504.000 2802.960 1885.335 2816.520 ;
      LAYER met3 ;
        RECT 1887.230 2815.705 1887.530 2816.920 ;
        RECT 1886.985 2815.390 1887.530 2815.705 ;
        RECT 1886.985 2815.375 1887.315 2815.390 ;
        RECT 1500.000 2802.280 1504.000 2802.560 ;
        RECT 1490.005 2802.090 1490.335 2802.105 ;
        RECT 1499.910 2802.090 1504.000 2802.280 ;
        RECT 1490.005 2801.960 1504.000 2802.090 ;
        RECT 1490.005 2801.790 1500.210 2801.960 ;
        RECT 1490.005 2801.775 1490.335 2801.790 ;
      LAYER met3 ;
        RECT 1504.400 2801.600 1885.335 2802.960 ;
        RECT 1504.400 2801.560 1884.935 2801.600 ;
        RECT 1504.000 2800.200 1884.935 2801.560 ;
      LAYER met3 ;
        RECT 1885.335 2801.070 1889.335 2801.200 ;
        RECT 1890.665 2801.070 1890.995 2801.085 ;
        RECT 1885.335 2800.770 1890.995 2801.070 ;
        RECT 1885.335 2800.600 1889.335 2800.770 ;
        RECT 1890.665 2800.755 1890.995 2800.770 ;
      LAYER met3 ;
        RECT 1504.000 2788.000 1885.335 2800.200 ;
        RECT 1004.000 2787.360 1096.000 2787.845 ;
      LAYER met3 ;
        RECT 1000.000 2786.360 1004.000 2786.960 ;
        RECT 992.950 2783.730 993.330 2783.740 ;
        RECT 1000.350 2783.730 1000.650 2786.360 ;
      LAYER met3 ;
        RECT 1004.400 2785.960 1096.000 2787.360 ;
      LAYER met3 ;
        RECT 1500.000 2787.320 1504.000 2787.600 ;
        RECT 992.950 2783.430 1000.650 2783.730 ;
      LAYER met3 ;
        RECT 1004.000 2784.640 1096.000 2785.960 ;
      LAYER met3 ;
        RECT 1499.910 2787.000 1504.000 2787.320 ;
        RECT 992.950 2783.420 993.330 2783.430 ;
      LAYER met3 ;
        RECT 1004.000 2783.240 1095.600 2784.640 ;
      LAYER met3 ;
        RECT 1485.405 2784.410 1485.735 2784.425 ;
        RECT 1499.910 2784.410 1500.210 2787.000 ;
      LAYER met3 ;
        RECT 1504.400 2786.640 1885.335 2788.000 ;
        RECT 1504.400 2786.600 1884.935 2786.640 ;
      LAYER met3 ;
        RECT 1096.000 2783.920 1100.000 2784.240 ;
        RECT 1485.405 2784.110 1500.210 2784.410 ;
      LAYER met3 ;
        RECT 1504.000 2785.240 1884.935 2786.600 ;
      LAYER met3 ;
        RECT 1885.335 2785.640 1889.335 2786.240 ;
        RECT 1485.405 2784.095 1485.735 2784.110 ;
        RECT 1096.000 2783.640 1100.010 2783.920 ;
      LAYER met3 ;
        RECT 1004.000 2764.240 1096.000 2783.240 ;
      LAYER met3 ;
        RECT 1099.710 2781.010 1100.010 2783.640 ;
        RECT 1110.965 2781.010 1111.295 2781.025 ;
        RECT 1099.710 2780.710 1111.295 2781.010 ;
        RECT 1110.965 2780.695 1111.295 2780.710 ;
      LAYER met3 ;
        RECT 1504.000 2771.680 1885.335 2785.240 ;
      LAYER met3 ;
        RECT 1887.230 2783.065 1887.530 2785.640 ;
        RECT 1887.230 2782.750 1887.775 2783.065 ;
        RECT 1887.445 2782.735 1887.775 2782.750 ;
        RECT 1500.000 2771.000 1504.000 2771.280 ;
        RECT 1499.910 2770.680 1504.000 2771.000 ;
        RECT 1489.545 2768.090 1489.875 2768.105 ;
        RECT 1499.910 2768.090 1500.210 2770.680 ;
      LAYER met3 ;
        RECT 1504.400 2770.320 1885.335 2771.680 ;
        RECT 1504.400 2770.280 1884.935 2770.320 ;
      LAYER met3 ;
        RECT 1489.545 2767.790 1500.210 2768.090 ;
      LAYER met3 ;
        RECT 1504.000 2768.920 1884.935 2770.280 ;
      LAYER met3 ;
        RECT 1885.335 2769.640 1889.335 2769.920 ;
        RECT 1885.335 2769.320 1889.370 2769.640 ;
        RECT 1489.545 2767.775 1489.875 2767.790 ;
        RECT 1000.000 2763.240 1004.000 2763.840 ;
        RECT 992.030 2760.610 992.410 2760.620 ;
        RECT 1000.350 2760.610 1000.650 2763.240 ;
      LAYER met3 ;
        RECT 1004.400 2762.840 1096.000 2764.240 ;
      LAYER met3 ;
        RECT 992.030 2760.310 1000.650 2760.610 ;
      LAYER met3 ;
        RECT 1004.000 2761.520 1096.000 2762.840 ;
      LAYER met3 ;
        RECT 992.030 2760.300 992.410 2760.310 ;
      LAYER met3 ;
        RECT 1004.000 2760.120 1095.600 2761.520 ;
      LAYER met3 ;
        RECT 1096.000 2760.800 1100.000 2761.120 ;
        RECT 1096.000 2760.610 1100.010 2760.800 ;
        RECT 1111.425 2760.610 1111.755 2760.625 ;
        RECT 1096.000 2760.520 1111.755 2760.610 ;
        RECT 1099.710 2760.310 1111.755 2760.520 ;
        RECT 1111.425 2760.295 1111.755 2760.310 ;
      LAYER met3 ;
        RECT 434.400 2751.960 574.800 2752.825 ;
        RECT 434.000 2734.320 574.800 2751.960 ;
        RECT 1004.000 2741.120 1096.000 2760.120 ;
        RECT 1504.000 2755.360 1885.335 2768.920 ;
      LAYER met3 ;
        RECT 1889.070 2767.410 1889.370 2769.320 ;
        RECT 1898.025 2767.410 1898.355 2767.425 ;
        RECT 1889.070 2767.110 1898.355 2767.410 ;
        RECT 1898.025 2767.095 1898.355 2767.110 ;
        RECT 1500.000 2754.680 1504.000 2754.960 ;
        RECT 1499.910 2754.360 1504.000 2754.680 ;
        RECT 1496.445 2753.810 1496.775 2753.825 ;
        RECT 1499.910 2753.810 1500.210 2754.360 ;
      LAYER met3 ;
        RECT 1504.400 2754.000 1885.335 2755.360 ;
        RECT 1504.400 2753.960 1884.935 2754.000 ;
      LAYER met3 ;
        RECT 1496.445 2753.510 1500.210 2753.810 ;
        RECT 1496.445 2753.495 1496.775 2753.510 ;
        RECT 1000.000 2740.120 1004.000 2740.720 ;
        RECT 991.110 2739.530 991.490 2739.540 ;
        RECT 1000.350 2739.530 1000.650 2740.120 ;
      LAYER met3 ;
        RECT 1004.400 2739.720 1096.000 2741.120 ;
        RECT 1504.000 2752.600 1884.935 2753.960 ;
      LAYER met3 ;
        RECT 1885.335 2753.470 1889.335 2753.600 ;
        RECT 1891.125 2753.470 1891.455 2753.485 ;
        RECT 1885.335 2753.170 1891.455 2753.470 ;
        RECT 1885.335 2753.000 1889.335 2753.170 ;
        RECT 1891.125 2753.155 1891.455 2753.170 ;
      LAYER met3 ;
        RECT 1504.000 2740.400 1885.335 2752.600 ;
      LAYER met3 ;
        RECT 1500.000 2739.720 1504.000 2740.000 ;
        RECT 991.110 2739.230 1000.650 2739.530 ;
        RECT 991.110 2739.220 991.490 2739.230 ;
      LAYER met3 ;
        RECT 1004.000 2738.400 1096.000 2739.720 ;
      LAYER met3 ;
        RECT 1495.985 2739.530 1496.315 2739.545 ;
        RECT 1499.910 2739.530 1504.000 2739.720 ;
        RECT 1495.985 2739.400 1504.000 2739.530 ;
        RECT 1495.985 2739.230 1500.210 2739.400 ;
        RECT 1495.985 2739.215 1496.315 2739.230 ;
      LAYER met3 ;
        RECT 1504.400 2739.040 1885.335 2740.400 ;
        RECT 1504.400 2739.000 1884.935 2739.040 ;
        RECT 1004.000 2737.000 1095.600 2738.400 ;
      LAYER met3 ;
        RECT 1096.000 2737.680 1100.000 2738.000 ;
        RECT 1096.000 2737.400 1100.010 2737.680 ;
      LAYER met3 ;
        RECT 434.000 2732.960 574.400 2734.320 ;
        RECT 434.400 2732.920 574.400 2732.960 ;
      LAYER met3 ;
        RECT 430.000 2732.240 434.000 2732.560 ;
        RECT 429.950 2731.960 434.000 2732.240 ;
        RECT 420.505 2729.330 420.835 2729.345 ;
        RECT 429.950 2729.330 430.250 2731.960 ;
      LAYER met3 ;
        RECT 434.400 2731.560 574.800 2732.920 ;
      LAYER met3 ;
        RECT 420.505 2729.030 430.250 2729.330 ;
        RECT 420.505 2729.015 420.835 2729.030 ;
      LAYER met3 ;
        RECT 434.000 2712.560 574.800 2731.560 ;
        RECT 1004.000 2719.360 1096.000 2737.000 ;
      LAYER met3 ;
        RECT 1099.710 2734.770 1100.010 2737.400 ;
      LAYER met3 ;
        RECT 1504.000 2737.640 1884.935 2739.000 ;
      LAYER met3 ;
        RECT 1885.335 2738.510 1889.335 2738.640 ;
        RECT 1891.585 2738.510 1891.915 2738.525 ;
        RECT 1885.335 2738.210 1891.915 2738.510 ;
        RECT 1885.335 2738.040 1889.335 2738.210 ;
        RECT 1891.585 2738.195 1891.915 2738.210 ;
        RECT 1112.805 2734.770 1113.135 2734.785 ;
        RECT 1099.710 2734.470 1113.135 2734.770 ;
        RECT 1112.805 2734.455 1113.135 2734.470 ;
      LAYER met3 ;
        RECT 1504.000 2724.080 1885.335 2737.640 ;
      LAYER met3 ;
        RECT 1500.000 2723.400 1504.000 2723.680 ;
        RECT 1499.910 2723.080 1504.000 2723.400 ;
        RECT 1489.085 2721.170 1489.415 2721.185 ;
        RECT 1499.910 2721.170 1500.210 2723.080 ;
      LAYER met3 ;
        RECT 1504.400 2722.720 1885.335 2724.080 ;
        RECT 1504.400 2722.680 1884.935 2722.720 ;
      LAYER met3 ;
        RECT 1489.085 2720.870 1500.210 2721.170 ;
      LAYER met3 ;
        RECT 1504.000 2721.320 1884.935 2722.680 ;
      LAYER met3 ;
        RECT 1885.335 2722.040 1889.335 2722.320 ;
        RECT 1885.335 2721.720 1889.370 2722.040 ;
        RECT 1489.085 2720.855 1489.415 2720.870 ;
        RECT 990.190 2719.130 990.570 2719.140 ;
        RECT 990.190 2718.960 1000.650 2719.130 ;
        RECT 990.190 2718.830 1004.000 2718.960 ;
        RECT 990.190 2718.820 990.570 2718.830 ;
        RECT 1000.000 2718.360 1004.000 2718.830 ;
      LAYER met3 ;
        RECT 1004.400 2717.960 1096.000 2719.360 ;
        RECT 1004.000 2716.640 1096.000 2717.960 ;
        RECT 1004.000 2715.240 1095.600 2716.640 ;
      LAYER met3 ;
        RECT 1096.000 2715.920 1100.000 2716.240 ;
        RECT 1096.000 2715.640 1100.010 2715.920 ;
      LAYER met3 ;
        RECT 434.000 2711.200 574.400 2712.560 ;
        RECT 434.400 2711.160 574.400 2711.200 ;
      LAYER met3 ;
        RECT 430.000 2710.480 434.000 2710.800 ;
        RECT 429.950 2710.200 434.000 2710.480 ;
        RECT 420.045 2707.570 420.375 2707.585 ;
        RECT 429.950 2707.570 430.250 2710.200 ;
      LAYER met3 ;
        RECT 434.400 2709.800 574.800 2711.160 ;
      LAYER met3 ;
        RECT 420.045 2707.270 430.250 2707.570 ;
        RECT 420.045 2707.255 420.375 2707.270 ;
      LAYER met3 ;
        RECT 434.000 2690.800 574.800 2709.800 ;
        RECT 1004.000 2696.240 1096.000 2715.240 ;
      LAYER met3 ;
        RECT 1099.710 2713.010 1100.010 2715.640 ;
        RECT 1112.345 2713.010 1112.675 2713.025 ;
        RECT 1099.710 2712.710 1112.675 2713.010 ;
        RECT 1112.345 2712.695 1112.675 2712.710 ;
      LAYER met3 ;
        RECT 1504.000 2709.120 1885.335 2721.320 ;
      LAYER met3 ;
        RECT 1889.070 2719.130 1889.370 2721.720 ;
        RECT 1898.485 2719.130 1898.815 2719.145 ;
        RECT 1889.070 2718.830 1898.815 2719.130 ;
        RECT 1898.485 2718.815 1898.815 2718.830 ;
      LAYER met3 ;
        RECT 1504.400 2707.760 1885.335 2709.120 ;
        RECT 1504.400 2707.720 1884.935 2707.760 ;
      LAYER met3 ;
        RECT 1000.000 2695.240 1004.000 2695.840 ;
        RECT 989.270 2692.610 989.650 2692.620 ;
        RECT 1000.350 2692.610 1000.650 2695.240 ;
      LAYER met3 ;
        RECT 1004.400 2694.840 1096.000 2696.240 ;
      LAYER met3 ;
        RECT 989.270 2692.310 1000.650 2692.610 ;
      LAYER met3 ;
        RECT 1004.000 2693.520 1096.000 2694.840 ;
        RECT 1504.000 2706.360 1884.935 2707.720 ;
      LAYER met3 ;
        RECT 989.270 2692.300 989.650 2692.310 ;
      LAYER met3 ;
        RECT 1004.000 2692.120 1095.600 2693.520 ;
      LAYER met3 ;
        RECT 1096.000 2692.800 1100.000 2693.120 ;
      LAYER met3 ;
        RECT 1504.000 2692.800 1885.335 2706.360 ;
      LAYER met3 ;
        RECT 1096.000 2692.520 1100.010 2692.800 ;
      LAYER met3 ;
        RECT 434.000 2689.440 574.400 2690.800 ;
      LAYER met3 ;
        RECT 574.800 2689.800 578.800 2690.400 ;
      LAYER met3 ;
        RECT 434.400 2689.400 574.400 2689.440 ;
        RECT 434.400 2688.040 574.800 2689.400 ;
        RECT 434.000 2670.400 574.800 2688.040 ;
      LAYER met3 ;
        RECT 578.070 2687.170 578.370 2689.800 ;
        RECT 586.565 2687.170 586.895 2687.185 ;
        RECT 578.070 2686.870 586.895 2687.170 ;
        RECT 586.565 2686.855 586.895 2686.870 ;
      LAYER met3 ;
        RECT 1004.000 2673.120 1096.000 2692.120 ;
      LAYER met3 ;
        RECT 1099.710 2691.930 1100.010 2692.520 ;
        RECT 1500.000 2692.120 1504.000 2692.400 ;
        RECT 1111.885 2691.930 1112.215 2691.945 ;
        RECT 1099.710 2691.630 1112.215 2691.930 ;
        RECT 1111.885 2691.615 1112.215 2691.630 ;
        RECT 1488.625 2691.930 1488.955 2691.945 ;
        RECT 1499.910 2691.930 1504.000 2692.120 ;
        RECT 1488.625 2691.800 1504.000 2691.930 ;
        RECT 1488.625 2691.630 1500.210 2691.800 ;
        RECT 1488.625 2691.615 1488.955 2691.630 ;
      LAYER met3 ;
        RECT 1504.400 2691.440 1885.335 2692.800 ;
        RECT 1504.400 2691.400 1884.935 2691.440 ;
        RECT 1504.000 2690.040 1884.935 2691.400 ;
      LAYER met3 ;
        RECT 1885.335 2690.760 1889.335 2691.040 ;
        RECT 1885.335 2690.440 1889.370 2690.760 ;
      LAYER met3 ;
        RECT 1504.000 2677.840 1885.335 2690.040 ;
      LAYER met3 ;
        RECT 1889.070 2687.850 1889.370 2690.440 ;
        RECT 1898.945 2687.850 1899.275 2687.865 ;
        RECT 1889.070 2687.550 1899.275 2687.850 ;
        RECT 1898.945 2687.535 1899.275 2687.550 ;
        RECT 1497.825 2677.310 1498.155 2677.325 ;
        RECT 1500.000 2677.310 1504.000 2677.440 ;
        RECT 1497.825 2677.010 1504.000 2677.310 ;
        RECT 1497.825 2676.995 1498.155 2677.010 ;
        RECT 1500.000 2676.840 1504.000 2677.010 ;
      LAYER met3 ;
        RECT 1504.400 2676.480 1885.335 2677.840 ;
        RECT 1504.400 2676.440 1884.935 2676.480 ;
      LAYER met3 ;
        RECT 1000.000 2672.120 1004.000 2672.720 ;
        RECT 993.205 2670.850 993.535 2670.865 ;
        RECT 1000.350 2670.850 1000.650 2672.120 ;
      LAYER met3 ;
        RECT 1004.400 2671.720 1096.000 2673.120 ;
      LAYER met3 ;
        RECT 993.205 2670.550 1000.650 2670.850 ;
        RECT 993.205 2670.535 993.535 2670.550 ;
      LAYER met3 ;
        RECT 1004.000 2670.400 1096.000 2671.720 ;
        RECT 1504.000 2675.080 1884.935 2676.440 ;
      LAYER met3 ;
        RECT 1885.335 2675.800 1889.335 2676.080 ;
        RECT 1885.335 2675.480 1889.370 2675.800 ;
      LAYER met3 ;
        RECT 434.000 2669.040 574.400 2670.400 ;
      LAYER met3 ;
        RECT 574.800 2669.400 578.800 2670.000 ;
      LAYER met3 ;
        RECT 434.400 2669.000 574.400 2669.040 ;
        RECT 434.400 2667.640 574.800 2669.000 ;
        RECT 434.000 2648.640 574.800 2667.640 ;
      LAYER met3 ;
        RECT 578.070 2666.770 578.370 2669.400 ;
      LAYER met3 ;
        RECT 1004.000 2669.000 1095.600 2670.400 ;
      LAYER met3 ;
        RECT 1096.000 2669.680 1100.000 2670.000 ;
        RECT 1096.000 2669.400 1100.010 2669.680 ;
        RECT 586.565 2666.770 586.895 2666.785 ;
        RECT 578.070 2666.470 586.895 2666.770 ;
        RECT 586.565 2666.455 586.895 2666.470 ;
      LAYER met3 ;
        RECT 1004.000 2650.000 1096.000 2669.000 ;
      LAYER met3 ;
        RECT 1099.710 2666.770 1100.010 2669.400 ;
        RECT 1113.265 2666.770 1113.595 2666.785 ;
        RECT 1099.710 2666.470 1113.595 2666.770 ;
        RECT 1113.265 2666.455 1113.595 2666.470 ;
      LAYER met3 ;
        RECT 1504.000 2661.520 1885.335 2675.080 ;
      LAYER met3 ;
        RECT 1889.070 2672.890 1889.370 2675.480 ;
        RECT 1899.405 2672.890 1899.735 2672.905 ;
        RECT 1889.070 2672.590 1899.735 2672.890 ;
        RECT 1899.405 2672.575 1899.735 2672.590 ;
        RECT 1500.000 2660.840 1504.000 2661.120 ;
        RECT 1499.910 2660.520 1504.000 2660.840 ;
        RECT 1482.645 2657.930 1482.975 2657.945 ;
        RECT 1499.910 2657.930 1500.210 2660.520 ;
      LAYER met3 ;
        RECT 1504.400 2660.160 1885.335 2661.520 ;
        RECT 1504.400 2660.120 1884.935 2660.160 ;
      LAYER met3 ;
        RECT 1482.645 2657.630 1500.210 2657.930 ;
      LAYER met3 ;
        RECT 1504.000 2658.760 1884.935 2660.120 ;
      LAYER met3 ;
        RECT 1885.335 2659.480 1889.335 2659.760 ;
        RECT 1885.335 2659.160 1889.370 2659.480 ;
        RECT 1482.645 2657.615 1482.975 2657.630 ;
        RECT 1000.000 2649.000 1004.000 2649.600 ;
      LAYER met3 ;
        RECT 434.000 2647.280 574.400 2648.640 ;
        RECT 434.400 2647.240 574.400 2647.280 ;
        RECT 434.400 2645.880 574.800 2647.240 ;
      LAYER met3 ;
        RECT 993.665 2646.370 993.995 2646.385 ;
        RECT 1000.350 2646.370 1000.650 2649.000 ;
      LAYER met3 ;
        RECT 1004.400 2648.600 1096.000 2650.000 ;
      LAYER met3 ;
        RECT 993.665 2646.070 1000.650 2646.370 ;
      LAYER met3 ;
        RECT 1004.000 2647.280 1096.000 2648.600 ;
      LAYER met3 ;
        RECT 993.665 2646.055 993.995 2646.070 ;
      LAYER met3 ;
        RECT 434.000 2626.880 574.800 2645.880 ;
        RECT 1004.000 2645.880 1095.600 2647.280 ;
      LAYER met3 ;
        RECT 1096.000 2646.560 1100.000 2646.880 ;
      LAYER met3 ;
        RECT 1504.000 2646.560 1885.335 2658.760 ;
      LAYER met3 ;
        RECT 1889.070 2657.250 1889.370 2659.160 ;
        RECT 1899.865 2657.250 1900.195 2657.265 ;
        RECT 1889.070 2656.950 1900.195 2657.250 ;
        RECT 1899.865 2656.935 1900.195 2656.950 ;
        RECT 1096.000 2646.280 1100.010 2646.560 ;
      LAYER met3 ;
        RECT 1004.000 2626.880 1096.000 2645.880 ;
      LAYER met3 ;
        RECT 1099.710 2645.010 1100.010 2646.280 ;
      LAYER met3 ;
        RECT 1504.400 2645.200 1885.335 2646.560 ;
        RECT 1504.400 2645.160 1884.935 2645.200 ;
      LAYER met3 ;
        RECT 1113.725 2645.010 1114.055 2645.025 ;
        RECT 1099.710 2644.710 1114.055 2645.010 ;
        RECT 1113.725 2644.695 1114.055 2644.710 ;
      LAYER met3 ;
        RECT 1504.000 2643.800 1884.935 2645.160 ;
        RECT 1504.000 2630.240 1885.335 2643.800 ;
      LAYER met3 ;
        RECT 1500.000 2629.560 1504.000 2629.840 ;
        RECT 1495.525 2629.370 1495.855 2629.385 ;
        RECT 1499.910 2629.370 1504.000 2629.560 ;
        RECT 1495.525 2629.240 1504.000 2629.370 ;
        RECT 1495.525 2629.070 1500.210 2629.240 ;
        RECT 1495.525 2629.055 1495.855 2629.070 ;
      LAYER met3 ;
        RECT 1504.400 2628.880 1885.335 2630.240 ;
        RECT 1504.400 2628.840 1884.935 2628.880 ;
        RECT 434.000 2625.520 574.400 2626.880 ;
      LAYER met3 ;
        RECT 1000.000 2625.880 1004.000 2626.480 ;
      LAYER met3 ;
        RECT 434.400 2625.480 574.400 2625.520 ;
        RECT 434.400 2624.120 574.800 2625.480 ;
        RECT 434.000 2606.480 574.800 2624.120 ;
      LAYER met3 ;
        RECT 992.745 2623.250 993.075 2623.265 ;
        RECT 1000.350 2623.250 1000.650 2625.880 ;
      LAYER met3 ;
        RECT 1004.400 2625.480 1096.000 2626.880 ;
      LAYER met3 ;
        RECT 992.745 2622.950 1000.650 2623.250 ;
      LAYER met3 ;
        RECT 1004.000 2624.160 1096.000 2625.480 ;
        RECT 1504.000 2627.480 1884.935 2628.840 ;
      LAYER met3 ;
        RECT 1885.335 2628.200 1889.335 2628.480 ;
        RECT 1885.335 2627.880 1889.370 2628.200 ;
        RECT 992.745 2622.935 993.075 2622.950 ;
      LAYER met3 ;
        RECT 1004.000 2622.760 1095.600 2624.160 ;
      LAYER met3 ;
        RECT 1096.000 2623.440 1100.000 2623.760 ;
        RECT 1096.000 2623.160 1100.010 2623.440 ;
      LAYER met3 ;
        RECT 1004.000 2610.715 1096.000 2622.760 ;
      LAYER met3 ;
        RECT 1099.710 2622.570 1100.010 2623.160 ;
        RECT 1114.185 2622.570 1114.515 2622.585 ;
        RECT 1099.710 2622.270 1114.515 2622.570 ;
        RECT 1114.185 2622.255 1114.515 2622.270 ;
      LAYER met3 ;
        RECT 1504.000 2613.920 1885.335 2627.480 ;
      LAYER met3 ;
        RECT 1889.070 2625.290 1889.370 2627.880 ;
        RECT 1900.325 2625.290 1900.655 2625.305 ;
        RECT 1889.070 2624.990 1900.655 2625.290 ;
        RECT 1900.325 2624.975 1900.655 2624.990 ;
        RECT 1500.000 2613.240 1504.000 2613.520 ;
        RECT 1499.910 2612.920 1504.000 2613.240 ;
        RECT 1485.405 2611.010 1485.735 2611.025 ;
        RECT 1499.910 2611.010 1500.210 2612.920 ;
      LAYER met3 ;
        RECT 1504.400 2612.560 1885.335 2613.920 ;
        RECT 1504.400 2612.520 1884.935 2612.560 ;
      LAYER met3 ;
        RECT 1485.405 2610.710 1500.210 2611.010 ;
      LAYER met3 ;
        RECT 1504.000 2611.160 1884.935 2612.520 ;
      LAYER met3 ;
        RECT 1885.335 2611.880 1889.335 2612.160 ;
        RECT 1885.335 2611.560 1889.370 2611.880 ;
        RECT 1485.405 2610.695 1485.735 2610.710 ;
      LAYER met3 ;
        RECT 434.000 2605.615 574.400 2606.480 ;
        RECT 1504.000 2598.960 1885.335 2611.160 ;
      LAYER met3 ;
        RECT 1889.070 2608.970 1889.370 2611.560 ;
      LAYER met3 ;
        RECT 2427.190 2610.715 2529.990 2760.645 ;
      LAYER met3 ;
        RECT 1900.785 2608.970 1901.115 2608.985 ;
        RECT 1889.070 2608.670 1901.115 2608.970 ;
        RECT 1900.785 2608.655 1901.115 2608.670 ;
        RECT 1500.000 2598.280 1504.000 2598.560 ;
        RECT 1499.910 2597.960 1504.000 2598.280 ;
        RECT 1488.625 2596.050 1488.955 2596.065 ;
        RECT 1499.910 2596.050 1500.210 2597.960 ;
      LAYER met3 ;
        RECT 1504.400 2597.600 1885.335 2598.960 ;
        RECT 1504.400 2597.560 1884.935 2597.600 ;
      LAYER met3 ;
        RECT 1488.625 2595.750 1500.210 2596.050 ;
      LAYER met3 ;
        RECT 1504.000 2596.200 1884.935 2597.560 ;
      LAYER met3 ;
        RECT 1488.625 2595.735 1488.955 2595.750 ;
      LAYER met3 ;
        RECT 1504.000 2582.640 1885.335 2596.200 ;
      LAYER met3 ;
        RECT 1500.000 2581.960 1504.000 2582.240 ;
        RECT 1499.910 2581.640 1504.000 2581.960 ;
        RECT 1488.625 2581.090 1488.955 2581.105 ;
        RECT 1499.910 2581.090 1500.210 2581.640 ;
      LAYER met3 ;
        RECT 1504.400 2581.280 1885.335 2582.640 ;
        RECT 1504.400 2581.240 1884.935 2581.280 ;
      LAYER met3 ;
        RECT 1488.625 2580.790 1500.210 2581.090 ;
        RECT 1488.625 2580.775 1488.955 2580.790 ;
      LAYER met3 ;
        RECT 1504.000 2579.880 1884.935 2581.240 ;
      LAYER met3 ;
        RECT 1885.335 2580.600 1889.335 2580.880 ;
        RECT 1885.335 2580.280 1889.370 2580.600 ;
      LAYER met3 ;
        RECT 1504.000 2567.680 1885.335 2579.880 ;
      LAYER met3 ;
        RECT 1889.070 2577.690 1889.370 2580.280 ;
        RECT 1894.805 2577.690 1895.135 2577.705 ;
        RECT 1889.070 2577.390 1895.135 2577.690 ;
        RECT 1894.805 2577.375 1895.135 2577.390 ;
        RECT 1488.625 2567.490 1488.955 2567.505 ;
        RECT 1488.625 2567.280 1500.210 2567.490 ;
        RECT 1488.625 2567.190 1504.000 2567.280 ;
        RECT 1488.625 2567.175 1488.955 2567.190 ;
        RECT 1499.910 2567.000 1504.000 2567.190 ;
        RECT 1500.000 2566.680 1504.000 2567.000 ;
      LAYER met3 ;
        RECT 1504.400 2566.320 1885.335 2567.680 ;
        RECT 1504.400 2566.280 1884.935 2566.320 ;
        RECT 1504.000 2564.920 1884.935 2566.280 ;
      LAYER met3 ;
        RECT 1885.335 2565.640 1889.335 2565.920 ;
        RECT 1885.335 2565.320 1889.370 2565.640 ;
        RECT 1501.965 2560.010 1502.295 2560.025 ;
        RECT 1501.965 2559.710 1502.970 2560.010 ;
        RECT 1501.965 2559.695 1502.295 2559.710 ;
        RECT 1500.125 2559.330 1500.455 2559.345 ;
        RECT 1502.670 2559.330 1502.970 2559.710 ;
        RECT 1500.125 2559.030 1502.970 2559.330 ;
        RECT 1500.125 2559.015 1500.455 2559.030 ;
      LAYER met3 ;
        RECT 1504.000 2551.360 1885.335 2564.920 ;
      LAYER met3 ;
        RECT 1889.070 2562.730 1889.370 2565.320 ;
        RECT 1901.245 2562.730 1901.575 2562.745 ;
        RECT 1889.070 2562.430 1901.575 2562.730 ;
        RECT 1901.245 2562.415 1901.575 2562.430 ;
        RECT 1500.000 2550.680 1504.000 2550.960 ;
        RECT 1499.910 2550.360 1504.000 2550.680 ;
        RECT 1483.565 2547.770 1483.895 2547.785 ;
        RECT 1499.910 2547.770 1500.210 2550.360 ;
      LAYER met3 ;
        RECT 1504.400 2550.000 1885.335 2551.360 ;
        RECT 1504.400 2549.960 1884.935 2550.000 ;
      LAYER met3 ;
        RECT 1483.565 2547.470 1500.210 2547.770 ;
      LAYER met3 ;
        RECT 1504.000 2548.600 1884.935 2549.960 ;
      LAYER met3 ;
        RECT 1885.335 2549.320 1889.335 2549.600 ;
        RECT 1885.335 2549.000 1889.370 2549.320 ;
        RECT 1483.565 2547.455 1483.895 2547.470 ;
      LAYER met3 ;
        RECT 1504.000 2536.400 1885.335 2548.600 ;
      LAYER met3 ;
        RECT 1889.070 2547.090 1889.370 2549.000 ;
        RECT 1901.705 2547.090 1902.035 2547.105 ;
        RECT 1889.070 2546.790 1902.035 2547.090 ;
        RECT 1901.705 2546.775 1902.035 2546.790 ;
      LAYER met3 ;
        RECT 1504.400 2535.040 1885.335 2536.400 ;
        RECT 1504.400 2535.000 1884.935 2535.040 ;
        RECT 1504.000 2533.640 1884.935 2535.000 ;
        RECT 1504.000 2520.080 1885.335 2533.640 ;
      LAYER met3 ;
        RECT 1498.285 2519.550 1498.615 2519.565 ;
        RECT 1500.000 2519.550 1504.000 2519.680 ;
        RECT 1498.285 2519.250 1504.000 2519.550 ;
        RECT 1498.285 2519.235 1498.615 2519.250 ;
        RECT 1500.000 2519.080 1504.000 2519.250 ;
      LAYER met3 ;
        RECT 1504.400 2518.720 1885.335 2520.080 ;
        RECT 1504.400 2518.680 1884.935 2518.720 ;
        RECT 1504.000 2517.320 1884.935 2518.680 ;
      LAYER met3 ;
        RECT 1885.335 2518.040 1889.335 2518.320 ;
        RECT 1885.335 2517.720 1889.370 2518.040 ;
      LAYER met3 ;
        RECT 1504.000 2504.255 1885.335 2517.320 ;
      LAYER met3 ;
        RECT 1889.070 2515.130 1889.370 2517.720 ;
        RECT 1903.545 2515.130 1903.875 2515.145 ;
        RECT 1889.070 2514.830 1903.875 2515.130 ;
        RECT 1903.545 2514.815 1903.875 2514.830 ;
        RECT 1441.705 2463.450 1442.035 2463.465 ;
        RECT 1442.625 2463.450 1442.955 2463.465 ;
        RECT 1441.705 2463.150 1442.955 2463.450 ;
        RECT 1441.705 2463.135 1442.035 2463.150 ;
        RECT 1442.625 2463.135 1442.955 2463.150 ;
        RECT 1520.825 2463.450 1521.155 2463.465 ;
        RECT 1530.025 2463.450 1530.355 2463.465 ;
        RECT 1520.825 2463.150 1530.355 2463.450 ;
        RECT 1520.825 2463.135 1521.155 2463.150 ;
        RECT 1530.025 2463.135 1530.355 2463.150 ;
        RECT 1519.905 2366.890 1520.235 2366.905 ;
        RECT 1520.825 2366.890 1521.155 2366.905 ;
        RECT 1519.905 2366.590 1521.155 2366.890 ;
        RECT 1519.905 2366.575 1520.235 2366.590 ;
        RECT 1520.825 2366.575 1521.155 2366.590 ;
        RECT 1439.405 2090.810 1439.735 2090.825 ;
        RECT 1440.325 2090.810 1440.655 2090.825 ;
        RECT 1439.405 2090.510 1440.655 2090.810 ;
        RECT 1439.405 2090.495 1439.735 2090.510 ;
        RECT 1440.325 2090.495 1440.655 2090.510 ;
        RECT 1016.665 2052.050 1016.995 2052.065 ;
        RECT 1334.270 2052.050 1334.650 2052.060 ;
        RECT 1016.665 2051.750 1334.650 2052.050 ;
        RECT 1016.665 2051.735 1016.995 2051.750 ;
        RECT 1334.270 2051.740 1334.650 2051.750 ;
        RECT 1159.265 2051.370 1159.595 2051.385 ;
        RECT 1339.790 2051.370 1340.170 2051.380 ;
        RECT 1159.265 2051.070 1340.170 2051.370 ;
        RECT 1159.265 2051.055 1159.595 2051.070 ;
        RECT 1339.790 2051.060 1340.170 2051.070 ;
        RECT 1130.745 2050.690 1131.075 2050.705 ;
        RECT 1338.870 2050.690 1339.250 2050.700 ;
        RECT 1130.745 2050.390 1339.250 2050.690 ;
        RECT 1130.745 2050.375 1131.075 2050.390 ;
        RECT 1338.870 2050.380 1339.250 2050.390 ;
        RECT 1315.665 2050.010 1315.995 2050.025 ;
        RECT 1340.710 2050.010 1341.090 2050.020 ;
        RECT 1315.665 2049.710 1341.090 2050.010 ;
        RECT 1315.665 2049.695 1315.995 2049.710 ;
        RECT 1340.710 2049.700 1341.090 2049.710 ;
        RECT 1439.865 2042.530 1440.195 2042.545 ;
        RECT 1441.705 2042.530 1442.035 2042.545 ;
        RECT 1439.865 2042.230 1442.035 2042.530 ;
        RECT 1439.865 2042.215 1440.195 2042.230 ;
        RECT 1441.705 2042.215 1442.035 2042.230 ;
      LAYER met3 ;
        RECT 1004.000 2019.280 1329.390 2032.005 ;
      LAYER met3 ;
        RECT 994.125 2018.730 994.455 2018.745 ;
        RECT 1000.000 2018.730 1004.000 2018.880 ;
        RECT 994.125 2018.430 1004.000 2018.730 ;
        RECT 994.125 2018.415 994.455 2018.430 ;
        RECT 1000.000 2018.280 1004.000 2018.430 ;
      LAYER met3 ;
        RECT 1004.400 2017.880 1328.990 2019.280 ;
      LAYER met3 ;
        RECT 1329.390 2018.730 1333.390 2018.880 ;
        RECT 1339.125 2018.730 1339.455 2018.745 ;
        RECT 1329.390 2018.430 1339.455 2018.730 ;
        RECT 1329.390 2018.280 1333.390 2018.430 ;
        RECT 1339.125 2018.415 1339.455 2018.430 ;
      LAYER met3 ;
        RECT 1004.000 1998.880 1329.390 2017.880 ;
      LAYER met3 ;
        RECT 992.285 1998.330 992.615 1998.345 ;
        RECT 1000.000 1998.330 1004.000 1998.480 ;
        RECT 992.285 1998.030 1004.000 1998.330 ;
        RECT 992.285 1998.015 992.615 1998.030 ;
        RECT 1000.000 1997.880 1004.000 1998.030 ;
      LAYER met3 ;
        RECT 1004.400 1997.480 1328.990 1998.880 ;
      LAYER met3 ;
        RECT 1329.390 1998.330 1333.390 1998.480 ;
        RECT 1335.905 1998.330 1336.235 1998.345 ;
        RECT 1329.390 1998.030 1336.235 1998.330 ;
        RECT 1329.390 1997.880 1333.390 1998.030 ;
        RECT 1335.905 1998.015 1336.235 1998.030 ;
      LAYER met3 ;
        RECT 1004.000 1977.120 1329.390 1997.480 ;
      LAYER met3 ;
        RECT 994.585 1976.570 994.915 1976.585 ;
        RECT 1000.000 1976.570 1004.000 1976.720 ;
        RECT 994.585 1976.270 1004.000 1976.570 ;
        RECT 994.585 1976.255 994.915 1976.270 ;
        RECT 1000.000 1976.120 1004.000 1976.270 ;
      LAYER met3 ;
        RECT 1004.400 1975.720 1328.990 1977.120 ;
      LAYER met3 ;
        RECT 1329.390 1976.570 1333.390 1976.720 ;
        RECT 1339.585 1976.570 1339.915 1976.585 ;
        RECT 1329.390 1976.270 1339.915 1976.570 ;
        RECT 1329.390 1976.120 1333.390 1976.270 ;
        RECT 1339.585 1976.255 1339.915 1976.270 ;
      LAYER met3 ;
        RECT 364.000 1963.520 627.030 1969.445 ;
        RECT 364.400 1962.120 627.030 1963.520 ;
        RECT 364.000 1940.400 627.030 1962.120 ;
        RECT 1004.000 1956.720 1329.390 1975.720 ;
      LAYER met3 ;
        RECT 995.045 1956.170 995.375 1956.185 ;
        RECT 1000.000 1956.170 1004.000 1956.320 ;
        RECT 995.045 1955.870 1004.000 1956.170 ;
        RECT 995.045 1955.855 995.375 1955.870 ;
        RECT 1000.000 1955.720 1004.000 1955.870 ;
      LAYER met3 ;
        RECT 1004.400 1955.320 1328.990 1956.720 ;
      LAYER met3 ;
        RECT 1329.390 1956.170 1333.390 1956.320 ;
        RECT 1340.045 1956.170 1340.375 1956.185 ;
        RECT 1329.390 1955.870 1340.375 1956.170 ;
        RECT 1329.390 1955.720 1333.390 1955.870 ;
        RECT 1340.045 1955.855 1340.375 1955.870 ;
      LAYER met3 ;
        RECT 364.000 1939.000 626.630 1940.400 ;
        RECT 364.000 1926.800 627.030 1939.000 ;
        RECT 1004.000 1936.320 1329.390 1955.320 ;
      LAYER met3 ;
        RECT 1441.705 1945.970 1442.035 1945.985 ;
        RECT 1442.625 1945.970 1442.955 1945.985 ;
        RECT 1441.705 1945.670 1442.955 1945.970 ;
        RECT 1441.705 1945.655 1442.035 1945.670 ;
        RECT 1442.625 1945.655 1442.955 1945.670 ;
        RECT 991.825 1935.770 992.155 1935.785 ;
        RECT 1000.000 1935.770 1004.000 1935.920 ;
        RECT 991.825 1935.470 1004.000 1935.770 ;
        RECT 991.825 1935.455 992.155 1935.470 ;
        RECT 1000.000 1935.320 1004.000 1935.470 ;
      LAYER met3 ;
        RECT 1004.400 1934.960 1329.390 1936.320 ;
        RECT 1004.400 1934.920 1328.990 1934.960 ;
        RECT 364.400 1925.400 627.030 1926.800 ;
        RECT 364.000 1903.680 627.030 1925.400 ;
        RECT 1004.000 1933.560 1328.990 1934.920 ;
      LAYER met3 ;
        RECT 1329.390 1934.410 1333.390 1934.560 ;
        RECT 1340.505 1934.410 1340.835 1934.425 ;
        RECT 1329.390 1934.110 1340.835 1934.410 ;
        RECT 1329.390 1933.960 1333.390 1934.110 ;
        RECT 1340.505 1934.095 1340.835 1934.110 ;
      LAYER met3 ;
        RECT 1004.000 1914.560 1329.390 1933.560 ;
      LAYER met3 ;
        RECT 995.505 1914.010 995.835 1914.025 ;
        RECT 1000.000 1914.010 1004.000 1914.160 ;
        RECT 995.505 1913.710 1004.000 1914.010 ;
        RECT 995.505 1913.695 995.835 1913.710 ;
        RECT 1000.000 1913.560 1004.000 1913.710 ;
      LAYER met3 ;
        RECT 1004.400 1913.160 1328.990 1914.560 ;
      LAYER met3 ;
        RECT 1329.390 1914.010 1333.390 1914.160 ;
        RECT 1340.965 1914.010 1341.295 1914.025 ;
        RECT 1329.390 1913.710 1341.295 1914.010 ;
        RECT 1329.390 1913.560 1333.390 1913.710 ;
        RECT 1340.965 1913.695 1341.295 1913.710 ;
      LAYER met3 ;
        RECT 364.000 1902.280 626.630 1903.680 ;
        RECT 364.000 1890.080 627.030 1902.280 ;
        RECT 1004.000 1894.160 1329.390 1913.160 ;
        RECT 1924.400 1906.040 2072.375 1906.905 ;
      LAYER met3 ;
        RECT 989.985 1893.610 990.315 1893.625 ;
        RECT 1000.000 1893.610 1004.000 1893.760 ;
        RECT 989.985 1893.310 1004.000 1893.610 ;
        RECT 989.985 1893.295 990.315 1893.310 ;
        RECT 1000.000 1893.160 1004.000 1893.310 ;
      LAYER met3 ;
        RECT 1004.400 1892.800 1329.390 1894.160 ;
        RECT 1924.000 1904.720 2072.375 1906.040 ;
        RECT 1924.000 1903.320 2071.975 1904.720 ;
        RECT 1004.400 1892.760 1328.990 1892.800 ;
        RECT 364.400 1888.680 627.030 1890.080 ;
        RECT 364.000 1866.960 627.030 1888.680 ;
        RECT 1004.000 1891.400 1328.990 1892.760 ;
      LAYER met3 ;
        RECT 1329.390 1892.250 1333.390 1892.400 ;
        RECT 1341.425 1892.250 1341.755 1892.265 ;
        RECT 1329.390 1891.950 1341.755 1892.250 ;
        RECT 1329.390 1891.800 1333.390 1891.950 ;
        RECT 1341.425 1891.935 1341.755 1891.950 ;
      LAYER met3 ;
        RECT 1004.000 1872.400 1329.390 1891.400 ;
        RECT 1924.000 1889.760 2072.375 1903.320 ;
      LAYER met3 ;
        RECT 1920.000 1888.760 1924.000 1889.360 ;
        RECT 1904.465 1886.130 1904.795 1886.145 ;
        RECT 1920.350 1886.130 1920.650 1888.760 ;
      LAYER met3 ;
        RECT 1924.400 1888.400 2072.375 1889.760 ;
        RECT 2304.000 1891.440 2523.025 1925.925 ;
      LAYER met3 ;
        RECT 2523.625 1892.250 2523.955 1892.265 ;
        RECT 2523.625 1891.935 2524.170 1892.250 ;
      LAYER met3 ;
        RECT 2304.000 1890.040 2522.625 1891.440 ;
      LAYER met3 ;
        RECT 2523.870 1891.040 2524.170 1891.935 ;
        RECT 2523.025 1890.440 2527.025 1891.040 ;
      LAYER met3 ;
        RECT 1924.400 1888.360 2071.975 1888.400 ;
      LAYER met3 ;
        RECT 1904.465 1885.830 1920.650 1886.130 ;
      LAYER met3 ;
        RECT 1924.000 1887.000 2071.975 1888.360 ;
      LAYER met3 ;
        RECT 2072.375 1887.400 2076.375 1888.000 ;
        RECT 1904.465 1885.815 1904.795 1885.830 ;
      LAYER met3 ;
        RECT 1924.000 1873.440 2072.375 1887.000 ;
      LAYER met3 ;
        RECT 2075.830 1884.770 2076.130 1887.400 ;
        RECT 2083.865 1884.770 2084.195 1884.785 ;
        RECT 2075.830 1884.470 2084.195 1884.770 ;
        RECT 2083.865 1884.455 2084.195 1884.470 ;
      LAYER met3 ;
        RECT 2304.000 1876.480 2523.025 1890.040 ;
      LAYER met3 ;
        RECT 2283.965 1875.930 2284.295 1875.945 ;
        RECT 2300.000 1875.930 2304.000 1876.080 ;
        RECT 2283.965 1875.630 2304.000 1875.930 ;
        RECT 2283.965 1875.615 2284.295 1875.630 ;
        RECT 2300.000 1875.480 2304.000 1875.630 ;
      LAYER met3 ;
        RECT 2304.400 1875.080 2523.025 1876.480 ;
      LAYER met3 ;
        RECT 1920.000 1872.440 1924.000 1873.040 ;
        RECT 989.525 1871.850 989.855 1871.865 ;
        RECT 1000.000 1871.850 1004.000 1872.000 ;
        RECT 989.525 1871.550 1004.000 1871.850 ;
        RECT 989.525 1871.535 989.855 1871.550 ;
        RECT 1000.000 1871.400 1004.000 1871.550 ;
      LAYER met3 ;
        RECT 1004.400 1871.000 1328.990 1872.400 ;
      LAYER met3 ;
        RECT 1329.390 1871.850 1333.390 1872.000 ;
        RECT 1341.885 1871.850 1342.215 1871.865 ;
        RECT 1329.390 1871.550 1342.215 1871.850 ;
        RECT 1329.390 1871.400 1333.390 1871.550 ;
        RECT 1341.885 1871.535 1342.215 1871.550 ;
      LAYER met3 ;
        RECT 364.000 1865.560 626.630 1866.960 ;
        RECT 364.000 1852.000 627.030 1865.560 ;
        RECT 1004.000 1852.000 1329.390 1871.000 ;
      LAYER met3 ;
        RECT 1904.465 1870.490 1904.795 1870.505 ;
        RECT 1920.350 1870.490 1920.650 1872.440 ;
      LAYER met3 ;
        RECT 1924.400 1872.040 2072.375 1873.440 ;
      LAYER met3 ;
        RECT 1904.465 1870.190 1920.650 1870.490 ;
      LAYER met3 ;
        RECT 1924.000 1870.720 2072.375 1872.040 ;
      LAYER met3 ;
        RECT 1904.465 1870.175 1904.795 1870.190 ;
      LAYER met3 ;
        RECT 1924.000 1869.320 2071.975 1870.720 ;
        RECT 1924.000 1855.760 2072.375 1869.320 ;
      LAYER met3 ;
        RECT 1920.000 1854.760 1924.000 1855.360 ;
      LAYER met3 ;
        RECT 364.400 1850.600 627.030 1852.000 ;
      LAYER met3 ;
        RECT 989.065 1851.450 989.395 1851.465 ;
        RECT 1000.000 1851.450 1004.000 1851.600 ;
        RECT 989.065 1851.150 1004.000 1851.450 ;
        RECT 989.065 1851.135 989.395 1851.150 ;
        RECT 1000.000 1851.000 1004.000 1851.150 ;
      LAYER met3 ;
        RECT 1004.400 1850.640 1329.390 1852.000 ;
      LAYER met3 ;
        RECT 1904.465 1852.130 1904.795 1852.145 ;
        RECT 1920.350 1852.130 1920.650 1854.760 ;
      LAYER met3 ;
        RECT 1924.400 1854.400 2072.375 1855.760 ;
        RECT 1924.400 1854.360 2071.975 1854.400 ;
      LAYER met3 ;
        RECT 1904.465 1851.830 1920.650 1852.130 ;
      LAYER met3 ;
        RECT 1924.000 1853.000 2071.975 1854.360 ;
      LAYER met3 ;
        RECT 2072.375 1853.400 2076.375 1854.000 ;
        RECT 1904.465 1851.815 1904.795 1851.830 ;
      LAYER met3 ;
        RECT 1004.400 1850.600 1328.990 1850.640 ;
        RECT 364.000 1830.240 627.030 1850.600 ;
        RECT 1004.000 1849.240 1328.990 1850.600 ;
      LAYER met3 ;
        RECT 1329.390 1850.090 1333.390 1850.240 ;
        RECT 1342.345 1850.090 1342.675 1850.105 ;
        RECT 1329.390 1849.790 1342.675 1850.090 ;
        RECT 1329.390 1849.640 1333.390 1849.790 ;
        RECT 1342.345 1849.775 1342.675 1849.790 ;
        RECT 1441.705 1849.410 1442.035 1849.425 ;
        RECT 1442.625 1849.410 1442.955 1849.425 ;
      LAYER met3 ;
        RECT 1004.000 1830.240 1329.390 1849.240 ;
      LAYER met3 ;
        RECT 1441.705 1849.110 1442.955 1849.410 ;
        RECT 1441.705 1849.095 1442.035 1849.110 ;
        RECT 1442.625 1849.095 1442.955 1849.110 ;
      LAYER met3 ;
        RECT 1924.000 1839.440 2072.375 1853.000 ;
      LAYER met3 ;
        RECT 2075.830 1850.770 2076.130 1853.400 ;
        RECT 2084.325 1850.770 2084.655 1850.785 ;
        RECT 2075.830 1850.470 2084.655 1850.770 ;
        RECT 2084.325 1850.455 2084.655 1850.470 ;
      LAYER met3 ;
        RECT 1924.400 1838.040 2072.375 1839.440 ;
        RECT 1924.000 1836.720 2072.375 1838.040 ;
        RECT 1924.000 1835.320 2071.975 1836.720 ;
      LAYER met3 ;
        RECT 2072.375 1835.810 2076.375 1836.320 ;
        RECT 2084.785 1835.810 2085.115 1835.825 ;
        RECT 2072.375 1835.720 2085.115 1835.810 ;
        RECT 2075.830 1835.510 2085.115 1835.720 ;
        RECT 2084.785 1835.495 2085.115 1835.510 ;
      LAYER met3 ;
        RECT 364.000 1828.840 626.630 1830.240 ;
      LAYER met3 ;
        RECT 995.965 1829.690 996.295 1829.705 ;
        RECT 1000.000 1829.690 1004.000 1829.840 ;
        RECT 995.965 1829.390 1004.000 1829.690 ;
        RECT 995.965 1829.375 996.295 1829.390 ;
        RECT 1000.000 1829.240 1004.000 1829.390 ;
      LAYER met3 ;
        RECT 1004.400 1828.840 1328.990 1830.240 ;
      LAYER met3 ;
        RECT 1329.390 1829.690 1333.390 1829.840 ;
        RECT 1342.805 1829.690 1343.135 1829.705 ;
        RECT 1329.390 1829.390 1343.135 1829.690 ;
        RECT 1329.390 1829.240 1333.390 1829.390 ;
        RECT 1342.805 1829.375 1343.135 1829.390 ;
      LAYER met3 ;
        RECT 364.000 1815.280 627.030 1828.840 ;
        RECT 364.400 1813.880 627.030 1815.280 ;
        RECT 364.000 1792.160 627.030 1813.880 ;
        RECT 1004.000 1809.840 1329.390 1828.840 ;
        RECT 1924.000 1821.760 2072.375 1835.320 ;
      LAYER met3 ;
        RECT 1920.000 1820.760 1924.000 1821.360 ;
        RECT 1904.465 1818.130 1904.795 1818.145 ;
        RECT 1920.350 1818.130 1920.650 1820.760 ;
      LAYER met3 ;
        RECT 1924.400 1820.400 2072.375 1821.760 ;
        RECT 1924.400 1820.360 2071.975 1820.400 ;
      LAYER met3 ;
        RECT 1904.465 1817.830 1920.650 1818.130 ;
      LAYER met3 ;
        RECT 1924.000 1819.000 2071.975 1820.360 ;
      LAYER met3 ;
        RECT 2072.375 1819.830 2076.375 1820.000 ;
        RECT 2076.965 1819.830 2077.295 1819.845 ;
        RECT 2072.375 1819.530 2077.295 1819.830 ;
        RECT 2072.375 1819.400 2076.375 1819.530 ;
        RECT 2076.965 1819.515 2077.295 1819.530 ;
        RECT 1904.465 1817.815 1904.795 1817.830 ;
        RECT 988.605 1809.290 988.935 1809.305 ;
        RECT 1000.000 1809.290 1004.000 1809.440 ;
        RECT 988.605 1808.990 1004.000 1809.290 ;
        RECT 988.605 1808.975 988.935 1808.990 ;
        RECT 1000.000 1808.840 1004.000 1808.990 ;
      LAYER met3 ;
        RECT 1004.400 1808.480 1329.390 1809.840 ;
        RECT 1004.400 1808.440 1328.990 1808.480 ;
        RECT 1004.000 1807.080 1328.990 1808.440 ;
      LAYER met3 ;
        RECT 1329.390 1807.930 1333.390 1808.080 ;
        RECT 1343.265 1807.930 1343.595 1807.945 ;
        RECT 1329.390 1807.630 1343.595 1807.930 ;
        RECT 1329.390 1807.480 1333.390 1807.630 ;
        RECT 1343.265 1807.615 1343.595 1807.630 ;
      LAYER met3 ;
        RECT 364.000 1790.760 626.630 1792.160 ;
        RECT 364.000 1778.560 627.030 1790.760 ;
        RECT 1004.000 1788.080 1329.390 1807.080 ;
        RECT 1924.000 1805.440 2072.375 1819.000 ;
        RECT 1924.400 1804.040 2072.375 1805.440 ;
        RECT 1924.000 1802.720 2072.375 1804.040 ;
        RECT 2304.000 1805.760 2523.025 1875.080 ;
        RECT 2304.000 1804.360 2522.625 1805.760 ;
      LAYER met3 ;
        RECT 2523.025 1804.760 2527.025 1805.360 ;
      LAYER met3 ;
        RECT 1924.000 1801.320 2071.975 1802.720 ;
      LAYER met3 ;
        RECT 2072.375 1801.720 2076.375 1802.320 ;
        RECT 987.685 1787.530 988.015 1787.545 ;
        RECT 1000.000 1787.530 1004.000 1787.680 ;
        RECT 987.685 1787.230 1004.000 1787.530 ;
        RECT 987.685 1787.215 988.015 1787.230 ;
        RECT 1000.000 1787.080 1004.000 1787.230 ;
      LAYER met3 ;
        RECT 1004.400 1786.680 1328.990 1788.080 ;
        RECT 1924.000 1787.760 2072.375 1801.320 ;
      LAYER met3 ;
        RECT 2075.830 1801.130 2076.130 1801.720 ;
        RECT 2085.245 1801.130 2085.575 1801.145 ;
        RECT 2075.830 1800.830 2085.575 1801.130 ;
        RECT 2085.245 1800.815 2085.575 1800.830 ;
      LAYER met3 ;
        RECT 2304.000 1790.800 2523.025 1804.360 ;
      LAYER met3 ;
        RECT 2523.870 1802.505 2524.170 1804.760 ;
        RECT 2523.625 1802.190 2524.170 1802.505 ;
        RECT 2523.625 1802.175 2523.955 1802.190 ;
        RECT 2287.185 1790.250 2287.515 1790.265 ;
        RECT 2300.000 1790.250 2304.000 1790.400 ;
        RECT 2287.185 1789.950 2304.000 1790.250 ;
        RECT 2287.185 1789.935 2287.515 1789.950 ;
        RECT 2300.000 1789.800 2304.000 1789.950 ;
      LAYER met3 ;
        RECT 2304.400 1789.400 2523.025 1790.800 ;
      LAYER met3 ;
        RECT 1329.390 1787.530 1333.390 1787.680 ;
        RECT 1336.365 1787.530 1336.695 1787.545 ;
        RECT 1329.390 1787.230 1336.695 1787.530 ;
        RECT 1329.390 1787.080 1333.390 1787.230 ;
        RECT 1336.365 1787.215 1336.695 1787.230 ;
      LAYER met3 ;
        RECT 364.400 1777.160 627.030 1778.560 ;
        RECT 364.000 1755.440 627.030 1777.160 ;
        RECT 1004.000 1767.680 1329.390 1786.680 ;
        RECT 1924.400 1786.400 2072.375 1787.760 ;
        RECT 1924.400 1786.360 2071.975 1786.400 ;
        RECT 1924.000 1785.000 2071.975 1786.360 ;
      LAYER met3 ;
        RECT 2072.375 1785.400 2076.375 1786.000 ;
      LAYER met3 ;
        RECT 1924.000 1771.440 2072.375 1785.000 ;
      LAYER met3 ;
        RECT 2075.830 1782.770 2076.130 1785.400 ;
        RECT 2085.705 1782.770 2086.035 1782.785 ;
        RECT 2075.830 1782.470 2086.035 1782.770 ;
        RECT 2085.705 1782.455 2086.035 1782.470 ;
        RECT 1920.000 1770.440 1924.000 1771.040 ;
        RECT 1904.465 1767.810 1904.795 1767.825 ;
        RECT 1920.350 1767.810 1920.650 1770.440 ;
      LAYER met3 ;
        RECT 1924.400 1770.040 2072.375 1771.440 ;
      LAYER met3 ;
        RECT 987.225 1767.130 987.555 1767.145 ;
        RECT 1000.000 1767.130 1004.000 1767.280 ;
        RECT 987.225 1766.830 1004.000 1767.130 ;
        RECT 987.225 1766.815 987.555 1766.830 ;
        RECT 1000.000 1766.680 1004.000 1766.830 ;
      LAYER met3 ;
        RECT 1004.400 1766.280 1328.990 1767.680 ;
      LAYER met3 ;
        RECT 1904.465 1767.510 1920.650 1767.810 ;
      LAYER met3 ;
        RECT 1924.000 1768.720 2072.375 1770.040 ;
      LAYER met3 ;
        RECT 1904.465 1767.495 1904.795 1767.510 ;
      LAYER met3 ;
        RECT 1924.000 1767.320 2071.975 1768.720 ;
      LAYER met3 ;
        RECT 2072.375 1767.720 2076.375 1768.320 ;
        RECT 1329.390 1767.130 1333.390 1767.280 ;
        RECT 1336.825 1767.130 1337.155 1767.145 ;
        RECT 1329.390 1766.830 1337.155 1767.130 ;
        RECT 1329.390 1766.680 1333.390 1766.830 ;
        RECT 1336.825 1766.815 1337.155 1766.830 ;
      LAYER met3 ;
        RECT 364.000 1754.040 626.630 1755.440 ;
        RECT 364.000 1741.840 627.030 1754.040 ;
        RECT 1004.000 1745.920 1329.390 1766.280 ;
        RECT 1924.000 1760.715 2072.375 1767.320 ;
      LAYER met3 ;
        RECT 2075.830 1767.130 2076.130 1767.720 ;
        RECT 2086.165 1767.130 2086.495 1767.145 ;
        RECT 2075.830 1766.830 2086.495 1767.130 ;
        RECT 2086.165 1766.815 2086.495 1766.830 ;
        RECT 986.765 1745.370 987.095 1745.385 ;
        RECT 1000.000 1745.370 1004.000 1745.520 ;
        RECT 986.765 1745.070 1004.000 1745.370 ;
        RECT 986.765 1745.055 987.095 1745.070 ;
        RECT 1000.000 1744.920 1004.000 1745.070 ;
      LAYER met3 ;
        RECT 1004.400 1744.520 1328.990 1745.920 ;
      LAYER met3 ;
        RECT 1329.390 1745.370 1333.390 1745.520 ;
        RECT 1337.285 1745.370 1337.615 1745.385 ;
        RECT 1329.390 1745.070 1337.615 1745.370 ;
        RECT 1329.390 1744.920 1333.390 1745.070 ;
        RECT 1337.285 1745.055 1337.615 1745.070 ;
      LAYER met3 ;
        RECT 364.400 1740.440 627.030 1741.840 ;
        RECT 364.000 1718.720 627.030 1740.440 ;
        RECT 1004.000 1725.520 1329.390 1744.520 ;
      LAYER met3 ;
        RECT 988.145 1724.970 988.475 1724.985 ;
        RECT 1000.000 1724.970 1004.000 1725.120 ;
        RECT 988.145 1724.670 1004.000 1724.970 ;
        RECT 988.145 1724.655 988.475 1724.670 ;
        RECT 1000.000 1724.520 1004.000 1724.670 ;
      LAYER met3 ;
        RECT 1004.400 1724.120 1328.990 1725.520 ;
      LAYER met3 ;
        RECT 1329.390 1724.970 1333.390 1725.120 ;
        RECT 1345.105 1724.970 1345.435 1724.985 ;
        RECT 1329.390 1724.670 1345.435 1724.970 ;
        RECT 1329.390 1724.520 1333.390 1724.670 ;
        RECT 1345.105 1724.655 1345.435 1724.670 ;
      LAYER met3 ;
        RECT 364.000 1717.320 626.630 1718.720 ;
        RECT 364.000 1710.715 627.030 1717.320 ;
        RECT 1004.000 1710.715 1329.390 1724.120 ;
        RECT 2304.000 1720.080 2523.025 1789.400 ;
        RECT 2304.000 1718.680 2522.625 1720.080 ;
      LAYER met3 ;
        RECT 2523.025 1719.080 2527.025 1719.680 ;
      LAYER met3 ;
        RECT 2304.000 1710.715 2523.025 1718.680 ;
      LAYER met3 ;
        RECT 2523.870 1718.185 2524.170 1719.080 ;
        RECT 2523.625 1717.870 2524.170 1718.185 ;
        RECT 2523.625 1717.855 2523.955 1717.870 ;
        RECT 2518.565 1704.570 2518.895 1704.585 ;
        RECT 2519.485 1704.570 2519.815 1704.585 ;
        RECT 2518.565 1704.270 2519.815 1704.570 ;
        RECT 2518.565 1704.255 2518.895 1704.270 ;
        RECT 2519.485 1704.255 2519.815 1704.270 ;
        RECT 1185.945 1693.690 1186.275 1693.705 ;
        RECT 1340.710 1693.690 1341.090 1693.700 ;
        RECT 1185.945 1693.390 1341.090 1693.690 ;
        RECT 1185.945 1693.375 1186.275 1693.390 ;
        RECT 1340.710 1693.380 1341.090 1693.390 ;
        RECT 1441.705 1663.090 1442.035 1663.105 ;
        RECT 1443.085 1663.090 1443.415 1663.105 ;
        RECT 1441.705 1662.790 1443.415 1663.090 ;
        RECT 1441.705 1662.775 1442.035 1662.790 ;
        RECT 1443.085 1662.775 1443.415 1662.790 ;
        RECT 2519.485 1608.690 2519.815 1608.705 ;
        RECT 2519.270 1608.375 2519.815 1608.690 ;
        RECT 2519.270 1607.345 2519.570 1608.375 ;
        RECT 2519.270 1607.030 2519.815 1607.345 ;
        RECT 2519.485 1607.015 2519.815 1607.030 ;
        RECT 1441.705 1338.730 1442.035 1338.745 ;
        RECT 1442.625 1338.730 1442.955 1338.745 ;
        RECT 1441.705 1338.430 1442.955 1338.730 ;
        RECT 1441.705 1338.415 1442.035 1338.430 ;
        RECT 1442.625 1338.415 1442.955 1338.430 ;
        RECT 1441.705 1290.450 1442.035 1290.465 ;
        RECT 1442.625 1290.450 1442.955 1290.465 ;
        RECT 1441.705 1290.150 1442.955 1290.450 ;
        RECT 1441.705 1290.135 1442.035 1290.150 ;
        RECT 1442.625 1290.135 1442.955 1290.150 ;
        RECT 1522.665 1257.130 1522.995 1257.145 ;
        RECT 1521.990 1256.830 1522.995 1257.130 ;
        RECT 1521.990 1255.785 1522.290 1256.830 ;
        RECT 1522.665 1256.815 1522.995 1256.830 ;
        RECT 1521.745 1255.470 1522.290 1255.785 ;
        RECT 1521.745 1255.455 1522.075 1255.470 ;
        RECT 1441.705 1159.210 1442.035 1159.225 ;
        RECT 1442.625 1159.210 1442.955 1159.225 ;
        RECT 1441.705 1158.910 1442.955 1159.210 ;
        RECT 1441.705 1158.895 1442.035 1158.910 ;
        RECT 1442.625 1158.895 1442.955 1158.910 ;
        RECT 1520.365 1055.850 1520.695 1055.865 ;
        RECT 1521.285 1055.850 1521.615 1055.865 ;
        RECT 1520.365 1055.550 1521.615 1055.850 ;
        RECT 1520.365 1055.535 1520.695 1055.550 ;
        RECT 1521.285 1055.535 1521.615 1055.550 ;
        RECT 985.385 1014.370 985.715 1014.385 ;
        RECT 1101.765 1014.370 1102.095 1014.385 ;
        RECT 985.385 1014.070 1102.095 1014.370 ;
        RECT 985.385 1014.055 985.715 1014.070 ;
        RECT 1101.765 1014.055 1102.095 1014.070 ;
        RECT 984.925 1013.690 985.255 1013.705 ;
        RECT 1119.245 1013.690 1119.575 1013.705 ;
        RECT 984.925 1013.390 1119.575 1013.690 ;
        RECT 984.925 1013.375 985.255 1013.390 ;
        RECT 1119.245 1013.375 1119.575 1013.390 ;
        RECT 989.270 1013.010 989.650 1013.020 ;
        RECT 1125.685 1013.010 1126.015 1013.025 ;
        RECT 989.270 1012.710 1126.015 1013.010 ;
        RECT 989.270 1012.700 989.650 1012.710 ;
        RECT 1125.685 1012.695 1126.015 1012.710 ;
        RECT 986.305 1012.330 986.635 1012.345 ;
        RECT 1131.665 1012.330 1131.995 1012.345 ;
        RECT 986.305 1012.030 1131.995 1012.330 ;
        RECT 986.305 1012.015 986.635 1012.030 ;
        RECT 1131.665 1012.015 1131.995 1012.030 ;
        RECT 1158.345 1012.330 1158.675 1012.345 ;
        RECT 1200.205 1012.330 1200.535 1012.345 ;
        RECT 1158.345 1012.030 1200.535 1012.330 ;
        RECT 1158.345 1012.015 1158.675 1012.030 ;
        RECT 1200.205 1012.015 1200.535 1012.030 ;
        RECT 991.110 1011.650 991.490 1011.660 ;
        RECT 1160.645 1011.650 1160.975 1011.665 ;
        RECT 991.110 1011.350 1160.975 1011.650 ;
        RECT 991.110 1011.340 991.490 1011.350 ;
        RECT 1160.645 1011.335 1160.975 1011.350 ;
        RECT 985.845 1010.970 986.175 1010.985 ;
        RECT 1167.085 1010.970 1167.415 1010.985 ;
        RECT 985.845 1010.670 1167.415 1010.970 ;
        RECT 985.845 1010.655 986.175 1010.670 ;
        RECT 1167.085 1010.655 1167.415 1010.670 ;
        RECT 1285.305 1010.970 1285.635 1010.985 ;
        RECT 1339.790 1010.970 1340.170 1010.980 ;
        RECT 1285.305 1010.670 1340.170 1010.970 ;
        RECT 1285.305 1010.655 1285.635 1010.670 ;
        RECT 1339.790 1010.660 1340.170 1010.670 ;
        RECT 998.470 1010.290 998.850 1010.300 ;
        RECT 1090.265 1010.290 1090.595 1010.305 ;
        RECT 998.470 1009.990 1090.595 1010.290 ;
        RECT 998.470 1009.980 998.850 1009.990 ;
        RECT 1090.265 1009.975 1090.595 1009.990 ;
        RECT 1160.185 1010.290 1160.515 1010.305 ;
        RECT 1191.465 1010.290 1191.795 1010.305 ;
        RECT 1160.185 1009.990 1191.795 1010.290 ;
        RECT 1160.185 1009.975 1160.515 1009.990 ;
        RECT 1191.465 1009.975 1191.795 1009.990 ;
        RECT 992.030 1009.610 992.410 1009.620 ;
        RECT 1062.665 1009.610 1062.995 1009.625 ;
        RECT 992.030 1009.310 1062.995 1009.610 ;
        RECT 992.030 1009.300 992.410 1009.310 ;
        RECT 1062.665 1009.295 1062.995 1009.310 ;
        RECT 1146.385 1009.610 1146.715 1009.625 ;
        RECT 1176.285 1009.610 1176.615 1009.625 ;
        RECT 1146.385 1009.310 1176.615 1009.610 ;
        RECT 1146.385 1009.295 1146.715 1009.310 ;
        RECT 1176.285 1009.295 1176.615 1009.310 ;
        RECT 992.950 1008.930 993.330 1008.940 ;
        RECT 1067.265 1008.930 1067.595 1008.945 ;
        RECT 992.950 1008.630 1067.595 1008.930 ;
        RECT 992.950 1008.620 993.330 1008.630 ;
        RECT 1067.265 1008.615 1067.595 1008.630 ;
        RECT 1111.425 1008.930 1111.755 1008.945 ;
        RECT 1158.345 1008.930 1158.675 1008.945 ;
        RECT 1111.425 1008.630 1158.675 1008.930 ;
        RECT 1111.425 1008.615 1111.755 1008.630 ;
        RECT 1158.345 1008.615 1158.675 1008.630 ;
        RECT 1159.265 1008.930 1159.595 1008.945 ;
        RECT 1161.105 1008.930 1161.435 1008.945 ;
        RECT 1159.265 1008.630 1161.435 1008.930 ;
        RECT 1159.265 1008.615 1159.595 1008.630 ;
        RECT 1161.105 1008.615 1161.435 1008.630 ;
        RECT 1207.565 1008.930 1207.895 1008.945 ;
        RECT 1209.405 1008.930 1209.735 1008.945 ;
        RECT 1207.565 1008.630 1209.735 1008.930 ;
        RECT 1207.565 1008.615 1207.895 1008.630 ;
        RECT 1209.405 1008.615 1209.735 1008.630 ;
        RECT 990.190 1008.250 990.570 1008.260 ;
        RECT 1055.765 1008.250 1056.095 1008.265 ;
        RECT 990.190 1007.950 1056.095 1008.250 ;
        RECT 990.190 1007.940 990.570 1007.950 ;
        RECT 1055.765 1007.935 1056.095 1007.950 ;
        RECT 1159.725 1008.250 1160.055 1008.265 ;
        RECT 1166.625 1008.250 1166.955 1008.265 ;
        RECT 1159.725 1007.950 1166.955 1008.250 ;
        RECT 1159.725 1007.935 1160.055 1007.950 ;
        RECT 1166.625 1007.935 1166.955 1007.950 ;
        RECT 1207.565 1008.250 1207.895 1008.265 ;
        RECT 1209.405 1008.250 1209.735 1008.265 ;
        RECT 1207.565 1007.950 1209.735 1008.250 ;
        RECT 1207.565 1007.935 1207.895 1007.950 ;
        RECT 1209.405 1007.935 1209.735 1007.950 ;
        RECT 1313.365 1008.250 1313.695 1008.265 ;
        RECT 1338.870 1008.250 1339.250 1008.260 ;
        RECT 1313.365 1007.950 1339.250 1008.250 ;
        RECT 1313.365 1007.935 1313.695 1007.950 ;
        RECT 1338.870 1007.940 1339.250 1007.950 ;
        RECT 1330.845 1007.570 1331.175 1007.585 ;
        RECT 1334.270 1007.570 1334.650 1007.580 ;
        RECT 1330.845 1007.270 1334.650 1007.570 ;
        RECT 1330.845 1007.255 1331.175 1007.270 ;
        RECT 1334.270 1007.260 1334.650 1007.270 ;
      LAYER met3 ;
        RECT 674.400 996.080 2166.000 996.945 ;
        RECT 674.000 994.760 2166.000 996.080 ;
        RECT 674.000 993.360 2165.600 994.760 ;
        RECT 674.000 992.040 2166.000 993.360 ;
        RECT 674.400 990.640 2166.000 992.040 ;
        RECT 674.000 986.600 2166.000 990.640 ;
        RECT 674.400 985.200 2166.000 986.600 ;
        RECT 674.000 984.560 2166.000 985.200 ;
        RECT 674.000 983.160 2165.600 984.560 ;
        RECT 674.000 981.840 2166.000 983.160 ;
        RECT 674.400 980.440 2166.000 981.840 ;
        RECT 674.000 976.400 2166.000 980.440 ;
        RECT 674.400 975.000 2166.000 976.400 ;
        RECT 674.000 973.680 2166.000 975.000 ;
        RECT 674.000 972.280 2165.600 973.680 ;
        RECT 674.000 970.960 2166.000 972.280 ;
        RECT 674.400 969.560 2166.000 970.960 ;
        RECT 674.000 965.520 2166.000 969.560 ;
        RECT 674.400 964.120 2166.000 965.520 ;
        RECT 674.000 963.480 2166.000 964.120 ;
        RECT 674.000 962.080 2165.600 963.480 ;
        RECT 674.000 960.760 2166.000 962.080 ;
        RECT 674.400 959.360 2166.000 960.760 ;
        RECT 674.000 955.320 2166.000 959.360 ;
        RECT 674.400 953.920 2166.000 955.320 ;
        RECT 674.000 952.600 2166.000 953.920 ;
        RECT 674.000 951.200 2165.600 952.600 ;
        RECT 674.000 949.880 2166.000 951.200 ;
        RECT 674.400 948.480 2166.000 949.880 ;
        RECT 674.000 944.440 2166.000 948.480 ;
        RECT 674.400 943.040 2166.000 944.440 ;
        RECT 674.000 942.400 2166.000 943.040 ;
        RECT 674.000 941.000 2165.600 942.400 ;
        RECT 674.000 939.680 2166.000 941.000 ;
        RECT 674.400 938.280 2166.000 939.680 ;
        RECT 674.000 934.240 2166.000 938.280 ;
        RECT 674.400 932.840 2166.000 934.240 ;
        RECT 674.000 931.520 2166.000 932.840 ;
        RECT 674.000 930.120 2165.600 931.520 ;
        RECT 674.000 928.800 2166.000 930.120 ;
        RECT 674.400 927.400 2166.000 928.800 ;
        RECT 674.000 923.360 2166.000 927.400 ;
        RECT 674.400 921.960 2166.000 923.360 ;
        RECT 674.000 921.320 2166.000 921.960 ;
        RECT 674.000 919.920 2165.600 921.320 ;
        RECT 674.000 918.600 2166.000 919.920 ;
        RECT 674.400 917.200 2166.000 918.600 ;
        RECT 674.000 913.160 2166.000 917.200 ;
        RECT 674.400 911.760 2166.000 913.160 ;
        RECT 674.000 910.440 2166.000 911.760 ;
        RECT 674.000 909.040 2165.600 910.440 ;
        RECT 674.000 907.720 2166.000 909.040 ;
        RECT 674.400 906.320 2166.000 907.720 ;
        RECT 674.000 902.960 2166.000 906.320 ;
        RECT 674.400 901.560 2166.000 902.960 ;
        RECT 674.000 900.240 2166.000 901.560 ;
        RECT 674.000 898.840 2165.600 900.240 ;
        RECT 674.000 897.520 2166.000 898.840 ;
        RECT 674.400 896.120 2166.000 897.520 ;
        RECT 674.000 892.080 2166.000 896.120 ;
        RECT 674.400 890.680 2166.000 892.080 ;
        RECT 674.000 889.360 2166.000 890.680 ;
        RECT 674.000 887.960 2165.600 889.360 ;
        RECT 674.000 886.640 2166.000 887.960 ;
        RECT 674.400 885.240 2166.000 886.640 ;
        RECT 674.000 881.880 2166.000 885.240 ;
        RECT 674.400 880.480 2166.000 881.880 ;
        RECT 674.000 879.160 2166.000 880.480 ;
        RECT 674.000 877.760 2165.600 879.160 ;
        RECT 674.000 876.440 2166.000 877.760 ;
        RECT 674.400 875.040 2166.000 876.440 ;
        RECT 674.000 871.000 2166.000 875.040 ;
        RECT 674.400 869.600 2166.000 871.000 ;
        RECT 674.000 868.280 2166.000 869.600 ;
        RECT 674.000 866.880 2165.600 868.280 ;
        RECT 674.000 865.560 2166.000 866.880 ;
        RECT 674.400 864.160 2166.000 865.560 ;
        RECT 674.000 860.800 2166.000 864.160 ;
        RECT 674.400 859.400 2166.000 860.800 ;
        RECT 674.000 858.080 2166.000 859.400 ;
        RECT 674.000 856.680 2165.600 858.080 ;
        RECT 674.000 855.360 2166.000 856.680 ;
        RECT 674.400 853.960 2166.000 855.360 ;
        RECT 674.000 849.920 2166.000 853.960 ;
        RECT 674.400 848.520 2166.000 849.920 ;
        RECT 674.000 847.200 2166.000 848.520 ;
        RECT 674.000 845.800 2165.600 847.200 ;
        RECT 674.000 844.480 2166.000 845.800 ;
        RECT 674.400 843.080 2166.000 844.480 ;
        RECT 674.000 839.720 2166.000 843.080 ;
        RECT 674.400 838.320 2166.000 839.720 ;
        RECT 674.000 837.000 2166.000 838.320 ;
        RECT 674.000 835.600 2165.600 837.000 ;
        RECT 674.000 834.280 2166.000 835.600 ;
        RECT 674.400 832.880 2166.000 834.280 ;
        RECT 674.000 828.840 2166.000 832.880 ;
        RECT 674.400 827.440 2166.000 828.840 ;
        RECT 674.000 826.120 2166.000 827.440 ;
        RECT 674.000 824.720 2165.600 826.120 ;
        RECT 674.000 823.400 2166.000 824.720 ;
        RECT 674.400 822.000 2166.000 823.400 ;
        RECT 674.000 818.640 2166.000 822.000 ;
        RECT 674.400 817.240 2166.000 818.640 ;
        RECT 674.000 815.920 2166.000 817.240 ;
        RECT 674.000 814.520 2165.600 815.920 ;
        RECT 674.000 813.200 2166.000 814.520 ;
        RECT 674.400 811.800 2166.000 813.200 ;
        RECT 674.000 807.760 2166.000 811.800 ;
        RECT 674.400 806.360 2166.000 807.760 ;
        RECT 674.000 805.720 2166.000 806.360 ;
        RECT 674.000 804.320 2165.600 805.720 ;
        RECT 674.000 803.000 2166.000 804.320 ;
        RECT 674.400 801.600 2166.000 803.000 ;
        RECT 674.000 797.560 2166.000 801.600 ;
        RECT 674.400 796.160 2166.000 797.560 ;
        RECT 674.000 794.840 2166.000 796.160 ;
        RECT 674.000 793.440 2165.600 794.840 ;
        RECT 674.000 792.120 2166.000 793.440 ;
        RECT 674.400 790.720 2166.000 792.120 ;
        RECT 674.000 786.680 2166.000 790.720 ;
        RECT 674.400 785.280 2166.000 786.680 ;
        RECT 674.000 784.640 2166.000 785.280 ;
        RECT 674.000 783.240 2165.600 784.640 ;
        RECT 674.000 781.920 2166.000 783.240 ;
        RECT 674.400 780.520 2166.000 781.920 ;
        RECT 674.000 776.480 2166.000 780.520 ;
        RECT 674.400 775.080 2166.000 776.480 ;
        RECT 674.000 773.760 2166.000 775.080 ;
        RECT 674.000 772.360 2165.600 773.760 ;
        RECT 674.000 771.040 2166.000 772.360 ;
        RECT 674.400 769.640 2166.000 771.040 ;
        RECT 674.000 765.600 2166.000 769.640 ;
        RECT 674.400 764.200 2166.000 765.600 ;
        RECT 674.000 763.560 2166.000 764.200 ;
        RECT 674.000 762.160 2165.600 763.560 ;
        RECT 674.000 760.840 2166.000 762.160 ;
        RECT 674.400 759.440 2166.000 760.840 ;
        RECT 674.000 755.400 2166.000 759.440 ;
        RECT 674.400 754.000 2166.000 755.400 ;
        RECT 674.000 752.680 2166.000 754.000 ;
        RECT 674.000 751.280 2165.600 752.680 ;
        RECT 674.000 749.960 2166.000 751.280 ;
        RECT 674.400 748.560 2166.000 749.960 ;
        RECT 674.000 744.520 2166.000 748.560 ;
        RECT 674.400 743.120 2166.000 744.520 ;
        RECT 674.000 742.480 2166.000 743.120 ;
        RECT 674.000 741.080 2165.600 742.480 ;
        RECT 674.000 739.760 2166.000 741.080 ;
        RECT 674.400 738.360 2166.000 739.760 ;
        RECT 674.000 734.320 2166.000 738.360 ;
        RECT 674.400 732.920 2166.000 734.320 ;
        RECT 674.000 731.600 2166.000 732.920 ;
        RECT 674.000 730.200 2165.600 731.600 ;
        RECT 674.000 728.880 2166.000 730.200 ;
        RECT 674.400 727.480 2166.000 728.880 ;
        RECT 674.000 723.440 2166.000 727.480 ;
        RECT 674.400 722.040 2166.000 723.440 ;
        RECT 674.000 721.400 2166.000 722.040 ;
        RECT 674.000 720.000 2165.600 721.400 ;
        RECT 674.000 718.680 2166.000 720.000 ;
        RECT 674.400 717.280 2166.000 718.680 ;
        RECT 674.000 713.240 2166.000 717.280 ;
        RECT 674.400 711.840 2166.000 713.240 ;
        RECT 674.000 710.520 2166.000 711.840 ;
        RECT 674.000 709.120 2165.600 710.520 ;
        RECT 674.000 707.800 2166.000 709.120 ;
        RECT 674.400 706.400 2166.000 707.800 ;
        RECT 674.000 703.040 2166.000 706.400 ;
        RECT 674.400 701.640 2166.000 703.040 ;
        RECT 674.000 700.320 2166.000 701.640 ;
        RECT 674.000 698.920 2165.600 700.320 ;
        RECT 674.000 697.600 2166.000 698.920 ;
        RECT 674.400 696.200 2166.000 697.600 ;
        RECT 674.000 692.160 2166.000 696.200 ;
        RECT 674.400 690.760 2166.000 692.160 ;
        RECT 674.000 689.440 2166.000 690.760 ;
        RECT 674.000 688.040 2165.600 689.440 ;
        RECT 674.000 686.720 2166.000 688.040 ;
        RECT 674.400 685.320 2166.000 686.720 ;
        RECT 674.000 681.960 2166.000 685.320 ;
        RECT 674.400 680.560 2166.000 681.960 ;
        RECT 674.000 679.240 2166.000 680.560 ;
        RECT 674.000 677.840 2165.600 679.240 ;
        RECT 674.000 676.520 2166.000 677.840 ;
        RECT 674.400 675.120 2166.000 676.520 ;
        RECT 674.000 671.080 2166.000 675.120 ;
        RECT 674.400 669.680 2166.000 671.080 ;
        RECT 674.000 668.360 2166.000 669.680 ;
        RECT 674.000 666.960 2165.600 668.360 ;
        RECT 674.000 665.640 2166.000 666.960 ;
        RECT 674.400 664.240 2166.000 665.640 ;
        RECT 674.000 660.880 2166.000 664.240 ;
        RECT 674.400 659.480 2166.000 660.880 ;
        RECT 674.000 658.160 2166.000 659.480 ;
        RECT 674.000 656.760 2165.600 658.160 ;
        RECT 674.000 655.440 2166.000 656.760 ;
        RECT 674.400 654.040 2166.000 655.440 ;
        RECT 674.000 650.000 2166.000 654.040 ;
        RECT 674.400 648.600 2166.000 650.000 ;
        RECT 674.000 647.280 2166.000 648.600 ;
        RECT 674.000 645.880 2165.600 647.280 ;
        RECT 674.000 644.560 2166.000 645.880 ;
        RECT 674.400 643.160 2166.000 644.560 ;
        RECT 674.000 639.800 2166.000 643.160 ;
        RECT 674.400 638.400 2166.000 639.800 ;
        RECT 674.000 637.080 2166.000 638.400 ;
        RECT 674.000 635.680 2165.600 637.080 ;
        RECT 674.000 634.360 2166.000 635.680 ;
        RECT 674.400 632.960 2166.000 634.360 ;
        RECT 674.000 628.920 2166.000 632.960 ;
        RECT 674.400 627.520 2166.000 628.920 ;
        RECT 674.000 626.200 2166.000 627.520 ;
        RECT 674.000 624.800 2165.600 626.200 ;
        RECT 674.000 623.480 2166.000 624.800 ;
        RECT 674.400 622.080 2166.000 623.480 ;
        RECT 674.000 618.720 2166.000 622.080 ;
        RECT 674.400 617.320 2166.000 618.720 ;
        RECT 674.000 616.000 2166.000 617.320 ;
        RECT 674.000 614.600 2165.600 616.000 ;
        RECT 674.000 613.280 2166.000 614.600 ;
        RECT 674.400 611.880 2166.000 613.280 ;
        RECT 674.000 607.840 2166.000 611.880 ;
        RECT 674.400 606.440 2166.000 607.840 ;
        RECT 674.000 605.800 2166.000 606.440 ;
        RECT 674.000 604.400 2165.600 605.800 ;
        RECT 674.000 603.080 2166.000 604.400 ;
        RECT 674.400 602.215 2166.000 603.080 ;
      LAYER via3 ;
        RECT 998.500 2808.580 998.820 2808.900 ;
        RECT 992.980 2783.420 993.300 2783.740 ;
        RECT 992.060 2760.300 992.380 2760.620 ;
        RECT 991.140 2739.220 991.460 2739.540 ;
        RECT 990.220 2718.820 990.540 2719.140 ;
        RECT 989.300 2692.300 989.620 2692.620 ;
        RECT 1334.300 2051.740 1334.620 2052.060 ;
        RECT 1339.820 2051.060 1340.140 2051.380 ;
        RECT 1338.900 2050.380 1339.220 2050.700 ;
        RECT 1340.740 2049.700 1341.060 2050.020 ;
        RECT 1340.740 1693.380 1341.060 1693.700 ;
        RECT 989.300 1012.700 989.620 1013.020 ;
        RECT 991.140 1011.340 991.460 1011.660 ;
        RECT 1339.820 1010.660 1340.140 1010.980 ;
        RECT 998.500 1009.980 998.820 1010.300 ;
        RECT 992.060 1009.300 992.380 1009.620 ;
        RECT 992.980 1008.620 993.300 1008.940 ;
        RECT 990.220 1007.940 990.540 1008.260 ;
        RECT 1338.900 1007.940 1339.220 1008.260 ;
        RECT 1334.300 1007.260 1334.620 1007.580 ;
      LAYER met4 ;
        RECT 998.495 2808.575 998.825 2808.905 ;
        RECT 992.975 2783.415 993.305 2783.745 ;
        RECT 992.055 2760.295 992.385 2760.625 ;
      LAYER met4 ;
        RECT 459.645 2610.640 480.165 2747.120 ;
        RECT 482.565 2610.640 550.935 2747.120 ;
      LAYER met4 ;
        RECT 991.135 2739.215 991.465 2739.545 ;
        RECT 990.215 2718.815 990.545 2719.145 ;
        RECT 989.295 2692.295 989.625 2692.625 ;
      LAYER met4 ;
        RECT 531.415 1710.640 613.040 1969.520 ;
      LAYER met4 ;
        RECT 989.310 1013.025 989.610 2692.295 ;
        RECT 989.295 1012.695 989.625 1013.025 ;
        RECT 990.230 1008.265 990.530 2718.815 ;
        RECT 991.150 1011.665 991.450 2739.215 ;
        RECT 991.135 1011.335 991.465 1011.665 ;
        RECT 992.070 1009.625 992.370 2760.295 ;
        RECT 992.055 1009.295 992.385 1009.625 ;
        RECT 992.990 1008.945 993.290 2783.415 ;
        RECT 998.510 1010.305 998.810 2808.575 ;
      LAYER met4 ;
        RECT 1036.375 2610.640 1080.450 2787.920 ;
        RECT 1674.640 2510.640 1829.840 2889.200 ;
        RECT 2477.790 2610.640 2529.990 2760.720 ;
      LAYER met4 ;
        RECT 1334.295 2051.735 1334.625 2052.065 ;
      LAYER met4 ;
        RECT 1174.640 1710.640 1253.040 2032.080 ;
      LAYER met4 ;
        RECT 998.495 1009.975 998.825 1010.305 ;
        RECT 992.975 1008.615 993.305 1008.945 ;
        RECT 990.215 1007.935 990.545 1008.265 ;
        RECT 1334.310 1007.585 1334.610 2051.735 ;
        RECT 1339.815 2051.055 1340.145 2051.385 ;
        RECT 1338.895 2050.375 1339.225 2050.705 ;
        RECT 1338.910 1008.265 1339.210 2050.375 ;
        RECT 1339.830 1010.985 1340.130 2051.055 ;
        RECT 1340.735 2049.695 1341.065 2050.025 ;
        RECT 1340.750 1693.705 1341.050 2049.695 ;
      LAYER met4 ;
        RECT 1997.170 1760.640 2047.070 1905.280 ;
        RECT 2474.640 1710.640 2476.240 1926.000 ;
      LAYER met4 ;
        RECT 1340.735 1693.375 1341.065 1693.705 ;
        RECT 1339.815 1010.655 1340.145 1010.985 ;
        RECT 1338.895 1007.935 1339.225 1008.265 ;
        RECT 1334.295 1007.255 1334.625 1007.585 ;
      LAYER met4 ;
        RECT 718.135 989.600 2151.840 995.585 ;
        RECT 718.135 610.640 767.440 989.600 ;
        RECT 769.840 610.640 2151.840 989.600 ;
      LAYER met5 ;
        RECT 855.500 966.380 1861.740 983.300 ;
        RECT 855.500 948.380 1861.740 963.380 ;
        RECT 855.500 944.300 1861.740 945.380 ;
  END
END user_project_wrapper
END LIBRARY

