VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multi_project_harness
  CLASS BLOCK ;
  FOREIGN multi_project_harness ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 400.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 4.800 1500.000 5.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 104.760 1500.000 105.360 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 114.280 1500.000 114.880 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 124.480 1500.000 125.080 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 134.680 1500.000 135.280 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 144.200 1500.000 144.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 154.400 1500.000 155.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 164.600 1500.000 165.200 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 174.120 1500.000 174.720 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 184.320 1500.000 184.920 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 194.520 1500.000 195.120 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 14.320 1500.000 14.920 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 204.720 1500.000 205.320 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 214.240 1500.000 214.840 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 224.440 1500.000 225.040 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 234.640 1500.000 235.240 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 244.160 1500.000 244.760 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 254.360 1500.000 254.960 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 264.560 1500.000 265.160 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 274.080 1500.000 274.680 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 284.280 1500.000 284.880 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 294.480 1500.000 295.080 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 24.520 1500.000 25.120 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 304.680 1500.000 305.280 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 314.200 1500.000 314.800 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 324.400 1500.000 325.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 334.600 1500.000 335.200 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 344.120 1500.000 344.720 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 354.320 1500.000 354.920 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 364.520 1500.000 365.120 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 374.040 1500.000 374.640 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 34.720 1500.000 35.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 44.240 1500.000 44.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 54.440 1500.000 55.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 64.640 1500.000 65.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 74.160 1500.000 74.760 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 84.360 1500.000 84.960 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 94.560 1500.000 95.160 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1241.630 0.000 1241.910 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1250.830 0.000 1251.110 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1260.030 0.000 1260.310 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.230 0.000 1269.510 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1278.430 0.000 1278.710 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.630 0.000 1287.910 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1296.830 0.000 1297.110 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1305.570 0.000 1305.850 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1314.770 0.000 1315.050 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1323.970 0.000 1324.250 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1351.570 0.000 1351.850 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1360.770 0.000 1361.050 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1369.970 0.000 1370.250 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1379.170 0.000 1379.450 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1388.370 0.000 1388.650 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1397.570 0.000 1397.850 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1406.770 0.000 1407.050 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1415.970 0.000 1416.250 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1424.710 0.000 1424.990 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1433.910 0.000 1434.190 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1443.110 0.000 1443.390 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1452.310 0.000 1452.590 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1461.510 0.000 1461.790 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1470.710 0.000 1470.990 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1479.910 0.000 1480.190 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.110 0.000 1489.390 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.130 0.000 609.410 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.130 0.000 655.410 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 691.470 0.000 691.750 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 709.870 0.000 710.150 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 746.670 0.000 746.950 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 755.870 0.000 756.150 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.070 0.000 765.350 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 774.270 0.000 774.550 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 792.670 0.000 792.950 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.010 0.000 829.290 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 847.410 0.000 847.690 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 865.810 0.000 866.090 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 911.810 0.000 912.090 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.210 0.000 930.490 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.950 0.000 939.230 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.150 0.000 948.430 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 957.350 0.000 957.630 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 966.550 0.000 966.830 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 994.150 0.000 994.430 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.350 0.000 1003.630 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1012.550 0.000 1012.830 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1021.750 0.000 1022.030 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1030.950 0.000 1031.230 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1049.350 0.000 1049.630 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1067.290 0.000 1067.570 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1076.490 0.000 1076.770 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1085.690 0.000 1085.970 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1113.290 0.000 1113.570 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1122.490 0.000 1122.770 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.690 0.000 1131.970 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1140.890 0.000 1141.170 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.090 0.000 1150.370 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.490 0.000 1168.770 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1177.230 0.000 1177.510 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1186.430 0.000 1186.710 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.630 0.000 1195.910 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1204.830 0.000 1205.110 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1223.230 0.000 1223.510 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1232.430 0.000 1232.710 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1244.850 0.000 1245.130 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1254.050 0.000 1254.330 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1262.790 0.000 1263.070 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.190 0.000 1281.470 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1290.390 0.000 1290.670 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1299.590 0.000 1299.870 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1308.790 0.000 1309.070 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1317.990 0.000 1318.270 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1327.190 0.000 1327.470 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1336.390 0.000 1336.670 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1345.590 0.000 1345.870 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1354.790 0.000 1355.070 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1363.990 0.000 1364.270 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1373.190 0.000 1373.470 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1381.930 0.000 1382.210 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1400.330 0.000 1400.610 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1409.530 0.000 1409.810 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1418.730 0.000 1419.010 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1427.930 0.000 1428.210 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1437.130 0.000 1437.410 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1446.330 0.000 1446.610 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1464.730 0.000 1465.010 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1473.930 0.000 1474.210 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1483.130 0.000 1483.410 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1492.330 0.000 1492.610 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 694.690 0.000 694.970 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 713.090 0.000 713.370 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 823.030 0.000 823.310 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 832.230 0.000 832.510 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 841.430 0.000 841.710 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 850.630 0.000 850.910 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 869.030 0.000 869.310 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 878.230 0.000 878.510 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 887.430 0.000 887.710 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 896.170 0.000 896.450 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 905.370 0.000 905.650 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 923.770 0.000 924.050 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 932.970 0.000 933.250 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 951.370 0.000 951.650 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.570 0.000 960.850 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 969.770 0.000 970.050 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 988.170 0.000 988.450 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.370 0.000 997.650 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1006.570 0.000 1006.850 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1015.310 0.000 1015.590 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.510 0.000 1024.790 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1042.910 0.000 1043.190 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1052.110 0.000 1052.390 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1061.310 0.000 1061.590 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1070.510 0.000 1070.790 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1088.910 0.000 1089.190 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1107.310 0.000 1107.590 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1116.510 0.000 1116.790 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1134.910 0.000 1135.190 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1162.050 0.000 1162.330 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1171.250 0.000 1171.530 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1180.450 0.000 1180.730 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1189.650 0.000 1189.930 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1198.850 0.000 1199.130 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1208.050 0.000 1208.330 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1217.250 0.000 1217.530 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1226.450 0.000 1226.730 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1235.650 0.000 1235.930 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1247.610 0.000 1247.890 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1256.810 0.000 1257.090 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.210 0.000 1275.490 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1284.410 0.000 1284.690 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.610 0.000 1293.890 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1302.810 0.000 1303.090 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1312.010 0.000 1312.290 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1321.210 0.000 1321.490 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1330.410 0.000 1330.690 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1339.150 0.000 1339.430 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1357.550 0.000 1357.830 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1366.750 0.000 1367.030 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1375.950 0.000 1376.230 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1403.550 0.000 1403.830 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.750 0.000 1413.030 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1421.950 0.000 1422.230 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1431.150 0.000 1431.430 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1440.350 0.000 1440.630 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1449.550 0.000 1449.830 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1458.750 0.000 1459.030 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1467.490 0.000 1467.770 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1476.690 0.000 1476.970 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1485.890 0.000 1486.170 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1495.090 0.000 1495.370 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 459.630 0.000 459.910 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 541.970 0.000 542.250 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.170 0.000 597.450 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 624.310 0.000 624.590 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 725.510 0.000 725.790 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 743.450 0.000 743.730 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 761.850 0.000 762.130 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 835.450 0.000 835.730 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 908.590 0.000 908.870 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 926.990 0.000 927.270 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.190 0.000 936.470 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 954.590 0.000 954.870 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 963.790 0.000 964.070 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 972.990 0.000 973.270 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 981.730 0.000 982.010 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 990.930 0.000 991.210 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1000.130 0.000 1000.410 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.530 0.000 1018.810 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1027.730 0.000 1028.010 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.930 0.000 1037.210 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.330 0.000 1055.610 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.730 0.000 1074.010 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1082.930 0.000 1083.210 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.130 0.000 1092.410 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1100.870 0.000 1101.150 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.070 0.000 1110.350 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1119.270 0.000 1119.550 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1128.470 0.000 1128.750 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1137.670 0.000 1137.950 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1146.870 0.000 1147.150 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1165.270 0.000 1165.550 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1174.470 0.000 1174.750 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1183.670 0.000 1183.950 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1192.870 0.000 1193.150 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1202.070 0.000 1202.350 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1211.270 0.000 1211.550 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1220.010 0.000 1220.290 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1229.210 0.000 1229.490 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1238.410 0.000 1238.690 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END la_oen[9]
  PIN proj0_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.130 396.000 172.410 400.000 ;
    END
  END proj0_clk
  PIN proj0_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 178.570 396.000 178.850 400.000 ;
    END
  END proj0_io_in[0]
  PIN proj0_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 221.810 396.000 222.090 400.000 ;
    END
  END proj0_io_in[10]
  PIN proj0_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 226.410 396.000 226.690 400.000 ;
    END
  END proj0_io_in[11]
  PIN proj0_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 230.550 396.000 230.830 400.000 ;
    END
  END proj0_io_in[12]
  PIN proj0_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.690 396.000 234.970 400.000 ;
    END
  END proj0_io_in[13]
  PIN proj0_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 239.290 396.000 239.570 400.000 ;
    END
  END proj0_io_in[14]
  PIN proj0_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.430 396.000 243.710 400.000 ;
    END
  END proj0_io_in[15]
  PIN proj0_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.030 396.000 248.310 400.000 ;
    END
  END proj0_io_in[16]
  PIN proj0_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.170 396.000 252.450 400.000 ;
    END
  END proj0_io_in[17]
  PIN proj0_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 256.770 396.000 257.050 400.000 ;
    END
  END proj0_io_in[18]
  PIN proj0_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 260.910 396.000 261.190 400.000 ;
    END
  END proj0_io_in[19]
  PIN proj0_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 182.710 396.000 182.990 400.000 ;
    END
  END proj0_io_in[1]
  PIN proj0_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 265.050 396.000 265.330 400.000 ;
    END
  END proj0_io_in[20]
  PIN proj0_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.650 396.000 269.930 400.000 ;
    END
  END proj0_io_in[21]
  PIN proj0_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.790 396.000 274.070 400.000 ;
    END
  END proj0_io_in[22]
  PIN proj0_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 278.390 396.000 278.670 400.000 ;
    END
  END proj0_io_in[23]
  PIN proj0_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 282.530 396.000 282.810 400.000 ;
    END
  END proj0_io_in[24]
  PIN proj0_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.130 396.000 287.410 400.000 ;
    END
  END proj0_io_in[25]
  PIN proj0_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.270 396.000 291.550 400.000 ;
    END
  END proj0_io_in[26]
  PIN proj0_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.410 396.000 295.690 400.000 ;
    END
  END proj0_io_in[27]
  PIN proj0_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.010 396.000 300.290 400.000 ;
    END
  END proj0_io_in[28]
  PIN proj0_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 304.150 396.000 304.430 400.000 ;
    END
  END proj0_io_in[29]
  PIN proj0_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 187.310 396.000 187.590 400.000 ;
    END
  END proj0_io_in[2]
  PIN proj0_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 308.750 396.000 309.030 400.000 ;
    END
  END proj0_io_in[30]
  PIN proj0_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 312.890 396.000 313.170 400.000 ;
    END
  END proj0_io_in[31]
  PIN proj0_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 317.490 396.000 317.770 400.000 ;
    END
  END proj0_io_in[32]
  PIN proj0_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.630 396.000 321.910 400.000 ;
    END
  END proj0_io_in[33]
  PIN proj0_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.770 396.000 326.050 400.000 ;
    END
  END proj0_io_in[34]
  PIN proj0_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 330.370 396.000 330.650 400.000 ;
    END
  END proj0_io_in[35]
  PIN proj0_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 334.510 396.000 334.790 400.000 ;
    END
  END proj0_io_in[36]
  PIN proj0_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 339.110 396.000 339.390 400.000 ;
    END
  END proj0_io_in[37]
  PIN proj0_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.450 396.000 191.730 400.000 ;
    END
  END proj0_io_in[3]
  PIN proj0_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.050 396.000 196.330 400.000 ;
    END
  END proj0_io_in[4]
  PIN proj0_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 200.190 396.000 200.470 400.000 ;
    END
  END proj0_io_in[5]
  PIN proj0_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 204.330 396.000 204.610 400.000 ;
    END
  END proj0_io_in[6]
  PIN proj0_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.930 396.000 209.210 400.000 ;
    END
  END proj0_io_in[7]
  PIN proj0_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.070 396.000 213.350 400.000 ;
    END
  END proj0_io_in[8]
  PIN proj0_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 217.670 396.000 217.950 400.000 ;
    END
  END proj0_io_in[9]
  PIN proj0_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.870 396.000 181.150 400.000 ;
    END
  END proj0_io_out[0]
  PIN proj0_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.110 396.000 224.390 400.000 ;
    END
  END proj0_io_out[10]
  PIN proj0_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.250 396.000 228.530 400.000 ;
    END
  END proj0_io_out[11]
  PIN proj0_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.850 396.000 233.130 400.000 ;
    END
  END proj0_io_out[12]
  PIN proj0_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.990 396.000 237.270 400.000 ;
    END
  END proj0_io_out[13]
  PIN proj0_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.590 396.000 241.870 400.000 ;
    END
  END proj0_io_out[14]
  PIN proj0_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 245.730 396.000 246.010 400.000 ;
    END
  END proj0_io_out[15]
  PIN proj0_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 249.870 396.000 250.150 400.000 ;
    END
  END proj0_io_out[16]
  PIN proj0_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.470 396.000 254.750 400.000 ;
    END
  END proj0_io_out[17]
  PIN proj0_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.610 396.000 258.890 400.000 ;
    END
  END proj0_io_out[18]
  PIN proj0_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.210 396.000 263.490 400.000 ;
    END
  END proj0_io_out[19]
  PIN proj0_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.010 396.000 185.290 400.000 ;
    END
  END proj0_io_out[1]
  PIN proj0_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 267.350 396.000 267.630 400.000 ;
    END
  END proj0_io_out[20]
  PIN proj0_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.950 396.000 272.230 400.000 ;
    END
  END proj0_io_out[21]
  PIN proj0_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.090 396.000 276.370 400.000 ;
    END
  END proj0_io_out[22]
  PIN proj0_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 280.230 396.000 280.510 400.000 ;
    END
  END proj0_io_out[23]
  PIN proj0_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 284.830 396.000 285.110 400.000 ;
    END
  END proj0_io_out[24]
  PIN proj0_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.970 396.000 289.250 400.000 ;
    END
  END proj0_io_out[25]
  PIN proj0_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.570 396.000 293.850 400.000 ;
    END
  END proj0_io_out[26]
  PIN proj0_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 297.710 396.000 297.990 400.000 ;
    END
  END proj0_io_out[27]
  PIN proj0_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.310 396.000 302.590 400.000 ;
    END
  END proj0_io_out[28]
  PIN proj0_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 306.450 396.000 306.730 400.000 ;
    END
  END proj0_io_out[29]
  PIN proj0_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.150 396.000 189.430 400.000 ;
    END
  END proj0_io_out[2]
  PIN proj0_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.590 396.000 310.870 400.000 ;
    END
  END proj0_io_out[30]
  PIN proj0_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.190 396.000 315.470 400.000 ;
    END
  END proj0_io_out[31]
  PIN proj0_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.330 396.000 319.610 400.000 ;
    END
  END proj0_io_out[32]
  PIN proj0_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 396.000 324.210 400.000 ;
    END
  END proj0_io_out[33]
  PIN proj0_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 328.070 396.000 328.350 400.000 ;
    END
  END proj0_io_out[34]
  PIN proj0_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 332.670 396.000 332.950 400.000 ;
    END
  END proj0_io_out[35]
  PIN proj0_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 336.810 396.000 337.090 400.000 ;
    END
  END proj0_io_out[36]
  PIN proj0_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.950 396.000 341.230 400.000 ;
    END
  END proj0_io_out[37]
  PIN proj0_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.750 396.000 194.030 400.000 ;
    END
  END proj0_io_out[3]
  PIN proj0_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.890 396.000 198.170 400.000 ;
    END
  END proj0_io_out[4]
  PIN proj0_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.490 396.000 202.770 400.000 ;
    END
  END proj0_io_out[5]
  PIN proj0_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.630 396.000 206.910 400.000 ;
    END
  END proj0_io_out[6]
  PIN proj0_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.230 396.000 211.510 400.000 ;
    END
  END proj0_io_out[7]
  PIN proj0_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.370 396.000 215.650 400.000 ;
    END
  END proj0_io_out[8]
  PIN proj0_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.510 396.000 219.790 400.000 ;
    END
  END proj0_io_out[9]
  PIN proj0_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.970 396.000 174.250 400.000 ;
    END
  END proj0_reset
  PIN proj0_wb_update
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.270 396.000 176.550 400.000 ;
    END
  END proj0_wb_update
  PIN proj1_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.010 396.000 1.290 400.000 ;
    END
  END proj1_clk
  PIN proj1_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 396.000 7.730 400.000 ;
    END
  END proj1_io_in[0]
  PIN proj1_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.690 396.000 50.970 400.000 ;
    END
  END proj1_io_in[10]
  PIN proj1_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.830 396.000 55.110 400.000 ;
    END
  END proj1_io_in[11]
  PIN proj1_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 396.000 59.710 400.000 ;
    END
  END proj1_io_in[12]
  PIN proj1_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 396.000 63.850 400.000 ;
    END
  END proj1_io_in[13]
  PIN proj1_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 396.000 68.450 400.000 ;
    END
  END proj1_io_in[14]
  PIN proj1_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.310 396.000 72.590 400.000 ;
    END
  END proj1_io_in[15]
  PIN proj1_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 396.000 76.730 400.000 ;
    END
  END proj1_io_in[16]
  PIN proj1_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 396.000 81.330 400.000 ;
    END
  END proj1_io_in[17]
  PIN proj1_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 396.000 85.470 400.000 ;
    END
  END proj1_io_in[18]
  PIN proj1_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 396.000 90.070 400.000 ;
    END
  END proj1_io_in[19]
  PIN proj1_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.590 396.000 11.870 400.000 ;
    END
  END proj1_io_in[1]
  PIN proj1_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 396.000 94.210 400.000 ;
    END
  END proj1_io_in[20]
  PIN proj1_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 396.000 98.810 400.000 ;
    END
  END proj1_io_in[21]
  PIN proj1_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.670 396.000 102.950 400.000 ;
    END
  END proj1_io_in[22]
  PIN proj1_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 396.000 107.090 400.000 ;
    END
  END proj1_io_in[23]
  PIN proj1_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.410 396.000 111.690 400.000 ;
    END
  END proj1_io_in[24]
  PIN proj1_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.550 396.000 115.830 400.000 ;
    END
  END proj1_io_in[25]
  PIN proj1_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.150 396.000 120.430 400.000 ;
    END
  END proj1_io_in[26]
  PIN proj1_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.290 396.000 124.570 400.000 ;
    END
  END proj1_io_in[27]
  PIN proj1_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.890 396.000 129.170 400.000 ;
    END
  END proj1_io_in[28]
  PIN proj1_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.030 396.000 133.310 400.000 ;
    END
  END proj1_io_in[29]
  PIN proj1_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 396.000 16.010 400.000 ;
    END
  END proj1_io_in[2]
  PIN proj1_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 396.000 137.450 400.000 ;
    END
  END proj1_io_in[30]
  PIN proj1_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.770 396.000 142.050 400.000 ;
    END
  END proj1_io_in[31]
  PIN proj1_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.910 396.000 146.190 400.000 ;
    END
  END proj1_io_in[32]
  PIN proj1_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.510 396.000 150.790 400.000 ;
    END
  END proj1_io_in[33]
  PIN proj1_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.650 396.000 154.930 400.000 ;
    END
  END proj1_io_in[34]
  PIN proj1_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 159.250 396.000 159.530 400.000 ;
    END
  END proj1_io_in[35]
  PIN proj1_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.390 396.000 163.670 400.000 ;
    END
  END proj1_io_in[36]
  PIN proj1_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.530 396.000 167.810 400.000 ;
    END
  END proj1_io_in[37]
  PIN proj1_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.330 396.000 20.610 400.000 ;
    END
  END proj1_io_in[3]
  PIN proj1_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.470 396.000 24.750 400.000 ;
    END
  END proj1_io_in[4]
  PIN proj1_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 396.000 29.350 400.000 ;
    END
  END proj1_io_in[5]
  PIN proj1_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.210 396.000 33.490 400.000 ;
    END
  END proj1_io_in[6]
  PIN proj1_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 396.000 38.090 400.000 ;
    END
  END proj1_io_in[7]
  PIN proj1_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 396.000 42.230 400.000 ;
    END
  END proj1_io_in[8]
  PIN proj1_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 396.000 46.370 400.000 ;
    END
  END proj1_io_in[9]
  PIN proj1_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 396.000 9.570 400.000 ;
    END
  END proj1_io_out[0]
  PIN proj1_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 396.000 53.270 400.000 ;
    END
  END proj1_io_out[10]
  PIN proj1_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 396.000 57.410 400.000 ;
    END
  END proj1_io_out[11]
  PIN proj1_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 396.000 61.550 400.000 ;
    END
  END proj1_io_out[12]
  PIN proj1_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 396.000 66.150 400.000 ;
    END
  END proj1_io_out[13]
  PIN proj1_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 396.000 70.290 400.000 ;
    END
  END proj1_io_out[14]
  PIN proj1_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 396.000 74.890 400.000 ;
    END
  END proj1_io_out[15]
  PIN proj1_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 396.000 79.030 400.000 ;
    END
  END proj1_io_out[16]
  PIN proj1_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.350 396.000 83.630 400.000 ;
    END
  END proj1_io_out[17]
  PIN proj1_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.490 396.000 87.770 400.000 ;
    END
  END proj1_io_out[18]
  PIN proj1_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 396.000 91.910 400.000 ;
    END
  END proj1_io_out[19]
  PIN proj1_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 396.000 14.170 400.000 ;
    END
  END proj1_io_out[1]
  PIN proj1_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.230 396.000 96.510 400.000 ;
    END
  END proj1_io_out[20]
  PIN proj1_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 396.000 100.650 400.000 ;
    END
  END proj1_io_out[21]
  PIN proj1_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 396.000 105.250 400.000 ;
    END
  END proj1_io_out[22]
  PIN proj1_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.110 396.000 109.390 400.000 ;
    END
  END proj1_io_out[23]
  PIN proj1_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 396.000 113.990 400.000 ;
    END
  END proj1_io_out[24]
  PIN proj1_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 396.000 118.130 400.000 ;
    END
  END proj1_io_out[25]
  PIN proj1_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 396.000 122.270 400.000 ;
    END
  END proj1_io_out[26]
  PIN proj1_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.590 396.000 126.870 400.000 ;
    END
  END proj1_io_out[27]
  PIN proj1_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.730 396.000 131.010 400.000 ;
    END
  END proj1_io_out[28]
  PIN proj1_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.330 396.000 135.610 400.000 ;
    END
  END proj1_io_out[29]
  PIN proj1_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 396.000 18.310 400.000 ;
    END
  END proj1_io_out[2]
  PIN proj1_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.470 396.000 139.750 400.000 ;
    END
  END proj1_io_out[30]
  PIN proj1_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.070 396.000 144.350 400.000 ;
    END
  END proj1_io_out[31]
  PIN proj1_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.210 396.000 148.490 400.000 ;
    END
  END proj1_io_out[32]
  PIN proj1_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.350 396.000 152.630 400.000 ;
    END
  END proj1_io_out[33]
  PIN proj1_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.950 396.000 157.230 400.000 ;
    END
  END proj1_io_out[34]
  PIN proj1_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.090 396.000 161.370 400.000 ;
    END
  END proj1_io_out[35]
  PIN proj1_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.690 396.000 165.970 400.000 ;
    END
  END proj1_io_out[36]
  PIN proj1_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.830 396.000 170.110 400.000 ;
    END
  END proj1_io_out[37]
  PIN proj1_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 396.000 22.910 400.000 ;
    END
  END proj1_io_out[3]
  PIN proj1_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 396.000 27.050 400.000 ;
    END
  END proj1_io_out[4]
  PIN proj1_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 396.000 31.190 400.000 ;
    END
  END proj1_io_out[5]
  PIN proj1_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 396.000 35.790 400.000 ;
    END
  END proj1_io_out[6]
  PIN proj1_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 396.000 39.930 400.000 ;
    END
  END proj1_io_out[7]
  PIN proj1_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 396.000 44.530 400.000 ;
    END
  END proj1_io_out[8]
  PIN proj1_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 396.000 48.670 400.000 ;
    END
  END proj1_io_out[9]
  PIN proj1_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 396.000 3.130 400.000 ;
    END
  END proj1_reset
  PIN proj1_wb_update
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.150 396.000 5.430 400.000 ;
    END
  END proj1_wb_update
  PIN proj2_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1327.650 396.000 1327.930 400.000 ;
    END
  END proj2_clk
  PIN proj2_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1331.790 396.000 1332.070 400.000 ;
    END
  END proj2_io_in[0]
  PIN proj2_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.030 396.000 1375.310 400.000 ;
    END
  END proj2_io_in[10]
  PIN proj2_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1379.630 396.000 1379.910 400.000 ;
    END
  END proj2_io_in[11]
  PIN proj2_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1383.770 396.000 1384.050 400.000 ;
    END
  END proj2_io_in[12]
  PIN proj2_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1387.910 396.000 1388.190 400.000 ;
    END
  END proj2_io_in[13]
  PIN proj2_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1392.510 396.000 1392.790 400.000 ;
    END
  END proj2_io_in[14]
  PIN proj2_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1396.650 396.000 1396.930 400.000 ;
    END
  END proj2_io_in[15]
  PIN proj2_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1401.250 396.000 1401.530 400.000 ;
    END
  END proj2_io_in[16]
  PIN proj2_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1405.390 396.000 1405.670 400.000 ;
    END
  END proj2_io_in[17]
  PIN proj2_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1409.990 396.000 1410.270 400.000 ;
    END
  END proj2_io_in[18]
  PIN proj2_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1414.130 396.000 1414.410 400.000 ;
    END
  END proj2_io_in[19]
  PIN proj2_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1335.930 396.000 1336.210 400.000 ;
    END
  END proj2_io_in[1]
  PIN proj2_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1418.270 396.000 1418.550 400.000 ;
    END
  END proj2_io_in[20]
  PIN proj2_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1422.870 396.000 1423.150 400.000 ;
    END
  END proj2_io_in[21]
  PIN proj2_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1427.010 396.000 1427.290 400.000 ;
    END
  END proj2_io_in[22]
  PIN proj2_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1431.610 396.000 1431.890 400.000 ;
    END
  END proj2_io_in[23]
  PIN proj2_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1435.750 396.000 1436.030 400.000 ;
    END
  END proj2_io_in[24]
  PIN proj2_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1440.350 396.000 1440.630 400.000 ;
    END
  END proj2_io_in[25]
  PIN proj2_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1444.490 396.000 1444.770 400.000 ;
    END
  END proj2_io_in[26]
  PIN proj2_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1448.630 396.000 1448.910 400.000 ;
    END
  END proj2_io_in[27]
  PIN proj2_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1453.230 396.000 1453.510 400.000 ;
    END
  END proj2_io_in[28]
  PIN proj2_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1457.370 396.000 1457.650 400.000 ;
    END
  END proj2_io_in[29]
  PIN proj2_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1340.530 396.000 1340.810 400.000 ;
    END
  END proj2_io_in[2]
  PIN proj2_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1461.970 396.000 1462.250 400.000 ;
    END
  END proj2_io_in[30]
  PIN proj2_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1466.110 396.000 1466.390 400.000 ;
    END
  END proj2_io_in[31]
  PIN proj2_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1470.710 396.000 1470.990 400.000 ;
    END
  END proj2_io_in[32]
  PIN proj2_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1474.850 396.000 1475.130 400.000 ;
    END
  END proj2_io_in[33]
  PIN proj2_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1478.990 396.000 1479.270 400.000 ;
    END
  END proj2_io_in[34]
  PIN proj2_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1483.590 396.000 1483.870 400.000 ;
    END
  END proj2_io_in[35]
  PIN proj2_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1487.730 396.000 1488.010 400.000 ;
    END
  END proj2_io_in[36]
  PIN proj2_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1492.330 396.000 1492.610 400.000 ;
    END
  END proj2_io_in[37]
  PIN proj2_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1344.670 396.000 1344.950 400.000 ;
    END
  END proj2_io_in[3]
  PIN proj2_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1349.270 396.000 1349.550 400.000 ;
    END
  END proj2_io_in[4]
  PIN proj2_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1353.410 396.000 1353.690 400.000 ;
    END
  END proj2_io_in[5]
  PIN proj2_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1357.550 396.000 1357.830 400.000 ;
    END
  END proj2_io_in[6]
  PIN proj2_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1362.150 396.000 1362.430 400.000 ;
    END
  END proj2_io_in[7]
  PIN proj2_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1366.290 396.000 1366.570 400.000 ;
    END
  END proj2_io_in[8]
  PIN proj2_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.890 396.000 1371.170 400.000 ;
    END
  END proj2_io_in[9]
  PIN proj2_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1334.090 396.000 1334.370 400.000 ;
    END
  END proj2_io_out[0]
  PIN proj2_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1377.330 396.000 1377.610 400.000 ;
    END
  END proj2_io_out[10]
  PIN proj2_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1381.470 396.000 1381.750 400.000 ;
    END
  END proj2_io_out[11]
  PIN proj2_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1386.070 396.000 1386.350 400.000 ;
    END
  END proj2_io_out[12]
  PIN proj2_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1390.210 396.000 1390.490 400.000 ;
    END
  END proj2_io_out[13]
  PIN proj2_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.810 396.000 1395.090 400.000 ;
    END
  END proj2_io_out[14]
  PIN proj2_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1398.950 396.000 1399.230 400.000 ;
    END
  END proj2_io_out[15]
  PIN proj2_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1403.090 396.000 1403.370 400.000 ;
    END
  END proj2_io_out[16]
  PIN proj2_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1407.690 396.000 1407.970 400.000 ;
    END
  END proj2_io_out[17]
  PIN proj2_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1411.830 396.000 1412.110 400.000 ;
    END
  END proj2_io_out[18]
  PIN proj2_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1416.430 396.000 1416.710 400.000 ;
    END
  END proj2_io_out[19]
  PIN proj2_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1338.230 396.000 1338.510 400.000 ;
    END
  END proj2_io_out[1]
  PIN proj2_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1420.570 396.000 1420.850 400.000 ;
    END
  END proj2_io_out[20]
  PIN proj2_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1425.170 396.000 1425.450 400.000 ;
    END
  END proj2_io_out[21]
  PIN proj2_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.310 396.000 1429.590 400.000 ;
    END
  END proj2_io_out[22]
  PIN proj2_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1433.450 396.000 1433.730 400.000 ;
    END
  END proj2_io_out[23]
  PIN proj2_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1438.050 396.000 1438.330 400.000 ;
    END
  END proj2_io_out[24]
  PIN proj2_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1442.190 396.000 1442.470 400.000 ;
    END
  END proj2_io_out[25]
  PIN proj2_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1446.790 396.000 1447.070 400.000 ;
    END
  END proj2_io_out[26]
  PIN proj2_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1450.930 396.000 1451.210 400.000 ;
    END
  END proj2_io_out[27]
  PIN proj2_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.530 396.000 1455.810 400.000 ;
    END
  END proj2_io_out[28]
  PIN proj2_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1459.670 396.000 1459.950 400.000 ;
    END
  END proj2_io_out[29]
  PIN proj2_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1342.370 396.000 1342.650 400.000 ;
    END
  END proj2_io_out[2]
  PIN proj2_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1463.810 396.000 1464.090 400.000 ;
    END
  END proj2_io_out[30]
  PIN proj2_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1468.410 396.000 1468.690 400.000 ;
    END
  END proj2_io_out[31]
  PIN proj2_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1472.550 396.000 1472.830 400.000 ;
    END
  END proj2_io_out[32]
  PIN proj2_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1477.150 396.000 1477.430 400.000 ;
    END
  END proj2_io_out[33]
  PIN proj2_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1481.290 396.000 1481.570 400.000 ;
    END
  END proj2_io_out[34]
  PIN proj2_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1485.890 396.000 1486.170 400.000 ;
    END
  END proj2_io_out[35]
  PIN proj2_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1490.030 396.000 1490.310 400.000 ;
    END
  END proj2_io_out[36]
  PIN proj2_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1494.170 396.000 1494.450 400.000 ;
    END
  END proj2_io_out[37]
  PIN proj2_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.970 396.000 1347.250 400.000 ;
    END
  END proj2_io_out[3]
  PIN proj2_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1351.110 396.000 1351.390 400.000 ;
    END
  END proj2_io_out[4]
  PIN proj2_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1355.710 396.000 1355.990 400.000 ;
    END
  END proj2_io_out[5]
  PIN proj2_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1359.850 396.000 1360.130 400.000 ;
    END
  END proj2_io_out[6]
  PIN proj2_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.450 396.000 1364.730 400.000 ;
    END
  END proj2_io_out[7]
  PIN proj2_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1368.590 396.000 1368.870 400.000 ;
    END
  END proj2_io_out[8]
  PIN proj2_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1372.730 396.000 1373.010 400.000 ;
    END
  END proj2_io_out[9]
  PIN proj2_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1329.490 396.000 1329.770 400.000 ;
    END
  END proj2_reset
  PIN proj3_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 510.230 396.000 510.510 400.000 ;
    END
  END proj3_clk
  PIN proj3_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 514.370 396.000 514.650 400.000 ;
    END
  END proj3_io_in[0]
  PIN proj3_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.070 396.000 558.350 400.000 ;
    END
  END proj3_io_in[10]
  PIN proj3_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 562.210 396.000 562.490 400.000 ;
    END
  END proj3_io_in[11]
  PIN proj3_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 566.350 396.000 566.630 400.000 ;
    END
  END proj3_io_in[12]
  PIN proj3_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.950 396.000 571.230 400.000 ;
    END
  END proj3_io_in[13]
  PIN proj3_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 575.090 396.000 575.370 400.000 ;
    END
  END proj3_io_in[14]
  PIN proj3_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 579.690 396.000 579.970 400.000 ;
    END
  END proj3_io_in[15]
  PIN proj3_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 583.830 396.000 584.110 400.000 ;
    END
  END proj3_io_in[16]
  PIN proj3_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 588.430 396.000 588.710 400.000 ;
    END
  END proj3_io_in[17]
  PIN proj3_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 592.570 396.000 592.850 400.000 ;
    END
  END proj3_io_in[18]
  PIN proj3_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 596.710 396.000 596.990 400.000 ;
    END
  END proj3_io_in[19]
  PIN proj3_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 518.970 396.000 519.250 400.000 ;
    END
  END proj3_io_in[1]
  PIN proj3_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 601.310 396.000 601.590 400.000 ;
    END
  END proj3_io_in[20]
  PIN proj3_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 605.450 396.000 605.730 400.000 ;
    END
  END proj3_io_in[21]
  PIN proj3_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.050 396.000 610.330 400.000 ;
    END
  END proj3_io_in[22]
  PIN proj3_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 614.190 396.000 614.470 400.000 ;
    END
  END proj3_io_in[23]
  PIN proj3_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 618.790 396.000 619.070 400.000 ;
    END
  END proj3_io_in[24]
  PIN proj3_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 622.930 396.000 623.210 400.000 ;
    END
  END proj3_io_in[25]
  PIN proj3_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.070 396.000 627.350 400.000 ;
    END
  END proj3_io_in[26]
  PIN proj3_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 631.670 396.000 631.950 400.000 ;
    END
  END proj3_io_in[27]
  PIN proj3_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 635.810 396.000 636.090 400.000 ;
    END
  END proj3_io_in[28]
  PIN proj3_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 640.410 396.000 640.690 400.000 ;
    END
  END proj3_io_in[29]
  PIN proj3_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 523.110 396.000 523.390 400.000 ;
    END
  END proj3_io_in[2]
  PIN proj3_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.550 396.000 644.830 400.000 ;
    END
  END proj3_io_in[30]
  PIN proj3_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 649.150 396.000 649.430 400.000 ;
    END
  END proj3_io_in[31]
  PIN proj3_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 653.290 396.000 653.570 400.000 ;
    END
  END proj3_io_in[32]
  PIN proj3_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 657.430 396.000 657.710 400.000 ;
    END
  END proj3_io_in[33]
  PIN proj3_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 662.030 396.000 662.310 400.000 ;
    END
  END proj3_io_in[34]
  PIN proj3_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 666.170 396.000 666.450 400.000 ;
    END
  END proj3_io_in[35]
  PIN proj3_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 670.770 396.000 671.050 400.000 ;
    END
  END proj3_io_in[36]
  PIN proj3_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.910 396.000 675.190 400.000 ;
    END
  END proj3_io_in[37]
  PIN proj3_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 527.710 396.000 527.990 400.000 ;
    END
  END proj3_io_in[3]
  PIN proj3_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 531.850 396.000 532.130 400.000 ;
    END
  END proj3_io_in[4]
  PIN proj3_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 535.990 396.000 536.270 400.000 ;
    END
  END proj3_io_in[5]
  PIN proj3_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 540.590 396.000 540.870 400.000 ;
    END
  END proj3_io_in[6]
  PIN proj3_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 544.730 396.000 545.010 400.000 ;
    END
  END proj3_io_in[7]
  PIN proj3_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 549.330 396.000 549.610 400.000 ;
    END
  END proj3_io_in[8]
  PIN proj3_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 553.470 396.000 553.750 400.000 ;
    END
  END proj3_io_in[9]
  PIN proj3_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 516.670 396.000 516.950 400.000 ;
    END
  END proj3_io_out[0]
  PIN proj3_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 559.910 396.000 560.190 400.000 ;
    END
  END proj3_io_out[10]
  PIN proj3_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 564.510 396.000 564.790 400.000 ;
    END
  END proj3_io_out[11]
  PIN proj3_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 568.650 396.000 568.930 400.000 ;
    END
  END proj3_io_out[12]
  PIN proj3_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 573.250 396.000 573.530 400.000 ;
    END
  END proj3_io_out[13]
  PIN proj3_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 577.390 396.000 577.670 400.000 ;
    END
  END proj3_io_out[14]
  PIN proj3_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.530 396.000 581.810 400.000 ;
    END
  END proj3_io_out[15]
  PIN proj3_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.130 396.000 586.410 400.000 ;
    END
  END proj3_io_out[16]
  PIN proj3_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 590.270 396.000 590.550 400.000 ;
    END
  END proj3_io_out[17]
  PIN proj3_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 594.870 396.000 595.150 400.000 ;
    END
  END proj3_io_out[18]
  PIN proj3_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 599.010 396.000 599.290 400.000 ;
    END
  END proj3_io_out[19]
  PIN proj3_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 520.810 396.000 521.090 400.000 ;
    END
  END proj3_io_out[1]
  PIN proj3_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.610 396.000 603.890 400.000 ;
    END
  END proj3_io_out[20]
  PIN proj3_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 607.750 396.000 608.030 400.000 ;
    END
  END proj3_io_out[21]
  PIN proj3_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 611.890 396.000 612.170 400.000 ;
    END
  END proj3_io_out[22]
  PIN proj3_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.490 396.000 616.770 400.000 ;
    END
  END proj3_io_out[23]
  PIN proj3_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.630 396.000 620.910 400.000 ;
    END
  END proj3_io_out[24]
  PIN proj3_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 625.230 396.000 625.510 400.000 ;
    END
  END proj3_io_out[25]
  PIN proj3_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 629.370 396.000 629.650 400.000 ;
    END
  END proj3_io_out[26]
  PIN proj3_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 633.970 396.000 634.250 400.000 ;
    END
  END proj3_io_out[27]
  PIN proj3_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 638.110 396.000 638.390 400.000 ;
    END
  END proj3_io_out[28]
  PIN proj3_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 642.250 396.000 642.530 400.000 ;
    END
  END proj3_io_out[29]
  PIN proj3_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.410 396.000 525.690 400.000 ;
    END
  END proj3_io_out[2]
  PIN proj3_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 646.850 396.000 647.130 400.000 ;
    END
  END proj3_io_out[30]
  PIN proj3_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.990 396.000 651.270 400.000 ;
    END
  END proj3_io_out[31]
  PIN proj3_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.590 396.000 655.870 400.000 ;
    END
  END proj3_io_out[32]
  PIN proj3_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 659.730 396.000 660.010 400.000 ;
    END
  END proj3_io_out[33]
  PIN proj3_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 664.330 396.000 664.610 400.000 ;
    END
  END proj3_io_out[34]
  PIN proj3_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.470 396.000 668.750 400.000 ;
    END
  END proj3_io_out[35]
  PIN proj3_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 672.610 396.000 672.890 400.000 ;
    END
  END proj3_io_out[36]
  PIN proj3_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 677.210 396.000 677.490 400.000 ;
    END
  END proj3_io_out[37]
  PIN proj3_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 529.550 396.000 529.830 400.000 ;
    END
  END proj3_io_out[3]
  PIN proj3_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 534.150 396.000 534.430 400.000 ;
    END
  END proj3_io_out[4]
  PIN proj3_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 538.290 396.000 538.570 400.000 ;
    END
  END proj3_io_out[5]
  PIN proj3_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 542.890 396.000 543.170 400.000 ;
    END
  END proj3_io_out[6]
  PIN proj3_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 547.030 396.000 547.310 400.000 ;
    END
  END proj3_io_out[7]
  PIN proj3_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 551.170 396.000 551.450 400.000 ;
    END
  END proj3_io_out[8]
  PIN proj3_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 555.770 396.000 556.050 400.000 ;
    END
  END proj3_io_out[9]
  PIN proj3_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 512.530 396.000 512.810 400.000 ;
    END
  END proj3_reset
  PIN proj4_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 679.050 396.000 679.330 400.000 ;
    END
  END proj4_clk
  PIN proj4_cnt[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 685.950 396.000 686.230 400.000 ;
    END
  END proj4_cnt[0]
  PIN proj4_cnt[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 772.430 396.000 772.710 400.000 ;
    END
  END proj4_cnt[10]
  PIN proj4_cnt[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.170 396.000 781.450 400.000 ;
    END
  END proj4_cnt[11]
  PIN proj4_cnt[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.910 396.000 790.190 400.000 ;
    END
  END proj4_cnt[12]
  PIN proj4_cnt[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 798.650 396.000 798.930 400.000 ;
    END
  END proj4_cnt[13]
  PIN proj4_cnt[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.390 396.000 807.670 400.000 ;
    END
  END proj4_cnt[14]
  PIN proj4_cnt[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 815.670 396.000 815.950 400.000 ;
    END
  END proj4_cnt[15]
  PIN proj4_cnt[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.410 396.000 824.690 400.000 ;
    END
  END proj4_cnt[16]
  PIN proj4_cnt[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 833.150 396.000 833.430 400.000 ;
    END
  END proj4_cnt[17]
  PIN proj4_cnt[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.890 396.000 842.170 400.000 ;
    END
  END proj4_cnt[18]
  PIN proj4_cnt[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 850.630 396.000 850.910 400.000 ;
    END
  END proj4_cnt[19]
  PIN proj4_cnt[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 694.230 396.000 694.510 400.000 ;
    END
  END proj4_cnt[1]
  PIN proj4_cnt[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 859.370 396.000 859.650 400.000 ;
    END
  END proj4_cnt[20]
  PIN proj4_cnt[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 867.650 396.000 867.930 400.000 ;
    END
  END proj4_cnt[21]
  PIN proj4_cnt[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.390 396.000 876.670 400.000 ;
    END
  END proj4_cnt[22]
  PIN proj4_cnt[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 885.130 396.000 885.410 400.000 ;
    END
  END proj4_cnt[23]
  PIN proj4_cnt[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 893.870 396.000 894.150 400.000 ;
    END
  END proj4_cnt[24]
  PIN proj4_cnt[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.610 396.000 902.890 400.000 ;
    END
  END proj4_cnt[25]
  PIN proj4_cnt[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 911.350 396.000 911.630 400.000 ;
    END
  END proj4_cnt[26]
  PIN proj4_cnt[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 920.090 396.000 920.370 400.000 ;
    END
  END proj4_cnt[27]
  PIN proj4_cnt[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 928.370 396.000 928.650 400.000 ;
    END
  END proj4_cnt[28]
  PIN proj4_cnt[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 937.110 396.000 937.390 400.000 ;
    END
  END proj4_cnt[29]
  PIN proj4_cnt[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.970 396.000 703.250 400.000 ;
    END
  END proj4_cnt[2]
  PIN proj4_cnt[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 945.850 396.000 946.130 400.000 ;
    END
  END proj4_cnt[30]
  PIN proj4_cnt[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 954.590 396.000 954.870 400.000 ;
    END
  END proj4_cnt[31]
  PIN proj4_cnt[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 711.710 396.000 711.990 400.000 ;
    END
  END proj4_cnt[3]
  PIN proj4_cnt[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.450 396.000 720.730 400.000 ;
    END
  END proj4_cnt[4]
  PIN proj4_cnt[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.190 396.000 729.470 400.000 ;
    END
  END proj4_cnt[5]
  PIN proj4_cnt[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 737.930 396.000 738.210 400.000 ;
    END
  END proj4_cnt[6]
  PIN proj4_cnt[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 746.670 396.000 746.950 400.000 ;
    END
  END proj4_cnt[7]
  PIN proj4_cnt[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.950 396.000 755.230 400.000 ;
    END
  END proj4_cnt[8]
  PIN proj4_cnt[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 763.690 396.000 763.970 400.000 ;
    END
  END proj4_cnt[9]
  PIN proj4_cnt_cont[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 687.790 396.000 688.070 400.000 ;
    END
  END proj4_cnt_cont[0]
  PIN proj4_cnt_cont[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 774.730 396.000 775.010 400.000 ;
    END
  END proj4_cnt_cont[10]
  PIN proj4_cnt_cont[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.470 396.000 783.750 400.000 ;
    END
  END proj4_cnt_cont[11]
  PIN proj4_cnt_cont[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 792.210 396.000 792.490 400.000 ;
    END
  END proj4_cnt_cont[12]
  PIN proj4_cnt_cont[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.490 396.000 800.770 400.000 ;
    END
  END proj4_cnt_cont[13]
  PIN proj4_cnt_cont[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 809.230 396.000 809.510 400.000 ;
    END
  END proj4_cnt_cont[14]
  PIN proj4_cnt_cont[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 817.970 396.000 818.250 400.000 ;
    END
  END proj4_cnt_cont[15]
  PIN proj4_cnt_cont[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 826.710 396.000 826.990 400.000 ;
    END
  END proj4_cnt_cont[16]
  PIN proj4_cnt_cont[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 835.450 396.000 835.730 400.000 ;
    END
  END proj4_cnt_cont[17]
  PIN proj4_cnt_cont[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 844.190 396.000 844.470 400.000 ;
    END
  END proj4_cnt_cont[18]
  PIN proj4_cnt_cont[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 852.470 396.000 852.750 400.000 ;
    END
  END proj4_cnt_cont[19]
  PIN proj4_cnt_cont[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 696.530 396.000 696.810 400.000 ;
    END
  END proj4_cnt_cont[1]
  PIN proj4_cnt_cont[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 861.210 396.000 861.490 400.000 ;
    END
  END proj4_cnt_cont[20]
  PIN proj4_cnt_cont[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 869.950 396.000 870.230 400.000 ;
    END
  END proj4_cnt_cont[21]
  PIN proj4_cnt_cont[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 878.690 396.000 878.970 400.000 ;
    END
  END proj4_cnt_cont[22]
  PIN proj4_cnt_cont[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 887.430 396.000 887.710 400.000 ;
    END
  END proj4_cnt_cont[23]
  PIN proj4_cnt_cont[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.170 396.000 896.450 400.000 ;
    END
  END proj4_cnt_cont[24]
  PIN proj4_cnt_cont[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 904.910 396.000 905.190 400.000 ;
    END
  END proj4_cnt_cont[25]
  PIN proj4_cnt_cont[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 913.190 396.000 913.470 400.000 ;
    END
  END proj4_cnt_cont[26]
  PIN proj4_cnt_cont[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 921.930 396.000 922.210 400.000 ;
    END
  END proj4_cnt_cont[27]
  PIN proj4_cnt_cont[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.670 396.000 930.950 400.000 ;
    END
  END proj4_cnt_cont[28]
  PIN proj4_cnt_cont[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 939.410 396.000 939.690 400.000 ;
    END
  END proj4_cnt_cont[29]
  PIN proj4_cnt_cont[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.270 396.000 705.550 400.000 ;
    END
  END proj4_cnt_cont[2]
  PIN proj4_cnt_cont[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.150 396.000 948.430 400.000 ;
    END
  END proj4_cnt_cont[30]
  PIN proj4_cnt_cont[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 956.890 396.000 957.170 400.000 ;
    END
  END proj4_cnt_cont[31]
  PIN proj4_cnt_cont[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.010 396.000 714.290 400.000 ;
    END
  END proj4_cnt_cont[3]
  PIN proj4_cnt_cont[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.750 396.000 723.030 400.000 ;
    END
  END proj4_cnt_cont[4]
  PIN proj4_cnt_cont[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 731.490 396.000 731.770 400.000 ;
    END
  END proj4_cnt_cont[5]
  PIN proj4_cnt_cont[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 739.770 396.000 740.050 400.000 ;
    END
  END proj4_cnt_cont[6]
  PIN proj4_cnt_cont[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 748.510 396.000 748.790 400.000 ;
    END
  END proj4_cnt_cont[7]
  PIN proj4_cnt_cont[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.250 396.000 757.530 400.000 ;
    END
  END proj4_cnt_cont[8]
  PIN proj4_cnt_cont[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.990 396.000 766.270 400.000 ;
    END
  END proj4_cnt_cont[9]
  PIN proj4_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 690.090 396.000 690.370 400.000 ;
    END
  END proj4_io_in[0]
  PIN proj4_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 777.030 396.000 777.310 400.000 ;
    END
  END proj4_io_in[10]
  PIN proj4_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 785.310 396.000 785.590 400.000 ;
    END
  END proj4_io_in[11]
  PIN proj4_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 794.050 396.000 794.330 400.000 ;
    END
  END proj4_io_in[12]
  PIN proj4_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 802.790 396.000 803.070 400.000 ;
    END
  END proj4_io_in[13]
  PIN proj4_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 811.530 396.000 811.810 400.000 ;
    END
  END proj4_io_in[14]
  PIN proj4_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 820.270 396.000 820.550 400.000 ;
    END
  END proj4_io_in[15]
  PIN proj4_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 829.010 396.000 829.290 400.000 ;
    END
  END proj4_io_in[16]
  PIN proj4_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 837.290 396.000 837.570 400.000 ;
    END
  END proj4_io_in[17]
  PIN proj4_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 846.030 396.000 846.310 400.000 ;
    END
  END proj4_io_in[18]
  PIN proj4_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 854.770 396.000 855.050 400.000 ;
    END
  END proj4_io_in[19]
  PIN proj4_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 698.830 396.000 699.110 400.000 ;
    END
  END proj4_io_in[1]
  PIN proj4_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 863.510 396.000 863.790 400.000 ;
    END
  END proj4_io_in[20]
  PIN proj4_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 872.250 396.000 872.530 400.000 ;
    END
  END proj4_io_in[21]
  PIN proj4_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.990 396.000 881.270 400.000 ;
    END
  END proj4_io_in[22]
  PIN proj4_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 889.730 396.000 890.010 400.000 ;
    END
  END proj4_io_in[23]
  PIN proj4_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 898.010 396.000 898.290 400.000 ;
    END
  END proj4_io_in[24]
  PIN proj4_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.750 396.000 907.030 400.000 ;
    END
  END proj4_io_in[25]
  PIN proj4_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 915.490 396.000 915.770 400.000 ;
    END
  END proj4_io_in[26]
  PIN proj4_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.230 396.000 924.510 400.000 ;
    END
  END proj4_io_in[27]
  PIN proj4_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 932.970 396.000 933.250 400.000 ;
    END
  END proj4_io_in[28]
  PIN proj4_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 941.710 396.000 941.990 400.000 ;
    END
  END proj4_io_in[29]
  PIN proj4_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 707.570 396.000 707.850 400.000 ;
    END
  END proj4_io_in[2]
  PIN proj4_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 950.450 396.000 950.730 400.000 ;
    END
  END proj4_io_in[30]
  PIN proj4_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 958.730 396.000 959.010 400.000 ;
    END
  END proj4_io_in[31]
  PIN proj4_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 963.330 396.000 963.610 400.000 ;
    END
  END proj4_io_in[32]
  PIN proj4_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.470 396.000 967.750 400.000 ;
    END
  END proj4_io_in[33]
  PIN proj4_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 972.070 396.000 972.350 400.000 ;
    END
  END proj4_io_in[34]
  PIN proj4_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 976.210 396.000 976.490 400.000 ;
    END
  END proj4_io_in[35]
  PIN proj4_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 980.810 396.000 981.090 400.000 ;
    END
  END proj4_io_in[36]
  PIN proj4_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 984.950 396.000 985.230 400.000 ;
    END
  END proj4_io_in[37]
  PIN proj4_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 716.310 396.000 716.590 400.000 ;
    END
  END proj4_io_in[3]
  PIN proj4_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.590 396.000 724.870 400.000 ;
    END
  END proj4_io_in[4]
  PIN proj4_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 733.330 396.000 733.610 400.000 ;
    END
  END proj4_io_in[5]
  PIN proj4_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 742.070 396.000 742.350 400.000 ;
    END
  END proj4_io_in[6]
  PIN proj4_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 750.810 396.000 751.090 400.000 ;
    END
  END proj4_io_in[7]
  PIN proj4_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 759.550 396.000 759.830 400.000 ;
    END
  END proj4_io_in[8]
  PIN proj4_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 768.290 396.000 768.570 400.000 ;
    END
  END proj4_io_in[9]
  PIN proj4_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 692.390 396.000 692.670 400.000 ;
    END
  END proj4_io_out[0]
  PIN proj4_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 778.870 396.000 779.150 400.000 ;
    END
  END proj4_io_out[10]
  PIN proj4_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.610 396.000 787.890 400.000 ;
    END
  END proj4_io_out[11]
  PIN proj4_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 796.350 396.000 796.630 400.000 ;
    END
  END proj4_io_out[12]
  PIN proj4_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.090 396.000 805.370 400.000 ;
    END
  END proj4_io_out[13]
  PIN proj4_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 813.830 396.000 814.110 400.000 ;
    END
  END proj4_io_out[14]
  PIN proj4_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 822.570 396.000 822.850 400.000 ;
    END
  END proj4_io_out[15]
  PIN proj4_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.850 396.000 831.130 400.000 ;
    END
  END proj4_io_out[16]
  PIN proj4_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 839.590 396.000 839.870 400.000 ;
    END
  END proj4_io_out[17]
  PIN proj4_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 848.330 396.000 848.610 400.000 ;
    END
  END proj4_io_out[18]
  PIN proj4_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 857.070 396.000 857.350 400.000 ;
    END
  END proj4_io_out[19]
  PIN proj4_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 701.130 396.000 701.410 400.000 ;
    END
  END proj4_io_out[1]
  PIN proj4_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 865.810 396.000 866.090 400.000 ;
    END
  END proj4_io_out[20]
  PIN proj4_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.550 396.000 874.830 400.000 ;
    END
  END proj4_io_out[21]
  PIN proj4_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.830 396.000 883.110 400.000 ;
    END
  END proj4_io_out[22]
  PIN proj4_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.570 396.000 891.850 400.000 ;
    END
  END proj4_io_out[23]
  PIN proj4_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.310 396.000 900.590 400.000 ;
    END
  END proj4_io_out[24]
  PIN proj4_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 909.050 396.000 909.330 400.000 ;
    END
  END proj4_io_out[25]
  PIN proj4_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 917.790 396.000 918.070 400.000 ;
    END
  END proj4_io_out[26]
  PIN proj4_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 926.530 396.000 926.810 400.000 ;
    END
  END proj4_io_out[27]
  PIN proj4_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 935.270 396.000 935.550 400.000 ;
    END
  END proj4_io_out[28]
  PIN proj4_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 943.550 396.000 943.830 400.000 ;
    END
  END proj4_io_out[29]
  PIN proj4_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 709.410 396.000 709.690 400.000 ;
    END
  END proj4_io_out[2]
  PIN proj4_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 952.290 396.000 952.570 400.000 ;
    END
  END proj4_io_out[30]
  PIN proj4_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 961.030 396.000 961.310 400.000 ;
    END
  END proj4_io_out[31]
  PIN proj4_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.630 396.000 965.910 400.000 ;
    END
  END proj4_io_out[32]
  PIN proj4_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.770 396.000 970.050 400.000 ;
    END
  END proj4_io_out[33]
  PIN proj4_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 973.910 396.000 974.190 400.000 ;
    END
  END proj4_io_out[34]
  PIN proj4_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.510 396.000 978.790 400.000 ;
    END
  END proj4_io_out[35]
  PIN proj4_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 982.650 396.000 982.930 400.000 ;
    END
  END proj4_io_out[36]
  PIN proj4_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 987.250 396.000 987.530 400.000 ;
    END
  END proj4_io_out[37]
  PIN proj4_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 718.150 396.000 718.430 400.000 ;
    END
  END proj4_io_out[3]
  PIN proj4_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 726.890 396.000 727.170 400.000 ;
    END
  END proj4_io_out[4]
  PIN proj4_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 735.630 396.000 735.910 400.000 ;
    END
  END proj4_io_out[5]
  PIN proj4_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 744.370 396.000 744.650 400.000 ;
    END
  END proj4_io_out[6]
  PIN proj4_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.110 396.000 753.390 400.000 ;
    END
  END proj4_io_out[7]
  PIN proj4_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 761.850 396.000 762.130 400.000 ;
    END
  END proj4_io_out[8]
  PIN proj4_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 770.130 396.000 770.410 400.000 ;
    END
  END proj4_io_out[9]
  PIN proj4_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 681.350 396.000 681.630 400.000 ;
    END
  END proj4_reset
  PIN proj4_wb_update
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 683.650 396.000 683.930 400.000 ;
    END
  END proj4_wb_update
  PIN proj5_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.090 396.000 989.370 400.000 ;
    END
  END proj5_clk
  PIN proj5_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.990 396.000 996.270 400.000 ;
    END
  END proj5_io_in[0]
  PIN proj5_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1039.230 396.000 1039.510 400.000 ;
    END
  END proj5_io_in[10]
  PIN proj5_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1043.370 396.000 1043.650 400.000 ;
    END
  END proj5_io_in[11]
  PIN proj5_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1047.970 396.000 1048.250 400.000 ;
    END
  END proj5_io_in[12]
  PIN proj5_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1052.110 396.000 1052.390 400.000 ;
    END
  END proj5_io_in[13]
  PIN proj5_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1056.250 396.000 1056.530 400.000 ;
    END
  END proj5_io_in[14]
  PIN proj5_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1060.850 396.000 1061.130 400.000 ;
    END
  END proj5_io_in[15]
  PIN proj5_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1064.990 396.000 1065.270 400.000 ;
    END
  END proj5_io_in[16]
  PIN proj5_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1069.590 396.000 1069.870 400.000 ;
    END
  END proj5_io_in[17]
  PIN proj5_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1073.730 396.000 1074.010 400.000 ;
    END
  END proj5_io_in[18]
  PIN proj5_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1078.330 396.000 1078.610 400.000 ;
    END
  END proj5_io_in[19]
  PIN proj5_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1000.130 396.000 1000.410 400.000 ;
    END
  END proj5_io_in[1]
  PIN proj5_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1082.470 396.000 1082.750 400.000 ;
    END
  END proj5_io_in[20]
  PIN proj5_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1086.610 396.000 1086.890 400.000 ;
    END
  END proj5_io_in[21]
  PIN proj5_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1091.210 396.000 1091.490 400.000 ;
    END
  END proj5_io_in[22]
  PIN proj5_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1095.350 396.000 1095.630 400.000 ;
    END
  END proj5_io_in[23]
  PIN proj5_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1099.950 396.000 1100.230 400.000 ;
    END
  END proj5_io_in[24]
  PIN proj5_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1104.090 396.000 1104.370 400.000 ;
    END
  END proj5_io_in[25]
  PIN proj5_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1108.690 396.000 1108.970 400.000 ;
    END
  END proj5_io_in[26]
  PIN proj5_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1112.830 396.000 1113.110 400.000 ;
    END
  END proj5_io_in[27]
  PIN proj5_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1116.970 396.000 1117.250 400.000 ;
    END
  END proj5_io_in[28]
  PIN proj5_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1121.570 396.000 1121.850 400.000 ;
    END
  END proj5_io_in[29]
  PIN proj5_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1004.270 396.000 1004.550 400.000 ;
    END
  END proj5_io_in[2]
  PIN proj5_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1125.710 396.000 1125.990 400.000 ;
    END
  END proj5_io_in[30]
  PIN proj5_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1130.310 396.000 1130.590 400.000 ;
    END
  END proj5_io_in[31]
  PIN proj5_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1134.450 396.000 1134.730 400.000 ;
    END
  END proj5_io_in[32]
  PIN proj5_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1139.050 396.000 1139.330 400.000 ;
    END
  END proj5_io_in[33]
  PIN proj5_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1143.190 396.000 1143.470 400.000 ;
    END
  END proj5_io_in[34]
  PIN proj5_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1147.330 396.000 1147.610 400.000 ;
    END
  END proj5_io_in[35]
  PIN proj5_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.930 396.000 1152.210 400.000 ;
    END
  END proj5_io_in[36]
  PIN proj5_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.070 396.000 1156.350 400.000 ;
    END
  END proj5_io_in[37]
  PIN proj5_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1008.870 396.000 1009.150 400.000 ;
    END
  END proj5_io_in[3]
  PIN proj5_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.010 396.000 1013.290 400.000 ;
    END
  END proj5_io_in[4]
  PIN proj5_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1017.610 396.000 1017.890 400.000 ;
    END
  END proj5_io_in[5]
  PIN proj5_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1021.750 396.000 1022.030 400.000 ;
    END
  END proj5_io_in[6]
  PIN proj5_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1025.890 396.000 1026.170 400.000 ;
    END
  END proj5_io_in[7]
  PIN proj5_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1030.490 396.000 1030.770 400.000 ;
    END
  END proj5_io_in[8]
  PIN proj5_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1034.630 396.000 1034.910 400.000 ;
    END
  END proj5_io_in[9]
  PIN proj5_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 997.830 396.000 998.110 400.000 ;
    END
  END proj5_io_out[0]
  PIN proj5_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1041.070 396.000 1041.350 400.000 ;
    END
  END proj5_io_out[10]
  PIN proj5_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.670 396.000 1045.950 400.000 ;
    END
  END proj5_io_out[11]
  PIN proj5_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1049.810 396.000 1050.090 400.000 ;
    END
  END proj5_io_out[12]
  PIN proj5_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1054.410 396.000 1054.690 400.000 ;
    END
  END proj5_io_out[13]
  PIN proj5_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.550 396.000 1058.830 400.000 ;
    END
  END proj5_io_out[14]
  PIN proj5_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.150 396.000 1063.430 400.000 ;
    END
  END proj5_io_out[15]
  PIN proj5_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1067.290 396.000 1067.570 400.000 ;
    END
  END proj5_io_out[16]
  PIN proj5_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1071.430 396.000 1071.710 400.000 ;
    END
  END proj5_io_out[17]
  PIN proj5_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1076.030 396.000 1076.310 400.000 ;
    END
  END proj5_io_out[18]
  PIN proj5_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.170 396.000 1080.450 400.000 ;
    END
  END proj5_io_out[19]
  PIN proj5_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1002.430 396.000 1002.710 400.000 ;
    END
  END proj5_io_out[1]
  PIN proj5_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1084.770 396.000 1085.050 400.000 ;
    END
  END proj5_io_out[20]
  PIN proj5_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1088.910 396.000 1089.190 400.000 ;
    END
  END proj5_io_out[21]
  PIN proj5_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1093.510 396.000 1093.790 400.000 ;
    END
  END proj5_io_out[22]
  PIN proj5_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.650 396.000 1097.930 400.000 ;
    END
  END proj5_io_out[23]
  PIN proj5_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1101.790 396.000 1102.070 400.000 ;
    END
  END proj5_io_out[24]
  PIN proj5_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1106.390 396.000 1106.670 400.000 ;
    END
  END proj5_io_out[25]
  PIN proj5_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.530 396.000 1110.810 400.000 ;
    END
  END proj5_io_out[26]
  PIN proj5_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1115.130 396.000 1115.410 400.000 ;
    END
  END proj5_io_out[27]
  PIN proj5_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1119.270 396.000 1119.550 400.000 ;
    END
  END proj5_io_out[28]
  PIN proj5_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1123.870 396.000 1124.150 400.000 ;
    END
  END proj5_io_out[29]
  PIN proj5_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1006.570 396.000 1006.850 400.000 ;
    END
  END proj5_io_out[2]
  PIN proj5_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1128.010 396.000 1128.290 400.000 ;
    END
  END proj5_io_out[30]
  PIN proj5_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.150 396.000 1132.430 400.000 ;
    END
  END proj5_io_out[31]
  PIN proj5_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1136.750 396.000 1137.030 400.000 ;
    END
  END proj5_io_out[32]
  PIN proj5_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1140.890 396.000 1141.170 400.000 ;
    END
  END proj5_io_out[33]
  PIN proj5_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1145.490 396.000 1145.770 400.000 ;
    END
  END proj5_io_out[34]
  PIN proj5_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1149.630 396.000 1149.910 400.000 ;
    END
  END proj5_io_out[35]
  PIN proj5_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1154.230 396.000 1154.510 400.000 ;
    END
  END proj5_io_out[36]
  PIN proj5_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1158.370 396.000 1158.650 400.000 ;
    END
  END proj5_io_out[37]
  PIN proj5_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1010.710 396.000 1010.990 400.000 ;
    END
  END proj5_io_out[3]
  PIN proj5_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.310 396.000 1015.590 400.000 ;
    END
  END proj5_io_out[4]
  PIN proj5_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.450 396.000 1019.730 400.000 ;
    END
  END proj5_io_out[5]
  PIN proj5_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1024.050 396.000 1024.330 400.000 ;
    END
  END proj5_io_out[6]
  PIN proj5_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1028.190 396.000 1028.470 400.000 ;
    END
  END proj5_io_out[7]
  PIN proj5_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.790 396.000 1033.070 400.000 ;
    END
  END proj5_io_out[8]
  PIN proj5_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.930 396.000 1037.210 400.000 ;
    END
  END proj5_io_out[9]
  PIN proj5_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 991.390 396.000 991.670 400.000 ;
    END
  END proj5_reset
  PIN proj5_wb_update
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 993.690 396.000 993.970 400.000 ;
    END
  END proj5_wb_update
  PIN proj6_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1160.670 396.000 1160.950 400.000 ;
    END
  END proj6_clk
  PIN proj6_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1162.510 396.000 1162.790 400.000 ;
    END
  END proj6_io_in[0]
  PIN proj6_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1206.210 396.000 1206.490 400.000 ;
    END
  END proj6_io_in[10]
  PIN proj6_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1210.350 396.000 1210.630 400.000 ;
    END
  END proj6_io_in[11]
  PIN proj6_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1214.490 396.000 1214.770 400.000 ;
    END
  END proj6_io_in[12]
  PIN proj6_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1219.090 396.000 1219.370 400.000 ;
    END
  END proj6_io_in[13]
  PIN proj6_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1223.230 396.000 1223.510 400.000 ;
    END
  END proj6_io_in[14]
  PIN proj6_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.830 396.000 1228.110 400.000 ;
    END
  END proj6_io_in[15]
  PIN proj6_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1231.970 396.000 1232.250 400.000 ;
    END
  END proj6_io_in[16]
  PIN proj6_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1236.570 396.000 1236.850 400.000 ;
    END
  END proj6_io_in[17]
  PIN proj6_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1240.710 396.000 1240.990 400.000 ;
    END
  END proj6_io_in[18]
  PIN proj6_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1244.850 396.000 1245.130 400.000 ;
    END
  END proj6_io_in[19]
  PIN proj6_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1167.110 396.000 1167.390 400.000 ;
    END
  END proj6_io_in[1]
  PIN proj6_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1249.450 396.000 1249.730 400.000 ;
    END
  END proj6_io_in[20]
  PIN proj6_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1253.590 396.000 1253.870 400.000 ;
    END
  END proj6_io_in[21]
  PIN proj6_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1258.190 396.000 1258.470 400.000 ;
    END
  END proj6_io_in[22]
  PIN proj6_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1262.330 396.000 1262.610 400.000 ;
    END
  END proj6_io_in[23]
  PIN proj6_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1266.930 396.000 1267.210 400.000 ;
    END
  END proj6_io_in[24]
  PIN proj6_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1271.070 396.000 1271.350 400.000 ;
    END
  END proj6_io_in[25]
  PIN proj6_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1275.210 396.000 1275.490 400.000 ;
    END
  END proj6_io_in[26]
  PIN proj6_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1279.810 396.000 1280.090 400.000 ;
    END
  END proj6_io_in[27]
  PIN proj6_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1283.950 396.000 1284.230 400.000 ;
    END
  END proj6_io_in[28]
  PIN proj6_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1288.550 396.000 1288.830 400.000 ;
    END
  END proj6_io_in[29]
  PIN proj6_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1171.250 396.000 1171.530 400.000 ;
    END
  END proj6_io_in[2]
  PIN proj6_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1292.690 396.000 1292.970 400.000 ;
    END
  END proj6_io_in[30]
  PIN proj6_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1297.290 396.000 1297.570 400.000 ;
    END
  END proj6_io_in[31]
  PIN proj6_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1301.430 396.000 1301.710 400.000 ;
    END
  END proj6_io_in[32]
  PIN proj6_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1305.570 396.000 1305.850 400.000 ;
    END
  END proj6_io_in[33]
  PIN proj6_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1310.170 396.000 1310.450 400.000 ;
    END
  END proj6_io_in[34]
  PIN proj6_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1314.310 396.000 1314.590 400.000 ;
    END
  END proj6_io_in[35]
  PIN proj6_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1318.910 396.000 1319.190 400.000 ;
    END
  END proj6_io_in[36]
  PIN proj6_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1323.050 396.000 1323.330 400.000 ;
    END
  END proj6_io_in[37]
  PIN proj6_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1175.850 396.000 1176.130 400.000 ;
    END
  END proj6_io_in[3]
  PIN proj6_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1179.990 396.000 1180.270 400.000 ;
    END
  END proj6_io_in[4]
  PIN proj6_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1184.130 396.000 1184.410 400.000 ;
    END
  END proj6_io_in[5]
  PIN proj6_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1188.730 396.000 1189.010 400.000 ;
    END
  END proj6_io_in[6]
  PIN proj6_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1192.870 396.000 1193.150 400.000 ;
    END
  END proj6_io_in[7]
  PIN proj6_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1197.470 396.000 1197.750 400.000 ;
    END
  END proj6_io_in[8]
  PIN proj6_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1201.610 396.000 1201.890 400.000 ;
    END
  END proj6_io_in[9]
  PIN proj6_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1164.810 396.000 1165.090 400.000 ;
    END
  END proj6_io_out[0]
  PIN proj6_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1208.050 396.000 1208.330 400.000 ;
    END
  END proj6_io_out[10]
  PIN proj6_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1212.650 396.000 1212.930 400.000 ;
    END
  END proj6_io_out[11]
  PIN proj6_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1216.790 396.000 1217.070 400.000 ;
    END
  END proj6_io_out[12]
  PIN proj6_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.390 396.000 1221.670 400.000 ;
    END
  END proj6_io_out[13]
  PIN proj6_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1225.530 396.000 1225.810 400.000 ;
    END
  END proj6_io_out[14]
  PIN proj6_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1229.670 396.000 1229.950 400.000 ;
    END
  END proj6_io_out[15]
  PIN proj6_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1234.270 396.000 1234.550 400.000 ;
    END
  END proj6_io_out[16]
  PIN proj6_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1238.410 396.000 1238.690 400.000 ;
    END
  END proj6_io_out[17]
  PIN proj6_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.010 396.000 1243.290 400.000 ;
    END
  END proj6_io_out[18]
  PIN proj6_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1247.150 396.000 1247.430 400.000 ;
    END
  END proj6_io_out[19]
  PIN proj6_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.950 396.000 1169.230 400.000 ;
    END
  END proj6_io_out[1]
  PIN proj6_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.750 396.000 1252.030 400.000 ;
    END
  END proj6_io_out[20]
  PIN proj6_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1255.890 396.000 1256.170 400.000 ;
    END
  END proj6_io_out[21]
  PIN proj6_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1260.030 396.000 1260.310 400.000 ;
    END
  END proj6_io_out[22]
  PIN proj6_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1264.630 396.000 1264.910 400.000 ;
    END
  END proj6_io_out[23]
  PIN proj6_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1268.770 396.000 1269.050 400.000 ;
    END
  END proj6_io_out[24]
  PIN proj6_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1273.370 396.000 1273.650 400.000 ;
    END
  END proj6_io_out[25]
  PIN proj6_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.510 396.000 1277.790 400.000 ;
    END
  END proj6_io_out[26]
  PIN proj6_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1282.110 396.000 1282.390 400.000 ;
    END
  END proj6_io_out[27]
  PIN proj6_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1286.250 396.000 1286.530 400.000 ;
    END
  END proj6_io_out[28]
  PIN proj6_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1290.390 396.000 1290.670 400.000 ;
    END
  END proj6_io_out[29]
  PIN proj6_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1173.550 396.000 1173.830 400.000 ;
    END
  END proj6_io_out[2]
  PIN proj6_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.990 396.000 1295.270 400.000 ;
    END
  END proj6_io_out[30]
  PIN proj6_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1299.130 396.000 1299.410 400.000 ;
    END
  END proj6_io_out[31]
  PIN proj6_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1303.730 396.000 1304.010 400.000 ;
    END
  END proj6_io_out[32]
  PIN proj6_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1307.870 396.000 1308.150 400.000 ;
    END
  END proj6_io_out[33]
  PIN proj6_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1312.470 396.000 1312.750 400.000 ;
    END
  END proj6_io_out[34]
  PIN proj6_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1316.610 396.000 1316.890 400.000 ;
    END
  END proj6_io_out[35]
  PIN proj6_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1320.750 396.000 1321.030 400.000 ;
    END
  END proj6_io_out[36]
  PIN proj6_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1325.350 396.000 1325.630 400.000 ;
    END
  END proj6_io_out[37]
  PIN proj6_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1177.690 396.000 1177.970 400.000 ;
    END
  END proj6_io_out[3]
  PIN proj6_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1182.290 396.000 1182.570 400.000 ;
    END
  END proj6_io_out[4]
  PIN proj6_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1186.430 396.000 1186.710 400.000 ;
    END
  END proj6_io_out[5]
  PIN proj6_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1191.030 396.000 1191.310 400.000 ;
    END
  END proj6_io_out[6]
  PIN proj6_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 396.000 1195.450 400.000 ;
    END
  END proj6_io_out[7]
  PIN proj6_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1199.310 396.000 1199.590 400.000 ;
    END
  END proj6_io_out[8]
  PIN proj6_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.910 396.000 1204.190 400.000 ;
    END
  END proj6_io_out[9]
  PIN proj7_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 345.550 396.000 345.830 400.000 ;
    END
  END proj7_io_in[0]
  PIN proj7_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.790 396.000 389.070 400.000 ;
    END
  END proj7_io_in[10]
  PIN proj7_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.930 396.000 393.210 400.000 ;
    END
  END proj7_io_in[11]
  PIN proj7_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 397.530 396.000 397.810 400.000 ;
    END
  END proj7_io_in[12]
  PIN proj7_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.670 396.000 401.950 400.000 ;
    END
  END proj7_io_in[13]
  PIN proj7_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 406.270 396.000 406.550 400.000 ;
    END
  END proj7_io_in[14]
  PIN proj7_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 410.410 396.000 410.690 400.000 ;
    END
  END proj7_io_in[15]
  PIN proj7_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 415.010 396.000 415.290 400.000 ;
    END
  END proj7_io_in[16]
  PIN proj7_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 419.150 396.000 419.430 400.000 ;
    END
  END proj7_io_in[17]
  PIN proj7_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.290 396.000 423.570 400.000 ;
    END
  END proj7_io_in[18]
  PIN proj7_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.890 396.000 428.170 400.000 ;
    END
  END proj7_io_in[19]
  PIN proj7_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 349.690 396.000 349.970 400.000 ;
    END
  END proj7_io_in[1]
  PIN proj7_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 432.030 396.000 432.310 400.000 ;
    END
  END proj7_io_in[20]
  PIN proj7_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 436.630 396.000 436.910 400.000 ;
    END
  END proj7_io_in[21]
  PIN proj7_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 440.770 396.000 441.050 400.000 ;
    END
  END proj7_io_in[22]
  PIN proj7_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.370 396.000 445.650 400.000 ;
    END
  END proj7_io_in[23]
  PIN proj7_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 449.510 396.000 449.790 400.000 ;
    END
  END proj7_io_in[24]
  PIN proj7_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 453.650 396.000 453.930 400.000 ;
    END
  END proj7_io_in[25]
  PIN proj7_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 458.250 396.000 458.530 400.000 ;
    END
  END proj7_io_in[26]
  PIN proj7_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 462.390 396.000 462.670 400.000 ;
    END
  END proj7_io_in[27]
  PIN proj7_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.990 396.000 467.270 400.000 ;
    END
  END proj7_io_in[28]
  PIN proj7_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 471.130 396.000 471.410 400.000 ;
    END
  END proj7_io_in[29]
  PIN proj7_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.290 396.000 354.570 400.000 ;
    END
  END proj7_io_in[2]
  PIN proj7_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.730 396.000 476.010 400.000 ;
    END
  END proj7_io_in[30]
  PIN proj7_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 479.870 396.000 480.150 400.000 ;
    END
  END proj7_io_in[31]
  PIN proj7_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.010 396.000 484.290 400.000 ;
    END
  END proj7_io_in[32]
  PIN proj7_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.610 396.000 488.890 400.000 ;
    END
  END proj7_io_in[33]
  PIN proj7_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.750 396.000 493.030 400.000 ;
    END
  END proj7_io_in[34]
  PIN proj7_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 497.350 396.000 497.630 400.000 ;
    END
  END proj7_io_in[35]
  PIN proj7_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 501.490 396.000 501.770 400.000 ;
    END
  END proj7_io_in[36]
  PIN proj7_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.630 396.000 505.910 400.000 ;
    END
  END proj7_io_in[37]
  PIN proj7_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 358.430 396.000 358.710 400.000 ;
    END
  END proj7_io_in[3]
  PIN proj7_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.570 396.000 362.850 400.000 ;
    END
  END proj7_io_in[4]
  PIN proj7_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 367.170 396.000 367.450 400.000 ;
    END
  END proj7_io_in[5]
  PIN proj7_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 371.310 396.000 371.590 400.000 ;
    END
  END proj7_io_in[6]
  PIN proj7_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 375.910 396.000 376.190 400.000 ;
    END
  END proj7_io_in[7]
  PIN proj7_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 380.050 396.000 380.330 400.000 ;
    END
  END proj7_io_in[8]
  PIN proj7_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 384.650 396.000 384.930 400.000 ;
    END
  END proj7_io_in[9]
  PIN proj7_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.390 396.000 347.670 400.000 ;
    END
  END proj7_io_out[0]
  PIN proj7_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 391.090 396.000 391.370 400.000 ;
    END
  END proj7_io_out[10]
  PIN proj7_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 395.230 396.000 395.510 400.000 ;
    END
  END proj7_io_out[11]
  PIN proj7_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.830 396.000 400.110 400.000 ;
    END
  END proj7_io_out[12]
  PIN proj7_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.970 396.000 404.250 400.000 ;
    END
  END proj7_io_out[13]
  PIN proj7_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.110 396.000 408.390 400.000 ;
    END
  END proj7_io_out[14]
  PIN proj7_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 412.710 396.000 412.990 400.000 ;
    END
  END proj7_io_out[15]
  PIN proj7_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 416.850 396.000 417.130 400.000 ;
    END
  END proj7_io_out[16]
  PIN proj7_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 421.450 396.000 421.730 400.000 ;
    END
  END proj7_io_out[17]
  PIN proj7_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.590 396.000 425.870 400.000 ;
    END
  END proj7_io_out[18]
  PIN proj7_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 430.190 396.000 430.470 400.000 ;
    END
  END proj7_io_out[19]
  PIN proj7_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.990 396.000 352.270 400.000 ;
    END
  END proj7_io_out[1]
  PIN proj7_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 434.330 396.000 434.610 400.000 ;
    END
  END proj7_io_out[20]
  PIN proj7_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.470 396.000 438.750 400.000 ;
    END
  END proj7_io_out[21]
  PIN proj7_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.070 396.000 443.350 400.000 ;
    END
  END proj7_io_out[22]
  PIN proj7_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 447.210 396.000 447.490 400.000 ;
    END
  END proj7_io_out[23]
  PIN proj7_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.810 396.000 452.090 400.000 ;
    END
  END proj7_io_out[24]
  PIN proj7_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.950 396.000 456.230 400.000 ;
    END
  END proj7_io_out[25]
  PIN proj7_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.550 396.000 460.830 400.000 ;
    END
  END proj7_io_out[26]
  PIN proj7_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 464.690 396.000 464.970 400.000 ;
    END
  END proj7_io_out[27]
  PIN proj7_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 468.830 396.000 469.110 400.000 ;
    END
  END proj7_io_out[28]
  PIN proj7_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 473.430 396.000 473.710 400.000 ;
    END
  END proj7_io_out[29]
  PIN proj7_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.130 396.000 356.410 400.000 ;
    END
  END proj7_io_out[2]
  PIN proj7_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.570 396.000 477.850 400.000 ;
    END
  END proj7_io_out[30]
  PIN proj7_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 482.170 396.000 482.450 400.000 ;
    END
  END proj7_io_out[31]
  PIN proj7_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 486.310 396.000 486.590 400.000 ;
    END
  END proj7_io_out[32]
  PIN proj7_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.910 396.000 491.190 400.000 ;
    END
  END proj7_io_out[33]
  PIN proj7_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.050 396.000 495.330 400.000 ;
    END
  END proj7_io_out[34]
  PIN proj7_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 499.190 396.000 499.470 400.000 ;
    END
  END proj7_io_out[35]
  PIN proj7_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 503.790 396.000 504.070 400.000 ;
    END
  END proj7_io_out[36]
  PIN proj7_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.930 396.000 508.210 400.000 ;
    END
  END proj7_io_out[37]
  PIN proj7_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 360.730 396.000 361.010 400.000 ;
    END
  END proj7_io_out[3]
  PIN proj7_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.870 396.000 365.150 400.000 ;
    END
  END proj7_io_out[4]
  PIN proj7_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 369.470 396.000 369.750 400.000 ;
    END
  END proj7_io_out[5]
  PIN proj7_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 373.610 396.000 373.890 400.000 ;
    END
  END proj7_io_out[6]
  PIN proj7_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 377.750 396.000 378.030 400.000 ;
    END
  END proj7_io_out[7]
  PIN proj7_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.350 396.000 382.630 400.000 ;
    END
  END proj7_io_out[8]
  PIN proj7_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.490 396.000 386.770 400.000 ;
    END
  END proj7_io_out[9]
  PIN proj7_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.250 396.000 343.530 400.000 ;
    END
  END proj7_reset
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 384.240 1500.000 384.840 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 394.440 1500.000 395.040 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1496.470 396.000 1496.750 400.000 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1498.310 0.000 1498.590 4.000 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1498.770 396.000 1499.050 400.000 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 398.055 ;
      LAYER met1 ;
        RECT 0.070 4.460 1494.080 398.440 ;
      LAYER met2 ;
        RECT 0.100 395.720 0.730 398.470 ;
        RECT 1.570 395.720 2.570 398.470 ;
        RECT 3.410 395.720 4.870 398.470 ;
        RECT 5.710 395.720 7.170 398.470 ;
        RECT 8.010 395.720 9.010 398.470 ;
        RECT 9.850 395.720 11.310 398.470 ;
        RECT 12.150 395.720 13.610 398.470 ;
        RECT 14.450 395.720 15.450 398.470 ;
        RECT 16.290 395.720 17.750 398.470 ;
        RECT 18.590 395.720 20.050 398.470 ;
        RECT 20.890 395.720 22.350 398.470 ;
        RECT 23.190 395.720 24.190 398.470 ;
        RECT 25.030 395.720 26.490 398.470 ;
        RECT 27.330 395.720 28.790 398.470 ;
        RECT 29.630 395.720 30.630 398.470 ;
        RECT 31.470 395.720 32.930 398.470 ;
        RECT 33.770 395.720 35.230 398.470 ;
        RECT 36.070 395.720 37.530 398.470 ;
        RECT 38.370 395.720 39.370 398.470 ;
        RECT 40.210 395.720 41.670 398.470 ;
        RECT 42.510 395.720 43.970 398.470 ;
        RECT 44.810 395.720 45.810 398.470 ;
        RECT 46.650 395.720 48.110 398.470 ;
        RECT 48.950 395.720 50.410 398.470 ;
        RECT 51.250 395.720 52.710 398.470 ;
        RECT 53.550 395.720 54.550 398.470 ;
        RECT 55.390 395.720 56.850 398.470 ;
        RECT 57.690 395.720 59.150 398.470 ;
        RECT 59.990 395.720 60.990 398.470 ;
        RECT 61.830 395.720 63.290 398.470 ;
        RECT 64.130 395.720 65.590 398.470 ;
        RECT 66.430 395.720 67.890 398.470 ;
        RECT 68.730 395.720 69.730 398.470 ;
        RECT 70.570 395.720 72.030 398.470 ;
        RECT 72.870 395.720 74.330 398.470 ;
        RECT 75.170 395.720 76.170 398.470 ;
        RECT 77.010 395.720 78.470 398.470 ;
        RECT 79.310 395.720 80.770 398.470 ;
        RECT 81.610 395.720 83.070 398.470 ;
        RECT 83.910 395.720 84.910 398.470 ;
        RECT 85.750 395.720 87.210 398.470 ;
        RECT 88.050 395.720 89.510 398.470 ;
        RECT 90.350 395.720 91.350 398.470 ;
        RECT 92.190 395.720 93.650 398.470 ;
        RECT 94.490 395.720 95.950 398.470 ;
        RECT 96.790 395.720 98.250 398.470 ;
        RECT 99.090 395.720 100.090 398.470 ;
        RECT 100.930 395.720 102.390 398.470 ;
        RECT 103.230 395.720 104.690 398.470 ;
        RECT 105.530 395.720 106.530 398.470 ;
        RECT 107.370 395.720 108.830 398.470 ;
        RECT 109.670 395.720 111.130 398.470 ;
        RECT 111.970 395.720 113.430 398.470 ;
        RECT 114.270 395.720 115.270 398.470 ;
        RECT 116.110 395.720 117.570 398.470 ;
        RECT 118.410 395.720 119.870 398.470 ;
        RECT 120.710 395.720 121.710 398.470 ;
        RECT 122.550 395.720 124.010 398.470 ;
        RECT 124.850 395.720 126.310 398.470 ;
        RECT 127.150 395.720 128.610 398.470 ;
        RECT 129.450 395.720 130.450 398.470 ;
        RECT 131.290 395.720 132.750 398.470 ;
        RECT 133.590 395.720 135.050 398.470 ;
        RECT 135.890 395.720 136.890 398.470 ;
        RECT 137.730 395.720 139.190 398.470 ;
        RECT 140.030 395.720 141.490 398.470 ;
        RECT 142.330 395.720 143.790 398.470 ;
        RECT 144.630 395.720 145.630 398.470 ;
        RECT 146.470 395.720 147.930 398.470 ;
        RECT 148.770 395.720 150.230 398.470 ;
        RECT 151.070 395.720 152.070 398.470 ;
        RECT 152.910 395.720 154.370 398.470 ;
        RECT 155.210 395.720 156.670 398.470 ;
        RECT 157.510 395.720 158.970 398.470 ;
        RECT 159.810 395.720 160.810 398.470 ;
        RECT 161.650 395.720 163.110 398.470 ;
        RECT 163.950 395.720 165.410 398.470 ;
        RECT 166.250 395.720 167.250 398.470 ;
        RECT 168.090 395.720 169.550 398.470 ;
        RECT 170.390 395.720 171.850 398.470 ;
        RECT 172.690 395.720 173.690 398.470 ;
        RECT 174.530 395.720 175.990 398.470 ;
        RECT 176.830 395.720 178.290 398.470 ;
        RECT 179.130 395.720 180.590 398.470 ;
        RECT 181.430 395.720 182.430 398.470 ;
        RECT 183.270 395.720 184.730 398.470 ;
        RECT 185.570 395.720 187.030 398.470 ;
        RECT 187.870 395.720 188.870 398.470 ;
        RECT 189.710 395.720 191.170 398.470 ;
        RECT 192.010 395.720 193.470 398.470 ;
        RECT 194.310 395.720 195.770 398.470 ;
        RECT 196.610 395.720 197.610 398.470 ;
        RECT 198.450 395.720 199.910 398.470 ;
        RECT 200.750 395.720 202.210 398.470 ;
        RECT 203.050 395.720 204.050 398.470 ;
        RECT 204.890 395.720 206.350 398.470 ;
        RECT 207.190 395.720 208.650 398.470 ;
        RECT 209.490 395.720 210.950 398.470 ;
        RECT 211.790 395.720 212.790 398.470 ;
        RECT 213.630 395.720 215.090 398.470 ;
        RECT 215.930 395.720 217.390 398.470 ;
        RECT 218.230 395.720 219.230 398.470 ;
        RECT 220.070 395.720 221.530 398.470 ;
        RECT 222.370 395.720 223.830 398.470 ;
        RECT 224.670 395.720 226.130 398.470 ;
        RECT 226.970 395.720 227.970 398.470 ;
        RECT 228.810 395.720 230.270 398.470 ;
        RECT 231.110 395.720 232.570 398.470 ;
        RECT 233.410 395.720 234.410 398.470 ;
        RECT 235.250 395.720 236.710 398.470 ;
        RECT 237.550 395.720 239.010 398.470 ;
        RECT 239.850 395.720 241.310 398.470 ;
        RECT 242.150 395.720 243.150 398.470 ;
        RECT 243.990 395.720 245.450 398.470 ;
        RECT 246.290 395.720 247.750 398.470 ;
        RECT 248.590 395.720 249.590 398.470 ;
        RECT 250.430 395.720 251.890 398.470 ;
        RECT 252.730 395.720 254.190 398.470 ;
        RECT 255.030 395.720 256.490 398.470 ;
        RECT 257.330 395.720 258.330 398.470 ;
        RECT 259.170 395.720 260.630 398.470 ;
        RECT 261.470 395.720 262.930 398.470 ;
        RECT 263.770 395.720 264.770 398.470 ;
        RECT 265.610 395.720 267.070 398.470 ;
        RECT 267.910 395.720 269.370 398.470 ;
        RECT 270.210 395.720 271.670 398.470 ;
        RECT 272.510 395.720 273.510 398.470 ;
        RECT 274.350 395.720 275.810 398.470 ;
        RECT 276.650 395.720 278.110 398.470 ;
        RECT 278.950 395.720 279.950 398.470 ;
        RECT 280.790 395.720 282.250 398.470 ;
        RECT 283.090 395.720 284.550 398.470 ;
        RECT 285.390 395.720 286.850 398.470 ;
        RECT 287.690 395.720 288.690 398.470 ;
        RECT 289.530 395.720 290.990 398.470 ;
        RECT 291.830 395.720 293.290 398.470 ;
        RECT 294.130 395.720 295.130 398.470 ;
        RECT 295.970 395.720 297.430 398.470 ;
        RECT 298.270 395.720 299.730 398.470 ;
        RECT 300.570 395.720 302.030 398.470 ;
        RECT 302.870 395.720 303.870 398.470 ;
        RECT 304.710 395.720 306.170 398.470 ;
        RECT 307.010 395.720 308.470 398.470 ;
        RECT 309.310 395.720 310.310 398.470 ;
        RECT 311.150 395.720 312.610 398.470 ;
        RECT 313.450 395.720 314.910 398.470 ;
        RECT 315.750 395.720 317.210 398.470 ;
        RECT 318.050 395.720 319.050 398.470 ;
        RECT 319.890 395.720 321.350 398.470 ;
        RECT 322.190 395.720 323.650 398.470 ;
        RECT 324.490 395.720 325.490 398.470 ;
        RECT 326.330 395.720 327.790 398.470 ;
        RECT 328.630 395.720 330.090 398.470 ;
        RECT 330.930 395.720 332.390 398.470 ;
        RECT 333.230 395.720 334.230 398.470 ;
        RECT 335.070 395.720 336.530 398.470 ;
        RECT 337.370 395.720 338.830 398.470 ;
        RECT 339.670 395.720 340.670 398.470 ;
        RECT 341.510 395.720 342.970 398.470 ;
        RECT 343.810 395.720 345.270 398.470 ;
        RECT 346.110 395.720 347.110 398.470 ;
        RECT 347.950 395.720 349.410 398.470 ;
        RECT 350.250 395.720 351.710 398.470 ;
        RECT 352.550 395.720 354.010 398.470 ;
        RECT 354.850 395.720 355.850 398.470 ;
        RECT 356.690 395.720 358.150 398.470 ;
        RECT 358.990 395.720 360.450 398.470 ;
        RECT 361.290 395.720 362.290 398.470 ;
        RECT 363.130 395.720 364.590 398.470 ;
        RECT 365.430 395.720 366.890 398.470 ;
        RECT 367.730 395.720 369.190 398.470 ;
        RECT 370.030 395.720 371.030 398.470 ;
        RECT 371.870 395.720 373.330 398.470 ;
        RECT 374.170 395.720 375.630 398.470 ;
        RECT 376.470 395.720 377.470 398.470 ;
        RECT 378.310 395.720 379.770 398.470 ;
        RECT 380.610 395.720 382.070 398.470 ;
        RECT 382.910 395.720 384.370 398.470 ;
        RECT 385.210 395.720 386.210 398.470 ;
        RECT 387.050 395.720 388.510 398.470 ;
        RECT 389.350 395.720 390.810 398.470 ;
        RECT 391.650 395.720 392.650 398.470 ;
        RECT 393.490 395.720 394.950 398.470 ;
        RECT 395.790 395.720 397.250 398.470 ;
        RECT 398.090 395.720 399.550 398.470 ;
        RECT 400.390 395.720 401.390 398.470 ;
        RECT 402.230 395.720 403.690 398.470 ;
        RECT 404.530 395.720 405.990 398.470 ;
        RECT 406.830 395.720 407.830 398.470 ;
        RECT 408.670 395.720 410.130 398.470 ;
        RECT 410.970 395.720 412.430 398.470 ;
        RECT 413.270 395.720 414.730 398.470 ;
        RECT 415.570 395.720 416.570 398.470 ;
        RECT 417.410 395.720 418.870 398.470 ;
        RECT 419.710 395.720 421.170 398.470 ;
        RECT 422.010 395.720 423.010 398.470 ;
        RECT 423.850 395.720 425.310 398.470 ;
        RECT 426.150 395.720 427.610 398.470 ;
        RECT 428.450 395.720 429.910 398.470 ;
        RECT 430.750 395.720 431.750 398.470 ;
        RECT 432.590 395.720 434.050 398.470 ;
        RECT 434.890 395.720 436.350 398.470 ;
        RECT 437.190 395.720 438.190 398.470 ;
        RECT 439.030 395.720 440.490 398.470 ;
        RECT 441.330 395.720 442.790 398.470 ;
        RECT 443.630 395.720 445.090 398.470 ;
        RECT 445.930 395.720 446.930 398.470 ;
        RECT 447.770 395.720 449.230 398.470 ;
        RECT 450.070 395.720 451.530 398.470 ;
        RECT 452.370 395.720 453.370 398.470 ;
        RECT 454.210 395.720 455.670 398.470 ;
        RECT 456.510 395.720 457.970 398.470 ;
        RECT 458.810 395.720 460.270 398.470 ;
        RECT 461.110 395.720 462.110 398.470 ;
        RECT 462.950 395.720 464.410 398.470 ;
        RECT 465.250 395.720 466.710 398.470 ;
        RECT 467.550 395.720 468.550 398.470 ;
        RECT 469.390 395.720 470.850 398.470 ;
        RECT 471.690 395.720 473.150 398.470 ;
        RECT 473.990 395.720 475.450 398.470 ;
        RECT 476.290 395.720 477.290 398.470 ;
        RECT 478.130 395.720 479.590 398.470 ;
        RECT 480.430 395.720 481.890 398.470 ;
        RECT 482.730 395.720 483.730 398.470 ;
        RECT 484.570 395.720 486.030 398.470 ;
        RECT 486.870 395.720 488.330 398.470 ;
        RECT 489.170 395.720 490.630 398.470 ;
        RECT 491.470 395.720 492.470 398.470 ;
        RECT 493.310 395.720 494.770 398.470 ;
        RECT 495.610 395.720 497.070 398.470 ;
        RECT 497.910 395.720 498.910 398.470 ;
        RECT 499.750 395.720 501.210 398.470 ;
        RECT 502.050 395.720 503.510 398.470 ;
        RECT 504.350 395.720 505.350 398.470 ;
        RECT 506.190 395.720 507.650 398.470 ;
        RECT 508.490 395.720 509.950 398.470 ;
        RECT 510.790 395.720 512.250 398.470 ;
        RECT 513.090 395.720 514.090 398.470 ;
        RECT 514.930 395.720 516.390 398.470 ;
        RECT 517.230 395.720 518.690 398.470 ;
        RECT 519.530 395.720 520.530 398.470 ;
        RECT 521.370 395.720 522.830 398.470 ;
        RECT 523.670 395.720 525.130 398.470 ;
        RECT 525.970 395.720 527.430 398.470 ;
        RECT 528.270 395.720 529.270 398.470 ;
        RECT 530.110 395.720 531.570 398.470 ;
        RECT 532.410 395.720 533.870 398.470 ;
        RECT 534.710 395.720 535.710 398.470 ;
        RECT 536.550 395.720 538.010 398.470 ;
        RECT 538.850 395.720 540.310 398.470 ;
        RECT 541.150 395.720 542.610 398.470 ;
        RECT 543.450 395.720 544.450 398.470 ;
        RECT 545.290 395.720 546.750 398.470 ;
        RECT 547.590 395.720 549.050 398.470 ;
        RECT 549.890 395.720 550.890 398.470 ;
        RECT 551.730 395.720 553.190 398.470 ;
        RECT 554.030 395.720 555.490 398.470 ;
        RECT 556.330 395.720 557.790 398.470 ;
        RECT 558.630 395.720 559.630 398.470 ;
        RECT 560.470 395.720 561.930 398.470 ;
        RECT 562.770 395.720 564.230 398.470 ;
        RECT 565.070 395.720 566.070 398.470 ;
        RECT 566.910 395.720 568.370 398.470 ;
        RECT 569.210 395.720 570.670 398.470 ;
        RECT 571.510 395.720 572.970 398.470 ;
        RECT 573.810 395.720 574.810 398.470 ;
        RECT 575.650 395.720 577.110 398.470 ;
        RECT 577.950 395.720 579.410 398.470 ;
        RECT 580.250 395.720 581.250 398.470 ;
        RECT 582.090 395.720 583.550 398.470 ;
        RECT 584.390 395.720 585.850 398.470 ;
        RECT 586.690 395.720 588.150 398.470 ;
        RECT 588.990 395.720 589.990 398.470 ;
        RECT 590.830 395.720 592.290 398.470 ;
        RECT 593.130 395.720 594.590 398.470 ;
        RECT 595.430 395.720 596.430 398.470 ;
        RECT 597.270 395.720 598.730 398.470 ;
        RECT 599.570 395.720 601.030 398.470 ;
        RECT 601.870 395.720 603.330 398.470 ;
        RECT 604.170 395.720 605.170 398.470 ;
        RECT 606.010 395.720 607.470 398.470 ;
        RECT 608.310 395.720 609.770 398.470 ;
        RECT 610.610 395.720 611.610 398.470 ;
        RECT 612.450 395.720 613.910 398.470 ;
        RECT 614.750 395.720 616.210 398.470 ;
        RECT 617.050 395.720 618.510 398.470 ;
        RECT 619.350 395.720 620.350 398.470 ;
        RECT 621.190 395.720 622.650 398.470 ;
        RECT 623.490 395.720 624.950 398.470 ;
        RECT 625.790 395.720 626.790 398.470 ;
        RECT 627.630 395.720 629.090 398.470 ;
        RECT 629.930 395.720 631.390 398.470 ;
        RECT 632.230 395.720 633.690 398.470 ;
        RECT 634.530 395.720 635.530 398.470 ;
        RECT 636.370 395.720 637.830 398.470 ;
        RECT 638.670 395.720 640.130 398.470 ;
        RECT 640.970 395.720 641.970 398.470 ;
        RECT 642.810 395.720 644.270 398.470 ;
        RECT 645.110 395.720 646.570 398.470 ;
        RECT 647.410 395.720 648.870 398.470 ;
        RECT 649.710 395.720 650.710 398.470 ;
        RECT 651.550 395.720 653.010 398.470 ;
        RECT 653.850 395.720 655.310 398.470 ;
        RECT 656.150 395.720 657.150 398.470 ;
        RECT 657.990 395.720 659.450 398.470 ;
        RECT 660.290 395.720 661.750 398.470 ;
        RECT 662.590 395.720 664.050 398.470 ;
        RECT 664.890 395.720 665.890 398.470 ;
        RECT 666.730 395.720 668.190 398.470 ;
        RECT 669.030 395.720 670.490 398.470 ;
        RECT 671.330 395.720 672.330 398.470 ;
        RECT 673.170 395.720 674.630 398.470 ;
        RECT 675.470 395.720 676.930 398.470 ;
        RECT 677.770 395.720 678.770 398.470 ;
        RECT 679.610 395.720 681.070 398.470 ;
        RECT 681.910 395.720 683.370 398.470 ;
        RECT 684.210 395.720 685.670 398.470 ;
        RECT 686.510 395.720 687.510 398.470 ;
        RECT 688.350 395.720 689.810 398.470 ;
        RECT 690.650 395.720 692.110 398.470 ;
        RECT 692.950 395.720 693.950 398.470 ;
        RECT 694.790 395.720 696.250 398.470 ;
        RECT 697.090 395.720 698.550 398.470 ;
        RECT 699.390 395.720 700.850 398.470 ;
        RECT 701.690 395.720 702.690 398.470 ;
        RECT 703.530 395.720 704.990 398.470 ;
        RECT 705.830 395.720 707.290 398.470 ;
        RECT 708.130 395.720 709.130 398.470 ;
        RECT 709.970 395.720 711.430 398.470 ;
        RECT 712.270 395.720 713.730 398.470 ;
        RECT 714.570 395.720 716.030 398.470 ;
        RECT 716.870 395.720 717.870 398.470 ;
        RECT 718.710 395.720 720.170 398.470 ;
        RECT 721.010 395.720 722.470 398.470 ;
        RECT 723.310 395.720 724.310 398.470 ;
        RECT 725.150 395.720 726.610 398.470 ;
        RECT 727.450 395.720 728.910 398.470 ;
        RECT 729.750 395.720 731.210 398.470 ;
        RECT 732.050 395.720 733.050 398.470 ;
        RECT 733.890 395.720 735.350 398.470 ;
        RECT 736.190 395.720 737.650 398.470 ;
        RECT 738.490 395.720 739.490 398.470 ;
        RECT 740.330 395.720 741.790 398.470 ;
        RECT 742.630 395.720 744.090 398.470 ;
        RECT 744.930 395.720 746.390 398.470 ;
        RECT 747.230 395.720 748.230 398.470 ;
        RECT 749.070 395.720 750.530 398.470 ;
        RECT 751.370 395.720 752.830 398.470 ;
        RECT 753.670 395.720 754.670 398.470 ;
        RECT 755.510 395.720 756.970 398.470 ;
        RECT 757.810 395.720 759.270 398.470 ;
        RECT 760.110 395.720 761.570 398.470 ;
        RECT 762.410 395.720 763.410 398.470 ;
        RECT 764.250 395.720 765.710 398.470 ;
        RECT 766.550 395.720 768.010 398.470 ;
        RECT 768.850 395.720 769.850 398.470 ;
        RECT 770.690 395.720 772.150 398.470 ;
        RECT 772.990 395.720 774.450 398.470 ;
        RECT 775.290 395.720 776.750 398.470 ;
        RECT 777.590 395.720 778.590 398.470 ;
        RECT 779.430 395.720 780.890 398.470 ;
        RECT 781.730 395.720 783.190 398.470 ;
        RECT 784.030 395.720 785.030 398.470 ;
        RECT 785.870 395.720 787.330 398.470 ;
        RECT 788.170 395.720 789.630 398.470 ;
        RECT 790.470 395.720 791.930 398.470 ;
        RECT 792.770 395.720 793.770 398.470 ;
        RECT 794.610 395.720 796.070 398.470 ;
        RECT 796.910 395.720 798.370 398.470 ;
        RECT 799.210 395.720 800.210 398.470 ;
        RECT 801.050 395.720 802.510 398.470 ;
        RECT 803.350 395.720 804.810 398.470 ;
        RECT 805.650 395.720 807.110 398.470 ;
        RECT 807.950 395.720 808.950 398.470 ;
        RECT 809.790 395.720 811.250 398.470 ;
        RECT 812.090 395.720 813.550 398.470 ;
        RECT 814.390 395.720 815.390 398.470 ;
        RECT 816.230 395.720 817.690 398.470 ;
        RECT 818.530 395.720 819.990 398.470 ;
        RECT 820.830 395.720 822.290 398.470 ;
        RECT 823.130 395.720 824.130 398.470 ;
        RECT 824.970 395.720 826.430 398.470 ;
        RECT 827.270 395.720 828.730 398.470 ;
        RECT 829.570 395.720 830.570 398.470 ;
        RECT 831.410 395.720 832.870 398.470 ;
        RECT 833.710 395.720 835.170 398.470 ;
        RECT 836.010 395.720 837.010 398.470 ;
        RECT 837.850 395.720 839.310 398.470 ;
        RECT 840.150 395.720 841.610 398.470 ;
        RECT 842.450 395.720 843.910 398.470 ;
        RECT 844.750 395.720 845.750 398.470 ;
        RECT 846.590 395.720 848.050 398.470 ;
        RECT 848.890 395.720 850.350 398.470 ;
        RECT 851.190 395.720 852.190 398.470 ;
        RECT 853.030 395.720 854.490 398.470 ;
        RECT 855.330 395.720 856.790 398.470 ;
        RECT 857.630 395.720 859.090 398.470 ;
        RECT 859.930 395.720 860.930 398.470 ;
        RECT 861.770 395.720 863.230 398.470 ;
        RECT 864.070 395.720 865.530 398.470 ;
        RECT 866.370 395.720 867.370 398.470 ;
        RECT 868.210 395.720 869.670 398.470 ;
        RECT 870.510 395.720 871.970 398.470 ;
        RECT 872.810 395.720 874.270 398.470 ;
        RECT 875.110 395.720 876.110 398.470 ;
        RECT 876.950 395.720 878.410 398.470 ;
        RECT 879.250 395.720 880.710 398.470 ;
        RECT 881.550 395.720 882.550 398.470 ;
        RECT 883.390 395.720 884.850 398.470 ;
        RECT 885.690 395.720 887.150 398.470 ;
        RECT 887.990 395.720 889.450 398.470 ;
        RECT 890.290 395.720 891.290 398.470 ;
        RECT 892.130 395.720 893.590 398.470 ;
        RECT 894.430 395.720 895.890 398.470 ;
        RECT 896.730 395.720 897.730 398.470 ;
        RECT 898.570 395.720 900.030 398.470 ;
        RECT 900.870 395.720 902.330 398.470 ;
        RECT 903.170 395.720 904.630 398.470 ;
        RECT 905.470 395.720 906.470 398.470 ;
        RECT 907.310 395.720 908.770 398.470 ;
        RECT 909.610 395.720 911.070 398.470 ;
        RECT 911.910 395.720 912.910 398.470 ;
        RECT 913.750 395.720 915.210 398.470 ;
        RECT 916.050 395.720 917.510 398.470 ;
        RECT 918.350 395.720 919.810 398.470 ;
        RECT 920.650 395.720 921.650 398.470 ;
        RECT 922.490 395.720 923.950 398.470 ;
        RECT 924.790 395.720 926.250 398.470 ;
        RECT 927.090 395.720 928.090 398.470 ;
        RECT 928.930 395.720 930.390 398.470 ;
        RECT 931.230 395.720 932.690 398.470 ;
        RECT 933.530 395.720 934.990 398.470 ;
        RECT 935.830 395.720 936.830 398.470 ;
        RECT 937.670 395.720 939.130 398.470 ;
        RECT 939.970 395.720 941.430 398.470 ;
        RECT 942.270 395.720 943.270 398.470 ;
        RECT 944.110 395.720 945.570 398.470 ;
        RECT 946.410 395.720 947.870 398.470 ;
        RECT 948.710 395.720 950.170 398.470 ;
        RECT 951.010 395.720 952.010 398.470 ;
        RECT 952.850 395.720 954.310 398.470 ;
        RECT 955.150 395.720 956.610 398.470 ;
        RECT 957.450 395.720 958.450 398.470 ;
        RECT 959.290 395.720 960.750 398.470 ;
        RECT 961.590 395.720 963.050 398.470 ;
        RECT 963.890 395.720 965.350 398.470 ;
        RECT 966.190 395.720 967.190 398.470 ;
        RECT 968.030 395.720 969.490 398.470 ;
        RECT 970.330 395.720 971.790 398.470 ;
        RECT 972.630 395.720 973.630 398.470 ;
        RECT 974.470 395.720 975.930 398.470 ;
        RECT 976.770 395.720 978.230 398.470 ;
        RECT 979.070 395.720 980.530 398.470 ;
        RECT 981.370 395.720 982.370 398.470 ;
        RECT 983.210 395.720 984.670 398.470 ;
        RECT 985.510 395.720 986.970 398.470 ;
        RECT 987.810 395.720 988.810 398.470 ;
        RECT 989.650 395.720 991.110 398.470 ;
        RECT 991.950 395.720 993.410 398.470 ;
        RECT 994.250 395.720 995.710 398.470 ;
        RECT 996.550 395.720 997.550 398.470 ;
        RECT 998.390 395.720 999.850 398.470 ;
        RECT 1000.690 395.720 1002.150 398.470 ;
        RECT 1002.990 395.720 1003.990 398.470 ;
        RECT 1004.830 395.720 1006.290 398.470 ;
        RECT 1007.130 395.720 1008.590 398.470 ;
        RECT 1009.430 395.720 1010.430 398.470 ;
        RECT 1011.270 395.720 1012.730 398.470 ;
        RECT 1013.570 395.720 1015.030 398.470 ;
        RECT 1015.870 395.720 1017.330 398.470 ;
        RECT 1018.170 395.720 1019.170 398.470 ;
        RECT 1020.010 395.720 1021.470 398.470 ;
        RECT 1022.310 395.720 1023.770 398.470 ;
        RECT 1024.610 395.720 1025.610 398.470 ;
        RECT 1026.450 395.720 1027.910 398.470 ;
        RECT 1028.750 395.720 1030.210 398.470 ;
        RECT 1031.050 395.720 1032.510 398.470 ;
        RECT 1033.350 395.720 1034.350 398.470 ;
        RECT 1035.190 395.720 1036.650 398.470 ;
        RECT 1037.490 395.720 1038.950 398.470 ;
        RECT 1039.790 395.720 1040.790 398.470 ;
        RECT 1041.630 395.720 1043.090 398.470 ;
        RECT 1043.930 395.720 1045.390 398.470 ;
        RECT 1046.230 395.720 1047.690 398.470 ;
        RECT 1048.530 395.720 1049.530 398.470 ;
        RECT 1050.370 395.720 1051.830 398.470 ;
        RECT 1052.670 395.720 1054.130 398.470 ;
        RECT 1054.970 395.720 1055.970 398.470 ;
        RECT 1056.810 395.720 1058.270 398.470 ;
        RECT 1059.110 395.720 1060.570 398.470 ;
        RECT 1061.410 395.720 1062.870 398.470 ;
        RECT 1063.710 395.720 1064.710 398.470 ;
        RECT 1065.550 395.720 1067.010 398.470 ;
        RECT 1067.850 395.720 1069.310 398.470 ;
        RECT 1070.150 395.720 1071.150 398.470 ;
        RECT 1071.990 395.720 1073.450 398.470 ;
        RECT 1074.290 395.720 1075.750 398.470 ;
        RECT 1076.590 395.720 1078.050 398.470 ;
        RECT 1078.890 395.720 1079.890 398.470 ;
        RECT 1080.730 395.720 1082.190 398.470 ;
        RECT 1083.030 395.720 1084.490 398.470 ;
        RECT 1085.330 395.720 1086.330 398.470 ;
        RECT 1087.170 395.720 1088.630 398.470 ;
        RECT 1089.470 395.720 1090.930 398.470 ;
        RECT 1091.770 395.720 1093.230 398.470 ;
        RECT 1094.070 395.720 1095.070 398.470 ;
        RECT 1095.910 395.720 1097.370 398.470 ;
        RECT 1098.210 395.720 1099.670 398.470 ;
        RECT 1100.510 395.720 1101.510 398.470 ;
        RECT 1102.350 395.720 1103.810 398.470 ;
        RECT 1104.650 395.720 1106.110 398.470 ;
        RECT 1106.950 395.720 1108.410 398.470 ;
        RECT 1109.250 395.720 1110.250 398.470 ;
        RECT 1111.090 395.720 1112.550 398.470 ;
        RECT 1113.390 395.720 1114.850 398.470 ;
        RECT 1115.690 395.720 1116.690 398.470 ;
        RECT 1117.530 395.720 1118.990 398.470 ;
        RECT 1119.830 395.720 1121.290 398.470 ;
        RECT 1122.130 395.720 1123.590 398.470 ;
        RECT 1124.430 395.720 1125.430 398.470 ;
        RECT 1126.270 395.720 1127.730 398.470 ;
        RECT 1128.570 395.720 1130.030 398.470 ;
        RECT 1130.870 395.720 1131.870 398.470 ;
        RECT 1132.710 395.720 1134.170 398.470 ;
        RECT 1135.010 395.720 1136.470 398.470 ;
        RECT 1137.310 395.720 1138.770 398.470 ;
        RECT 1139.610 395.720 1140.610 398.470 ;
        RECT 1141.450 395.720 1142.910 398.470 ;
        RECT 1143.750 395.720 1145.210 398.470 ;
        RECT 1146.050 395.720 1147.050 398.470 ;
        RECT 1147.890 395.720 1149.350 398.470 ;
        RECT 1150.190 395.720 1151.650 398.470 ;
        RECT 1152.490 395.720 1153.950 398.470 ;
        RECT 1154.790 395.720 1155.790 398.470 ;
        RECT 1156.630 395.720 1158.090 398.470 ;
        RECT 1158.930 395.720 1160.390 398.470 ;
        RECT 1161.230 395.720 1162.230 398.470 ;
        RECT 1163.070 395.720 1164.530 398.470 ;
        RECT 1165.370 395.720 1166.830 398.470 ;
        RECT 1167.670 395.720 1168.670 398.470 ;
        RECT 1169.510 395.720 1170.970 398.470 ;
        RECT 1171.810 395.720 1173.270 398.470 ;
        RECT 1174.110 395.720 1175.570 398.470 ;
        RECT 1176.410 395.720 1177.410 398.470 ;
        RECT 1178.250 395.720 1179.710 398.470 ;
        RECT 1180.550 395.720 1182.010 398.470 ;
        RECT 1182.850 395.720 1183.850 398.470 ;
        RECT 1184.690 395.720 1186.150 398.470 ;
        RECT 1186.990 395.720 1188.450 398.470 ;
        RECT 1189.290 395.720 1190.750 398.470 ;
        RECT 1191.590 395.720 1192.590 398.470 ;
        RECT 1193.430 395.720 1194.890 398.470 ;
        RECT 1195.730 395.720 1197.190 398.470 ;
        RECT 1198.030 395.720 1199.030 398.470 ;
        RECT 1199.870 395.720 1201.330 398.470 ;
        RECT 1202.170 395.720 1203.630 398.470 ;
        RECT 1204.470 395.720 1205.930 398.470 ;
        RECT 1206.770 395.720 1207.770 398.470 ;
        RECT 1208.610 395.720 1210.070 398.470 ;
        RECT 1210.910 395.720 1212.370 398.470 ;
        RECT 1213.210 395.720 1214.210 398.470 ;
        RECT 1215.050 395.720 1216.510 398.470 ;
        RECT 1217.350 395.720 1218.810 398.470 ;
        RECT 1219.650 395.720 1221.110 398.470 ;
        RECT 1221.950 395.720 1222.950 398.470 ;
        RECT 1223.790 395.720 1225.250 398.470 ;
        RECT 1226.090 395.720 1227.550 398.470 ;
        RECT 1228.390 395.720 1229.390 398.470 ;
        RECT 1230.230 395.720 1231.690 398.470 ;
        RECT 1232.530 395.720 1233.990 398.470 ;
        RECT 1234.830 395.720 1236.290 398.470 ;
        RECT 1237.130 395.720 1238.130 398.470 ;
        RECT 1238.970 395.720 1240.430 398.470 ;
        RECT 1241.270 395.720 1242.730 398.470 ;
        RECT 1243.570 395.720 1244.570 398.470 ;
        RECT 1245.410 395.720 1246.870 398.470 ;
        RECT 1247.710 395.720 1249.170 398.470 ;
        RECT 1250.010 395.720 1251.470 398.470 ;
        RECT 1252.310 395.720 1253.310 398.470 ;
        RECT 1254.150 395.720 1255.610 398.470 ;
        RECT 1256.450 395.720 1257.910 398.470 ;
        RECT 1258.750 395.720 1259.750 398.470 ;
        RECT 1260.590 395.720 1262.050 398.470 ;
        RECT 1262.890 395.720 1264.350 398.470 ;
        RECT 1265.190 395.720 1266.650 398.470 ;
        RECT 1267.490 395.720 1268.490 398.470 ;
        RECT 1269.330 395.720 1270.790 398.470 ;
        RECT 1271.630 395.720 1273.090 398.470 ;
        RECT 1273.930 395.720 1274.930 398.470 ;
        RECT 1275.770 395.720 1277.230 398.470 ;
        RECT 1278.070 395.720 1279.530 398.470 ;
        RECT 1280.370 395.720 1281.830 398.470 ;
        RECT 1282.670 395.720 1283.670 398.470 ;
        RECT 1284.510 395.720 1285.970 398.470 ;
        RECT 1286.810 395.720 1288.270 398.470 ;
        RECT 1289.110 395.720 1290.110 398.470 ;
        RECT 1290.950 395.720 1292.410 398.470 ;
        RECT 1293.250 395.720 1294.710 398.470 ;
        RECT 1295.550 395.720 1297.010 398.470 ;
        RECT 1297.850 395.720 1298.850 398.470 ;
        RECT 1299.690 395.720 1301.150 398.470 ;
        RECT 1301.990 395.720 1303.450 398.470 ;
        RECT 1304.290 395.720 1305.290 398.470 ;
        RECT 1306.130 395.720 1307.590 398.470 ;
        RECT 1308.430 395.720 1309.890 398.470 ;
        RECT 1310.730 395.720 1312.190 398.470 ;
        RECT 1313.030 395.720 1314.030 398.470 ;
        RECT 1314.870 395.720 1316.330 398.470 ;
        RECT 1317.170 395.720 1318.630 398.470 ;
        RECT 1319.470 395.720 1320.470 398.470 ;
        RECT 1321.310 395.720 1322.770 398.470 ;
        RECT 1323.610 395.720 1325.070 398.470 ;
        RECT 1325.910 395.720 1327.370 398.470 ;
        RECT 1328.210 395.720 1329.210 398.470 ;
        RECT 1330.050 395.720 1331.510 398.470 ;
        RECT 1332.350 395.720 1333.810 398.470 ;
        RECT 1334.650 395.720 1335.650 398.470 ;
        RECT 1336.490 395.720 1337.950 398.470 ;
        RECT 1338.790 395.720 1340.250 398.470 ;
        RECT 1341.090 395.720 1342.090 398.470 ;
        RECT 1342.930 395.720 1344.390 398.470 ;
        RECT 1345.230 395.720 1346.690 398.470 ;
        RECT 1347.530 395.720 1348.990 398.470 ;
        RECT 1349.830 395.720 1350.830 398.470 ;
        RECT 1351.670 395.720 1353.130 398.470 ;
        RECT 1353.970 395.720 1355.430 398.470 ;
        RECT 1356.270 395.720 1357.270 398.470 ;
        RECT 1358.110 395.720 1359.570 398.470 ;
        RECT 1360.410 395.720 1361.870 398.470 ;
        RECT 1362.710 395.720 1364.170 398.470 ;
        RECT 1365.010 395.720 1366.010 398.470 ;
        RECT 1366.850 395.720 1368.310 398.470 ;
        RECT 1369.150 395.720 1370.610 398.470 ;
        RECT 1371.450 395.720 1372.450 398.470 ;
        RECT 1373.290 395.720 1374.750 398.470 ;
        RECT 1375.590 395.720 1377.050 398.470 ;
        RECT 1377.890 395.720 1379.350 398.470 ;
        RECT 1380.190 395.720 1381.190 398.470 ;
        RECT 1382.030 395.720 1383.490 398.470 ;
        RECT 1384.330 395.720 1385.790 398.470 ;
        RECT 1386.630 395.720 1387.630 398.470 ;
        RECT 1388.470 395.720 1389.930 398.470 ;
        RECT 1390.770 395.720 1392.230 398.470 ;
        RECT 1393.070 395.720 1394.530 398.470 ;
        RECT 1395.370 395.720 1396.370 398.470 ;
        RECT 1397.210 395.720 1398.670 398.470 ;
        RECT 1399.510 395.720 1400.970 398.470 ;
        RECT 1401.810 395.720 1402.810 398.470 ;
        RECT 1403.650 395.720 1405.110 398.470 ;
        RECT 1405.950 395.720 1407.410 398.470 ;
        RECT 1408.250 395.720 1409.710 398.470 ;
        RECT 1410.550 395.720 1411.550 398.470 ;
        RECT 1412.390 395.720 1413.850 398.470 ;
        RECT 1414.690 395.720 1416.150 398.470 ;
        RECT 1416.990 395.720 1417.990 398.470 ;
        RECT 1418.830 395.720 1420.290 398.470 ;
        RECT 1421.130 395.720 1422.590 398.470 ;
        RECT 1423.430 395.720 1424.890 398.470 ;
        RECT 1425.730 395.720 1426.730 398.470 ;
        RECT 1427.570 395.720 1429.030 398.470 ;
        RECT 1429.870 395.720 1431.330 398.470 ;
        RECT 1432.170 395.720 1433.170 398.470 ;
        RECT 1434.010 395.720 1435.470 398.470 ;
        RECT 1436.310 395.720 1437.770 398.470 ;
        RECT 1438.610 395.720 1440.070 398.470 ;
        RECT 1440.910 395.720 1441.910 398.470 ;
        RECT 1442.750 395.720 1444.210 398.470 ;
        RECT 1445.050 395.720 1446.510 398.470 ;
        RECT 1447.350 395.720 1448.350 398.470 ;
        RECT 1449.190 395.720 1450.650 398.470 ;
        RECT 1451.490 395.720 1452.950 398.470 ;
        RECT 1453.790 395.720 1455.250 398.470 ;
        RECT 1456.090 395.720 1457.090 398.470 ;
        RECT 1457.930 395.720 1459.390 398.470 ;
        RECT 1460.230 395.720 1461.690 398.470 ;
        RECT 1462.530 395.720 1463.530 398.470 ;
        RECT 1464.370 395.720 1465.830 398.470 ;
        RECT 1466.670 395.720 1468.130 398.470 ;
        RECT 1468.970 395.720 1470.430 398.470 ;
        RECT 1471.270 395.720 1472.270 398.470 ;
        RECT 1473.110 395.720 1474.570 398.470 ;
        RECT 1475.410 395.720 1476.870 398.470 ;
        RECT 1477.710 395.720 1478.710 398.470 ;
        RECT 1479.550 395.720 1481.010 398.470 ;
        RECT 1481.850 395.720 1483.310 398.470 ;
        RECT 1484.150 395.720 1485.610 398.470 ;
        RECT 1486.450 395.720 1487.450 398.470 ;
        RECT 1488.290 395.720 1489.750 398.470 ;
        RECT 1490.590 395.720 1492.050 398.470 ;
        RECT 1492.890 395.720 1493.890 398.470 ;
        RECT 0.100 4.280 1494.380 395.720 ;
        RECT 0.100 2.195 1.190 4.280 ;
        RECT 2.030 2.195 3.950 4.280 ;
        RECT 4.790 2.195 7.170 4.280 ;
        RECT 8.010 2.195 9.930 4.280 ;
        RECT 10.770 2.195 13.150 4.280 ;
        RECT 13.990 2.195 16.370 4.280 ;
        RECT 17.210 2.195 19.130 4.280 ;
        RECT 19.970 2.195 22.350 4.280 ;
        RECT 23.190 2.195 25.570 4.280 ;
        RECT 26.410 2.195 28.330 4.280 ;
        RECT 29.170 2.195 31.550 4.280 ;
        RECT 32.390 2.195 34.770 4.280 ;
        RECT 35.610 2.195 37.530 4.280 ;
        RECT 38.370 2.195 40.750 4.280 ;
        RECT 41.590 2.195 43.510 4.280 ;
        RECT 44.350 2.195 46.730 4.280 ;
        RECT 47.570 2.195 49.950 4.280 ;
        RECT 50.790 2.195 52.710 4.280 ;
        RECT 53.550 2.195 55.930 4.280 ;
        RECT 56.770 2.195 59.150 4.280 ;
        RECT 59.990 2.195 61.910 4.280 ;
        RECT 62.750 2.195 65.130 4.280 ;
        RECT 65.970 2.195 68.350 4.280 ;
        RECT 69.190 2.195 71.110 4.280 ;
        RECT 71.950 2.195 74.330 4.280 ;
        RECT 75.170 2.195 77.550 4.280 ;
        RECT 78.390 2.195 80.310 4.280 ;
        RECT 81.150 2.195 83.530 4.280 ;
        RECT 84.370 2.195 86.290 4.280 ;
        RECT 87.130 2.195 89.510 4.280 ;
        RECT 90.350 2.195 92.730 4.280 ;
        RECT 93.570 2.195 95.490 4.280 ;
        RECT 96.330 2.195 98.710 4.280 ;
        RECT 99.550 2.195 101.930 4.280 ;
        RECT 102.770 2.195 104.690 4.280 ;
        RECT 105.530 2.195 107.910 4.280 ;
        RECT 108.750 2.195 111.130 4.280 ;
        RECT 111.970 2.195 113.890 4.280 ;
        RECT 114.730 2.195 117.110 4.280 ;
        RECT 117.950 2.195 120.330 4.280 ;
        RECT 121.170 2.195 123.090 4.280 ;
        RECT 123.930 2.195 126.310 4.280 ;
        RECT 127.150 2.195 129.070 4.280 ;
        RECT 129.910 2.195 132.290 4.280 ;
        RECT 133.130 2.195 135.510 4.280 ;
        RECT 136.350 2.195 138.270 4.280 ;
        RECT 139.110 2.195 141.490 4.280 ;
        RECT 142.330 2.195 144.710 4.280 ;
        RECT 145.550 2.195 147.470 4.280 ;
        RECT 148.310 2.195 150.690 4.280 ;
        RECT 151.530 2.195 153.910 4.280 ;
        RECT 154.750 2.195 156.670 4.280 ;
        RECT 157.510 2.195 159.890 4.280 ;
        RECT 160.730 2.195 163.110 4.280 ;
        RECT 163.950 2.195 165.870 4.280 ;
        RECT 166.710 2.195 169.090 4.280 ;
        RECT 169.930 2.195 171.850 4.280 ;
        RECT 172.690 2.195 175.070 4.280 ;
        RECT 175.910 2.195 178.290 4.280 ;
        RECT 179.130 2.195 181.050 4.280 ;
        RECT 181.890 2.195 184.270 4.280 ;
        RECT 185.110 2.195 187.490 4.280 ;
        RECT 188.330 2.195 190.250 4.280 ;
        RECT 191.090 2.195 193.470 4.280 ;
        RECT 194.310 2.195 196.690 4.280 ;
        RECT 197.530 2.195 199.450 4.280 ;
        RECT 200.290 2.195 202.670 4.280 ;
        RECT 203.510 2.195 205.430 4.280 ;
        RECT 206.270 2.195 208.650 4.280 ;
        RECT 209.490 2.195 211.870 4.280 ;
        RECT 212.710 2.195 214.630 4.280 ;
        RECT 215.470 2.195 217.850 4.280 ;
        RECT 218.690 2.195 221.070 4.280 ;
        RECT 221.910 2.195 223.830 4.280 ;
        RECT 224.670 2.195 227.050 4.280 ;
        RECT 227.890 2.195 230.270 4.280 ;
        RECT 231.110 2.195 233.030 4.280 ;
        RECT 233.870 2.195 236.250 4.280 ;
        RECT 237.090 2.195 239.470 4.280 ;
        RECT 240.310 2.195 242.230 4.280 ;
        RECT 243.070 2.195 245.450 4.280 ;
        RECT 246.290 2.195 248.210 4.280 ;
        RECT 249.050 2.195 251.430 4.280 ;
        RECT 252.270 2.195 254.650 4.280 ;
        RECT 255.490 2.195 257.410 4.280 ;
        RECT 258.250 2.195 260.630 4.280 ;
        RECT 261.470 2.195 263.850 4.280 ;
        RECT 264.690 2.195 266.610 4.280 ;
        RECT 267.450 2.195 269.830 4.280 ;
        RECT 270.670 2.195 273.050 4.280 ;
        RECT 273.890 2.195 275.810 4.280 ;
        RECT 276.650 2.195 279.030 4.280 ;
        RECT 279.870 2.195 282.250 4.280 ;
        RECT 283.090 2.195 285.010 4.280 ;
        RECT 285.850 2.195 288.230 4.280 ;
        RECT 289.070 2.195 290.990 4.280 ;
        RECT 291.830 2.195 294.210 4.280 ;
        RECT 295.050 2.195 297.430 4.280 ;
        RECT 298.270 2.195 300.190 4.280 ;
        RECT 301.030 2.195 303.410 4.280 ;
        RECT 304.250 2.195 306.630 4.280 ;
        RECT 307.470 2.195 309.390 4.280 ;
        RECT 310.230 2.195 312.610 4.280 ;
        RECT 313.450 2.195 315.830 4.280 ;
        RECT 316.670 2.195 318.590 4.280 ;
        RECT 319.430 2.195 321.810 4.280 ;
        RECT 322.650 2.195 325.030 4.280 ;
        RECT 325.870 2.195 327.790 4.280 ;
        RECT 328.630 2.195 331.010 4.280 ;
        RECT 331.850 2.195 333.770 4.280 ;
        RECT 334.610 2.195 336.990 4.280 ;
        RECT 337.830 2.195 340.210 4.280 ;
        RECT 341.050 2.195 342.970 4.280 ;
        RECT 343.810 2.195 346.190 4.280 ;
        RECT 347.030 2.195 349.410 4.280 ;
        RECT 350.250 2.195 352.170 4.280 ;
        RECT 353.010 2.195 355.390 4.280 ;
        RECT 356.230 2.195 358.610 4.280 ;
        RECT 359.450 2.195 361.370 4.280 ;
        RECT 362.210 2.195 364.590 4.280 ;
        RECT 365.430 2.195 367.350 4.280 ;
        RECT 368.190 2.195 370.570 4.280 ;
        RECT 371.410 2.195 373.790 4.280 ;
        RECT 374.630 2.195 376.550 4.280 ;
        RECT 377.390 2.195 379.770 4.280 ;
        RECT 380.610 2.195 382.990 4.280 ;
        RECT 383.830 2.195 385.750 4.280 ;
        RECT 386.590 2.195 388.970 4.280 ;
        RECT 389.810 2.195 392.190 4.280 ;
        RECT 393.030 2.195 394.950 4.280 ;
        RECT 395.790 2.195 398.170 4.280 ;
        RECT 399.010 2.195 401.390 4.280 ;
        RECT 402.230 2.195 404.150 4.280 ;
        RECT 404.990 2.195 407.370 4.280 ;
        RECT 408.210 2.195 410.130 4.280 ;
        RECT 410.970 2.195 413.350 4.280 ;
        RECT 414.190 2.195 416.570 4.280 ;
        RECT 417.410 2.195 419.330 4.280 ;
        RECT 420.170 2.195 422.550 4.280 ;
        RECT 423.390 2.195 425.770 4.280 ;
        RECT 426.610 2.195 428.530 4.280 ;
        RECT 429.370 2.195 431.750 4.280 ;
        RECT 432.590 2.195 434.970 4.280 ;
        RECT 435.810 2.195 437.730 4.280 ;
        RECT 438.570 2.195 440.950 4.280 ;
        RECT 441.790 2.195 444.170 4.280 ;
        RECT 445.010 2.195 446.930 4.280 ;
        RECT 447.770 2.195 450.150 4.280 ;
        RECT 450.990 2.195 452.910 4.280 ;
        RECT 453.750 2.195 456.130 4.280 ;
        RECT 456.970 2.195 459.350 4.280 ;
        RECT 460.190 2.195 462.110 4.280 ;
        RECT 462.950 2.195 465.330 4.280 ;
        RECT 466.170 2.195 468.550 4.280 ;
        RECT 469.390 2.195 471.310 4.280 ;
        RECT 472.150 2.195 474.530 4.280 ;
        RECT 475.370 2.195 477.750 4.280 ;
        RECT 478.590 2.195 480.510 4.280 ;
        RECT 481.350 2.195 483.730 4.280 ;
        RECT 484.570 2.195 486.950 4.280 ;
        RECT 487.790 2.195 489.710 4.280 ;
        RECT 490.550 2.195 492.930 4.280 ;
        RECT 493.770 2.195 495.690 4.280 ;
        RECT 496.530 2.195 498.910 4.280 ;
        RECT 499.750 2.195 502.130 4.280 ;
        RECT 502.970 2.195 504.890 4.280 ;
        RECT 505.730 2.195 508.110 4.280 ;
        RECT 508.950 2.195 511.330 4.280 ;
        RECT 512.170 2.195 514.090 4.280 ;
        RECT 514.930 2.195 517.310 4.280 ;
        RECT 518.150 2.195 520.530 4.280 ;
        RECT 521.370 2.195 523.290 4.280 ;
        RECT 524.130 2.195 526.510 4.280 ;
        RECT 527.350 2.195 529.270 4.280 ;
        RECT 530.110 2.195 532.490 4.280 ;
        RECT 533.330 2.195 535.710 4.280 ;
        RECT 536.550 2.195 538.470 4.280 ;
        RECT 539.310 2.195 541.690 4.280 ;
        RECT 542.530 2.195 544.910 4.280 ;
        RECT 545.750 2.195 547.670 4.280 ;
        RECT 548.510 2.195 550.890 4.280 ;
        RECT 551.730 2.195 554.110 4.280 ;
        RECT 554.950 2.195 556.870 4.280 ;
        RECT 557.710 2.195 560.090 4.280 ;
        RECT 560.930 2.195 563.310 4.280 ;
        RECT 564.150 2.195 566.070 4.280 ;
        RECT 566.910 2.195 569.290 4.280 ;
        RECT 570.130 2.195 572.050 4.280 ;
        RECT 572.890 2.195 575.270 4.280 ;
        RECT 576.110 2.195 578.490 4.280 ;
        RECT 579.330 2.195 581.250 4.280 ;
        RECT 582.090 2.195 584.470 4.280 ;
        RECT 585.310 2.195 587.690 4.280 ;
        RECT 588.530 2.195 590.450 4.280 ;
        RECT 591.290 2.195 593.670 4.280 ;
        RECT 594.510 2.195 596.890 4.280 ;
        RECT 597.730 2.195 599.650 4.280 ;
        RECT 600.490 2.195 602.870 4.280 ;
        RECT 603.710 2.195 606.090 4.280 ;
        RECT 606.930 2.195 608.850 4.280 ;
        RECT 609.690 2.195 612.070 4.280 ;
        RECT 612.910 2.195 614.830 4.280 ;
        RECT 615.670 2.195 618.050 4.280 ;
        RECT 618.890 2.195 621.270 4.280 ;
        RECT 622.110 2.195 624.030 4.280 ;
        RECT 624.870 2.195 627.250 4.280 ;
        RECT 628.090 2.195 630.470 4.280 ;
        RECT 631.310 2.195 633.230 4.280 ;
        RECT 634.070 2.195 636.450 4.280 ;
        RECT 637.290 2.195 639.670 4.280 ;
        RECT 640.510 2.195 642.430 4.280 ;
        RECT 643.270 2.195 645.650 4.280 ;
        RECT 646.490 2.195 648.870 4.280 ;
        RECT 649.710 2.195 651.630 4.280 ;
        RECT 652.470 2.195 654.850 4.280 ;
        RECT 655.690 2.195 657.610 4.280 ;
        RECT 658.450 2.195 660.830 4.280 ;
        RECT 661.670 2.195 664.050 4.280 ;
        RECT 664.890 2.195 666.810 4.280 ;
        RECT 667.650 2.195 670.030 4.280 ;
        RECT 670.870 2.195 673.250 4.280 ;
        RECT 674.090 2.195 676.010 4.280 ;
        RECT 676.850 2.195 679.230 4.280 ;
        RECT 680.070 2.195 682.450 4.280 ;
        RECT 683.290 2.195 685.210 4.280 ;
        RECT 686.050 2.195 688.430 4.280 ;
        RECT 689.270 2.195 691.190 4.280 ;
        RECT 692.030 2.195 694.410 4.280 ;
        RECT 695.250 2.195 697.630 4.280 ;
        RECT 698.470 2.195 700.390 4.280 ;
        RECT 701.230 2.195 703.610 4.280 ;
        RECT 704.450 2.195 706.830 4.280 ;
        RECT 707.670 2.195 709.590 4.280 ;
        RECT 710.430 2.195 712.810 4.280 ;
        RECT 713.650 2.195 716.030 4.280 ;
        RECT 716.870 2.195 718.790 4.280 ;
        RECT 719.630 2.195 722.010 4.280 ;
        RECT 722.850 2.195 725.230 4.280 ;
        RECT 726.070 2.195 727.990 4.280 ;
        RECT 728.830 2.195 731.210 4.280 ;
        RECT 732.050 2.195 733.970 4.280 ;
        RECT 734.810 2.195 737.190 4.280 ;
        RECT 738.030 2.195 740.410 4.280 ;
        RECT 741.250 2.195 743.170 4.280 ;
        RECT 744.010 2.195 746.390 4.280 ;
        RECT 747.230 2.195 749.610 4.280 ;
        RECT 750.450 2.195 752.370 4.280 ;
        RECT 753.210 2.195 755.590 4.280 ;
        RECT 756.430 2.195 758.810 4.280 ;
        RECT 759.650 2.195 761.570 4.280 ;
        RECT 762.410 2.195 764.790 4.280 ;
        RECT 765.630 2.195 768.010 4.280 ;
        RECT 768.850 2.195 770.770 4.280 ;
        RECT 771.610 2.195 773.990 4.280 ;
        RECT 774.830 2.195 776.750 4.280 ;
        RECT 777.590 2.195 779.970 4.280 ;
        RECT 780.810 2.195 783.190 4.280 ;
        RECT 784.030 2.195 785.950 4.280 ;
        RECT 786.790 2.195 789.170 4.280 ;
        RECT 790.010 2.195 792.390 4.280 ;
        RECT 793.230 2.195 795.150 4.280 ;
        RECT 795.990 2.195 798.370 4.280 ;
        RECT 799.210 2.195 801.590 4.280 ;
        RECT 802.430 2.195 804.350 4.280 ;
        RECT 805.190 2.195 807.570 4.280 ;
        RECT 808.410 2.195 810.790 4.280 ;
        RECT 811.630 2.195 813.550 4.280 ;
        RECT 814.390 2.195 816.770 4.280 ;
        RECT 817.610 2.195 819.530 4.280 ;
        RECT 820.370 2.195 822.750 4.280 ;
        RECT 823.590 2.195 825.970 4.280 ;
        RECT 826.810 2.195 828.730 4.280 ;
        RECT 829.570 2.195 831.950 4.280 ;
        RECT 832.790 2.195 835.170 4.280 ;
        RECT 836.010 2.195 837.930 4.280 ;
        RECT 838.770 2.195 841.150 4.280 ;
        RECT 841.990 2.195 844.370 4.280 ;
        RECT 845.210 2.195 847.130 4.280 ;
        RECT 847.970 2.195 850.350 4.280 ;
        RECT 851.190 2.195 853.110 4.280 ;
        RECT 853.950 2.195 856.330 4.280 ;
        RECT 857.170 2.195 859.550 4.280 ;
        RECT 860.390 2.195 862.310 4.280 ;
        RECT 863.150 2.195 865.530 4.280 ;
        RECT 866.370 2.195 868.750 4.280 ;
        RECT 869.590 2.195 871.510 4.280 ;
        RECT 872.350 2.195 874.730 4.280 ;
        RECT 875.570 2.195 877.950 4.280 ;
        RECT 878.790 2.195 880.710 4.280 ;
        RECT 881.550 2.195 883.930 4.280 ;
        RECT 884.770 2.195 887.150 4.280 ;
        RECT 887.990 2.195 889.910 4.280 ;
        RECT 890.750 2.195 893.130 4.280 ;
        RECT 893.970 2.195 895.890 4.280 ;
        RECT 896.730 2.195 899.110 4.280 ;
        RECT 899.950 2.195 902.330 4.280 ;
        RECT 903.170 2.195 905.090 4.280 ;
        RECT 905.930 2.195 908.310 4.280 ;
        RECT 909.150 2.195 911.530 4.280 ;
        RECT 912.370 2.195 914.290 4.280 ;
        RECT 915.130 2.195 917.510 4.280 ;
        RECT 918.350 2.195 920.730 4.280 ;
        RECT 921.570 2.195 923.490 4.280 ;
        RECT 924.330 2.195 926.710 4.280 ;
        RECT 927.550 2.195 929.930 4.280 ;
        RECT 930.770 2.195 932.690 4.280 ;
        RECT 933.530 2.195 935.910 4.280 ;
        RECT 936.750 2.195 938.670 4.280 ;
        RECT 939.510 2.195 941.890 4.280 ;
        RECT 942.730 2.195 945.110 4.280 ;
        RECT 945.950 2.195 947.870 4.280 ;
        RECT 948.710 2.195 951.090 4.280 ;
        RECT 951.930 2.195 954.310 4.280 ;
        RECT 955.150 2.195 957.070 4.280 ;
        RECT 957.910 2.195 960.290 4.280 ;
        RECT 961.130 2.195 963.510 4.280 ;
        RECT 964.350 2.195 966.270 4.280 ;
        RECT 967.110 2.195 969.490 4.280 ;
        RECT 970.330 2.195 972.710 4.280 ;
        RECT 973.550 2.195 975.470 4.280 ;
        RECT 976.310 2.195 978.690 4.280 ;
        RECT 979.530 2.195 981.450 4.280 ;
        RECT 982.290 2.195 984.670 4.280 ;
        RECT 985.510 2.195 987.890 4.280 ;
        RECT 988.730 2.195 990.650 4.280 ;
        RECT 991.490 2.195 993.870 4.280 ;
        RECT 994.710 2.195 997.090 4.280 ;
        RECT 997.930 2.195 999.850 4.280 ;
        RECT 1000.690 2.195 1003.070 4.280 ;
        RECT 1003.910 2.195 1006.290 4.280 ;
        RECT 1007.130 2.195 1009.050 4.280 ;
        RECT 1009.890 2.195 1012.270 4.280 ;
        RECT 1013.110 2.195 1015.030 4.280 ;
        RECT 1015.870 2.195 1018.250 4.280 ;
        RECT 1019.090 2.195 1021.470 4.280 ;
        RECT 1022.310 2.195 1024.230 4.280 ;
        RECT 1025.070 2.195 1027.450 4.280 ;
        RECT 1028.290 2.195 1030.670 4.280 ;
        RECT 1031.510 2.195 1033.430 4.280 ;
        RECT 1034.270 2.195 1036.650 4.280 ;
        RECT 1037.490 2.195 1039.870 4.280 ;
        RECT 1040.710 2.195 1042.630 4.280 ;
        RECT 1043.470 2.195 1045.850 4.280 ;
        RECT 1046.690 2.195 1049.070 4.280 ;
        RECT 1049.910 2.195 1051.830 4.280 ;
        RECT 1052.670 2.195 1055.050 4.280 ;
        RECT 1055.890 2.195 1057.810 4.280 ;
        RECT 1058.650 2.195 1061.030 4.280 ;
        RECT 1061.870 2.195 1064.250 4.280 ;
        RECT 1065.090 2.195 1067.010 4.280 ;
        RECT 1067.850 2.195 1070.230 4.280 ;
        RECT 1071.070 2.195 1073.450 4.280 ;
        RECT 1074.290 2.195 1076.210 4.280 ;
        RECT 1077.050 2.195 1079.430 4.280 ;
        RECT 1080.270 2.195 1082.650 4.280 ;
        RECT 1083.490 2.195 1085.410 4.280 ;
        RECT 1086.250 2.195 1088.630 4.280 ;
        RECT 1089.470 2.195 1091.850 4.280 ;
        RECT 1092.690 2.195 1094.610 4.280 ;
        RECT 1095.450 2.195 1097.830 4.280 ;
        RECT 1098.670 2.195 1100.590 4.280 ;
        RECT 1101.430 2.195 1103.810 4.280 ;
        RECT 1104.650 2.195 1107.030 4.280 ;
        RECT 1107.870 2.195 1109.790 4.280 ;
        RECT 1110.630 2.195 1113.010 4.280 ;
        RECT 1113.850 2.195 1116.230 4.280 ;
        RECT 1117.070 2.195 1118.990 4.280 ;
        RECT 1119.830 2.195 1122.210 4.280 ;
        RECT 1123.050 2.195 1125.430 4.280 ;
        RECT 1126.270 2.195 1128.190 4.280 ;
        RECT 1129.030 2.195 1131.410 4.280 ;
        RECT 1132.250 2.195 1134.630 4.280 ;
        RECT 1135.470 2.195 1137.390 4.280 ;
        RECT 1138.230 2.195 1140.610 4.280 ;
        RECT 1141.450 2.195 1143.370 4.280 ;
        RECT 1144.210 2.195 1146.590 4.280 ;
        RECT 1147.430 2.195 1149.810 4.280 ;
        RECT 1150.650 2.195 1152.570 4.280 ;
        RECT 1153.410 2.195 1155.790 4.280 ;
        RECT 1156.630 2.195 1159.010 4.280 ;
        RECT 1159.850 2.195 1161.770 4.280 ;
        RECT 1162.610 2.195 1164.990 4.280 ;
        RECT 1165.830 2.195 1168.210 4.280 ;
        RECT 1169.050 2.195 1170.970 4.280 ;
        RECT 1171.810 2.195 1174.190 4.280 ;
        RECT 1175.030 2.195 1176.950 4.280 ;
        RECT 1177.790 2.195 1180.170 4.280 ;
        RECT 1181.010 2.195 1183.390 4.280 ;
        RECT 1184.230 2.195 1186.150 4.280 ;
        RECT 1186.990 2.195 1189.370 4.280 ;
        RECT 1190.210 2.195 1192.590 4.280 ;
        RECT 1193.430 2.195 1195.350 4.280 ;
        RECT 1196.190 2.195 1198.570 4.280 ;
        RECT 1199.410 2.195 1201.790 4.280 ;
        RECT 1202.630 2.195 1204.550 4.280 ;
        RECT 1205.390 2.195 1207.770 4.280 ;
        RECT 1208.610 2.195 1210.990 4.280 ;
        RECT 1211.830 2.195 1213.750 4.280 ;
        RECT 1214.590 2.195 1216.970 4.280 ;
        RECT 1217.810 2.195 1219.730 4.280 ;
        RECT 1220.570 2.195 1222.950 4.280 ;
        RECT 1223.790 2.195 1226.170 4.280 ;
        RECT 1227.010 2.195 1228.930 4.280 ;
        RECT 1229.770 2.195 1232.150 4.280 ;
        RECT 1232.990 2.195 1235.370 4.280 ;
        RECT 1236.210 2.195 1238.130 4.280 ;
        RECT 1238.970 2.195 1241.350 4.280 ;
        RECT 1242.190 2.195 1244.570 4.280 ;
        RECT 1245.410 2.195 1247.330 4.280 ;
        RECT 1248.170 2.195 1250.550 4.280 ;
        RECT 1251.390 2.195 1253.770 4.280 ;
        RECT 1254.610 2.195 1256.530 4.280 ;
        RECT 1257.370 2.195 1259.750 4.280 ;
        RECT 1260.590 2.195 1262.510 4.280 ;
        RECT 1263.350 2.195 1265.730 4.280 ;
        RECT 1266.570 2.195 1268.950 4.280 ;
        RECT 1269.790 2.195 1271.710 4.280 ;
        RECT 1272.550 2.195 1274.930 4.280 ;
        RECT 1275.770 2.195 1278.150 4.280 ;
        RECT 1278.990 2.195 1280.910 4.280 ;
        RECT 1281.750 2.195 1284.130 4.280 ;
        RECT 1284.970 2.195 1287.350 4.280 ;
        RECT 1288.190 2.195 1290.110 4.280 ;
        RECT 1290.950 2.195 1293.330 4.280 ;
        RECT 1294.170 2.195 1296.550 4.280 ;
        RECT 1297.390 2.195 1299.310 4.280 ;
        RECT 1300.150 2.195 1302.530 4.280 ;
        RECT 1303.370 2.195 1305.290 4.280 ;
        RECT 1306.130 2.195 1308.510 4.280 ;
        RECT 1309.350 2.195 1311.730 4.280 ;
        RECT 1312.570 2.195 1314.490 4.280 ;
        RECT 1315.330 2.195 1317.710 4.280 ;
        RECT 1318.550 2.195 1320.930 4.280 ;
        RECT 1321.770 2.195 1323.690 4.280 ;
        RECT 1324.530 2.195 1326.910 4.280 ;
        RECT 1327.750 2.195 1330.130 4.280 ;
        RECT 1330.970 2.195 1332.890 4.280 ;
        RECT 1333.730 2.195 1336.110 4.280 ;
        RECT 1336.950 2.195 1338.870 4.280 ;
        RECT 1339.710 2.195 1342.090 4.280 ;
        RECT 1342.930 2.195 1345.310 4.280 ;
        RECT 1346.150 2.195 1348.070 4.280 ;
        RECT 1348.910 2.195 1351.290 4.280 ;
        RECT 1352.130 2.195 1354.510 4.280 ;
        RECT 1355.350 2.195 1357.270 4.280 ;
        RECT 1358.110 2.195 1360.490 4.280 ;
        RECT 1361.330 2.195 1363.710 4.280 ;
        RECT 1364.550 2.195 1366.470 4.280 ;
        RECT 1367.310 2.195 1369.690 4.280 ;
        RECT 1370.530 2.195 1372.910 4.280 ;
        RECT 1373.750 2.195 1375.670 4.280 ;
        RECT 1376.510 2.195 1378.890 4.280 ;
        RECT 1379.730 2.195 1381.650 4.280 ;
        RECT 1382.490 2.195 1384.870 4.280 ;
        RECT 1385.710 2.195 1388.090 4.280 ;
        RECT 1388.930 2.195 1390.850 4.280 ;
        RECT 1391.690 2.195 1394.070 4.280 ;
        RECT 1394.910 2.195 1397.290 4.280 ;
        RECT 1398.130 2.195 1400.050 4.280 ;
        RECT 1400.890 2.195 1403.270 4.280 ;
        RECT 1404.110 2.195 1406.490 4.280 ;
        RECT 1407.330 2.195 1409.250 4.280 ;
        RECT 1410.090 2.195 1412.470 4.280 ;
        RECT 1413.310 2.195 1415.690 4.280 ;
        RECT 1416.530 2.195 1418.450 4.280 ;
        RECT 1419.290 2.195 1421.670 4.280 ;
        RECT 1422.510 2.195 1424.430 4.280 ;
        RECT 1425.270 2.195 1427.650 4.280 ;
        RECT 1428.490 2.195 1430.870 4.280 ;
        RECT 1431.710 2.195 1433.630 4.280 ;
        RECT 1434.470 2.195 1436.850 4.280 ;
        RECT 1437.690 2.195 1440.070 4.280 ;
        RECT 1440.910 2.195 1442.830 4.280 ;
        RECT 1443.670 2.195 1446.050 4.280 ;
        RECT 1446.890 2.195 1449.270 4.280 ;
        RECT 1450.110 2.195 1452.030 4.280 ;
        RECT 1452.870 2.195 1455.250 4.280 ;
        RECT 1456.090 2.195 1458.470 4.280 ;
        RECT 1459.310 2.195 1461.230 4.280 ;
        RECT 1462.070 2.195 1464.450 4.280 ;
        RECT 1465.290 2.195 1467.210 4.280 ;
        RECT 1468.050 2.195 1470.430 4.280 ;
        RECT 1471.270 2.195 1473.650 4.280 ;
        RECT 1474.490 2.195 1476.410 4.280 ;
        RECT 1477.250 2.195 1479.630 4.280 ;
        RECT 1480.470 2.195 1482.850 4.280 ;
        RECT 1483.690 2.195 1485.610 4.280 ;
        RECT 1486.450 2.195 1488.830 4.280 ;
        RECT 1489.670 2.195 1492.050 4.280 ;
        RECT 1492.890 2.195 1494.380 4.280 ;
      LAYER met3 ;
        RECT 4.000 392.720 1496.000 392.865 ;
        RECT 4.400 391.320 1496.000 392.720 ;
        RECT 4.000 387.280 1496.000 391.320 ;
        RECT 4.400 385.880 1496.000 387.280 ;
        RECT 4.000 385.240 1496.000 385.880 ;
        RECT 4.000 383.840 1495.600 385.240 ;
        RECT 4.000 382.520 1496.000 383.840 ;
        RECT 4.400 381.120 1496.000 382.520 ;
        RECT 4.000 377.080 1496.000 381.120 ;
        RECT 4.400 375.680 1496.000 377.080 ;
        RECT 4.000 375.040 1496.000 375.680 ;
        RECT 4.000 373.640 1495.600 375.040 ;
        RECT 4.000 372.320 1496.000 373.640 ;
        RECT 4.400 370.920 1496.000 372.320 ;
        RECT 4.000 366.880 1496.000 370.920 ;
        RECT 4.400 365.520 1496.000 366.880 ;
        RECT 4.400 365.480 1495.600 365.520 ;
        RECT 4.000 364.120 1495.600 365.480 ;
        RECT 4.000 362.120 1496.000 364.120 ;
        RECT 4.400 360.720 1496.000 362.120 ;
        RECT 4.000 357.360 1496.000 360.720 ;
        RECT 4.400 355.960 1496.000 357.360 ;
        RECT 4.000 355.320 1496.000 355.960 ;
        RECT 4.000 353.920 1495.600 355.320 ;
        RECT 4.000 351.920 1496.000 353.920 ;
        RECT 4.400 350.520 1496.000 351.920 ;
        RECT 4.000 347.160 1496.000 350.520 ;
        RECT 4.400 345.760 1496.000 347.160 ;
        RECT 4.000 345.120 1496.000 345.760 ;
        RECT 4.000 343.720 1495.600 345.120 ;
        RECT 4.000 341.720 1496.000 343.720 ;
        RECT 4.400 340.320 1496.000 341.720 ;
        RECT 4.000 336.960 1496.000 340.320 ;
        RECT 4.400 335.600 1496.000 336.960 ;
        RECT 4.400 335.560 1495.600 335.600 ;
        RECT 4.000 334.200 1495.600 335.560 ;
        RECT 4.000 331.520 1496.000 334.200 ;
        RECT 4.400 330.120 1496.000 331.520 ;
        RECT 4.000 326.760 1496.000 330.120 ;
        RECT 4.400 325.400 1496.000 326.760 ;
        RECT 4.400 325.360 1495.600 325.400 ;
        RECT 4.000 324.000 1495.600 325.360 ;
        RECT 4.000 321.320 1496.000 324.000 ;
        RECT 4.400 319.920 1496.000 321.320 ;
        RECT 4.000 316.560 1496.000 319.920 ;
        RECT 4.400 315.200 1496.000 316.560 ;
        RECT 4.400 315.160 1495.600 315.200 ;
        RECT 4.000 313.800 1495.600 315.160 ;
        RECT 4.000 311.800 1496.000 313.800 ;
        RECT 4.400 310.400 1496.000 311.800 ;
        RECT 4.000 306.360 1496.000 310.400 ;
        RECT 4.400 305.680 1496.000 306.360 ;
        RECT 4.400 304.960 1495.600 305.680 ;
        RECT 4.000 304.280 1495.600 304.960 ;
        RECT 4.000 301.600 1496.000 304.280 ;
        RECT 4.400 300.200 1496.000 301.600 ;
        RECT 4.000 296.160 1496.000 300.200 ;
        RECT 4.400 295.480 1496.000 296.160 ;
        RECT 4.400 294.760 1495.600 295.480 ;
        RECT 4.000 294.080 1495.600 294.760 ;
        RECT 4.000 291.400 1496.000 294.080 ;
        RECT 4.400 290.000 1496.000 291.400 ;
        RECT 4.000 285.960 1496.000 290.000 ;
        RECT 4.400 285.280 1496.000 285.960 ;
        RECT 4.400 284.560 1495.600 285.280 ;
        RECT 4.000 283.880 1495.600 284.560 ;
        RECT 4.000 281.200 1496.000 283.880 ;
        RECT 4.400 279.800 1496.000 281.200 ;
        RECT 4.000 275.760 1496.000 279.800 ;
        RECT 4.400 275.080 1496.000 275.760 ;
        RECT 4.400 274.360 1495.600 275.080 ;
        RECT 4.000 273.680 1495.600 274.360 ;
        RECT 4.000 271.000 1496.000 273.680 ;
        RECT 4.400 269.600 1496.000 271.000 ;
        RECT 4.000 266.240 1496.000 269.600 ;
        RECT 4.400 265.560 1496.000 266.240 ;
        RECT 4.400 264.840 1495.600 265.560 ;
        RECT 4.000 264.160 1495.600 264.840 ;
        RECT 4.000 260.800 1496.000 264.160 ;
        RECT 4.400 259.400 1496.000 260.800 ;
        RECT 4.000 256.040 1496.000 259.400 ;
        RECT 4.400 255.360 1496.000 256.040 ;
        RECT 4.400 254.640 1495.600 255.360 ;
        RECT 4.000 253.960 1495.600 254.640 ;
        RECT 4.000 250.600 1496.000 253.960 ;
        RECT 4.400 249.200 1496.000 250.600 ;
        RECT 4.000 245.840 1496.000 249.200 ;
        RECT 4.400 245.160 1496.000 245.840 ;
        RECT 4.400 244.440 1495.600 245.160 ;
        RECT 4.000 243.760 1495.600 244.440 ;
        RECT 4.000 240.400 1496.000 243.760 ;
        RECT 4.400 239.000 1496.000 240.400 ;
        RECT 4.000 235.640 1496.000 239.000 ;
        RECT 4.400 234.240 1495.600 235.640 ;
        RECT 4.000 230.200 1496.000 234.240 ;
        RECT 4.400 228.800 1496.000 230.200 ;
        RECT 4.000 225.440 1496.000 228.800 ;
        RECT 4.400 224.040 1495.600 225.440 ;
        RECT 4.000 220.680 1496.000 224.040 ;
        RECT 4.400 219.280 1496.000 220.680 ;
        RECT 4.000 215.240 1496.000 219.280 ;
        RECT 4.400 213.840 1495.600 215.240 ;
        RECT 4.000 210.480 1496.000 213.840 ;
        RECT 4.400 209.080 1496.000 210.480 ;
        RECT 4.000 205.720 1496.000 209.080 ;
        RECT 4.000 205.040 1495.600 205.720 ;
        RECT 4.400 204.320 1495.600 205.040 ;
        RECT 4.400 203.640 1496.000 204.320 ;
        RECT 4.000 200.280 1496.000 203.640 ;
        RECT 4.400 198.880 1496.000 200.280 ;
        RECT 4.000 195.520 1496.000 198.880 ;
        RECT 4.000 194.840 1495.600 195.520 ;
        RECT 4.400 194.120 1495.600 194.840 ;
        RECT 4.400 193.440 1496.000 194.120 ;
        RECT 4.000 190.080 1496.000 193.440 ;
        RECT 4.400 188.680 1496.000 190.080 ;
        RECT 4.000 185.320 1496.000 188.680 ;
        RECT 4.000 184.640 1495.600 185.320 ;
        RECT 4.400 183.920 1495.600 184.640 ;
        RECT 4.400 183.240 1496.000 183.920 ;
        RECT 4.000 179.880 1496.000 183.240 ;
        RECT 4.400 178.480 1496.000 179.880 ;
        RECT 4.000 175.120 1496.000 178.480 ;
        RECT 4.400 173.720 1495.600 175.120 ;
        RECT 4.000 169.680 1496.000 173.720 ;
        RECT 4.400 168.280 1496.000 169.680 ;
        RECT 4.000 165.600 1496.000 168.280 ;
        RECT 4.000 164.920 1495.600 165.600 ;
        RECT 4.400 164.200 1495.600 164.920 ;
        RECT 4.400 163.520 1496.000 164.200 ;
        RECT 4.000 159.480 1496.000 163.520 ;
        RECT 4.400 158.080 1496.000 159.480 ;
        RECT 4.000 155.400 1496.000 158.080 ;
        RECT 4.000 154.720 1495.600 155.400 ;
        RECT 4.400 154.000 1495.600 154.720 ;
        RECT 4.400 153.320 1496.000 154.000 ;
        RECT 4.000 149.280 1496.000 153.320 ;
        RECT 4.400 147.880 1496.000 149.280 ;
        RECT 4.000 145.200 1496.000 147.880 ;
        RECT 4.000 144.520 1495.600 145.200 ;
        RECT 4.400 143.800 1495.600 144.520 ;
        RECT 4.400 143.120 1496.000 143.800 ;
        RECT 4.000 139.080 1496.000 143.120 ;
        RECT 4.400 137.680 1496.000 139.080 ;
        RECT 4.000 135.680 1496.000 137.680 ;
        RECT 4.000 134.320 1495.600 135.680 ;
        RECT 4.400 134.280 1495.600 134.320 ;
        RECT 4.400 132.920 1496.000 134.280 ;
        RECT 4.000 129.560 1496.000 132.920 ;
        RECT 4.400 128.160 1496.000 129.560 ;
        RECT 4.000 125.480 1496.000 128.160 ;
        RECT 4.000 124.120 1495.600 125.480 ;
        RECT 4.400 124.080 1495.600 124.120 ;
        RECT 4.400 122.720 1496.000 124.080 ;
        RECT 4.000 119.360 1496.000 122.720 ;
        RECT 4.400 117.960 1496.000 119.360 ;
        RECT 4.000 115.280 1496.000 117.960 ;
        RECT 4.000 113.920 1495.600 115.280 ;
        RECT 4.400 113.880 1495.600 113.920 ;
        RECT 4.400 112.520 1496.000 113.880 ;
        RECT 4.000 109.160 1496.000 112.520 ;
        RECT 4.400 107.760 1496.000 109.160 ;
        RECT 4.000 105.760 1496.000 107.760 ;
        RECT 4.000 104.360 1495.600 105.760 ;
        RECT 4.000 103.720 1496.000 104.360 ;
        RECT 4.400 102.320 1496.000 103.720 ;
        RECT 4.000 98.960 1496.000 102.320 ;
        RECT 4.400 97.560 1496.000 98.960 ;
        RECT 4.000 95.560 1496.000 97.560 ;
        RECT 4.000 94.160 1495.600 95.560 ;
        RECT 4.000 93.520 1496.000 94.160 ;
        RECT 4.400 92.120 1496.000 93.520 ;
        RECT 4.000 88.760 1496.000 92.120 ;
        RECT 4.400 87.360 1496.000 88.760 ;
        RECT 4.000 85.360 1496.000 87.360 ;
        RECT 4.000 84.000 1495.600 85.360 ;
        RECT 4.400 83.960 1495.600 84.000 ;
        RECT 4.400 82.600 1496.000 83.960 ;
        RECT 4.000 78.560 1496.000 82.600 ;
        RECT 4.400 77.160 1496.000 78.560 ;
        RECT 4.000 75.160 1496.000 77.160 ;
        RECT 4.000 73.800 1495.600 75.160 ;
        RECT 4.400 73.760 1495.600 73.800 ;
        RECT 4.400 72.400 1496.000 73.760 ;
        RECT 4.000 68.360 1496.000 72.400 ;
        RECT 4.400 66.960 1496.000 68.360 ;
        RECT 4.000 65.640 1496.000 66.960 ;
        RECT 4.000 64.240 1495.600 65.640 ;
        RECT 4.000 63.600 1496.000 64.240 ;
        RECT 4.400 62.200 1496.000 63.600 ;
        RECT 4.000 58.160 1496.000 62.200 ;
        RECT 4.400 56.760 1496.000 58.160 ;
        RECT 4.000 55.440 1496.000 56.760 ;
        RECT 4.000 54.040 1495.600 55.440 ;
        RECT 4.000 53.400 1496.000 54.040 ;
        RECT 4.400 52.000 1496.000 53.400 ;
        RECT 4.000 47.960 1496.000 52.000 ;
        RECT 4.400 46.560 1496.000 47.960 ;
        RECT 4.000 45.240 1496.000 46.560 ;
        RECT 4.000 43.840 1495.600 45.240 ;
        RECT 4.000 43.200 1496.000 43.840 ;
        RECT 4.400 41.800 1496.000 43.200 ;
        RECT 4.000 38.440 1496.000 41.800 ;
        RECT 4.400 37.040 1496.000 38.440 ;
        RECT 4.000 35.720 1496.000 37.040 ;
        RECT 4.000 34.320 1495.600 35.720 ;
        RECT 4.000 33.000 1496.000 34.320 ;
        RECT 4.400 31.600 1496.000 33.000 ;
        RECT 4.000 28.240 1496.000 31.600 ;
        RECT 4.400 26.840 1496.000 28.240 ;
        RECT 4.000 25.520 1496.000 26.840 ;
        RECT 4.000 24.120 1495.600 25.520 ;
        RECT 4.000 22.800 1496.000 24.120 ;
        RECT 4.400 21.400 1496.000 22.800 ;
        RECT 4.000 18.040 1496.000 21.400 ;
        RECT 4.400 16.640 1496.000 18.040 ;
        RECT 4.000 15.320 1496.000 16.640 ;
        RECT 4.000 13.920 1495.600 15.320 ;
        RECT 4.000 12.600 1496.000 13.920 ;
        RECT 4.400 11.200 1496.000 12.600 ;
        RECT 4.000 7.840 1496.000 11.200 ;
        RECT 4.400 6.440 1496.000 7.840 ;
        RECT 4.000 5.800 1496.000 6.440 ;
        RECT 4.000 4.400 1495.600 5.800 ;
        RECT 4.000 3.080 1496.000 4.400 ;
        RECT 4.400 2.215 1496.000 3.080 ;
      LAYER met4 ;
        RECT 138.295 10.640 1481.840 390.825 ;
  END
END multi_project_harness
END LIBRARY

