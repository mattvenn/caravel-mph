VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vga_clock
  CLASS BLOCK ;
  FOREIGN vga_clock ;
  ORIGIN 0.000 0.000 ;
  SIZE 227.025 BY 237.745 ;
  PIN adj_hrs
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END adj_hrs
  PIN adj_min
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 223.025 190.440 227.025 191.040 ;
    END
  END adj_min
  PIN adj_sec
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END adj_sec
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END clk
  PIN hsync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 223.025 104.760 227.025 105.360 ;
    END
  END hsync
  PIN reset_n
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 233.745 79.490 237.745 ;
    END
  END reset_n
  PIN rrggbb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END rrggbb[0]
  PIN rrggbb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END rrggbb[1]
  PIN rrggbb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 223.025 19.080 227.025 19.680 ;
    END
  END rrggbb[2]
  PIN rrggbb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.250 233.745 21.530 237.745 ;
    END
  END rrggbb[3]
  PIN rrggbb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.130 233.745 195.410 237.745 ;
    END
  END rrggbb[4]
  PIN rrggbb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 233.745 137.450 237.745 ;
    END
  END rrggbb[5]
  PIN vsync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END vsync
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 226.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 226.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 221.260 225.845 ;
      LAYER met1 ;
        RECT 2.830 10.640 221.260 226.000 ;
      LAYER met2 ;
        RECT 2.860 233.465 20.970 233.745 ;
        RECT 21.810 233.465 78.930 233.745 ;
        RECT 79.770 233.465 136.890 233.745 ;
        RECT 137.730 233.465 194.850 233.745 ;
        RECT 195.690 233.465 214.720 233.745 ;
        RECT 2.860 4.280 214.720 233.465 ;
        RECT 3.410 4.000 60.530 4.280 ;
        RECT 61.370 4.000 118.490 4.280 ;
        RECT 119.330 4.000 176.450 4.280 ;
        RECT 177.290 4.000 214.720 4.280 ;
      LAYER met3 ;
        RECT 4.000 191.440 223.025 225.925 ;
        RECT 4.000 190.040 222.625 191.440 ;
        RECT 4.000 176.480 223.025 190.040 ;
        RECT 4.400 175.080 223.025 176.480 ;
        RECT 4.000 105.760 223.025 175.080 ;
        RECT 4.000 104.360 222.625 105.760 ;
        RECT 4.000 90.800 223.025 104.360 ;
        RECT 4.400 89.400 223.025 90.800 ;
        RECT 4.000 20.080 223.025 89.400 ;
        RECT 4.000 18.680 222.625 20.080 ;
        RECT 4.000 10.715 223.025 18.680 ;
      LAYER met4 ;
        RECT 174.640 10.640 176.240 226.000 ;
  END
END vga_clock
END LIBRARY

