VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2183.690 89.660 2184.010 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2183.690 89.520 2899.310 89.660 ;
        RECT 2183.690 89.460 2184.010 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2183.720 89.460 2183.980 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2183.710 601.955 2183.990 602.325 ;
        RECT 2183.780 89.750 2183.920 601.955 ;
        RECT 2183.720 89.430 2183.980 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2183.710 602.000 2183.990 602.280 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2166.000 604.800 2170.000 605.400 ;
        RECT 2169.670 602.290 2169.970 604.800 ;
        RECT 2183.685 602.290 2184.015 602.305 ;
        RECT 2169.670 601.990 2184.015 602.290 ;
        RECT 2183.685 601.975 2184.015 601.990 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2191.970 2429.200 2192.290 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 2191.970 2429.060 2901.150 2429.200 ;
        RECT 2191.970 2429.000 2192.290 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 2180.470 707.780 2180.790 707.840 ;
        RECT 2191.970 707.780 2192.290 707.840 ;
        RECT 2180.470 707.640 2192.290 707.780 ;
        RECT 2180.470 707.580 2180.790 707.640 ;
        RECT 2191.970 707.580 2192.290 707.640 ;
      LAYER via ;
        RECT 2192.000 2429.000 2192.260 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 2180.500 707.580 2180.760 707.840 ;
        RECT 2192.000 707.580 2192.260 707.840 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 2192.000 2428.970 2192.260 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 2192.060 707.870 2192.200 2428.970 ;
        RECT 2180.500 707.550 2180.760 707.870 ;
        RECT 2192.000 707.550 2192.260 707.870 ;
        RECT 2180.560 706.365 2180.700 707.550 ;
        RECT 2180.490 705.995 2180.770 706.365 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 2180.490 706.040 2180.770 706.320 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2180.465 706.330 2180.795 706.345 ;
        RECT 2169.670 706.030 2180.795 706.330 ;
        RECT 2169.670 705.360 2169.970 706.030 ;
        RECT 2180.465 706.015 2180.795 706.030 ;
        RECT 2166.000 704.760 2170.000 705.360 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.470 717.640 2180.790 717.700 ;
        RECT 2901.290 717.640 2901.610 717.700 ;
        RECT 2180.470 717.500 2901.610 717.640 ;
        RECT 2180.470 717.440 2180.790 717.500 ;
        RECT 2901.290 717.440 2901.610 717.500 ;
      LAYER via ;
        RECT 2180.500 717.440 2180.760 717.700 ;
        RECT 2901.320 717.440 2901.580 717.700 ;
      LAYER met2 ;
        RECT 2901.310 2669.155 2901.590 2669.525 ;
        RECT 2901.380 717.730 2901.520 2669.155 ;
        RECT 2180.500 717.410 2180.760 717.730 ;
        RECT 2901.320 717.410 2901.580 717.730 ;
        RECT 2180.560 715.885 2180.700 717.410 ;
        RECT 2180.490 715.515 2180.770 715.885 ;
      LAYER via2 ;
        RECT 2901.310 2669.200 2901.590 2669.480 ;
        RECT 2180.490 715.560 2180.770 715.840 ;
      LAYER met3 ;
        RECT 2901.285 2669.490 2901.615 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2901.285 2669.190 2924.800 2669.490 ;
        RECT 2901.285 2669.175 2901.615 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2180.465 715.850 2180.795 715.865 ;
        RECT 2169.670 715.550 2180.795 715.850 ;
        RECT 2169.670 714.880 2169.970 715.550 ;
        RECT 2180.465 715.535 2180.795 715.550 ;
        RECT 2166.000 714.280 2170.000 714.880 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2191.510 2898.400 2191.830 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2191.510 2898.260 2901.150 2898.400 ;
        RECT 2191.510 2898.200 2191.830 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2180.470 729.200 2180.790 729.260 ;
        RECT 2191.510 729.200 2191.830 729.260 ;
        RECT 2180.470 729.060 2191.830 729.200 ;
        RECT 2180.470 729.000 2180.790 729.060 ;
        RECT 2191.510 729.000 2191.830 729.060 ;
      LAYER via ;
        RECT 2191.540 2898.200 2191.800 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2180.500 729.000 2180.760 729.260 ;
        RECT 2191.540 729.000 2191.800 729.260 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2191.540 2898.170 2191.800 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2191.600 729.290 2191.740 2898.170 ;
        RECT 2180.500 728.970 2180.760 729.290 ;
        RECT 2191.540 728.970 2191.800 729.290 ;
        RECT 2180.560 726.765 2180.700 728.970 ;
        RECT 2180.490 726.395 2180.770 726.765 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 2180.490 726.440 2180.770 726.720 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2180.465 726.730 2180.795 726.745 ;
        RECT 2169.670 726.430 2180.795 726.730 ;
        RECT 2169.670 725.080 2169.970 726.430 ;
        RECT 2180.465 726.415 2180.795 726.430 ;
        RECT 2166.000 724.480 2170.000 725.080 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2191.050 3133.000 2191.370 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2191.050 3132.860 2901.150 3133.000 ;
        RECT 2191.050 3132.800 2191.370 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 2180.470 737.700 2180.790 737.760 ;
        RECT 2191.050 737.700 2191.370 737.760 ;
        RECT 2180.470 737.560 2191.370 737.700 ;
        RECT 2180.470 737.500 2180.790 737.560 ;
        RECT 2191.050 737.500 2191.370 737.560 ;
      LAYER via ;
        RECT 2191.080 3132.800 2191.340 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 2180.500 737.500 2180.760 737.760 ;
        RECT 2191.080 737.500 2191.340 737.760 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2191.080 3132.770 2191.340 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 2191.140 737.790 2191.280 3132.770 ;
        RECT 2180.500 737.470 2180.760 737.790 ;
        RECT 2191.080 737.470 2191.340 737.790 ;
        RECT 2180.560 736.285 2180.700 737.470 ;
        RECT 2180.490 735.915 2180.770 736.285 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 2180.490 735.960 2180.770 736.240 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2180.465 736.250 2180.795 736.265 ;
        RECT 2169.670 735.950 2180.795 736.250 ;
        RECT 2169.670 735.280 2169.970 735.950 ;
        RECT 2180.465 735.935 2180.795 735.950 ;
        RECT 2166.000 734.680 2170.000 735.280 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2197.490 3367.600 2197.810 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2197.490 3367.460 2901.150 3367.600 ;
        RECT 2197.490 3367.400 2197.810 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 2180.470 745.180 2180.790 745.240 ;
        RECT 2197.490 745.180 2197.810 745.240 ;
        RECT 2180.470 745.040 2197.810 745.180 ;
        RECT 2180.470 744.980 2180.790 745.040 ;
        RECT 2197.490 744.980 2197.810 745.040 ;
      LAYER via ;
        RECT 2197.520 3367.400 2197.780 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 2180.500 744.980 2180.760 745.240 ;
        RECT 2197.520 744.980 2197.780 745.240 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2197.520 3367.370 2197.780 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 2197.580 745.270 2197.720 3367.370 ;
        RECT 2180.500 745.125 2180.760 745.270 ;
        RECT 2180.490 744.755 2180.770 745.125 ;
        RECT 2197.520 744.950 2197.780 745.270 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 2180.490 744.800 2180.770 745.080 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2180.465 745.090 2180.795 745.105 ;
        RECT 2169.670 744.800 2180.795 745.090 ;
        RECT 2166.000 744.790 2180.795 744.800 ;
        RECT 2166.000 744.200 2170.000 744.790 ;
        RECT 2180.465 744.775 2180.795 744.790 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2204.390 3502.240 2204.710 3502.300 ;
        RECT 2798.250 3502.240 2798.570 3502.300 ;
        RECT 2204.390 3502.100 2798.570 3502.240 ;
        RECT 2204.390 3502.040 2204.710 3502.100 ;
        RECT 2798.250 3502.040 2798.570 3502.100 ;
        RECT 2180.470 757.080 2180.790 757.140 ;
        RECT 2204.390 757.080 2204.710 757.140 ;
        RECT 2180.470 756.940 2204.710 757.080 ;
        RECT 2180.470 756.880 2180.790 756.940 ;
        RECT 2204.390 756.880 2204.710 756.940 ;
      LAYER via ;
        RECT 2204.420 3502.040 2204.680 3502.300 ;
        RECT 2798.280 3502.040 2798.540 3502.300 ;
        RECT 2180.500 756.880 2180.760 757.140 ;
        RECT 2204.420 756.880 2204.680 757.140 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3502.330 2798.480 3517.600 ;
        RECT 2204.420 3502.010 2204.680 3502.330 ;
        RECT 2798.280 3502.010 2798.540 3502.330 ;
        RECT 2204.480 757.170 2204.620 3502.010 ;
        RECT 2180.500 756.850 2180.760 757.170 ;
        RECT 2204.420 756.850 2204.680 757.170 ;
        RECT 2180.560 756.005 2180.700 756.850 ;
        RECT 2180.490 755.635 2180.770 756.005 ;
      LAYER via2 ;
        RECT 2180.490 755.680 2180.770 755.960 ;
      LAYER met3 ;
        RECT 2180.465 755.970 2180.795 755.985 ;
        RECT 2169.670 755.670 2180.795 755.970 ;
        RECT 2169.670 755.000 2169.970 755.670 ;
        RECT 2180.465 755.655 2180.795 755.670 ;
        RECT 2166.000 754.400 2170.000 755.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2190.590 3502.920 2190.910 3502.980 ;
        RECT 2473.950 3502.920 2474.270 3502.980 ;
        RECT 2190.590 3502.780 2474.270 3502.920 ;
        RECT 2190.590 3502.720 2190.910 3502.780 ;
        RECT 2473.950 3502.720 2474.270 3502.780 ;
        RECT 2180.470 765.580 2180.790 765.640 ;
        RECT 2190.590 765.580 2190.910 765.640 ;
        RECT 2180.470 765.440 2190.910 765.580 ;
        RECT 2180.470 765.380 2180.790 765.440 ;
        RECT 2190.590 765.380 2190.910 765.440 ;
      LAYER via ;
        RECT 2190.620 3502.720 2190.880 3502.980 ;
        RECT 2473.980 3502.720 2474.240 3502.980 ;
        RECT 2180.500 765.380 2180.760 765.640 ;
        RECT 2190.620 765.380 2190.880 765.640 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3503.010 2474.180 3517.600 ;
        RECT 2190.620 3502.690 2190.880 3503.010 ;
        RECT 2473.980 3502.690 2474.240 3503.010 ;
        RECT 2190.680 765.670 2190.820 3502.690 ;
        RECT 2180.500 765.525 2180.760 765.670 ;
        RECT 2180.490 765.155 2180.770 765.525 ;
        RECT 2190.620 765.350 2190.880 765.670 ;
      LAYER via2 ;
        RECT 2180.490 765.200 2180.770 765.480 ;
      LAYER met3 ;
        RECT 2180.465 765.490 2180.795 765.505 ;
        RECT 2169.670 765.200 2180.795 765.490 ;
        RECT 2166.000 765.190 2180.795 765.200 ;
        RECT 2166.000 764.600 2170.000 765.190 ;
        RECT 2180.465 765.175 2180.795 765.190 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2149.190 3498.500 2149.510 3498.560 ;
        RECT 2164.830 3498.500 2165.150 3498.560 ;
        RECT 2149.190 3498.360 2165.150 3498.500 ;
        RECT 2149.190 3498.300 2149.510 3498.360 ;
        RECT 2164.830 3498.300 2165.150 3498.360 ;
      LAYER via ;
        RECT 2149.220 3498.300 2149.480 3498.560 ;
        RECT 2164.860 3498.300 2165.120 3498.560 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3498.590 2149.420 3517.600 ;
        RECT 2149.220 3498.270 2149.480 3498.590 ;
        RECT 2164.860 3498.270 2165.120 3498.590 ;
        RECT 2164.920 776.970 2165.060 3498.270 ;
        RECT 2166.690 776.970 2166.970 777.085 ;
        RECT 2164.920 776.830 2166.970 776.970 ;
        RECT 2166.690 776.715 2166.970 776.830 ;
      LAYER via2 ;
        RECT 2166.690 776.760 2166.970 777.040 ;
      LAYER met3 ;
        RECT 2166.665 777.050 2166.995 777.065 ;
        RECT 2166.665 776.735 2167.210 777.050 ;
        RECT 2166.910 774.720 2167.210 776.735 ;
        RECT 2166.000 774.120 2170.000 774.720 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3504.620 1825.210 3504.680 ;
        RECT 2170.810 3504.620 2171.130 3504.680 ;
        RECT 1824.890 3504.480 2171.130 3504.620 ;
        RECT 1824.890 3504.420 1825.210 3504.480 ;
        RECT 2170.810 3504.420 2171.130 3504.480 ;
      LAYER via ;
        RECT 1824.920 3504.420 1825.180 3504.680 ;
        RECT 2170.840 3504.420 2171.100 3504.680 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3504.710 1825.120 3517.600 ;
        RECT 1824.920 3504.390 1825.180 3504.710 ;
        RECT 2170.840 3504.390 2171.100 3504.710 ;
        RECT 2170.900 785.925 2171.040 3504.390 ;
        RECT 2170.830 785.555 2171.110 785.925 ;
      LAYER via2 ;
        RECT 2170.830 785.600 2171.110 785.880 ;
      LAYER met3 ;
        RECT 2170.805 785.890 2171.135 785.905 ;
        RECT 2169.670 785.590 2171.135 785.890 ;
        RECT 2169.670 784.920 2169.970 785.590 ;
        RECT 2170.805 785.575 2171.135 785.590 ;
        RECT 2166.000 784.320 2170.000 784.920 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3500.880 1500.910 3500.940 ;
        RECT 2167.130 3500.880 2167.450 3500.940 ;
        RECT 1500.590 3500.740 2167.450 3500.880 ;
        RECT 1500.590 3500.680 1500.910 3500.740 ;
        RECT 2167.130 3500.680 2167.450 3500.740 ;
      LAYER via ;
        RECT 1500.620 3500.680 1500.880 3500.940 ;
        RECT 2167.160 3500.680 2167.420 3500.940 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3500.970 1500.820 3517.600 ;
        RECT 1500.620 3500.650 1500.880 3500.970 ;
        RECT 2167.160 3500.650 2167.420 3500.970 ;
        RECT 2167.220 797.485 2167.360 3500.650 ;
        RECT 2167.150 797.115 2167.430 797.485 ;
      LAYER via2 ;
        RECT 2167.150 797.160 2167.430 797.440 ;
      LAYER met3 ;
        RECT 2167.125 797.450 2167.455 797.465 ;
        RECT 2166.910 797.135 2167.455 797.450 ;
        RECT 2166.910 795.120 2167.210 797.135 ;
        RECT 2166.000 794.520 2170.000 795.120 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2184.150 324.260 2184.470 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2184.150 324.120 2899.310 324.260 ;
        RECT 2184.150 324.060 2184.470 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2184.180 324.060 2184.440 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2184.170 614.875 2184.450 615.245 ;
        RECT 2184.240 324.350 2184.380 614.875 ;
        RECT 2184.180 324.030 2184.440 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2184.170 614.920 2184.450 615.200 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2184.145 615.210 2184.475 615.225 ;
        RECT 2169.670 614.920 2184.475 615.210 ;
        RECT 2166.000 614.910 2184.475 614.920 ;
        RECT 2166.000 614.320 2170.000 614.910 ;
        RECT 2184.145 614.895 2184.475 614.910 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3504.960 1176.150 3505.020 ;
        RECT 2167.590 3504.960 2167.910 3505.020 ;
        RECT 1175.830 3504.820 2167.910 3504.960 ;
        RECT 1175.830 3504.760 1176.150 3504.820 ;
        RECT 2167.590 3504.760 2167.910 3504.820 ;
      LAYER via ;
        RECT 1175.860 3504.760 1176.120 3505.020 ;
        RECT 2167.620 3504.760 2167.880 3505.020 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3505.050 1176.060 3517.600 ;
        RECT 1175.860 3504.730 1176.120 3505.050 ;
        RECT 2167.620 3504.730 2167.880 3505.050 ;
        RECT 2167.680 807.005 2167.820 3504.730 ;
        RECT 2167.610 806.635 2167.890 807.005 ;
      LAYER via2 ;
        RECT 2167.610 806.680 2167.890 806.960 ;
      LAYER met3 ;
        RECT 2167.585 806.970 2167.915 806.985 ;
        RECT 2167.585 806.655 2168.130 806.970 ;
        RECT 2167.830 805.320 2168.130 806.655 ;
        RECT 2166.000 804.720 2170.000 805.320 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3504.280 851.850 3504.340 ;
        RECT 2165.290 3504.280 2165.610 3504.340 ;
        RECT 851.530 3504.140 2165.610 3504.280 ;
        RECT 851.530 3504.080 851.850 3504.140 ;
        RECT 2165.290 3504.080 2165.610 3504.140 ;
        RECT 2165.290 883.220 2165.610 883.280 ;
        RECT 2168.510 883.220 2168.830 883.280 ;
        RECT 2165.290 883.080 2168.830 883.220 ;
        RECT 2165.290 883.020 2165.610 883.080 ;
        RECT 2168.510 883.020 2168.830 883.080 ;
        RECT 2166.210 846.500 2166.530 846.560 ;
        RECT 2168.510 846.500 2168.830 846.560 ;
        RECT 2166.210 846.360 2168.830 846.500 ;
        RECT 2166.210 846.300 2166.530 846.360 ;
        RECT 2168.510 846.300 2168.830 846.360 ;
      LAYER via ;
        RECT 851.560 3504.080 851.820 3504.340 ;
        RECT 2165.320 3504.080 2165.580 3504.340 ;
        RECT 2165.320 883.020 2165.580 883.280 ;
        RECT 2168.540 883.020 2168.800 883.280 ;
        RECT 2166.240 846.300 2166.500 846.560 ;
        RECT 2168.540 846.300 2168.800 846.560 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3504.370 851.760 3517.600 ;
        RECT 851.560 3504.050 851.820 3504.370 ;
        RECT 2165.320 3504.050 2165.580 3504.370 ;
        RECT 2165.380 883.310 2165.520 3504.050 ;
        RECT 2165.320 882.990 2165.580 883.310 ;
        RECT 2168.540 882.990 2168.800 883.310 ;
        RECT 2168.600 846.590 2168.740 882.990 ;
        RECT 2166.240 846.270 2166.500 846.590 ;
        RECT 2168.540 846.270 2168.800 846.590 ;
        RECT 2166.300 817.090 2166.440 846.270 ;
        RECT 2166.690 817.090 2166.970 817.205 ;
        RECT 2166.300 816.950 2166.970 817.090 ;
        RECT 2166.690 816.835 2166.970 816.950 ;
      LAYER via2 ;
        RECT 2166.690 816.880 2166.970 817.160 ;
      LAYER met3 ;
        RECT 2166.665 817.170 2166.995 817.185 ;
        RECT 2166.665 816.855 2167.210 817.170 ;
        RECT 2166.910 814.840 2167.210 816.855 ;
        RECT 2166.000 814.240 2170.000 814.840 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3502.920 527.550 3502.980 ;
        RECT 2168.050 3502.920 2168.370 3502.980 ;
        RECT 527.230 3502.780 2168.370 3502.920 ;
        RECT 527.230 3502.720 527.550 3502.780 ;
        RECT 2168.050 3502.720 2168.370 3502.780 ;
      LAYER via ;
        RECT 527.260 3502.720 527.520 3502.980 ;
        RECT 2168.080 3502.720 2168.340 3502.980 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.010 527.460 3517.600 ;
        RECT 527.260 3502.690 527.520 3503.010 ;
        RECT 2168.080 3502.690 2168.340 3503.010 ;
        RECT 2168.140 827.405 2168.280 3502.690 ;
        RECT 2168.070 827.035 2168.350 827.405 ;
      LAYER via2 ;
        RECT 2168.070 827.080 2168.350 827.360 ;
      LAYER met3 ;
        RECT 2168.045 827.370 2168.375 827.385 ;
        RECT 2167.830 827.055 2168.375 827.370 ;
        RECT 2167.830 825.040 2168.130 827.055 ;
        RECT 2166.000 824.440 2170.000 825.040 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.240 202.790 3502.300 ;
        RECT 2165.750 3502.240 2166.070 3502.300 ;
        RECT 202.470 3502.100 2166.070 3502.240 ;
        RECT 202.470 3502.040 202.790 3502.100 ;
        RECT 2165.750 3502.040 2166.070 3502.100 ;
        RECT 2165.290 834.260 2165.610 834.320 ;
        RECT 2166.670 834.260 2166.990 834.320 ;
        RECT 2165.290 834.120 2166.990 834.260 ;
        RECT 2165.290 834.060 2165.610 834.120 ;
        RECT 2166.670 834.060 2166.990 834.120 ;
      LAYER via ;
        RECT 202.500 3502.040 202.760 3502.300 ;
        RECT 2165.780 3502.040 2166.040 3502.300 ;
        RECT 2165.320 834.060 2165.580 834.320 ;
        RECT 2166.700 834.060 2166.960 834.320 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.330 202.700 3517.600 ;
        RECT 202.500 3502.010 202.760 3502.330 ;
        RECT 2165.780 3502.010 2166.040 3502.330 ;
        RECT 2165.840 845.650 2165.980 3502.010 ;
        RECT 2165.380 845.510 2165.980 845.650 ;
        RECT 2165.380 834.350 2165.520 845.510 ;
        RECT 2165.320 834.030 2165.580 834.350 ;
        RECT 2166.700 834.205 2166.960 834.350 ;
        RECT 2166.690 833.835 2166.970 834.205 ;
      LAYER via2 ;
        RECT 2166.690 833.880 2166.970 834.160 ;
      LAYER met3 ;
        RECT 2166.000 834.640 2170.000 835.240 ;
        RECT 2166.910 834.185 2167.210 834.640 ;
        RECT 2166.665 833.870 2167.210 834.185 ;
        RECT 2166.665 833.855 2166.995 833.870 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.930 3408.740 19.250 3408.800 ;
        RECT 2166.210 3408.740 2166.530 3408.800 ;
        RECT 18.930 3408.600 2166.530 3408.740 ;
        RECT 18.930 3408.540 19.250 3408.600 ;
        RECT 2166.210 3408.540 2166.530 3408.600 ;
        RECT 2166.210 1001.200 2166.530 1001.260 ;
        RECT 2171.730 1001.200 2172.050 1001.260 ;
        RECT 2166.210 1001.060 2172.050 1001.200 ;
        RECT 2166.210 1001.000 2166.530 1001.060 ;
        RECT 2171.730 1001.000 2172.050 1001.060 ;
        RECT 2166.210 990.320 2166.530 990.380 ;
        RECT 2171.730 990.320 2172.050 990.380 ;
        RECT 2166.210 990.180 2172.050 990.320 ;
        RECT 2166.210 990.120 2166.530 990.180 ;
        RECT 2171.730 990.120 2172.050 990.180 ;
      LAYER via ;
        RECT 18.960 3408.540 19.220 3408.800 ;
        RECT 2166.240 3408.540 2166.500 3408.800 ;
        RECT 2166.240 1001.000 2166.500 1001.260 ;
        RECT 2171.760 1001.000 2172.020 1001.260 ;
        RECT 2166.240 990.120 2166.500 990.380 ;
        RECT 2171.760 990.120 2172.020 990.380 ;
      LAYER met2 ;
        RECT 18.950 3411.035 19.230 3411.405 ;
        RECT 19.020 3408.830 19.160 3411.035 ;
        RECT 18.960 3408.510 19.220 3408.830 ;
        RECT 2166.240 3408.510 2166.500 3408.830 ;
        RECT 2166.300 1001.290 2166.440 3408.510 ;
        RECT 2166.240 1000.970 2166.500 1001.290 ;
        RECT 2171.760 1000.970 2172.020 1001.290 ;
        RECT 2171.820 990.410 2171.960 1000.970 ;
        RECT 2166.240 990.090 2166.500 990.410 ;
        RECT 2171.760 990.090 2172.020 990.410 ;
        RECT 2166.300 847.010 2166.440 990.090 ;
        RECT 2166.690 847.010 2166.970 847.125 ;
        RECT 2166.300 846.870 2166.970 847.010 ;
        RECT 2166.690 846.755 2166.970 846.870 ;
      LAYER via2 ;
        RECT 18.950 3411.080 19.230 3411.360 ;
        RECT 2166.690 846.800 2166.970 847.080 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 18.925 3411.370 19.255 3411.385 ;
        RECT -4.800 3411.070 19.255 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 18.925 3411.055 19.255 3411.070 ;
        RECT 2166.665 847.090 2166.995 847.105 ;
        RECT 2166.665 846.775 2167.210 847.090 ;
        RECT 2166.910 844.760 2167.210 846.775 ;
        RECT 2166.000 844.160 2170.000 844.760 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 3119.060 16.490 3119.120 ;
        RECT 2162.990 3119.060 2163.310 3119.120 ;
        RECT 16.170 3118.920 2163.310 3119.060 ;
        RECT 16.170 3118.860 16.490 3118.920 ;
        RECT 2162.990 3118.860 2163.310 3118.920 ;
        RECT 2162.990 1001.540 2163.310 1001.600 ;
        RECT 2172.190 1001.540 2172.510 1001.600 ;
        RECT 2162.990 1001.400 2172.510 1001.540 ;
        RECT 2162.990 1001.340 2163.310 1001.400 ;
        RECT 2172.190 1001.340 2172.510 1001.400 ;
        RECT 2166.670 989.980 2166.990 990.040 ;
        RECT 2172.190 989.980 2172.510 990.040 ;
        RECT 2166.670 989.840 2172.510 989.980 ;
        RECT 2166.670 989.780 2166.990 989.840 ;
        RECT 2172.190 989.780 2172.510 989.840 ;
        RECT 2165.290 882.540 2165.610 882.600 ;
        RECT 2166.670 882.540 2166.990 882.600 ;
        RECT 2165.290 882.400 2166.990 882.540 ;
        RECT 2165.290 882.340 2165.610 882.400 ;
        RECT 2166.670 882.340 2166.990 882.400 ;
        RECT 2165.290 853.980 2165.610 854.040 ;
        RECT 2166.670 853.980 2166.990 854.040 ;
        RECT 2165.290 853.840 2166.990 853.980 ;
        RECT 2165.290 853.780 2165.610 853.840 ;
        RECT 2166.670 853.780 2166.990 853.840 ;
      LAYER via ;
        RECT 16.200 3118.860 16.460 3119.120 ;
        RECT 2163.020 3118.860 2163.280 3119.120 ;
        RECT 2163.020 1001.340 2163.280 1001.600 ;
        RECT 2172.220 1001.340 2172.480 1001.600 ;
        RECT 2166.700 989.780 2166.960 990.040 ;
        RECT 2172.220 989.780 2172.480 990.040 ;
        RECT 2165.320 882.340 2165.580 882.600 ;
        RECT 2166.700 882.340 2166.960 882.600 ;
        RECT 2165.320 853.780 2165.580 854.040 ;
        RECT 2166.700 853.780 2166.960 854.040 ;
      LAYER met2 ;
        RECT 16.190 3124.075 16.470 3124.445 ;
        RECT 16.260 3119.150 16.400 3124.075 ;
        RECT 16.200 3118.830 16.460 3119.150 ;
        RECT 2163.020 3118.830 2163.280 3119.150 ;
        RECT 2163.080 1001.630 2163.220 3118.830 ;
        RECT 2163.020 1001.310 2163.280 1001.630 ;
        RECT 2172.220 1001.310 2172.480 1001.630 ;
        RECT 2172.280 990.070 2172.420 1001.310 ;
        RECT 2166.700 989.750 2166.960 990.070 ;
        RECT 2172.220 989.750 2172.480 990.070 ;
        RECT 2166.760 882.630 2166.900 989.750 ;
        RECT 2165.320 882.310 2165.580 882.630 ;
        RECT 2166.700 882.310 2166.960 882.630 ;
        RECT 2165.380 854.070 2165.520 882.310 ;
        RECT 2165.320 853.750 2165.580 854.070 ;
        RECT 2166.700 853.925 2166.960 854.070 ;
        RECT 2166.690 853.555 2166.970 853.925 ;
      LAYER via2 ;
        RECT 16.190 3124.120 16.470 3124.400 ;
        RECT 2166.690 853.600 2166.970 853.880 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 16.165 3124.410 16.495 3124.425 ;
        RECT -4.800 3124.110 16.495 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 16.165 3124.095 16.495 3124.110 ;
        RECT 2166.000 854.360 2170.000 854.960 ;
        RECT 2166.910 853.905 2167.210 854.360 ;
        RECT 2166.665 853.590 2167.210 853.905 ;
        RECT 2166.665 853.575 2166.995 853.590 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2836.180 20.630 2836.240 ;
        RECT 831.750 2836.180 832.070 2836.240 ;
        RECT 20.310 2836.040 832.070 2836.180 ;
        RECT 20.310 2835.980 20.630 2836.040 ;
        RECT 831.750 2835.980 832.070 2836.040 ;
        RECT 831.750 1003.580 832.070 1003.640 ;
        RECT 860.730 1003.580 861.050 1003.640 ;
        RECT 831.750 1003.440 861.050 1003.580 ;
        RECT 831.750 1003.380 832.070 1003.440 ;
        RECT 860.730 1003.380 861.050 1003.440 ;
        RECT 1762.330 1000.860 1762.650 1000.920 ;
        RECT 1766.010 1000.860 1766.330 1000.920 ;
        RECT 1762.330 1000.720 1766.330 1000.860 ;
        RECT 1762.330 1000.660 1762.650 1000.720 ;
        RECT 1766.010 1000.660 1766.330 1000.720 ;
        RECT 1766.470 1000.860 1766.790 1000.920 ;
        RECT 1788.550 1000.860 1788.870 1000.920 ;
        RECT 1766.470 1000.720 1788.870 1000.860 ;
        RECT 1766.470 1000.660 1766.790 1000.720 ;
        RECT 1788.550 1000.660 1788.870 1000.720 ;
        RECT 1220.450 1000.520 1220.770 1000.580 ;
        RECT 1232.870 1000.520 1233.190 1000.580 ;
        RECT 1220.450 1000.380 1233.190 1000.520 ;
        RECT 1220.450 1000.320 1220.770 1000.380 ;
        RECT 1232.870 1000.320 1233.190 1000.380 ;
        RECT 1398.470 1000.520 1398.790 1000.580 ;
        RECT 1421.470 1000.520 1421.790 1000.580 ;
        RECT 1398.470 1000.380 1421.790 1000.520 ;
        RECT 1398.470 1000.320 1398.790 1000.380 ;
        RECT 1421.470 1000.320 1421.790 1000.380 ;
        RECT 1563.150 1000.520 1563.470 1000.580 ;
        RECT 1577.870 1000.520 1578.190 1000.580 ;
        RECT 1563.150 1000.380 1578.190 1000.520 ;
        RECT 1563.150 1000.320 1563.470 1000.380 ;
        RECT 1577.870 1000.320 1578.190 1000.380 ;
        RECT 1885.150 1000.520 1885.470 1000.580 ;
        RECT 1885.150 1000.380 1932.300 1000.520 ;
        RECT 1885.150 1000.320 1885.470 1000.380 ;
        RECT 1276.570 1000.180 1276.890 1000.240 ;
        RECT 1435.270 1000.180 1435.590 1000.240 ;
        RECT 1666.650 1000.180 1666.970 1000.240 ;
        RECT 935.340 1000.040 959.400 1000.180 ;
        RECT 860.730 999.500 861.050 999.560 ;
        RECT 935.340 999.500 935.480 1000.040 ;
        RECT 860.730 999.360 935.480 999.500 ;
        RECT 959.260 999.500 959.400 1000.040 ;
        RECT 1276.570 1000.040 1290.140 1000.180 ;
        RECT 1276.570 999.980 1276.890 1000.040 ;
        RECT 1159.270 999.640 1159.590 999.900 ;
        RECT 1007.470 999.500 1007.790 999.560 ;
        RECT 959.260 999.360 1007.790 999.500 ;
        RECT 860.730 999.300 861.050 999.360 ;
        RECT 1007.470 999.300 1007.790 999.360 ;
        RECT 1008.390 999.500 1008.710 999.560 ;
        RECT 1070.490 999.500 1070.810 999.560 ;
        RECT 1008.390 999.360 1070.810 999.500 ;
        RECT 1008.390 999.300 1008.710 999.360 ;
        RECT 1070.490 999.300 1070.810 999.360 ;
        RECT 1096.710 999.500 1097.030 999.560 ;
        RECT 1159.360 999.500 1159.500 999.640 ;
        RECT 1096.710 999.360 1159.500 999.500 ;
        RECT 1174.910 999.500 1175.230 999.560 ;
        RECT 1220.450 999.500 1220.770 999.560 ;
        RECT 1174.910 999.360 1220.770 999.500 ;
        RECT 1096.710 999.300 1097.030 999.360 ;
        RECT 1174.910 999.300 1175.230 999.360 ;
        RECT 1220.450 999.300 1220.770 999.360 ;
        RECT 1232.870 999.500 1233.190 999.560 ;
        RECT 1242.070 999.500 1242.390 999.560 ;
        RECT 1232.870 999.360 1242.390 999.500 ;
        RECT 1290.000 999.500 1290.140 1000.040 ;
        RECT 1362.220 1000.040 1375.700 1000.180 ;
        RECT 1362.220 999.500 1362.360 1000.040 ;
        RECT 1290.000 999.360 1362.360 999.500 ;
        RECT 1375.560 999.500 1375.700 1000.040 ;
        RECT 1435.270 1000.040 1435.960 1000.180 ;
        RECT 1435.270 999.980 1435.590 1000.040 ;
        RECT 1435.820 999.840 1435.960 1000.040 ;
        RECT 1642.360 1000.040 1666.970 1000.180 ;
        RECT 1435.820 999.700 1463.560 999.840 ;
        RECT 1398.470 999.500 1398.790 999.560 ;
        RECT 1375.560 999.360 1398.790 999.500 ;
        RECT 1232.870 999.300 1233.190 999.360 ;
        RECT 1242.070 999.300 1242.390 999.360 ;
        RECT 1398.470 999.300 1398.790 999.360 ;
        RECT 1421.470 999.500 1421.790 999.560 ;
        RECT 1435.270 999.500 1435.590 999.560 ;
        RECT 1421.470 999.360 1435.590 999.500 ;
        RECT 1463.420 999.500 1463.560 999.700 ;
        RECT 1563.150 999.500 1563.470 999.560 ;
        RECT 1463.420 999.360 1563.470 999.500 ;
        RECT 1421.470 999.300 1421.790 999.360 ;
        RECT 1435.270 999.300 1435.590 999.360 ;
        RECT 1563.150 999.300 1563.470 999.360 ;
        RECT 1577.870 999.500 1578.190 999.560 ;
        RECT 1642.360 999.500 1642.500 1000.040 ;
        RECT 1666.650 999.980 1666.970 1000.040 ;
        RECT 1766.470 999.980 1766.790 1000.240 ;
        RECT 1814.400 1000.040 1815.460 1000.180 ;
        RECT 1766.010 999.840 1766.330 999.900 ;
        RECT 1766.560 999.840 1766.700 999.980 ;
        RECT 1766.010 999.700 1766.700 999.840 ;
        RECT 1788.550 999.840 1788.870 999.900 ;
        RECT 1814.400 999.840 1814.540 1000.040 ;
        RECT 1788.550 999.700 1814.540 999.840 ;
        RECT 1815.320 999.840 1815.460 1000.040 ;
        RECT 1932.160 999.840 1932.300 1000.380 ;
        RECT 1950.930 1000.180 1951.250 1000.240 ;
        RECT 1933.540 1000.040 1951.250 1000.180 ;
        RECT 1933.540 999.840 1933.680 1000.040 ;
        RECT 1950.930 999.980 1951.250 1000.040 ;
        RECT 2149.650 1000.180 2149.970 1000.240 ;
        RECT 2149.650 1000.040 2167.820 1000.180 ;
        RECT 2149.650 999.980 2149.970 1000.040 ;
        RECT 1815.320 999.700 1815.920 999.840 ;
        RECT 1932.160 999.700 1933.680 999.840 ;
        RECT 1766.010 999.640 1766.330 999.700 ;
        RECT 1788.550 999.640 1788.870 999.700 ;
        RECT 1577.870 999.360 1642.500 999.500 ;
        RECT 1666.650 999.500 1666.970 999.560 ;
        RECT 1762.330 999.500 1762.650 999.560 ;
        RECT 1666.650 999.360 1762.650 999.500 ;
        RECT 1815.780 999.500 1815.920 999.700 ;
        RECT 1950.930 999.500 1951.250 999.560 ;
        RECT 2149.650 999.500 2149.970 999.560 ;
        RECT 1815.780 999.360 1884.460 999.500 ;
        RECT 1577.870 999.300 1578.190 999.360 ;
        RECT 1666.650 999.300 1666.970 999.360 ;
        RECT 1762.330 999.300 1762.650 999.360 ;
        RECT 1884.320 999.160 1884.460 999.360 ;
        RECT 1950.930 999.360 2149.970 999.500 ;
        RECT 1950.930 999.300 1951.250 999.360 ;
        RECT 2149.650 999.300 2149.970 999.360 ;
        RECT 1885.150 999.160 1885.470 999.220 ;
        RECT 1884.320 999.020 1885.470 999.160 ;
        RECT 1885.150 998.960 1885.470 999.020 ;
        RECT 2167.680 998.480 2167.820 1000.040 ;
        RECT 2181.390 998.480 2181.710 998.540 ;
        RECT 2167.680 998.340 2181.710 998.480 ;
        RECT 2181.390 998.280 2181.710 998.340 ;
      LAYER via ;
        RECT 20.340 2835.980 20.600 2836.240 ;
        RECT 831.780 2835.980 832.040 2836.240 ;
        RECT 831.780 1003.380 832.040 1003.640 ;
        RECT 860.760 1003.380 861.020 1003.640 ;
        RECT 1762.360 1000.660 1762.620 1000.920 ;
        RECT 1766.040 1000.660 1766.300 1000.920 ;
        RECT 1766.500 1000.660 1766.760 1000.920 ;
        RECT 1788.580 1000.660 1788.840 1000.920 ;
        RECT 1220.480 1000.320 1220.740 1000.580 ;
        RECT 1232.900 1000.320 1233.160 1000.580 ;
        RECT 1398.500 1000.320 1398.760 1000.580 ;
        RECT 1421.500 1000.320 1421.760 1000.580 ;
        RECT 1563.180 1000.320 1563.440 1000.580 ;
        RECT 1577.900 1000.320 1578.160 1000.580 ;
        RECT 1885.180 1000.320 1885.440 1000.580 ;
        RECT 860.760 999.300 861.020 999.560 ;
        RECT 1276.600 999.980 1276.860 1000.240 ;
        RECT 1159.300 999.640 1159.560 999.900 ;
        RECT 1007.500 999.300 1007.760 999.560 ;
        RECT 1008.420 999.300 1008.680 999.560 ;
        RECT 1070.520 999.300 1070.780 999.560 ;
        RECT 1096.740 999.300 1097.000 999.560 ;
        RECT 1174.940 999.300 1175.200 999.560 ;
        RECT 1220.480 999.300 1220.740 999.560 ;
        RECT 1232.900 999.300 1233.160 999.560 ;
        RECT 1242.100 999.300 1242.360 999.560 ;
        RECT 1435.300 999.980 1435.560 1000.240 ;
        RECT 1398.500 999.300 1398.760 999.560 ;
        RECT 1421.500 999.300 1421.760 999.560 ;
        RECT 1435.300 999.300 1435.560 999.560 ;
        RECT 1563.180 999.300 1563.440 999.560 ;
        RECT 1577.900 999.300 1578.160 999.560 ;
        RECT 1666.680 999.980 1666.940 1000.240 ;
        RECT 1766.500 999.980 1766.760 1000.240 ;
        RECT 1766.040 999.640 1766.300 999.900 ;
        RECT 1788.580 999.640 1788.840 999.900 ;
        RECT 1950.960 999.980 1951.220 1000.240 ;
        RECT 2149.680 999.980 2149.940 1000.240 ;
        RECT 1666.680 999.300 1666.940 999.560 ;
        RECT 1762.360 999.300 1762.620 999.560 ;
        RECT 1950.960 999.300 1951.220 999.560 ;
        RECT 2149.680 999.300 2149.940 999.560 ;
        RECT 1885.180 998.960 1885.440 999.220 ;
        RECT 2181.420 998.280 2181.680 998.540 ;
      LAYER met2 ;
        RECT 20.330 2836.435 20.610 2836.805 ;
        RECT 20.400 2836.270 20.540 2836.435 ;
        RECT 20.340 2835.950 20.600 2836.270 ;
        RECT 831.780 2835.950 832.040 2836.270 ;
        RECT 831.840 1003.670 831.980 2835.950 ;
        RECT 831.780 1003.350 832.040 1003.670 ;
        RECT 860.760 1003.350 861.020 1003.670 ;
        RECT 860.820 999.590 860.960 1003.350 ;
        RECT 1762.360 1000.630 1762.620 1000.950 ;
        RECT 1766.040 1000.630 1766.300 1000.950 ;
        RECT 1766.500 1000.630 1766.760 1000.950 ;
        RECT 1788.580 1000.630 1788.840 1000.950 ;
        RECT 1220.480 1000.290 1220.740 1000.610 ;
        RECT 1232.900 1000.290 1233.160 1000.610 ;
        RECT 1398.500 1000.290 1398.760 1000.610 ;
        RECT 1421.500 1000.290 1421.760 1000.610 ;
        RECT 1563.180 1000.290 1563.440 1000.610 ;
        RECT 1577.900 1000.290 1578.160 1000.610 ;
        RECT 1070.510 999.755 1070.790 1000.125 ;
        RECT 1096.730 999.755 1097.010 1000.125 ;
        RECT 1159.290 999.755 1159.570 1000.125 ;
        RECT 1174.930 999.755 1175.210 1000.125 ;
        RECT 1070.580 999.590 1070.720 999.755 ;
        RECT 1096.800 999.590 1096.940 999.755 ;
        RECT 1159.300 999.610 1159.560 999.755 ;
        RECT 1175.000 999.590 1175.140 999.755 ;
        RECT 1220.540 999.590 1220.680 1000.290 ;
        RECT 1232.960 999.590 1233.100 1000.290 ;
        RECT 1276.600 1000.125 1276.860 1000.270 ;
        RECT 1276.590 999.755 1276.870 1000.125 ;
        RECT 1398.560 999.590 1398.700 1000.290 ;
        RECT 1421.560 999.590 1421.700 1000.290 ;
        RECT 1435.300 999.950 1435.560 1000.270 ;
        RECT 1435.360 999.590 1435.500 999.950 ;
        RECT 1563.240 999.590 1563.380 1000.290 ;
        RECT 1577.960 999.590 1578.100 1000.290 ;
        RECT 1666.680 999.950 1666.940 1000.270 ;
        RECT 1666.740 999.590 1666.880 999.950 ;
        RECT 1762.420 999.590 1762.560 1000.630 ;
        RECT 1766.100 999.930 1766.240 1000.630 ;
        RECT 1766.560 1000.270 1766.700 1000.630 ;
        RECT 1766.500 999.950 1766.760 1000.270 ;
        RECT 1788.640 999.930 1788.780 1000.630 ;
        RECT 1885.180 1000.290 1885.440 1000.610 ;
        RECT 1766.040 999.610 1766.300 999.930 ;
        RECT 1788.580 999.610 1788.840 999.930 ;
        RECT 860.760 999.270 861.020 999.590 ;
        RECT 1007.500 999.445 1007.760 999.590 ;
        RECT 1008.420 999.445 1008.680 999.590 ;
        RECT 1007.490 999.075 1007.770 999.445 ;
        RECT 1008.410 999.075 1008.690 999.445 ;
        RECT 1070.520 999.270 1070.780 999.590 ;
        RECT 1096.740 999.270 1097.000 999.590 ;
        RECT 1174.940 999.270 1175.200 999.590 ;
        RECT 1220.480 999.270 1220.740 999.590 ;
        RECT 1232.900 999.270 1233.160 999.590 ;
        RECT 1242.100 999.445 1242.360 999.590 ;
        RECT 1242.090 999.075 1242.370 999.445 ;
        RECT 1398.500 999.270 1398.760 999.590 ;
        RECT 1421.500 999.270 1421.760 999.590 ;
        RECT 1435.300 999.270 1435.560 999.590 ;
        RECT 1563.180 999.270 1563.440 999.590 ;
        RECT 1577.900 999.270 1578.160 999.590 ;
        RECT 1666.680 999.270 1666.940 999.590 ;
        RECT 1762.360 999.270 1762.620 999.590 ;
        RECT 1885.240 999.250 1885.380 1000.290 ;
        RECT 1950.960 999.950 1951.220 1000.270 ;
        RECT 2149.680 999.950 2149.940 1000.270 ;
        RECT 1951.020 999.590 1951.160 999.950 ;
        RECT 2149.740 999.590 2149.880 999.950 ;
        RECT 1950.960 999.270 1951.220 999.590 ;
        RECT 2149.680 999.270 2149.940 999.590 ;
        RECT 1885.180 998.930 1885.440 999.250 ;
        RECT 2181.420 998.250 2181.680 998.570 ;
        RECT 2181.480 867.525 2181.620 998.250 ;
        RECT 2181.410 867.155 2181.690 867.525 ;
      LAYER via2 ;
        RECT 20.330 2836.480 20.610 2836.760 ;
        RECT 1070.510 999.800 1070.790 1000.080 ;
        RECT 1096.730 999.800 1097.010 1000.080 ;
        RECT 1159.290 999.800 1159.570 1000.080 ;
        RECT 1174.930 999.800 1175.210 1000.080 ;
        RECT 1276.590 999.800 1276.870 1000.080 ;
        RECT 1007.490 999.120 1007.770 999.400 ;
        RECT 1008.410 999.120 1008.690 999.400 ;
        RECT 1242.090 999.120 1242.370 999.400 ;
        RECT 2181.410 867.200 2181.690 867.480 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 20.305 2836.770 20.635 2836.785 ;
        RECT -4.800 2836.470 20.635 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 20.305 2836.455 20.635 2836.470 ;
        RECT 1070.485 1000.090 1070.815 1000.105 ;
        RECT 1096.705 1000.090 1097.035 1000.105 ;
        RECT 1070.485 999.790 1097.035 1000.090 ;
        RECT 1070.485 999.775 1070.815 999.790 ;
        RECT 1096.705 999.775 1097.035 999.790 ;
        RECT 1159.265 1000.090 1159.595 1000.105 ;
        RECT 1174.905 1000.090 1175.235 1000.105 ;
        RECT 1276.565 1000.090 1276.895 1000.105 ;
        RECT 1159.265 999.790 1175.235 1000.090 ;
        RECT 1159.265 999.775 1159.595 999.790 ;
        RECT 1174.905 999.775 1175.235 999.790 ;
        RECT 1242.310 999.790 1276.895 1000.090 ;
        RECT 1242.310 999.425 1242.610 999.790 ;
        RECT 1276.565 999.775 1276.895 999.790 ;
        RECT 1007.465 999.410 1007.795 999.425 ;
        RECT 1008.385 999.410 1008.715 999.425 ;
        RECT 1007.465 999.110 1008.715 999.410 ;
        RECT 1007.465 999.095 1007.795 999.110 ;
        RECT 1008.385 999.095 1008.715 999.110 ;
        RECT 1242.065 999.110 1242.610 999.425 ;
        RECT 1242.065 999.095 1242.395 999.110 ;
        RECT 2181.385 867.490 2181.715 867.505 ;
        RECT 2169.670 867.190 2181.715 867.490 ;
        RECT 2169.670 865.160 2169.970 867.190 ;
        RECT 2181.385 867.175 2181.715 867.190 ;
        RECT 2166.000 864.560 2170.000 865.160 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 1005.620 19.710 1005.680 ;
        RECT 2181.850 1005.620 2182.170 1005.680 ;
        RECT 19.390 1005.480 2182.170 1005.620 ;
        RECT 19.390 1005.420 19.710 1005.480 ;
        RECT 2181.850 1005.420 2182.170 1005.480 ;
      LAYER via ;
        RECT 19.420 1005.420 19.680 1005.680 ;
        RECT 2181.880 1005.420 2182.140 1005.680 ;
      LAYER met2 ;
        RECT 19.410 2549.475 19.690 2549.845 ;
        RECT 19.480 1005.710 19.620 2549.475 ;
        RECT 19.420 1005.390 19.680 1005.710 ;
        RECT 2181.880 1005.390 2182.140 1005.710 ;
        RECT 2181.940 876.365 2182.080 1005.390 ;
        RECT 2181.870 875.995 2182.150 876.365 ;
      LAYER via2 ;
        RECT 19.410 2549.520 19.690 2549.800 ;
        RECT 2181.870 876.040 2182.150 876.320 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 19.385 2549.810 19.715 2549.825 ;
        RECT -4.800 2549.510 19.715 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 19.385 2549.495 19.715 2549.510 ;
        RECT 2181.845 876.330 2182.175 876.345 ;
        RECT 2169.670 876.030 2182.175 876.330 ;
        RECT 2169.670 874.680 2169.970 876.030 ;
        RECT 2181.845 876.015 2182.175 876.030 ;
        RECT 2166.000 874.080 2170.000 874.680 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2256.820 20.630 2256.880 ;
        RECT 2170.350 2256.820 2170.670 2256.880 ;
        RECT 20.310 2256.680 2170.670 2256.820 ;
        RECT 20.310 2256.620 20.630 2256.680 ;
        RECT 2170.350 2256.620 2170.670 2256.680 ;
      LAYER via ;
        RECT 20.340 2256.620 20.600 2256.880 ;
        RECT 2170.380 2256.620 2170.640 2256.880 ;
      LAYER met2 ;
        RECT 20.330 2261.835 20.610 2262.205 ;
        RECT 20.400 2256.910 20.540 2261.835 ;
        RECT 20.340 2256.590 20.600 2256.910 ;
        RECT 2170.380 2256.590 2170.640 2256.910 ;
        RECT 2170.440 887.245 2170.580 2256.590 ;
        RECT 2170.370 886.875 2170.650 887.245 ;
      LAYER via2 ;
        RECT 20.330 2261.880 20.610 2262.160 ;
        RECT 2170.370 886.920 2170.650 887.200 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 20.305 2262.170 20.635 2262.185 ;
        RECT -4.800 2261.870 20.635 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 20.305 2261.855 20.635 2261.870 ;
        RECT 2170.345 887.210 2170.675 887.225 ;
        RECT 2169.670 886.910 2170.675 887.210 ;
        RECT 2169.670 884.880 2169.970 886.910 ;
        RECT 2170.345 886.895 2170.675 886.910 ;
        RECT 2166.000 884.280 2170.000 884.880 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 14.330 1052.200 14.650 1052.260 ;
        RECT 16.170 1052.200 16.490 1052.260 ;
        RECT 14.330 1052.060 16.490 1052.200 ;
        RECT 14.330 1052.000 14.650 1052.060 ;
        RECT 16.170 1052.000 16.490 1052.060 ;
        RECT 14.330 1005.280 14.650 1005.340 ;
        RECT 2182.310 1005.280 2182.630 1005.340 ;
        RECT 14.330 1005.140 2182.630 1005.280 ;
        RECT 14.330 1005.080 14.650 1005.140 ;
        RECT 2182.310 1005.080 2182.630 1005.140 ;
      LAYER via ;
        RECT 14.360 1052.000 14.620 1052.260 ;
        RECT 16.200 1052.000 16.460 1052.260 ;
        RECT 14.360 1005.080 14.620 1005.340 ;
        RECT 2182.340 1005.080 2182.600 1005.340 ;
      LAYER met2 ;
        RECT 16.190 1974.875 16.470 1975.245 ;
        RECT 16.260 1052.290 16.400 1974.875 ;
        RECT 14.360 1051.970 14.620 1052.290 ;
        RECT 16.200 1051.970 16.460 1052.290 ;
        RECT 14.420 1005.370 14.560 1051.970 ;
        RECT 14.360 1005.050 14.620 1005.370 ;
        RECT 2182.340 1005.050 2182.600 1005.370 ;
        RECT 2182.400 896.765 2182.540 1005.050 ;
        RECT 2182.330 896.395 2182.610 896.765 ;
      LAYER via2 ;
        RECT 16.190 1974.920 16.470 1975.200 ;
        RECT 2182.330 896.440 2182.610 896.720 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 16.165 1975.210 16.495 1975.225 ;
        RECT -4.800 1974.910 16.495 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 16.165 1974.895 16.495 1974.910 ;
        RECT 2182.305 896.730 2182.635 896.745 ;
        RECT 2169.670 896.430 2182.635 896.730 ;
        RECT 2169.670 895.080 2169.970 896.430 ;
        RECT 2182.305 896.415 2182.635 896.430 ;
        RECT 2166.000 894.480 2170.000 895.080 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2184.610 558.860 2184.930 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2184.610 558.720 2899.310 558.860 ;
        RECT 2184.610 558.660 2184.930 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2184.640 558.660 2184.900 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2184.630 621.675 2184.910 622.045 ;
        RECT 2184.700 558.950 2184.840 621.675 ;
        RECT 2184.640 558.630 2184.900 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2184.630 621.720 2184.910 622.000 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2166.000 624.520 2170.000 625.120 ;
        RECT 2169.670 622.010 2169.970 624.520 ;
        RECT 2184.605 622.010 2184.935 622.025 ;
        RECT 2169.670 621.710 2184.935 622.010 ;
        RECT 2184.605 621.695 2184.935 621.710 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 1683.920 16.030 1683.980 ;
        RECT 2169.890 1683.920 2170.210 1683.980 ;
        RECT 15.710 1683.780 2170.210 1683.920 ;
        RECT 15.710 1683.720 16.030 1683.780 ;
        RECT 2169.890 1683.720 2170.210 1683.780 ;
      LAYER via ;
        RECT 15.740 1683.720 16.000 1683.980 ;
        RECT 2169.920 1683.720 2170.180 1683.980 ;
      LAYER met2 ;
        RECT 15.730 1687.235 16.010 1687.605 ;
        RECT 15.800 1684.010 15.940 1687.235 ;
        RECT 15.740 1683.690 16.000 1684.010 ;
        RECT 2169.920 1683.690 2170.180 1684.010 ;
        RECT 2169.980 907.645 2170.120 1683.690 ;
        RECT 2169.910 907.275 2170.190 907.645 ;
      LAYER via2 ;
        RECT 15.730 1687.280 16.010 1687.560 ;
        RECT 2169.910 907.320 2170.190 907.600 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 15.705 1687.570 16.035 1687.585 ;
        RECT -4.800 1687.270 16.035 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 15.705 1687.255 16.035 1687.270 ;
        RECT 2169.885 907.610 2170.215 907.625 ;
        RECT 2169.670 907.295 2170.215 907.610 ;
        RECT 2169.670 905.280 2169.970 907.295 ;
        RECT 2166.000 904.680 2170.000 905.280 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 1470.060 15.570 1470.120 ;
        RECT 2174.030 1470.060 2174.350 1470.120 ;
        RECT 15.250 1469.920 2174.350 1470.060 ;
        RECT 15.250 1469.860 15.570 1469.920 ;
        RECT 2174.030 1469.860 2174.350 1469.920 ;
      LAYER via ;
        RECT 15.280 1469.860 15.540 1470.120 ;
        RECT 2174.060 1469.860 2174.320 1470.120 ;
      LAYER met2 ;
        RECT 15.270 1471.675 15.550 1472.045 ;
        RECT 15.340 1470.150 15.480 1471.675 ;
        RECT 15.280 1469.830 15.540 1470.150 ;
        RECT 2174.060 1469.830 2174.320 1470.150 ;
        RECT 2174.120 917.165 2174.260 1469.830 ;
        RECT 2174.050 916.795 2174.330 917.165 ;
      LAYER via2 ;
        RECT 15.270 1471.720 15.550 1472.000 ;
        RECT 2174.050 916.840 2174.330 917.120 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 15.245 1472.010 15.575 1472.025 ;
        RECT -4.800 1471.710 15.575 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 15.245 1471.695 15.575 1471.710 ;
        RECT 2174.025 917.130 2174.355 917.145 ;
        RECT 2169.670 916.830 2174.355 917.130 ;
        RECT 2169.670 914.800 2169.970 916.830 ;
        RECT 2174.025 916.815 2174.355 916.830 ;
        RECT 2166.000 914.200 2170.000 914.800 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1328.090 1257.220 1328.410 1257.280 ;
        RECT 1352.010 1257.220 1352.330 1257.280 ;
        RECT 1328.090 1257.080 1352.330 1257.220 ;
        RECT 1328.090 1257.020 1328.410 1257.080 ;
        RECT 1352.010 1257.020 1352.330 1257.080 ;
        RECT 14.790 1256.200 15.110 1256.260 ;
        RECT 1328.090 1256.200 1328.410 1256.260 ;
        RECT 14.790 1256.060 1328.410 1256.200 ;
        RECT 14.790 1256.000 15.110 1256.060 ;
        RECT 1328.090 1256.000 1328.410 1256.060 ;
        RECT 1352.010 1256.200 1352.330 1256.260 ;
        RECT 2169.430 1256.200 2169.750 1256.260 ;
        RECT 1352.010 1256.060 2169.750 1256.200 ;
        RECT 1352.010 1256.000 1352.330 1256.060 ;
        RECT 2169.430 1256.000 2169.750 1256.060 ;
      LAYER via ;
        RECT 1328.120 1257.020 1328.380 1257.280 ;
        RECT 1352.040 1257.020 1352.300 1257.280 ;
        RECT 14.820 1256.000 15.080 1256.260 ;
        RECT 1328.120 1256.000 1328.380 1256.260 ;
        RECT 1352.040 1256.000 1352.300 1256.260 ;
        RECT 2169.460 1256.000 2169.720 1256.260 ;
      LAYER met2 ;
        RECT 1328.120 1256.990 1328.380 1257.310 ;
        RECT 1352.040 1256.990 1352.300 1257.310 ;
        RECT 14.810 1256.115 15.090 1256.485 ;
        RECT 1328.180 1256.290 1328.320 1256.990 ;
        RECT 1352.100 1256.290 1352.240 1256.990 ;
        RECT 14.820 1255.970 15.080 1256.115 ;
        RECT 1328.120 1255.970 1328.380 1256.290 ;
        RECT 1352.040 1255.970 1352.300 1256.290 ;
        RECT 2169.460 1255.970 2169.720 1256.290 ;
        RECT 2169.520 923.965 2169.660 1255.970 ;
        RECT 2169.450 923.595 2169.730 923.965 ;
      LAYER via2 ;
        RECT 14.810 1256.160 15.090 1256.440 ;
        RECT 2169.450 923.640 2169.730 923.920 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 14.785 1256.450 15.115 1256.465 ;
        RECT -4.800 1256.150 15.115 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 14.785 1256.135 15.115 1256.150 ;
        RECT 2166.000 924.400 2170.000 925.000 ;
        RECT 2169.670 923.945 2169.970 924.400 ;
        RECT 2169.425 923.630 2169.970 923.945 ;
        RECT 2169.425 923.615 2169.755 923.630 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 1035.200 16.490 1035.260 ;
        RECT 2174.490 1035.200 2174.810 1035.260 ;
        RECT 16.170 1035.060 2174.810 1035.200 ;
        RECT 16.170 1035.000 16.490 1035.060 ;
        RECT 2174.490 1035.000 2174.810 1035.060 ;
      LAYER via ;
        RECT 16.200 1035.000 16.460 1035.260 ;
        RECT 2174.520 1035.000 2174.780 1035.260 ;
      LAYER met2 ;
        RECT 16.190 1040.555 16.470 1040.925 ;
        RECT 16.260 1035.290 16.400 1040.555 ;
        RECT 16.200 1034.970 16.460 1035.290 ;
        RECT 2174.520 1034.970 2174.780 1035.290 ;
        RECT 2174.580 937.565 2174.720 1034.970 ;
        RECT 2174.510 937.195 2174.790 937.565 ;
      LAYER via2 ;
        RECT 16.190 1040.600 16.470 1040.880 ;
        RECT 2174.510 937.240 2174.790 937.520 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 16.165 1040.890 16.495 1040.905 ;
        RECT -4.800 1040.590 16.495 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 16.165 1040.575 16.495 1040.590 ;
        RECT 2174.485 937.530 2174.815 937.545 ;
        RECT 2169.670 937.230 2174.815 937.530 ;
        RECT 2169.670 935.200 2169.970 937.230 ;
        RECT 2174.485 937.215 2174.815 937.230 ;
        RECT 2166.000 934.600 2170.000 935.200 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.770 1000.860 1815.090 1000.920 ;
        RECT 1838.230 1000.860 1838.550 1000.920 ;
        RECT 1814.770 1000.720 1838.550 1000.860 ;
        RECT 1814.770 1000.660 1815.090 1000.720 ;
        RECT 1838.230 1000.660 1838.550 1000.720 ;
        RECT 2165.840 1000.720 2166.900 1000.860 ;
        RECT 2091.230 1000.520 2091.550 1000.580 ;
        RECT 2165.840 1000.520 2165.980 1000.720 ;
        RECT 2091.230 1000.380 2165.980 1000.520 ;
        RECT 2166.760 1000.520 2166.900 1000.720 ;
        RECT 2180.930 1000.520 2181.250 1000.580 ;
        RECT 2166.760 1000.380 2181.250 1000.520 ;
        RECT 2091.230 1000.320 2091.550 1000.380 ;
        RECT 2180.930 1000.320 2181.250 1000.380 ;
        RECT 1069.110 1000.180 1069.430 1000.240 ;
        RECT 1069.110 1000.040 1073.940 1000.180 ;
        RECT 1069.110 999.980 1069.430 1000.040 ;
        RECT 13.870 999.160 14.190 999.220 ;
        RECT 834.510 999.160 834.830 999.220 ;
        RECT 13.870 999.020 834.830 999.160 ;
        RECT 13.870 998.960 14.190 999.020 ;
        RECT 834.510 998.960 834.830 999.020 ;
        RECT 838.190 999.160 838.510 999.220 ;
        RECT 862.570 999.160 862.890 999.220 ;
        RECT 838.190 999.020 862.890 999.160 ;
        RECT 838.190 998.960 838.510 999.020 ;
        RECT 862.570 998.960 862.890 999.020 ;
        RECT 883.730 999.160 884.050 999.220 ;
        RECT 933.870 999.160 934.190 999.220 ;
        RECT 883.730 999.020 934.190 999.160 ;
        RECT 883.730 998.960 884.050 999.020 ;
        RECT 933.870 998.960 934.190 999.020 ;
        RECT 935.710 999.160 936.030 999.220 ;
        RECT 957.790 999.160 958.110 999.220 ;
        RECT 935.710 999.020 958.110 999.160 ;
        RECT 935.710 998.960 936.030 999.020 ;
        RECT 957.790 998.960 958.110 999.020 ;
        RECT 959.630 999.160 959.950 999.220 ;
        RECT 1069.110 999.160 1069.430 999.220 ;
        RECT 959.630 999.020 1069.430 999.160 ;
        RECT 1073.800 999.160 1073.940 1000.040 ;
        RECT 1253.660 999.700 1270.360 999.840 ;
        RECT 1172.150 999.500 1172.470 999.560 ;
        RECT 1159.820 999.360 1172.470 999.500 ;
        RECT 1159.820 999.160 1159.960 999.360 ;
        RECT 1172.150 999.300 1172.470 999.360 ;
        RECT 1253.110 999.500 1253.430 999.560 ;
        RECT 1253.660 999.500 1253.800 999.700 ;
        RECT 1253.110 999.360 1253.800 999.500 ;
        RECT 1253.110 999.300 1253.430 999.360 ;
        RECT 1073.800 999.020 1159.960 999.160 ;
        RECT 1173.070 999.160 1173.390 999.220 ;
        RECT 1219.990 999.160 1220.310 999.220 ;
        RECT 1173.070 999.020 1220.310 999.160 ;
        RECT 959.630 998.960 959.950 999.020 ;
        RECT 1069.110 998.960 1069.430 999.020 ;
        RECT 1173.070 998.960 1173.390 999.020 ;
        RECT 1219.990 998.960 1220.310 999.020 ;
        RECT 1222.750 999.160 1223.070 999.220 ;
        RECT 1252.190 999.160 1252.510 999.220 ;
        RECT 1222.750 999.020 1252.510 999.160 ;
        RECT 1270.220 999.160 1270.360 999.700 ;
        RECT 1362.680 999.700 1371.560 999.840 ;
        RECT 1352.470 999.160 1352.790 999.220 ;
        RECT 1270.220 999.020 1352.790 999.160 ;
        RECT 1222.750 998.960 1223.070 999.020 ;
        RECT 1252.190 998.960 1252.510 999.020 ;
        RECT 1352.470 998.960 1352.790 999.020 ;
        RECT 1352.930 999.160 1353.250 999.220 ;
        RECT 1362.680 999.160 1362.820 999.700 ;
        RECT 1352.930 999.020 1362.820 999.160 ;
        RECT 1371.420 999.160 1371.560 999.700 ;
        RECT 1400.310 999.160 1400.630 999.220 ;
        RECT 1371.420 999.020 1400.630 999.160 ;
        RECT 1352.930 998.960 1353.250 999.020 ;
        RECT 1400.310 998.960 1400.630 999.020 ;
        RECT 1415.030 999.160 1415.350 999.220 ;
        RECT 1452.750 999.160 1453.070 999.220 ;
        RECT 1415.030 999.020 1453.070 999.160 ;
        RECT 1415.030 998.960 1415.350 999.020 ;
        RECT 1452.750 998.960 1453.070 999.020 ;
        RECT 1464.710 999.160 1465.030 999.220 ;
        RECT 1559.010 999.160 1559.330 999.220 ;
        RECT 1464.710 999.020 1559.330 999.160 ;
        RECT 1464.710 998.960 1465.030 999.020 ;
        RECT 1559.010 998.960 1559.330 999.020 ;
        RECT 1578.330 999.160 1578.650 999.220 ;
        RECT 1642.730 999.160 1643.050 999.220 ;
        RECT 1578.330 999.020 1643.050 999.160 ;
        RECT 1578.330 998.960 1578.650 999.020 ;
        RECT 1642.730 998.960 1643.050 999.020 ;
        RECT 1657.910 999.160 1658.230 999.220 ;
        RECT 1762.790 999.160 1763.110 999.220 ;
        RECT 1657.910 999.020 1763.110 999.160 ;
        RECT 1657.910 998.960 1658.230 999.020 ;
        RECT 1762.790 998.960 1763.110 999.020 ;
        RECT 1786.250 999.160 1786.570 999.220 ;
        RECT 1814.770 999.160 1815.090 999.220 ;
        RECT 1786.250 999.020 1815.090 999.160 ;
        RECT 1786.250 998.960 1786.570 999.020 ;
        RECT 1814.770 998.960 1815.090 999.020 ;
        RECT 1838.230 999.160 1838.550 999.220 ;
        RECT 1883.770 999.160 1884.090 999.220 ;
        RECT 1838.230 999.020 1884.090 999.160 ;
        RECT 1838.230 998.960 1838.550 999.020 ;
        RECT 1883.770 998.960 1884.090 999.020 ;
        RECT 1909.530 999.160 1909.850 999.220 ;
        RECT 1931.610 999.160 1931.930 999.220 ;
        RECT 1909.530 999.020 1931.930 999.160 ;
        RECT 1909.530 998.960 1909.850 999.020 ;
        RECT 1931.610 998.960 1931.930 999.020 ;
        RECT 1950.470 999.160 1950.790 999.220 ;
        RECT 2091.230 999.160 2091.550 999.220 ;
        RECT 1950.470 999.020 2091.550 999.160 ;
        RECT 1950.470 998.960 1950.790 999.020 ;
        RECT 2091.230 998.960 2091.550 999.020 ;
      LAYER via ;
        RECT 1814.800 1000.660 1815.060 1000.920 ;
        RECT 1838.260 1000.660 1838.520 1000.920 ;
        RECT 2091.260 1000.320 2091.520 1000.580 ;
        RECT 2180.960 1000.320 2181.220 1000.580 ;
        RECT 1069.140 999.980 1069.400 1000.240 ;
        RECT 13.900 998.960 14.160 999.220 ;
        RECT 834.540 998.960 834.800 999.220 ;
        RECT 838.220 998.960 838.480 999.220 ;
        RECT 862.600 998.960 862.860 999.220 ;
        RECT 883.760 998.960 884.020 999.220 ;
        RECT 933.900 998.960 934.160 999.220 ;
        RECT 935.740 998.960 936.000 999.220 ;
        RECT 957.820 998.960 958.080 999.220 ;
        RECT 959.660 998.960 959.920 999.220 ;
        RECT 1069.140 998.960 1069.400 999.220 ;
        RECT 1172.180 999.300 1172.440 999.560 ;
        RECT 1253.140 999.300 1253.400 999.560 ;
        RECT 1173.100 998.960 1173.360 999.220 ;
        RECT 1220.020 998.960 1220.280 999.220 ;
        RECT 1222.780 998.960 1223.040 999.220 ;
        RECT 1252.220 998.960 1252.480 999.220 ;
        RECT 1352.500 998.960 1352.760 999.220 ;
        RECT 1352.960 998.960 1353.220 999.220 ;
        RECT 1400.340 998.960 1400.600 999.220 ;
        RECT 1415.060 998.960 1415.320 999.220 ;
        RECT 1452.780 998.960 1453.040 999.220 ;
        RECT 1464.740 998.960 1465.000 999.220 ;
        RECT 1559.040 998.960 1559.300 999.220 ;
        RECT 1578.360 998.960 1578.620 999.220 ;
        RECT 1642.760 998.960 1643.020 999.220 ;
        RECT 1657.940 998.960 1658.200 999.220 ;
        RECT 1762.820 998.960 1763.080 999.220 ;
        RECT 1786.280 998.960 1786.540 999.220 ;
        RECT 1814.800 998.960 1815.060 999.220 ;
        RECT 1838.260 998.960 1838.520 999.220 ;
        RECT 1883.800 998.960 1884.060 999.220 ;
        RECT 1909.560 998.960 1909.820 999.220 ;
        RECT 1931.640 998.960 1931.900 999.220 ;
        RECT 1950.500 998.960 1950.760 999.220 ;
        RECT 2091.260 998.960 2091.520 999.220 ;
      LAYER met2 ;
        RECT 1814.800 1000.630 1815.060 1000.950 ;
        RECT 1838.260 1000.630 1838.520 1000.950 ;
        RECT 1069.140 999.950 1069.400 1000.270 ;
        RECT 13.900 998.930 14.160 999.250 ;
        RECT 834.530 999.075 834.810 999.445 ;
        RECT 838.210 999.075 838.490 999.445 ;
        RECT 862.590 999.075 862.870 999.445 ;
        RECT 883.750 999.075 884.030 999.445 ;
        RECT 933.890 999.075 934.170 999.445 ;
        RECT 935.730 999.075 936.010 999.445 ;
        RECT 957.810 999.075 958.090 999.445 ;
        RECT 959.650 999.075 959.930 999.445 ;
        RECT 1069.200 999.250 1069.340 999.950 ;
        RECT 1172.180 999.330 1172.440 999.590 ;
        RECT 1172.180 999.270 1173.300 999.330 ;
        RECT 1172.240 999.250 1173.300 999.270 ;
        RECT 834.540 998.930 834.800 999.075 ;
        RECT 838.220 998.930 838.480 999.075 ;
        RECT 862.600 998.930 862.860 999.075 ;
        RECT 883.760 998.930 884.020 999.075 ;
        RECT 933.900 998.930 934.160 999.075 ;
        RECT 935.740 998.930 936.000 999.075 ;
        RECT 957.820 998.930 958.080 999.075 ;
        RECT 959.660 998.930 959.920 999.075 ;
        RECT 1069.140 998.930 1069.400 999.250 ;
        RECT 1172.240 999.190 1173.360 999.250 ;
        RECT 1173.100 998.930 1173.360 999.190 ;
        RECT 1220.010 999.075 1220.290 999.445 ;
        RECT 1222.770 999.075 1223.050 999.445 ;
        RECT 1253.140 999.330 1253.400 999.590 ;
        RECT 1252.280 999.270 1253.400 999.330 ;
        RECT 1252.280 999.250 1253.340 999.270 ;
        RECT 1352.560 999.250 1353.160 999.330 ;
        RECT 1252.220 999.190 1253.340 999.250 ;
        RECT 1352.500 999.190 1353.220 999.250 ;
        RECT 1220.020 998.930 1220.280 999.075 ;
        RECT 1222.780 998.930 1223.040 999.075 ;
        RECT 1252.220 998.930 1252.480 999.190 ;
        RECT 1352.500 998.930 1352.760 999.190 ;
        RECT 1352.960 998.930 1353.220 999.190 ;
        RECT 1400.330 999.075 1400.610 999.445 ;
        RECT 1415.050 999.075 1415.330 999.445 ;
        RECT 1452.770 999.075 1453.050 999.445 ;
        RECT 1464.730 999.075 1465.010 999.445 ;
        RECT 1559.030 999.075 1559.310 999.445 ;
        RECT 1578.350 999.075 1578.630 999.445 ;
        RECT 1642.750 999.075 1643.030 999.445 ;
        RECT 1657.930 999.075 1658.210 999.445 ;
        RECT 1762.810 999.075 1763.090 999.445 ;
        RECT 1786.270 999.075 1786.550 999.445 ;
        RECT 1814.860 999.250 1815.000 1000.630 ;
        RECT 1838.320 999.250 1838.460 1000.630 ;
        RECT 2091.260 1000.290 2091.520 1000.610 ;
        RECT 2180.960 1000.290 2181.220 1000.610 ;
        RECT 1400.340 998.930 1400.600 999.075 ;
        RECT 1415.060 998.930 1415.320 999.075 ;
        RECT 1452.780 998.930 1453.040 999.075 ;
        RECT 1464.740 998.930 1465.000 999.075 ;
        RECT 1559.040 998.930 1559.300 999.075 ;
        RECT 1578.360 998.930 1578.620 999.075 ;
        RECT 1642.760 998.930 1643.020 999.075 ;
        RECT 1657.940 998.930 1658.200 999.075 ;
        RECT 1762.820 998.930 1763.080 999.075 ;
        RECT 1786.280 998.930 1786.540 999.075 ;
        RECT 1814.800 998.930 1815.060 999.250 ;
        RECT 1838.260 998.930 1838.520 999.250 ;
        RECT 1883.790 999.075 1884.070 999.445 ;
        RECT 1909.550 999.075 1909.830 999.445 ;
        RECT 1931.630 999.075 1931.910 999.445 ;
        RECT 1950.490 999.075 1950.770 999.445 ;
        RECT 2091.320 999.250 2091.460 1000.290 ;
        RECT 1883.800 998.930 1884.060 999.075 ;
        RECT 1909.560 998.930 1909.820 999.075 ;
        RECT 1931.640 998.930 1931.900 999.075 ;
        RECT 1950.500 998.930 1950.760 999.075 ;
        RECT 2091.260 998.930 2091.520 999.250 ;
        RECT 13.960 825.365 14.100 998.930 ;
        RECT 2181.020 945.045 2181.160 1000.290 ;
        RECT 2180.950 944.675 2181.230 945.045 ;
        RECT 13.890 824.995 14.170 825.365 ;
      LAYER via2 ;
        RECT 834.530 999.120 834.810 999.400 ;
        RECT 838.210 999.120 838.490 999.400 ;
        RECT 862.590 999.120 862.870 999.400 ;
        RECT 883.750 999.120 884.030 999.400 ;
        RECT 933.890 999.120 934.170 999.400 ;
        RECT 935.730 999.120 936.010 999.400 ;
        RECT 957.810 999.120 958.090 999.400 ;
        RECT 959.650 999.120 959.930 999.400 ;
        RECT 1220.010 999.120 1220.290 999.400 ;
        RECT 1222.770 999.120 1223.050 999.400 ;
        RECT 1400.330 999.120 1400.610 999.400 ;
        RECT 1415.050 999.120 1415.330 999.400 ;
        RECT 1452.770 999.120 1453.050 999.400 ;
        RECT 1464.730 999.120 1465.010 999.400 ;
        RECT 1559.030 999.120 1559.310 999.400 ;
        RECT 1578.350 999.120 1578.630 999.400 ;
        RECT 1642.750 999.120 1643.030 999.400 ;
        RECT 1657.930 999.120 1658.210 999.400 ;
        RECT 1762.810 999.120 1763.090 999.400 ;
        RECT 1786.270 999.120 1786.550 999.400 ;
        RECT 1883.790 999.120 1884.070 999.400 ;
        RECT 1909.550 999.120 1909.830 999.400 ;
        RECT 1931.630 999.120 1931.910 999.400 ;
        RECT 1950.490 999.120 1950.770 999.400 ;
        RECT 2180.950 944.720 2181.230 945.000 ;
        RECT 13.890 825.040 14.170 825.320 ;
      LAYER met3 ;
        RECT 834.505 999.410 834.835 999.425 ;
        RECT 838.185 999.410 838.515 999.425 ;
        RECT 834.505 999.110 838.515 999.410 ;
        RECT 834.505 999.095 834.835 999.110 ;
        RECT 838.185 999.095 838.515 999.110 ;
        RECT 862.565 999.410 862.895 999.425 ;
        RECT 883.725 999.410 884.055 999.425 ;
        RECT 862.565 999.110 884.055 999.410 ;
        RECT 862.565 999.095 862.895 999.110 ;
        RECT 883.725 999.095 884.055 999.110 ;
        RECT 933.865 999.410 934.195 999.425 ;
        RECT 935.705 999.410 936.035 999.425 ;
        RECT 933.865 999.110 936.035 999.410 ;
        RECT 933.865 999.095 934.195 999.110 ;
        RECT 935.705 999.095 936.035 999.110 ;
        RECT 957.785 999.410 958.115 999.425 ;
        RECT 959.625 999.410 959.955 999.425 ;
        RECT 957.785 999.110 959.955 999.410 ;
        RECT 957.785 999.095 958.115 999.110 ;
        RECT 959.625 999.095 959.955 999.110 ;
        RECT 1219.985 999.410 1220.315 999.425 ;
        RECT 1222.745 999.410 1223.075 999.425 ;
        RECT 1219.985 999.110 1223.075 999.410 ;
        RECT 1219.985 999.095 1220.315 999.110 ;
        RECT 1222.745 999.095 1223.075 999.110 ;
        RECT 1400.305 999.410 1400.635 999.425 ;
        RECT 1415.025 999.410 1415.355 999.425 ;
        RECT 1400.305 999.110 1415.355 999.410 ;
        RECT 1400.305 999.095 1400.635 999.110 ;
        RECT 1415.025 999.095 1415.355 999.110 ;
        RECT 1452.745 999.410 1453.075 999.425 ;
        RECT 1464.705 999.410 1465.035 999.425 ;
        RECT 1452.745 999.110 1465.035 999.410 ;
        RECT 1452.745 999.095 1453.075 999.110 ;
        RECT 1464.705 999.095 1465.035 999.110 ;
        RECT 1559.005 999.410 1559.335 999.425 ;
        RECT 1578.325 999.410 1578.655 999.425 ;
        RECT 1559.005 999.110 1578.655 999.410 ;
        RECT 1559.005 999.095 1559.335 999.110 ;
        RECT 1578.325 999.095 1578.655 999.110 ;
        RECT 1642.725 999.410 1643.055 999.425 ;
        RECT 1657.905 999.410 1658.235 999.425 ;
        RECT 1642.725 999.110 1658.235 999.410 ;
        RECT 1642.725 999.095 1643.055 999.110 ;
        RECT 1657.905 999.095 1658.235 999.110 ;
        RECT 1762.785 999.410 1763.115 999.425 ;
        RECT 1786.245 999.410 1786.575 999.425 ;
        RECT 1883.765 999.410 1884.095 999.425 ;
        RECT 1909.525 999.410 1909.855 999.425 ;
        RECT 1762.785 999.110 1786.575 999.410 ;
        RECT 1762.785 999.095 1763.115 999.110 ;
        RECT 1786.245 999.095 1786.575 999.110 ;
        RECT 1883.550 999.095 1884.095 999.410 ;
        RECT 1909.310 999.095 1909.855 999.410 ;
        RECT 1931.605 999.410 1931.935 999.425 ;
        RECT 1950.465 999.410 1950.795 999.425 ;
        RECT 1931.605 999.110 1950.795 999.410 ;
        RECT 1931.605 999.095 1931.935 999.110 ;
        RECT 1950.465 999.095 1950.795 999.110 ;
        RECT 1883.550 998.730 1883.850 999.095 ;
        RECT 1909.310 998.730 1909.610 999.095 ;
        RECT 1883.550 998.430 1909.610 998.730 ;
        RECT 2180.925 945.010 2181.255 945.025 ;
        RECT 2169.670 944.720 2181.255 945.010 ;
        RECT 2166.000 944.710 2181.255 944.720 ;
        RECT 2166.000 944.120 2170.000 944.710 ;
        RECT 2180.925 944.695 2181.255 944.710 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 13.865 825.330 14.195 825.345 ;
        RECT -4.800 825.030 14.195 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 13.865 825.015 14.195 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 603.060 17.870 603.120 ;
        RECT 669.370 603.060 669.690 603.120 ;
        RECT 2183.230 603.060 2183.550 603.120 ;
        RECT 17.550 602.920 669.690 603.060 ;
        RECT 17.550 602.860 17.870 602.920 ;
        RECT 669.370 602.860 669.690 602.920 ;
        RECT 695.220 602.920 2183.550 603.060 ;
        RECT 695.220 601.760 695.360 602.920 ;
        RECT 2183.230 602.860 2183.550 602.920 ;
        RECT 695.130 601.500 695.450 601.760 ;
      LAYER via ;
        RECT 17.580 602.860 17.840 603.120 ;
        RECT 669.400 602.860 669.660 603.120 ;
        RECT 2183.260 602.860 2183.520 603.120 ;
        RECT 695.160 601.500 695.420 601.760 ;
      LAYER met2 ;
        RECT 2183.250 952.835 2183.530 953.205 ;
        RECT 17.570 610.115 17.850 610.485 ;
        RECT 17.640 603.150 17.780 610.115 ;
        RECT 2183.320 603.150 2183.460 952.835 ;
        RECT 17.580 602.830 17.840 603.150 ;
        RECT 669.400 602.830 669.660 603.150 ;
        RECT 2183.260 602.830 2183.520 603.150 ;
        RECT 669.460 601.645 669.600 602.830 ;
        RECT 695.160 601.645 695.420 601.790 ;
        RECT 669.390 601.275 669.670 601.645 ;
        RECT 695.150 601.275 695.430 601.645 ;
      LAYER via2 ;
        RECT 2183.250 952.880 2183.530 953.160 ;
        RECT 17.570 610.160 17.850 610.440 ;
        RECT 669.390 601.320 669.670 601.600 ;
        RECT 695.150 601.320 695.430 601.600 ;
      LAYER met3 ;
        RECT 2166.000 954.320 2170.000 954.920 ;
        RECT 2169.670 953.170 2169.970 954.320 ;
        RECT 2183.225 953.170 2183.555 953.185 ;
        RECT 2169.670 952.870 2183.555 953.170 ;
        RECT 2183.225 952.855 2183.555 952.870 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.545 610.450 17.875 610.465 ;
        RECT -4.800 610.150 17.875 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.545 610.135 17.875 610.150 ;
        RECT 669.365 601.610 669.695 601.625 ;
        RECT 695.125 601.610 695.455 601.625 ;
        RECT 669.365 601.310 695.455 601.610 ;
        RECT 669.365 601.295 669.695 601.310 ;
        RECT 695.125 601.295 695.455 601.310 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2173.570 903.760 2173.890 904.020 ;
        RECT 2173.660 903.620 2173.800 903.760 ;
        RECT 2174.030 903.620 2174.350 903.680 ;
        RECT 2173.660 903.480 2174.350 903.620 ;
        RECT 2174.030 903.420 2174.350 903.480 ;
        RECT 2173.570 821.000 2173.890 821.060 ;
        RECT 2174.950 821.000 2175.270 821.060 ;
        RECT 2173.570 820.860 2175.270 821.000 ;
        RECT 2173.570 820.800 2173.890 820.860 ;
        RECT 2174.950 820.800 2175.270 820.860 ;
        RECT 2174.490 642.160 2174.810 642.220 ;
        RECT 2174.120 642.020 2174.810 642.160 ;
        RECT 2174.120 641.540 2174.260 642.020 ;
        RECT 2174.490 641.960 2174.810 642.020 ;
        RECT 2174.030 641.280 2174.350 641.540 ;
        RECT 2174.030 600.340 2174.350 600.400 ;
        RECT 2174.950 600.340 2175.270 600.400 ;
        RECT 2174.030 600.200 2175.270 600.340 ;
        RECT 2174.030 600.140 2174.350 600.200 ;
        RECT 2174.950 600.140 2175.270 600.200 ;
        RECT 2174.950 545.400 2175.270 545.660 ;
        RECT 2175.040 544.980 2175.180 545.400 ;
        RECT 2174.950 544.720 2175.270 544.980 ;
        RECT 2174.950 496.980 2175.270 497.040 ;
        RECT 2174.580 496.840 2175.270 496.980 ;
        RECT 2174.580 496.700 2174.720 496.840 ;
        RECT 2174.950 496.780 2175.270 496.840 ;
        RECT 2174.490 496.440 2174.810 496.700 ;
        RECT 2174.490 483.040 2174.810 483.100 ;
        RECT 2175.410 483.040 2175.730 483.100 ;
        RECT 2174.490 482.900 2175.730 483.040 ;
        RECT 2174.490 482.840 2174.810 482.900 ;
        RECT 2175.410 482.840 2175.730 482.900 ;
        RECT 2174.030 435.100 2174.350 435.160 ;
        RECT 2175.410 435.100 2175.730 435.160 ;
        RECT 2174.030 434.960 2175.730 435.100 ;
        RECT 2174.030 434.900 2174.350 434.960 ;
        RECT 2175.410 434.900 2175.730 434.960 ;
        RECT 2174.030 400.760 2174.350 400.820 ;
        RECT 2174.030 400.620 2175.180 400.760 ;
        RECT 2174.030 400.560 2174.350 400.620 ;
        RECT 1932.160 400.280 1952.080 400.420 ;
        RECT 15.250 400.080 15.570 400.140 ;
        RECT 1932.160 400.080 1932.300 400.280 ;
        RECT 15.250 399.940 1932.300 400.080 ;
        RECT 1951.940 400.080 1952.080 400.280 ;
        RECT 2028.760 400.280 2055.120 400.420 ;
        RECT 2028.760 400.080 2028.900 400.280 ;
        RECT 1951.940 399.940 2028.900 400.080 ;
        RECT 2054.980 400.080 2055.120 400.280 ;
        RECT 2175.040 400.080 2175.180 400.620 ;
        RECT 2054.980 399.940 2175.180 400.080 ;
        RECT 15.250 399.880 15.570 399.940 ;
      LAYER via ;
        RECT 2173.600 903.760 2173.860 904.020 ;
        RECT 2174.060 903.420 2174.320 903.680 ;
        RECT 2173.600 820.800 2173.860 821.060 ;
        RECT 2174.980 820.800 2175.240 821.060 ;
        RECT 2174.520 641.960 2174.780 642.220 ;
        RECT 2174.060 641.280 2174.320 641.540 ;
        RECT 2174.060 600.140 2174.320 600.400 ;
        RECT 2174.980 600.140 2175.240 600.400 ;
        RECT 2174.980 545.400 2175.240 545.660 ;
        RECT 2174.980 544.720 2175.240 544.980 ;
        RECT 2174.980 496.780 2175.240 497.040 ;
        RECT 2174.520 496.440 2174.780 496.700 ;
        RECT 2174.520 482.840 2174.780 483.100 ;
        RECT 2175.440 482.840 2175.700 483.100 ;
        RECT 2174.060 434.900 2174.320 435.160 ;
        RECT 2175.440 434.900 2175.700 435.160 ;
        RECT 2174.060 400.560 2174.320 400.820 ;
        RECT 15.280 399.880 15.540 400.140 ;
      LAYER met2 ;
        RECT 2173.590 961.675 2173.870 962.045 ;
        RECT 2173.660 904.050 2173.800 961.675 ;
        RECT 2173.600 903.730 2173.860 904.050 ;
        RECT 2174.060 903.390 2174.320 903.710 ;
        RECT 2174.120 883.050 2174.260 903.390 ;
        RECT 2174.120 882.910 2174.720 883.050 ;
        RECT 2174.580 834.770 2174.720 882.910 ;
        RECT 2173.660 834.630 2174.720 834.770 ;
        RECT 2173.660 821.090 2173.800 834.630 ;
        RECT 2173.600 820.770 2173.860 821.090 ;
        RECT 2174.980 820.770 2175.240 821.090 ;
        RECT 2175.040 773.005 2175.180 820.770 ;
        RECT 2174.050 772.635 2174.330 773.005 ;
        RECT 2174.970 772.635 2175.250 773.005 ;
        RECT 2174.120 738.210 2174.260 772.635 ;
        RECT 2174.120 738.070 2174.720 738.210 ;
        RECT 2174.580 642.250 2174.720 738.070 ;
        RECT 2174.520 641.930 2174.780 642.250 ;
        RECT 2174.060 641.250 2174.320 641.570 ;
        RECT 2174.120 600.430 2174.260 641.250 ;
        RECT 2174.060 600.110 2174.320 600.430 ;
        RECT 2174.980 600.110 2175.240 600.430 ;
        RECT 2175.040 545.690 2175.180 600.110 ;
        RECT 2174.980 545.370 2175.240 545.690 ;
        RECT 2174.980 544.690 2175.240 545.010 ;
        RECT 2175.040 497.070 2175.180 544.690 ;
        RECT 2174.980 496.750 2175.240 497.070 ;
        RECT 2174.520 496.410 2174.780 496.730 ;
        RECT 2174.580 483.130 2174.720 496.410 ;
        RECT 2174.520 482.810 2174.780 483.130 ;
        RECT 2175.440 482.810 2175.700 483.130 ;
        RECT 2175.500 435.190 2175.640 482.810 ;
        RECT 2174.060 434.870 2174.320 435.190 ;
        RECT 2175.440 434.870 2175.700 435.190 ;
        RECT 2174.120 400.850 2174.260 434.870 ;
        RECT 2174.060 400.530 2174.320 400.850 ;
        RECT 15.280 399.850 15.540 400.170 ;
        RECT 15.340 394.925 15.480 399.850 ;
        RECT 15.270 394.555 15.550 394.925 ;
      LAYER via2 ;
        RECT 2173.590 961.720 2173.870 962.000 ;
        RECT 2174.050 772.680 2174.330 772.960 ;
        RECT 2174.970 772.680 2175.250 772.960 ;
        RECT 15.270 394.600 15.550 394.880 ;
      LAYER met3 ;
        RECT 2166.000 964.520 2170.000 965.120 ;
        RECT 2169.670 962.010 2169.970 964.520 ;
        RECT 2173.565 962.010 2173.895 962.025 ;
        RECT 2169.670 961.710 2173.895 962.010 ;
        RECT 2173.565 961.695 2173.895 961.710 ;
        RECT 2174.025 772.970 2174.355 772.985 ;
        RECT 2174.945 772.970 2175.275 772.985 ;
        RECT 2174.025 772.670 2175.275 772.970 ;
        RECT 2174.025 772.655 2174.355 772.670 ;
        RECT 2174.945 772.655 2175.275 772.670 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 15.245 394.890 15.575 394.905 ;
        RECT -4.800 394.590 15.575 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 15.245 394.575 15.575 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 2182.770 179.420 2183.090 179.480 ;
        RECT 17.090 179.280 2087.320 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 2087.180 179.080 2087.320 179.280 ;
        RECT 2110.180 179.280 2183.090 179.420 ;
        RECT 2110.180 179.080 2110.320 179.280 ;
        RECT 2182.770 179.220 2183.090 179.280 ;
        RECT 2087.180 178.940 2110.320 179.080 ;
      LAYER via ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 2182.800 179.220 2183.060 179.480 ;
      LAYER met2 ;
        RECT 2182.790 973.235 2183.070 973.605 ;
        RECT 2182.860 179.510 2183.000 973.235 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 2182.800 179.190 2183.060 179.510 ;
      LAYER via2 ;
        RECT 2182.790 973.280 2183.070 973.560 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 2166.000 974.040 2170.000 974.640 ;
        RECT 2169.670 973.570 2169.970 974.040 ;
        RECT 2182.765 973.570 2183.095 973.585 ;
        RECT 2169.670 973.270 2183.095 973.570 ;
        RECT 2182.765 973.255 2183.095 973.270 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2184.610 672.760 2184.930 672.820 ;
        RECT 2903.590 672.760 2903.910 672.820 ;
        RECT 2184.610 672.620 2903.910 672.760 ;
        RECT 2184.610 672.560 2184.930 672.620 ;
        RECT 2903.590 672.560 2903.910 672.620 ;
      LAYER via ;
        RECT 2184.640 672.560 2184.900 672.820 ;
        RECT 2903.620 672.560 2903.880 672.820 ;
      LAYER met2 ;
        RECT 2903.610 791.675 2903.890 792.045 ;
        RECT 2903.680 672.850 2903.820 791.675 ;
        RECT 2184.640 672.530 2184.900 672.850 ;
        RECT 2903.620 672.530 2903.880 672.850 ;
        RECT 2184.700 634.285 2184.840 672.530 ;
        RECT 2184.630 633.915 2184.910 634.285 ;
      LAYER via2 ;
        RECT 2903.610 791.720 2903.890 792.000 ;
        RECT 2184.630 633.960 2184.910 634.240 ;
      LAYER met3 ;
        RECT 2903.585 792.010 2903.915 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2903.585 791.710 2924.800 792.010 ;
        RECT 2903.585 791.695 2903.915 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2166.000 634.720 2170.000 635.320 ;
        RECT 2169.670 634.250 2169.970 634.720 ;
        RECT 2184.605 634.250 2184.935 634.265 ;
        RECT 2169.670 633.950 2184.935 634.250 ;
        RECT 2184.605 633.935 2184.935 633.950 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.470 648.620 2180.790 648.680 ;
        RECT 2899.910 648.620 2900.230 648.680 ;
        RECT 2180.470 648.480 2900.230 648.620 ;
        RECT 2180.470 648.420 2180.790 648.480 ;
        RECT 2899.910 648.420 2900.230 648.480 ;
      LAYER via ;
        RECT 2180.500 648.420 2180.760 648.680 ;
        RECT 2899.940 648.420 2900.200 648.680 ;
      LAYER met2 ;
        RECT 2899.930 1026.275 2900.210 1026.645 ;
        RECT 2900.000 648.710 2900.140 1026.275 ;
        RECT 2180.500 648.390 2180.760 648.710 ;
        RECT 2899.940 648.390 2900.200 648.710 ;
        RECT 2180.560 646.525 2180.700 648.390 ;
        RECT 2180.490 646.155 2180.770 646.525 ;
      LAYER via2 ;
        RECT 2899.930 1026.320 2900.210 1026.600 ;
        RECT 2180.490 646.200 2180.770 646.480 ;
      LAYER met3 ;
        RECT 2899.905 1026.610 2900.235 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2899.905 1026.310 2924.800 1026.610 ;
        RECT 2899.905 1026.295 2900.235 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2180.465 646.490 2180.795 646.505 ;
        RECT 2169.670 646.190 2180.795 646.490 ;
        RECT 2169.670 644.840 2169.970 646.190 ;
        RECT 2180.465 646.175 2180.795 646.190 ;
        RECT 2166.000 644.240 2170.000 644.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.470 655.420 2180.790 655.480 ;
        RECT 2900.370 655.420 2900.690 655.480 ;
        RECT 2180.470 655.280 2900.690 655.420 ;
        RECT 2180.470 655.220 2180.790 655.280 ;
        RECT 2900.370 655.220 2900.690 655.280 ;
      LAYER via ;
        RECT 2180.500 655.220 2180.760 655.480 ;
        RECT 2900.400 655.220 2900.660 655.480 ;
      LAYER met2 ;
        RECT 2900.390 1260.875 2900.670 1261.245 ;
        RECT 2900.460 655.510 2900.600 1260.875 ;
        RECT 2180.500 655.365 2180.760 655.510 ;
        RECT 2180.490 654.995 2180.770 655.365 ;
        RECT 2900.400 655.190 2900.660 655.510 ;
      LAYER via2 ;
        RECT 2900.390 1260.920 2900.670 1261.200 ;
        RECT 2180.490 655.040 2180.770 655.320 ;
      LAYER met3 ;
        RECT 2900.365 1261.210 2900.695 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.365 1260.910 2924.800 1261.210 ;
        RECT 2900.365 1260.895 2900.695 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2180.465 655.330 2180.795 655.345 ;
        RECT 2169.670 655.040 2180.795 655.330 ;
        RECT 2166.000 655.030 2180.795 655.040 ;
        RECT 2166.000 654.440 2170.000 655.030 ;
        RECT 2180.465 655.015 2180.795 655.030 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.470 669.360 2180.790 669.420 ;
        RECT 2904.510 669.360 2904.830 669.420 ;
        RECT 2180.470 669.220 2904.830 669.360 ;
        RECT 2180.470 669.160 2180.790 669.220 ;
        RECT 2904.510 669.160 2904.830 669.220 ;
      LAYER via ;
        RECT 2180.500 669.160 2180.760 669.420 ;
        RECT 2904.540 669.160 2904.800 669.420 ;
      LAYER met2 ;
        RECT 2904.530 1495.475 2904.810 1495.845 ;
        RECT 2904.600 669.450 2904.740 1495.475 ;
        RECT 2180.500 669.130 2180.760 669.450 ;
        RECT 2904.540 669.130 2904.800 669.450 ;
        RECT 2180.560 666.925 2180.700 669.130 ;
        RECT 2180.490 666.555 2180.770 666.925 ;
      LAYER via2 ;
        RECT 2904.530 1495.520 2904.810 1495.800 ;
        RECT 2180.490 666.600 2180.770 666.880 ;
      LAYER met3 ;
        RECT 2904.505 1495.810 2904.835 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2904.505 1495.510 2924.800 1495.810 ;
        RECT 2904.505 1495.495 2904.835 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2180.465 666.890 2180.795 666.905 ;
        RECT 2169.670 666.590 2180.795 666.890 ;
        RECT 2169.670 665.240 2169.970 666.590 ;
        RECT 2180.465 666.575 2180.795 666.590 ;
        RECT 2166.000 664.640 2170.000 665.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.470 676.160 2180.790 676.220 ;
        RECT 2903.130 676.160 2903.450 676.220 ;
        RECT 2180.470 676.020 2903.450 676.160 ;
        RECT 2180.470 675.960 2180.790 676.020 ;
        RECT 2903.130 675.960 2903.450 676.020 ;
      LAYER via ;
        RECT 2180.500 675.960 2180.760 676.220 ;
        RECT 2903.160 675.960 2903.420 676.220 ;
      LAYER met2 ;
        RECT 2903.150 1730.075 2903.430 1730.445 ;
        RECT 2903.220 676.250 2903.360 1730.075 ;
        RECT 2180.500 675.930 2180.760 676.250 ;
        RECT 2903.160 675.930 2903.420 676.250 ;
        RECT 2180.560 675.085 2180.700 675.930 ;
        RECT 2180.490 674.715 2180.770 675.085 ;
      LAYER via2 ;
        RECT 2903.150 1730.120 2903.430 1730.400 ;
        RECT 2180.490 674.760 2180.770 675.040 ;
      LAYER met3 ;
        RECT 2903.125 1730.410 2903.455 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2903.125 1730.110 2924.800 1730.410 ;
        RECT 2903.125 1730.095 2903.455 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2180.465 675.050 2180.795 675.065 ;
        RECT 2169.670 674.760 2180.795 675.050 ;
        RECT 2166.000 674.750 2180.795 674.760 ;
        RECT 2166.000 674.160 2170.000 674.750 ;
        RECT 2180.465 674.735 2180.795 674.750 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.470 689.760 2180.790 689.820 ;
        RECT 2902.670 689.760 2902.990 689.820 ;
        RECT 2180.470 689.620 2902.990 689.760 ;
        RECT 2180.470 689.560 2180.790 689.620 ;
        RECT 2902.670 689.560 2902.990 689.620 ;
      LAYER via ;
        RECT 2180.500 689.560 2180.760 689.820 ;
        RECT 2902.700 689.560 2902.960 689.820 ;
      LAYER met2 ;
        RECT 2902.690 1964.675 2902.970 1965.045 ;
        RECT 2902.760 689.850 2902.900 1964.675 ;
        RECT 2180.500 689.530 2180.760 689.850 ;
        RECT 2902.700 689.530 2902.960 689.850 ;
        RECT 2180.560 687.325 2180.700 689.530 ;
        RECT 2180.490 686.955 2180.770 687.325 ;
      LAYER via2 ;
        RECT 2902.690 1964.720 2902.970 1965.000 ;
        RECT 2180.490 687.000 2180.770 687.280 ;
      LAYER met3 ;
        RECT 2902.665 1965.010 2902.995 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2902.665 1964.710 2924.800 1965.010 ;
        RECT 2902.665 1964.695 2902.995 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2180.465 687.290 2180.795 687.305 ;
        RECT 2169.670 686.990 2180.795 687.290 ;
        RECT 2169.670 684.960 2169.970 686.990 ;
        RECT 2180.465 686.975 2180.795 686.990 ;
        RECT 2166.000 684.360 2170.000 684.960 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.470 696.900 2180.790 696.960 ;
        RECT 2902.210 696.900 2902.530 696.960 ;
        RECT 2180.470 696.760 2902.530 696.900 ;
        RECT 2180.470 696.700 2180.790 696.760 ;
        RECT 2902.210 696.700 2902.530 696.760 ;
      LAYER via ;
        RECT 2180.500 696.700 2180.760 696.960 ;
        RECT 2902.240 696.700 2902.500 696.960 ;
      LAYER met2 ;
        RECT 2902.230 2199.275 2902.510 2199.645 ;
        RECT 2902.300 696.990 2902.440 2199.275 ;
        RECT 2180.500 696.670 2180.760 696.990 ;
        RECT 2902.240 696.670 2902.500 696.990 ;
        RECT 2180.560 696.165 2180.700 696.670 ;
        RECT 2180.490 695.795 2180.770 696.165 ;
      LAYER via2 ;
        RECT 2902.230 2199.320 2902.510 2199.600 ;
        RECT 2180.490 695.840 2180.770 696.120 ;
      LAYER met3 ;
        RECT 2902.205 2199.610 2902.535 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2902.205 2199.310 2924.800 2199.610 ;
        RECT 2902.205 2199.295 2902.535 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2180.465 696.130 2180.795 696.145 ;
        RECT 2169.670 695.830 2180.795 696.130 ;
        RECT 2169.670 695.160 2169.970 695.830 ;
        RECT 2180.465 695.815 2180.795 695.830 ;
        RECT 2166.000 694.560 2170.000 695.160 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.070 206.960 667.390 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 667.070 206.820 2901.150 206.960 ;
        RECT 667.070 206.760 667.390 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 667.100 206.760 667.360 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 667.090 793.715 667.370 794.085 ;
        RECT 667.160 207.050 667.300 793.715 ;
        RECT 667.100 206.730 667.360 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 667.090 793.760 667.370 794.040 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 667.065 794.050 667.395 794.065 ;
        RECT 670.000 794.050 674.000 794.440 ;
        RECT 667.065 793.840 674.000 794.050 ;
        RECT 667.065 793.750 670.220 793.840 ;
        RECT 667.065 793.735 667.395 793.750 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 653.270 2501.280 653.590 2501.340 ;
        RECT 2902.670 2501.280 2902.990 2501.340 ;
        RECT 653.270 2501.140 2902.990 2501.280 ;
        RECT 653.270 2501.080 653.590 2501.140 ;
        RECT 2902.670 2501.080 2902.990 2501.140 ;
      LAYER via ;
        RECT 653.300 2501.080 653.560 2501.340 ;
        RECT 2902.700 2501.080 2902.960 2501.340 ;
      LAYER met2 ;
        RECT 2902.690 2551.515 2902.970 2551.885 ;
        RECT 2902.760 2501.370 2902.900 2551.515 ;
        RECT 653.300 2501.050 653.560 2501.370 ;
        RECT 2902.700 2501.050 2902.960 2501.370 ;
        RECT 653.360 845.085 653.500 2501.050 ;
        RECT 653.290 844.715 653.570 845.085 ;
      LAYER via2 ;
        RECT 2902.690 2551.560 2902.970 2551.840 ;
        RECT 653.290 844.760 653.570 845.040 ;
      LAYER met3 ;
        RECT 2902.665 2551.850 2902.995 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2902.665 2551.550 2924.800 2551.850 ;
        RECT 2902.665 2551.535 2902.995 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 653.265 845.050 653.595 845.065 ;
        RECT 670.000 845.050 674.000 845.440 ;
        RECT 653.265 844.840 674.000 845.050 ;
        RECT 653.265 844.750 670.220 844.840 ;
        RECT 653.265 844.735 653.595 844.750 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 652.810 2501.620 653.130 2501.680 ;
        RECT 2902.210 2501.620 2902.530 2501.680 ;
        RECT 652.810 2501.480 2902.530 2501.620 ;
        RECT 652.810 2501.420 653.130 2501.480 ;
        RECT 2902.210 2501.420 2902.530 2501.480 ;
      LAYER via ;
        RECT 652.840 2501.420 653.100 2501.680 ;
        RECT 2902.240 2501.420 2902.500 2501.680 ;
      LAYER met2 ;
        RECT 2902.230 2786.115 2902.510 2786.485 ;
        RECT 2902.300 2501.710 2902.440 2786.115 ;
        RECT 652.840 2501.390 653.100 2501.710 ;
        RECT 2902.240 2501.390 2902.500 2501.710 ;
        RECT 652.900 849.845 653.040 2501.390 ;
        RECT 652.830 849.475 653.110 849.845 ;
      LAYER via2 ;
        RECT 2902.230 2786.160 2902.510 2786.440 ;
        RECT 652.830 849.520 653.110 849.800 ;
      LAYER met3 ;
        RECT 2902.205 2786.450 2902.535 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2902.205 2786.150 2924.800 2786.450 ;
        RECT 2902.205 2786.135 2902.535 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 652.805 849.810 653.135 849.825 ;
        RECT 670.000 849.810 674.000 850.200 ;
        RECT 652.805 849.600 674.000 849.810 ;
        RECT 652.805 849.510 670.220 849.600 ;
        RECT 652.805 849.495 653.135 849.510 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 659.250 3015.700 659.570 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 659.250 3015.560 2901.150 3015.700 ;
        RECT 659.250 3015.500 659.570 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 659.280 3015.500 659.540 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 659.280 3015.470 659.540 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 659.340 855.285 659.480 3015.470 ;
        RECT 659.270 854.915 659.550 855.285 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 659.270 854.960 659.550 855.240 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 659.245 855.250 659.575 855.265 ;
        RECT 670.000 855.250 674.000 855.640 ;
        RECT 659.245 855.040 674.000 855.250 ;
        RECT 659.245 854.950 670.220 855.040 ;
        RECT 659.245 854.935 659.575 854.950 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 655.110 3250.300 655.430 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 655.110 3250.160 2901.150 3250.300 ;
        RECT 655.110 3250.100 655.430 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 655.140 3250.100 655.400 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 655.140 3250.070 655.400 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 655.200 860.045 655.340 3250.070 ;
        RECT 655.130 859.675 655.410 860.045 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 655.130 859.720 655.410 860.000 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 655.105 860.010 655.435 860.025 ;
        RECT 670.000 860.010 674.000 860.400 ;
        RECT 655.105 859.800 674.000 860.010 ;
        RECT 655.105 859.710 670.220 859.800 ;
        RECT 655.105 859.695 655.435 859.710 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 647.750 3484.900 648.070 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 647.750 3484.760 2901.150 3484.900 ;
        RECT 647.750 3484.700 648.070 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 647.750 869.280 648.070 869.340 ;
        RECT 656.490 869.280 656.810 869.340 ;
        RECT 647.750 869.140 656.810 869.280 ;
        RECT 647.750 869.080 648.070 869.140 ;
        RECT 656.490 869.080 656.810 869.140 ;
      LAYER via ;
        RECT 647.780 3484.700 648.040 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 647.780 869.080 648.040 869.340 ;
        RECT 656.520 869.080 656.780 869.340 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 647.780 3484.670 648.040 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 647.840 869.370 647.980 3484.670 ;
        RECT 647.780 869.050 648.040 869.370 ;
        RECT 656.520 869.050 656.780 869.370 ;
        RECT 656.580 865.485 656.720 869.050 ;
        RECT 656.510 865.115 656.790 865.485 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 656.510 865.160 656.790 865.440 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 656.485 865.450 656.815 865.465 ;
        RECT 670.000 865.450 674.000 865.840 ;
        RECT 656.485 865.240 674.000 865.450 ;
        RECT 656.485 865.150 670.220 865.240 ;
        RECT 656.485 865.135 656.815 865.150 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.990 3501.900 668.310 3501.960 ;
        RECT 2635.870 3501.900 2636.190 3501.960 ;
        RECT 667.990 3501.760 2636.190 3501.900 ;
        RECT 667.990 3501.700 668.310 3501.760 ;
        RECT 2635.870 3501.700 2636.190 3501.760 ;
      LAYER via ;
        RECT 668.020 3501.700 668.280 3501.960 ;
        RECT 2635.900 3501.700 2636.160 3501.960 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.990 2636.100 3517.600 ;
        RECT 668.020 3501.670 668.280 3501.990 ;
        RECT 2635.900 3501.670 2636.160 3501.990 ;
        RECT 668.080 870.245 668.220 3501.670 ;
        RECT 668.010 869.875 668.290 870.245 ;
      LAYER via2 ;
        RECT 668.010 869.920 668.290 870.200 ;
      LAYER met3 ;
        RECT 667.985 870.210 668.315 870.225 ;
        RECT 670.000 870.210 674.000 870.600 ;
        RECT 667.985 870.000 674.000 870.210 ;
        RECT 667.985 869.910 670.220 870.000 ;
        RECT 667.985 869.895 668.315 869.910 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.930 3503.260 663.250 3503.320 ;
        RECT 2311.570 3503.260 2311.890 3503.320 ;
        RECT 662.930 3503.120 2311.890 3503.260 ;
        RECT 662.930 3503.060 663.250 3503.120 ;
        RECT 2311.570 3503.060 2311.890 3503.120 ;
      LAYER via ;
        RECT 662.960 3503.060 663.220 3503.320 ;
        RECT 2311.600 3503.060 2311.860 3503.320 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3503.350 2311.800 3517.600 ;
        RECT 662.960 3503.030 663.220 3503.350 ;
        RECT 2311.600 3503.030 2311.860 3503.350 ;
        RECT 663.020 875.005 663.160 3503.030 ;
        RECT 662.950 874.635 663.230 875.005 ;
      LAYER via2 ;
        RECT 662.950 874.680 663.230 874.960 ;
      LAYER met3 ;
        RECT 662.925 874.970 663.255 874.985 ;
        RECT 670.000 874.970 674.000 875.360 ;
        RECT 662.925 874.760 674.000 874.970 ;
        RECT 662.925 874.670 670.220 874.760 ;
        RECT 662.925 874.655 663.255 874.670 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.530 3503.940 667.850 3504.000 ;
        RECT 1987.270 3503.940 1987.590 3504.000 ;
        RECT 667.530 3503.800 1987.590 3503.940 ;
        RECT 667.530 3503.740 667.850 3503.800 ;
        RECT 1987.270 3503.740 1987.590 3503.800 ;
      LAYER via ;
        RECT 667.560 3503.740 667.820 3504.000 ;
        RECT 1987.300 3503.740 1987.560 3504.000 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3504.030 1987.500 3517.600 ;
        RECT 667.560 3503.710 667.820 3504.030 ;
        RECT 1987.300 3503.710 1987.560 3504.030 ;
        RECT 667.620 880.445 667.760 3503.710 ;
        RECT 667.550 880.075 667.830 880.445 ;
      LAYER via2 ;
        RECT 667.550 880.120 667.830 880.400 ;
      LAYER met3 ;
        RECT 667.525 880.410 667.855 880.425 ;
        RECT 670.000 880.410 674.000 880.800 ;
        RECT 667.525 880.200 674.000 880.410 ;
        RECT 667.525 880.110 670.220 880.200 ;
        RECT 667.525 880.095 667.855 880.110 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.070 3501.220 667.390 3501.280 ;
        RECT 1662.510 3501.220 1662.830 3501.280 ;
        RECT 667.070 3501.080 1662.830 3501.220 ;
        RECT 667.070 3501.020 667.390 3501.080 ;
        RECT 1662.510 3501.020 1662.830 3501.080 ;
      LAYER via ;
        RECT 667.100 3501.020 667.360 3501.280 ;
        RECT 1662.540 3501.020 1662.800 3501.280 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3501.310 1662.740 3517.600 ;
        RECT 667.100 3500.990 667.360 3501.310 ;
        RECT 1662.540 3500.990 1662.800 3501.310 ;
        RECT 667.160 885.205 667.300 3500.990 ;
        RECT 667.090 884.835 667.370 885.205 ;
      LAYER via2 ;
        RECT 667.090 884.880 667.370 885.160 ;
      LAYER met3 ;
        RECT 667.065 885.170 667.395 885.185 ;
        RECT 670.000 885.170 674.000 885.560 ;
        RECT 667.065 884.960 674.000 885.170 ;
        RECT 667.065 884.870 670.220 884.960 ;
        RECT 667.065 884.855 667.395 884.870 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1331.770 3487.960 1332.090 3488.020 ;
        RECT 1338.210 3487.960 1338.530 3488.020 ;
        RECT 1331.770 3487.820 1338.530 3487.960 ;
        RECT 1331.770 3487.760 1332.090 3487.820 ;
        RECT 1338.210 3487.760 1338.530 3487.820 ;
        RECT 662.470 1005.960 662.790 1006.020 ;
        RECT 1331.770 1005.960 1332.090 1006.020 ;
        RECT 662.470 1005.820 1332.090 1005.960 ;
        RECT 662.470 1005.760 662.790 1005.820 ;
        RECT 1331.770 1005.760 1332.090 1005.820 ;
        RECT 658.330 999.500 658.650 999.560 ;
        RECT 662.470 999.500 662.790 999.560 ;
        RECT 658.330 999.360 662.790 999.500 ;
        RECT 658.330 999.300 658.650 999.360 ;
        RECT 662.470 999.300 662.790 999.360 ;
        RECT 658.330 979.780 658.650 979.840 ;
        RECT 662.470 979.780 662.790 979.840 ;
        RECT 658.330 979.640 662.790 979.780 ;
        RECT 658.330 979.580 658.650 979.640 ;
        RECT 662.470 979.580 662.790 979.640 ;
      LAYER via ;
        RECT 1331.800 3487.760 1332.060 3488.020 ;
        RECT 1338.240 3487.760 1338.500 3488.020 ;
        RECT 662.500 1005.760 662.760 1006.020 ;
        RECT 1331.800 1005.760 1332.060 1006.020 ;
        RECT 658.360 999.300 658.620 999.560 ;
        RECT 662.500 999.300 662.760 999.560 ;
        RECT 658.360 979.580 658.620 979.840 ;
        RECT 662.500 979.580 662.760 979.840 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3488.050 1338.440 3517.600 ;
        RECT 1331.800 3487.730 1332.060 3488.050 ;
        RECT 1338.240 3487.730 1338.500 3488.050 ;
        RECT 1331.860 1006.050 1332.000 3487.730 ;
        RECT 662.500 1005.730 662.760 1006.050 ;
        RECT 1331.800 1005.730 1332.060 1006.050 ;
        RECT 662.560 999.590 662.700 1005.730 ;
        RECT 658.360 999.270 658.620 999.590 ;
        RECT 662.500 999.270 662.760 999.590 ;
        RECT 658.420 979.870 658.560 999.270 ;
        RECT 658.360 979.550 658.620 979.870 ;
        RECT 662.500 979.550 662.760 979.870 ;
        RECT 662.560 890.645 662.700 979.550 ;
        RECT 662.490 890.275 662.770 890.645 ;
      LAYER via2 ;
        RECT 662.490 890.320 662.770 890.600 ;
      LAYER met3 ;
        RECT 662.465 890.610 662.795 890.625 ;
        RECT 670.000 890.610 674.000 891.000 ;
        RECT 662.465 890.400 674.000 890.610 ;
        RECT 662.465 890.310 670.220 890.400 ;
        RECT 662.465 890.295 662.795 890.310 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.990 441.560 668.310 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 667.990 441.420 2901.150 441.560 ;
        RECT 667.990 441.360 668.310 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 668.020 441.360 668.280 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 668.010 799.155 668.290 799.525 ;
        RECT 668.080 441.650 668.220 799.155 ;
        RECT 668.020 441.330 668.280 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 668.010 799.200 668.290 799.480 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 667.985 799.490 668.315 799.505 ;
        RECT 670.000 799.490 674.000 799.880 ;
        RECT 667.985 799.280 674.000 799.490 ;
        RECT 667.985 799.190 670.220 799.280 ;
        RECT 667.985 799.175 668.315 799.190 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 666.610 3504.960 666.930 3505.020 ;
        RECT 1013.910 3504.960 1014.230 3505.020 ;
        RECT 666.610 3504.820 1014.230 3504.960 ;
        RECT 666.610 3504.760 666.930 3504.820 ;
        RECT 1013.910 3504.760 1014.230 3504.820 ;
      LAYER via ;
        RECT 666.640 3504.760 666.900 3505.020 ;
        RECT 1013.940 3504.760 1014.200 3505.020 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3505.050 1014.140 3517.600 ;
        RECT 666.640 3504.730 666.900 3505.050 ;
        RECT 1013.940 3504.730 1014.200 3505.050 ;
        RECT 666.700 895.405 666.840 3504.730 ;
        RECT 666.630 895.035 666.910 895.405 ;
      LAYER via2 ;
        RECT 666.630 895.080 666.910 895.360 ;
      LAYER met3 ;
        RECT 666.605 895.370 666.935 895.385 ;
        RECT 670.000 895.370 674.000 895.760 ;
        RECT 666.605 895.160 674.000 895.370 ;
        RECT 666.605 895.070 670.220 895.160 ;
        RECT 666.605 895.055 666.935 895.070 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 666.150 3498.500 666.470 3498.560 ;
        RECT 689.150 3498.500 689.470 3498.560 ;
        RECT 666.150 3498.360 689.470 3498.500 ;
        RECT 666.150 3498.300 666.470 3498.360 ;
        RECT 689.150 3498.300 689.470 3498.360 ;
      LAYER via ;
        RECT 666.180 3498.300 666.440 3498.560 ;
        RECT 689.180 3498.300 689.440 3498.560 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3498.590 689.380 3517.600 ;
        RECT 666.180 3498.270 666.440 3498.590 ;
        RECT 689.180 3498.270 689.440 3498.590 ;
        RECT 666.240 900.845 666.380 3498.270 ;
        RECT 666.170 900.475 666.450 900.845 ;
      LAYER via2 ;
        RECT 666.170 900.520 666.450 900.800 ;
      LAYER met3 ;
        RECT 666.145 900.810 666.475 900.825 ;
        RECT 670.000 900.810 674.000 901.200 ;
        RECT 666.145 900.600 674.000 900.810 ;
        RECT 666.145 900.510 670.220 900.600 ;
        RECT 666.145 900.495 666.475 900.510 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 362.090 3498.500 362.410 3498.560 ;
        RECT 364.850 3498.500 365.170 3498.560 ;
        RECT 362.090 3498.360 365.170 3498.500 ;
        RECT 362.090 3498.300 362.410 3498.360 ;
        RECT 364.850 3498.300 365.170 3498.360 ;
        RECT 362.090 910.760 362.410 910.820 ;
        RECT 656.030 910.760 656.350 910.820 ;
        RECT 362.090 910.620 656.350 910.760 ;
        RECT 362.090 910.560 362.410 910.620 ;
        RECT 656.030 910.560 656.350 910.620 ;
      LAYER via ;
        RECT 362.120 3498.300 362.380 3498.560 ;
        RECT 364.880 3498.300 365.140 3498.560 ;
        RECT 362.120 910.560 362.380 910.820 ;
        RECT 656.060 910.560 656.320 910.820 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3498.590 365.080 3517.600 ;
        RECT 362.120 3498.270 362.380 3498.590 ;
        RECT 364.880 3498.270 365.140 3498.590 ;
        RECT 362.180 910.850 362.320 3498.270 ;
        RECT 362.120 910.530 362.380 910.850 ;
        RECT 656.060 910.530 656.320 910.850 ;
        RECT 656.120 905.605 656.260 910.530 ;
        RECT 656.050 905.235 656.330 905.605 ;
      LAYER via2 ;
        RECT 656.050 905.280 656.330 905.560 ;
      LAYER met3 ;
        RECT 656.025 905.570 656.355 905.585 ;
        RECT 670.000 905.570 674.000 905.960 ;
        RECT 656.025 905.360 674.000 905.570 ;
        RECT 656.025 905.270 670.220 905.360 ;
        RECT 656.025 905.255 656.355 905.270 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 39.630 3477.420 39.950 3477.480 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 39.630 3477.280 41.330 3477.420 ;
        RECT 39.630 3477.220 39.950 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 39.630 3429.480 39.950 3429.540 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 39.630 3429.340 40.870 3429.480 ;
        RECT 39.630 3429.280 39.950 3429.340 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3270.700 40.410 3270.760 ;
        RECT 41.010 3270.700 41.330 3270.760 ;
        RECT 40.090 3270.560 41.330 3270.700 ;
        RECT 40.090 3270.500 40.410 3270.560 ;
        RECT 41.010 3270.500 41.330 3270.560 ;
        RECT 40.090 3174.140 40.410 3174.200 ;
        RECT 41.010 3174.140 41.330 3174.200 ;
        RECT 40.090 3174.000 41.330 3174.140 ;
        RECT 40.090 3173.940 40.410 3174.000 ;
        RECT 41.010 3173.940 41.330 3174.000 ;
        RECT 40.090 3077.580 40.410 3077.640 ;
        RECT 41.010 3077.580 41.330 3077.640 ;
        RECT 40.090 3077.440 41.330 3077.580 ;
        RECT 40.090 3077.380 40.410 3077.440 ;
        RECT 41.010 3077.380 41.330 3077.440 ;
        RECT 40.090 2981.020 40.410 2981.080 ;
        RECT 41.010 2981.020 41.330 2981.080 ;
        RECT 40.090 2980.880 41.330 2981.020 ;
        RECT 40.090 2980.820 40.410 2980.880 ;
        RECT 41.010 2980.820 41.330 2980.880 ;
        RECT 38.250 2898.060 38.570 2898.120 ;
        RECT 39.630 2898.060 39.950 2898.120 ;
        RECT 38.250 2897.920 39.950 2898.060 ;
        RECT 38.250 2897.860 38.570 2897.920 ;
        RECT 39.630 2897.860 39.950 2897.920 ;
        RECT 38.250 2849.780 38.570 2849.840 ;
        RECT 39.170 2849.780 39.490 2849.840 ;
        RECT 38.250 2849.640 39.490 2849.780 ;
        RECT 38.250 2849.580 38.570 2849.640 ;
        RECT 39.170 2849.580 39.490 2849.640 ;
        RECT 39.170 2815.240 39.490 2815.500 ;
        RECT 39.260 2814.760 39.400 2815.240 ;
        RECT 39.630 2814.760 39.950 2814.820 ;
        RECT 39.260 2814.620 39.950 2814.760 ;
        RECT 39.630 2814.560 39.950 2814.620 ;
        RECT 40.090 2752.880 40.410 2752.940 ;
        RECT 40.550 2752.880 40.870 2752.940 ;
        RECT 40.090 2752.740 40.870 2752.880 ;
        RECT 40.090 2752.680 40.410 2752.740 ;
        RECT 40.550 2752.680 40.870 2752.740 ;
        RECT 40.550 2704.940 40.870 2705.000 ;
        RECT 41.010 2704.940 41.330 2705.000 ;
        RECT 40.550 2704.800 41.330 2704.940 ;
        RECT 40.550 2704.740 40.870 2704.800 ;
        RECT 41.010 2704.740 41.330 2704.800 ;
        RECT 41.010 2608.380 41.330 2608.440 ;
        RECT 41.930 2608.380 42.250 2608.440 ;
        RECT 41.010 2608.240 42.250 2608.380 ;
        RECT 41.010 2608.180 41.330 2608.240 ;
        RECT 41.930 2608.180 42.250 2608.240 ;
        RECT 41.010 2511.820 41.330 2511.880 ;
        RECT 41.930 2511.820 42.250 2511.880 ;
        RECT 41.010 2511.680 42.250 2511.820 ;
        RECT 41.010 2511.620 41.330 2511.680 ;
        RECT 41.930 2511.620 42.250 2511.680 ;
        RECT 40.550 2429.000 40.870 2429.260 ;
        RECT 40.640 2428.860 40.780 2429.000 ;
        RECT 41.010 2428.860 41.330 2428.920 ;
        RECT 40.640 2428.720 41.330 2428.860 ;
        RECT 41.010 2428.660 41.330 2428.720 ;
        RECT 39.630 2414.920 39.950 2414.980 ;
        RECT 41.010 2414.920 41.330 2414.980 ;
        RECT 39.630 2414.780 41.330 2414.920 ;
        RECT 39.630 2414.720 39.950 2414.780 ;
        RECT 41.010 2414.720 41.330 2414.780 ;
        RECT 40.550 2332.100 40.870 2332.360 ;
        RECT 40.640 2331.960 40.780 2332.100 ;
        RECT 41.010 2331.960 41.330 2332.020 ;
        RECT 40.640 2331.820 41.330 2331.960 ;
        RECT 41.010 2331.760 41.330 2331.820 ;
        RECT 39.170 2270.080 39.490 2270.140 ;
        RECT 40.090 2270.080 40.410 2270.140 ;
        RECT 39.170 2269.940 40.410 2270.080 ;
        RECT 39.170 2269.880 39.490 2269.940 ;
        RECT 40.090 2269.880 40.410 2269.940 ;
        RECT 39.170 2222.140 39.490 2222.200 ;
        RECT 39.630 2222.140 39.950 2222.200 ;
        RECT 39.170 2222.000 39.950 2222.140 ;
        RECT 39.170 2221.940 39.490 2222.000 ;
        RECT 39.630 2221.940 39.950 2222.000 ;
        RECT 40.550 2138.980 40.870 2139.240 ;
        RECT 40.640 2138.840 40.780 2138.980 ;
        RECT 41.010 2138.840 41.330 2138.900 ;
        RECT 40.640 2138.700 41.330 2138.840 ;
        RECT 41.010 2138.640 41.330 2138.700 ;
        RECT 39.630 2125.240 39.950 2125.300 ;
        RECT 41.010 2125.240 41.330 2125.300 ;
        RECT 39.630 2125.100 41.330 2125.240 ;
        RECT 39.630 2125.040 39.950 2125.100 ;
        RECT 41.010 2125.040 41.330 2125.100 ;
        RECT 39.630 2077.300 39.950 2077.360 ;
        RECT 40.550 2077.300 40.870 2077.360 ;
        RECT 39.630 2077.160 40.870 2077.300 ;
        RECT 39.630 2077.100 39.950 2077.160 ;
        RECT 40.550 2077.100 40.870 2077.160 ;
        RECT 40.550 2042.420 40.870 2042.680 ;
        RECT 40.640 2041.940 40.780 2042.420 ;
        RECT 41.010 2041.940 41.330 2042.000 ;
        RECT 40.640 2041.800 41.330 2041.940 ;
        RECT 41.010 2041.740 41.330 2041.800 ;
        RECT 41.010 2004.540 41.330 2004.600 ;
        RECT 41.930 2004.540 42.250 2004.600 ;
        RECT 41.010 2004.400 42.250 2004.540 ;
        RECT 41.010 2004.340 41.330 2004.400 ;
        RECT 41.930 2004.340 42.250 2004.400 ;
        RECT 40.090 1980.400 40.410 1980.460 ;
        RECT 41.930 1980.400 42.250 1980.460 ;
        RECT 40.090 1980.260 42.250 1980.400 ;
        RECT 40.090 1980.200 40.410 1980.260 ;
        RECT 41.930 1980.200 42.250 1980.260 ;
        RECT 40.090 1973.600 40.410 1973.660 ;
        RECT 40.550 1973.600 40.870 1973.660 ;
        RECT 40.090 1973.460 40.870 1973.600 ;
        RECT 40.090 1973.400 40.410 1973.460 ;
        RECT 40.550 1973.400 40.870 1973.460 ;
        RECT 40.550 1945.860 40.870 1946.120 ;
        RECT 40.640 1945.380 40.780 1945.860 ;
        RECT 41.010 1945.380 41.330 1945.440 ;
        RECT 40.640 1945.240 41.330 1945.380 ;
        RECT 41.010 1945.180 41.330 1945.240 ;
        RECT 41.010 1897.780 41.330 1897.840 ;
        RECT 40.180 1897.640 41.330 1897.780 ;
        RECT 40.180 1897.500 40.320 1897.640 ;
        RECT 41.010 1897.580 41.330 1897.640 ;
        RECT 40.090 1897.240 40.410 1897.500 ;
        RECT 39.170 1876.700 39.490 1876.760 ;
        RECT 40.090 1876.700 40.410 1876.760 ;
        RECT 39.170 1876.560 40.410 1876.700 ;
        RECT 39.170 1876.500 39.490 1876.560 ;
        RECT 40.090 1876.500 40.410 1876.560 ;
        RECT 39.170 1828.760 39.490 1828.820 ;
        RECT 40.550 1828.760 40.870 1828.820 ;
        RECT 39.170 1828.620 40.870 1828.760 ;
        RECT 39.170 1828.560 39.490 1828.620 ;
        RECT 40.550 1828.560 40.870 1828.620 ;
        RECT 40.550 1801.020 40.870 1801.280 ;
        RECT 40.640 1800.880 40.780 1801.020 ;
        RECT 41.010 1800.880 41.330 1800.940 ;
        RECT 40.640 1800.740 41.330 1800.880 ;
        RECT 41.010 1800.680 41.330 1800.740 ;
        RECT 41.010 1773.340 41.330 1773.400 ;
        RECT 41.930 1773.340 42.250 1773.400 ;
        RECT 41.010 1773.200 42.250 1773.340 ;
        RECT 41.010 1773.140 41.330 1773.200 ;
        RECT 41.930 1773.140 42.250 1773.200 ;
        RECT 41.010 1725.400 41.330 1725.460 ;
        RECT 41.930 1725.400 42.250 1725.460 ;
        RECT 41.010 1725.260 42.250 1725.400 ;
        RECT 41.010 1725.200 41.330 1725.260 ;
        RECT 41.930 1725.200 42.250 1725.260 ;
        RECT 40.090 1628.500 40.410 1628.560 ;
        RECT 41.010 1628.500 41.330 1628.560 ;
        RECT 40.090 1628.360 41.330 1628.500 ;
        RECT 40.090 1628.300 40.410 1628.360 ;
        RECT 41.010 1628.300 41.330 1628.360 ;
        RECT 40.090 1531.940 40.410 1532.000 ;
        RECT 41.010 1531.940 41.330 1532.000 ;
        RECT 40.090 1531.800 41.330 1531.940 ;
        RECT 40.090 1531.740 40.410 1531.800 ;
        RECT 41.010 1531.740 41.330 1531.800 ;
        RECT 40.090 1435.380 40.410 1435.440 ;
        RECT 41.010 1435.380 41.330 1435.440 ;
        RECT 40.090 1435.240 41.330 1435.380 ;
        RECT 40.090 1435.180 40.410 1435.240 ;
        RECT 41.010 1435.180 41.330 1435.240 ;
        RECT 40.090 1338.820 40.410 1338.880 ;
        RECT 41.010 1338.820 41.330 1338.880 ;
        RECT 40.090 1338.680 41.330 1338.820 ;
        RECT 40.090 1338.620 40.410 1338.680 ;
        RECT 41.010 1338.620 41.330 1338.680 ;
        RECT 38.710 1255.860 39.030 1255.920 ;
        RECT 39.630 1255.860 39.950 1255.920 ;
        RECT 38.710 1255.720 39.950 1255.860 ;
        RECT 38.710 1255.660 39.030 1255.720 ;
        RECT 39.630 1255.660 39.950 1255.720 ;
        RECT 38.710 1207.580 39.030 1207.640 ;
        RECT 40.090 1207.580 40.410 1207.640 ;
        RECT 38.710 1207.440 40.410 1207.580 ;
        RECT 38.710 1207.380 39.030 1207.440 ;
        RECT 40.090 1207.380 40.410 1207.440 ;
        RECT 40.090 1173.580 40.410 1173.640 ;
        RECT 39.720 1173.440 40.410 1173.580 ;
        RECT 39.720 1172.960 39.860 1173.440 ;
        RECT 40.090 1173.380 40.410 1173.440 ;
        RECT 39.630 1172.700 39.950 1172.960 ;
        RECT 38.710 1158.960 39.030 1159.020 ;
        RECT 39.630 1158.960 39.950 1159.020 ;
        RECT 38.710 1158.820 39.950 1158.960 ;
        RECT 38.710 1158.760 39.030 1158.820 ;
        RECT 39.630 1158.760 39.950 1158.820 ;
        RECT 38.710 1111.020 39.030 1111.080 ;
        RECT 40.090 1111.020 40.410 1111.080 ;
        RECT 38.710 1110.880 40.410 1111.020 ;
        RECT 38.710 1110.820 39.030 1110.880 ;
        RECT 40.090 1110.820 40.410 1110.880 ;
        RECT 40.090 1077.020 40.410 1077.080 ;
        RECT 39.720 1076.880 40.410 1077.020 ;
        RECT 39.720 1076.400 39.860 1076.880 ;
        RECT 40.090 1076.820 40.410 1076.880 ;
        RECT 39.630 1076.140 39.950 1076.400 ;
        RECT 39.170 979.780 39.490 979.840 ;
        RECT 40.550 979.780 40.870 979.840 ;
        RECT 39.170 979.640 40.870 979.780 ;
        RECT 39.170 979.580 39.490 979.640 ;
        RECT 40.550 979.580 40.870 979.640 ;
        RECT 96.300 917.080 96.900 917.220 ;
        RECT 40.090 916.540 40.410 916.600 ;
        RECT 48.370 916.540 48.690 916.600 ;
        RECT 40.090 916.400 48.690 916.540 ;
        RECT 40.090 916.340 40.410 916.400 ;
        RECT 48.370 916.340 48.690 916.400 ;
        RECT 62.170 916.540 62.490 916.600 ;
        RECT 96.300 916.540 96.440 917.080 ;
        RECT 96.760 916.880 96.900 917.080 ;
        RECT 241.570 916.880 241.890 916.940 ;
        RECT 338.170 916.880 338.490 916.940 ;
        RECT 448.110 916.880 448.430 916.940 ;
        RECT 96.760 916.740 158.540 916.880 ;
        RECT 62.170 916.400 96.440 916.540 ;
        RECT 158.400 916.540 158.540 916.740 ;
        RECT 213.140 916.740 241.890 916.880 ;
        RECT 206.610 916.540 206.930 916.600 ;
        RECT 158.400 916.400 206.930 916.540 ;
        RECT 62.170 916.340 62.490 916.400 ;
        RECT 206.610 916.340 206.930 916.400 ;
        RECT 207.070 916.540 207.390 916.600 ;
        RECT 213.140 916.540 213.280 916.740 ;
        RECT 241.570 916.680 241.890 916.740 ;
        RECT 309.740 916.740 338.490 916.880 ;
        RECT 207.070 916.400 213.280 916.540 ;
        RECT 289.410 916.540 289.730 916.600 ;
        RECT 303.210 916.540 303.530 916.600 ;
        RECT 289.410 916.400 303.530 916.540 ;
        RECT 207.070 916.340 207.390 916.400 ;
        RECT 289.410 916.340 289.730 916.400 ;
        RECT 303.210 916.340 303.530 916.400 ;
        RECT 303.670 916.540 303.990 916.600 ;
        RECT 309.740 916.540 309.880 916.740 ;
        RECT 338.170 916.680 338.490 916.740 ;
        RECT 406.340 916.740 448.430 916.880 ;
        RECT 303.670 916.400 309.880 916.540 ;
        RECT 386.010 916.540 386.330 916.600 ;
        RECT 399.810 916.540 400.130 916.600 ;
        RECT 386.010 916.400 400.130 916.540 ;
        RECT 303.670 916.340 303.990 916.400 ;
        RECT 386.010 916.340 386.330 916.400 ;
        RECT 399.810 916.340 400.130 916.400 ;
        RECT 400.270 916.540 400.590 916.600 ;
        RECT 406.340 916.540 406.480 916.740 ;
        RECT 448.110 916.680 448.430 916.740 ;
        RECT 400.270 916.400 406.480 916.540 ;
        RECT 448.570 916.540 448.890 916.600 ;
        RECT 476.170 916.540 476.490 916.600 ;
        RECT 448.570 916.400 476.490 916.540 ;
        RECT 400.270 916.340 400.590 916.400 ;
        RECT 448.570 916.340 448.890 916.400 ;
        RECT 476.170 916.340 476.490 916.400 ;
        RECT 524.010 916.540 524.330 916.600 ;
        RECT 572.770 916.540 573.090 916.600 ;
        RECT 524.010 916.400 573.090 916.540 ;
        RECT 524.010 916.340 524.330 916.400 ;
        RECT 572.770 916.340 573.090 916.400 ;
        RECT 620.610 916.200 620.930 916.260 ;
        RECT 620.610 916.060 641.540 916.200 ;
        RECT 620.610 916.000 620.930 916.060 ;
        RECT 641.400 915.860 641.540 916.060 ;
        RECT 641.400 915.720 656.260 915.860 ;
        RECT 572.770 915.520 573.090 915.580 ;
        RECT 620.610 915.520 620.930 915.580 ;
        RECT 572.770 915.380 620.930 915.520 ;
        RECT 572.770 915.320 573.090 915.380 ;
        RECT 620.610 915.320 620.930 915.380 ;
        RECT 656.120 915.240 656.260 915.720 ;
        RECT 656.030 914.980 656.350 915.240 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 39.660 3477.220 39.920 3477.480 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 39.660 3429.280 39.920 3429.540 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3270.500 40.380 3270.760 ;
        RECT 41.040 3270.500 41.300 3270.760 ;
        RECT 40.120 3173.940 40.380 3174.200 ;
        RECT 41.040 3173.940 41.300 3174.200 ;
        RECT 40.120 3077.380 40.380 3077.640 ;
        RECT 41.040 3077.380 41.300 3077.640 ;
        RECT 40.120 2980.820 40.380 2981.080 ;
        RECT 41.040 2980.820 41.300 2981.080 ;
        RECT 38.280 2897.860 38.540 2898.120 ;
        RECT 39.660 2897.860 39.920 2898.120 ;
        RECT 38.280 2849.580 38.540 2849.840 ;
        RECT 39.200 2849.580 39.460 2849.840 ;
        RECT 39.200 2815.240 39.460 2815.500 ;
        RECT 39.660 2814.560 39.920 2814.820 ;
        RECT 40.120 2752.680 40.380 2752.940 ;
        RECT 40.580 2752.680 40.840 2752.940 ;
        RECT 40.580 2704.740 40.840 2705.000 ;
        RECT 41.040 2704.740 41.300 2705.000 ;
        RECT 41.040 2608.180 41.300 2608.440 ;
        RECT 41.960 2608.180 42.220 2608.440 ;
        RECT 41.040 2511.620 41.300 2511.880 ;
        RECT 41.960 2511.620 42.220 2511.880 ;
        RECT 40.580 2429.000 40.840 2429.260 ;
        RECT 41.040 2428.660 41.300 2428.920 ;
        RECT 39.660 2414.720 39.920 2414.980 ;
        RECT 41.040 2414.720 41.300 2414.980 ;
        RECT 40.580 2332.100 40.840 2332.360 ;
        RECT 41.040 2331.760 41.300 2332.020 ;
        RECT 39.200 2269.880 39.460 2270.140 ;
        RECT 40.120 2269.880 40.380 2270.140 ;
        RECT 39.200 2221.940 39.460 2222.200 ;
        RECT 39.660 2221.940 39.920 2222.200 ;
        RECT 40.580 2138.980 40.840 2139.240 ;
        RECT 41.040 2138.640 41.300 2138.900 ;
        RECT 39.660 2125.040 39.920 2125.300 ;
        RECT 41.040 2125.040 41.300 2125.300 ;
        RECT 39.660 2077.100 39.920 2077.360 ;
        RECT 40.580 2077.100 40.840 2077.360 ;
        RECT 40.580 2042.420 40.840 2042.680 ;
        RECT 41.040 2041.740 41.300 2042.000 ;
        RECT 41.040 2004.340 41.300 2004.600 ;
        RECT 41.960 2004.340 42.220 2004.600 ;
        RECT 40.120 1980.200 40.380 1980.460 ;
        RECT 41.960 1980.200 42.220 1980.460 ;
        RECT 40.120 1973.400 40.380 1973.660 ;
        RECT 40.580 1973.400 40.840 1973.660 ;
        RECT 40.580 1945.860 40.840 1946.120 ;
        RECT 41.040 1945.180 41.300 1945.440 ;
        RECT 41.040 1897.580 41.300 1897.840 ;
        RECT 40.120 1897.240 40.380 1897.500 ;
        RECT 39.200 1876.500 39.460 1876.760 ;
        RECT 40.120 1876.500 40.380 1876.760 ;
        RECT 39.200 1828.560 39.460 1828.820 ;
        RECT 40.580 1828.560 40.840 1828.820 ;
        RECT 40.580 1801.020 40.840 1801.280 ;
        RECT 41.040 1800.680 41.300 1800.940 ;
        RECT 41.040 1773.140 41.300 1773.400 ;
        RECT 41.960 1773.140 42.220 1773.400 ;
        RECT 41.040 1725.200 41.300 1725.460 ;
        RECT 41.960 1725.200 42.220 1725.460 ;
        RECT 40.120 1628.300 40.380 1628.560 ;
        RECT 41.040 1628.300 41.300 1628.560 ;
        RECT 40.120 1531.740 40.380 1532.000 ;
        RECT 41.040 1531.740 41.300 1532.000 ;
        RECT 40.120 1435.180 40.380 1435.440 ;
        RECT 41.040 1435.180 41.300 1435.440 ;
        RECT 40.120 1338.620 40.380 1338.880 ;
        RECT 41.040 1338.620 41.300 1338.880 ;
        RECT 38.740 1255.660 39.000 1255.920 ;
        RECT 39.660 1255.660 39.920 1255.920 ;
        RECT 38.740 1207.380 39.000 1207.640 ;
        RECT 40.120 1207.380 40.380 1207.640 ;
        RECT 40.120 1173.380 40.380 1173.640 ;
        RECT 39.660 1172.700 39.920 1172.960 ;
        RECT 38.740 1158.760 39.000 1159.020 ;
        RECT 39.660 1158.760 39.920 1159.020 ;
        RECT 38.740 1110.820 39.000 1111.080 ;
        RECT 40.120 1110.820 40.380 1111.080 ;
        RECT 40.120 1076.820 40.380 1077.080 ;
        RECT 39.660 1076.140 39.920 1076.400 ;
        RECT 39.200 979.580 39.460 979.840 ;
        RECT 40.580 979.580 40.840 979.840 ;
        RECT 40.120 916.340 40.380 916.600 ;
        RECT 48.400 916.340 48.660 916.600 ;
        RECT 62.200 916.340 62.460 916.600 ;
        RECT 206.640 916.340 206.900 916.600 ;
        RECT 207.100 916.340 207.360 916.600 ;
        RECT 241.600 916.680 241.860 916.940 ;
        RECT 289.440 916.340 289.700 916.600 ;
        RECT 303.240 916.340 303.500 916.600 ;
        RECT 303.700 916.340 303.960 916.600 ;
        RECT 338.200 916.680 338.460 916.940 ;
        RECT 386.040 916.340 386.300 916.600 ;
        RECT 399.840 916.340 400.100 916.600 ;
        RECT 400.300 916.340 400.560 916.600 ;
        RECT 448.140 916.680 448.400 916.940 ;
        RECT 448.600 916.340 448.860 916.600 ;
        RECT 476.200 916.340 476.460 916.600 ;
        RECT 524.040 916.340 524.300 916.600 ;
        RECT 572.800 916.340 573.060 916.600 ;
        RECT 620.640 916.000 620.900 916.260 ;
        RECT 572.800 915.320 573.060 915.580 ;
        RECT 620.640 915.320 620.900 915.580 ;
        RECT 656.060 914.980 656.320 915.240 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 39.660 3477.190 39.920 3477.510 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 39.720 3429.570 39.860 3477.190 ;
        RECT 39.660 3429.250 39.920 3429.570 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3270.790 40.320 3318.670 ;
        RECT 40.120 3270.470 40.380 3270.790 ;
        RECT 41.040 3270.470 41.300 3270.790 ;
        RECT 41.100 3222.250 41.240 3270.470 ;
        RECT 40.180 3222.110 41.240 3222.250 ;
        RECT 40.180 3174.230 40.320 3222.110 ;
        RECT 40.120 3173.910 40.380 3174.230 ;
        RECT 41.040 3173.910 41.300 3174.230 ;
        RECT 41.100 3125.690 41.240 3173.910 ;
        RECT 40.180 3125.550 41.240 3125.690 ;
        RECT 40.180 3077.670 40.320 3125.550 ;
        RECT 40.120 3077.350 40.380 3077.670 ;
        RECT 41.040 3077.350 41.300 3077.670 ;
        RECT 41.100 3029.130 41.240 3077.350 ;
        RECT 40.180 3028.990 41.240 3029.130 ;
        RECT 40.180 2981.110 40.320 3028.990 ;
        RECT 40.120 2980.790 40.380 2981.110 ;
        RECT 41.040 2980.850 41.300 2981.110 ;
        RECT 40.640 2980.790 41.300 2980.850 ;
        RECT 40.640 2980.710 41.240 2980.790 ;
        RECT 40.640 2959.770 40.780 2980.710 ;
        RECT 40.180 2959.630 40.780 2959.770 ;
        RECT 40.180 2912.170 40.320 2959.630 ;
        RECT 39.720 2912.030 40.320 2912.170 ;
        RECT 39.720 2898.150 39.860 2912.030 ;
        RECT 38.280 2897.830 38.540 2898.150 ;
        RECT 39.660 2897.830 39.920 2898.150 ;
        RECT 38.340 2849.870 38.480 2897.830 ;
        RECT 38.280 2849.550 38.540 2849.870 ;
        RECT 39.200 2849.550 39.460 2849.870 ;
        RECT 39.260 2815.530 39.400 2849.550 ;
        RECT 39.200 2815.210 39.460 2815.530 ;
        RECT 39.660 2814.530 39.920 2814.850 ;
        RECT 39.720 2766.650 39.860 2814.530 ;
        RECT 39.720 2766.510 40.320 2766.650 ;
        RECT 40.180 2752.970 40.320 2766.510 ;
        RECT 40.120 2752.650 40.380 2752.970 ;
        RECT 40.580 2752.650 40.840 2752.970 ;
        RECT 40.640 2705.030 40.780 2752.650 ;
        RECT 40.580 2704.710 40.840 2705.030 ;
        RECT 41.040 2704.710 41.300 2705.030 ;
        RECT 41.100 2670.090 41.240 2704.710 ;
        RECT 40.640 2669.950 41.240 2670.090 ;
        RECT 40.640 2656.605 40.780 2669.950 ;
        RECT 40.570 2656.235 40.850 2656.605 ;
        RECT 41.950 2656.235 42.230 2656.605 ;
        RECT 42.020 2608.470 42.160 2656.235 ;
        RECT 41.040 2608.150 41.300 2608.470 ;
        RECT 41.960 2608.150 42.220 2608.470 ;
        RECT 41.100 2573.530 41.240 2608.150 ;
        RECT 40.640 2573.390 41.240 2573.530 ;
        RECT 40.640 2560.045 40.780 2573.390 ;
        RECT 40.570 2559.675 40.850 2560.045 ;
        RECT 41.950 2559.675 42.230 2560.045 ;
        RECT 42.020 2511.910 42.160 2559.675 ;
        RECT 41.040 2511.590 41.300 2511.910 ;
        RECT 41.960 2511.590 42.220 2511.910 ;
        RECT 41.100 2476.970 41.240 2511.590 ;
        RECT 40.640 2476.830 41.240 2476.970 ;
        RECT 40.640 2429.290 40.780 2476.830 ;
        RECT 40.580 2428.970 40.840 2429.290 ;
        RECT 41.040 2428.630 41.300 2428.950 ;
        RECT 41.100 2415.010 41.240 2428.630 ;
        RECT 39.660 2414.690 39.920 2415.010 ;
        RECT 41.040 2414.690 41.300 2415.010 ;
        RECT 39.720 2366.925 39.860 2414.690 ;
        RECT 39.650 2366.555 39.930 2366.925 ;
        RECT 40.570 2366.555 40.850 2366.925 ;
        RECT 40.640 2332.390 40.780 2366.555 ;
        RECT 40.580 2332.070 40.840 2332.390 ;
        RECT 41.040 2331.730 41.300 2332.050 ;
        RECT 41.100 2283.850 41.240 2331.730 ;
        RECT 40.180 2283.710 41.240 2283.850 ;
        RECT 40.180 2270.170 40.320 2283.710 ;
        RECT 39.200 2269.850 39.460 2270.170 ;
        RECT 40.120 2269.850 40.380 2270.170 ;
        RECT 39.260 2222.230 39.400 2269.850 ;
        RECT 39.200 2221.910 39.460 2222.230 ;
        RECT 39.660 2221.910 39.920 2222.230 ;
        RECT 39.720 2187.290 39.860 2221.910 ;
        RECT 39.720 2187.150 40.780 2187.290 ;
        RECT 40.640 2139.270 40.780 2187.150 ;
        RECT 40.580 2138.950 40.840 2139.270 ;
        RECT 41.040 2138.610 41.300 2138.930 ;
        RECT 41.100 2125.330 41.240 2138.610 ;
        RECT 39.660 2125.010 39.920 2125.330 ;
        RECT 41.040 2125.010 41.300 2125.330 ;
        RECT 39.720 2077.390 39.860 2125.010 ;
        RECT 39.660 2077.070 39.920 2077.390 ;
        RECT 40.580 2077.070 40.840 2077.390 ;
        RECT 40.640 2042.710 40.780 2077.070 ;
        RECT 40.580 2042.390 40.840 2042.710 ;
        RECT 41.040 2041.710 41.300 2042.030 ;
        RECT 41.100 2004.630 41.240 2041.710 ;
        RECT 41.040 2004.310 41.300 2004.630 ;
        RECT 41.960 2004.310 42.220 2004.630 ;
        RECT 42.020 1980.490 42.160 2004.310 ;
        RECT 40.120 1980.170 40.380 1980.490 ;
        RECT 41.960 1980.170 42.220 1980.490 ;
        RECT 40.180 1973.690 40.320 1980.170 ;
        RECT 40.120 1973.370 40.380 1973.690 ;
        RECT 40.580 1973.370 40.840 1973.690 ;
        RECT 40.640 1946.150 40.780 1973.370 ;
        RECT 40.580 1945.830 40.840 1946.150 ;
        RECT 41.040 1945.150 41.300 1945.470 ;
        RECT 41.100 1897.870 41.240 1945.150 ;
        RECT 41.040 1897.550 41.300 1897.870 ;
        RECT 40.120 1897.210 40.380 1897.530 ;
        RECT 40.180 1876.790 40.320 1897.210 ;
        RECT 39.200 1876.470 39.460 1876.790 ;
        RECT 40.120 1876.470 40.380 1876.790 ;
        RECT 39.260 1828.850 39.400 1876.470 ;
        RECT 39.200 1828.530 39.460 1828.850 ;
        RECT 40.580 1828.530 40.840 1828.850 ;
        RECT 40.640 1801.310 40.780 1828.530 ;
        RECT 40.580 1800.990 40.840 1801.310 ;
        RECT 41.040 1800.650 41.300 1800.970 ;
        RECT 41.100 1773.430 41.240 1800.650 ;
        RECT 41.040 1773.110 41.300 1773.430 ;
        RECT 41.960 1773.110 42.220 1773.430 ;
        RECT 42.020 1725.490 42.160 1773.110 ;
        RECT 41.040 1725.170 41.300 1725.490 ;
        RECT 41.960 1725.170 42.220 1725.490 ;
        RECT 41.100 1676.610 41.240 1725.170 ;
        RECT 40.180 1676.470 41.240 1676.610 ;
        RECT 40.180 1628.590 40.320 1676.470 ;
        RECT 40.120 1628.270 40.380 1628.590 ;
        RECT 41.040 1628.270 41.300 1628.590 ;
        RECT 41.100 1580.050 41.240 1628.270 ;
        RECT 40.180 1579.910 41.240 1580.050 ;
        RECT 40.180 1532.030 40.320 1579.910 ;
        RECT 40.120 1531.710 40.380 1532.030 ;
        RECT 41.040 1531.710 41.300 1532.030 ;
        RECT 41.100 1483.490 41.240 1531.710 ;
        RECT 40.180 1483.350 41.240 1483.490 ;
        RECT 40.180 1435.470 40.320 1483.350 ;
        RECT 40.120 1435.150 40.380 1435.470 ;
        RECT 41.040 1435.150 41.300 1435.470 ;
        RECT 41.100 1386.930 41.240 1435.150 ;
        RECT 40.180 1386.790 41.240 1386.930 ;
        RECT 40.180 1338.910 40.320 1386.790 ;
        RECT 40.120 1338.590 40.380 1338.910 ;
        RECT 41.040 1338.650 41.300 1338.910 ;
        RECT 40.640 1338.590 41.300 1338.650 ;
        RECT 40.640 1338.510 41.240 1338.590 ;
        RECT 40.640 1317.570 40.780 1338.510 ;
        RECT 40.180 1317.430 40.780 1317.570 ;
        RECT 40.180 1269.970 40.320 1317.430 ;
        RECT 39.720 1269.830 40.320 1269.970 ;
        RECT 39.720 1255.950 39.860 1269.830 ;
        RECT 38.740 1255.630 39.000 1255.950 ;
        RECT 39.660 1255.630 39.920 1255.950 ;
        RECT 38.800 1207.670 38.940 1255.630 ;
        RECT 38.740 1207.350 39.000 1207.670 ;
        RECT 40.120 1207.350 40.380 1207.670 ;
        RECT 40.180 1173.670 40.320 1207.350 ;
        RECT 40.120 1173.350 40.380 1173.670 ;
        RECT 39.660 1172.670 39.920 1172.990 ;
        RECT 39.720 1159.050 39.860 1172.670 ;
        RECT 38.740 1158.730 39.000 1159.050 ;
        RECT 39.660 1158.730 39.920 1159.050 ;
        RECT 38.800 1111.110 38.940 1158.730 ;
        RECT 38.740 1110.790 39.000 1111.110 ;
        RECT 40.120 1110.790 40.380 1111.110 ;
        RECT 40.180 1077.110 40.320 1110.790 ;
        RECT 40.120 1076.790 40.380 1077.110 ;
        RECT 39.660 1076.110 39.920 1076.430 ;
        RECT 39.720 1027.890 39.860 1076.110 ;
        RECT 39.720 1027.750 40.320 1027.890 ;
        RECT 40.180 1014.405 40.320 1027.750 ;
        RECT 39.190 1014.035 39.470 1014.405 ;
        RECT 40.110 1014.035 40.390 1014.405 ;
        RECT 39.260 979.870 39.400 1014.035 ;
        RECT 39.200 979.550 39.460 979.870 ;
        RECT 40.580 979.550 40.840 979.870 ;
        RECT 40.640 932.125 40.780 979.550 ;
        RECT 40.570 931.755 40.850 932.125 ;
        RECT 40.110 931.075 40.390 931.445 ;
        RECT 40.180 916.630 40.320 931.075 ;
        RECT 241.590 916.795 241.870 917.165 ;
        RECT 289.430 916.795 289.710 917.165 ;
        RECT 338.190 916.795 338.470 917.165 ;
        RECT 386.030 916.795 386.310 917.165 ;
        RECT 448.200 916.970 448.800 917.050 ;
        RECT 448.140 916.910 448.800 916.970 ;
        RECT 241.600 916.650 241.860 916.795 ;
        RECT 289.500 916.630 289.640 916.795 ;
        RECT 338.200 916.650 338.460 916.795 ;
        RECT 386.100 916.630 386.240 916.795 ;
        RECT 448.140 916.650 448.400 916.910 ;
        RECT 448.660 916.630 448.800 916.910 ;
        RECT 524.030 916.795 524.310 917.165 ;
        RECT 524.100 916.630 524.240 916.795 ;
        RECT 40.120 916.310 40.380 916.630 ;
        RECT 48.400 916.485 48.660 916.630 ;
        RECT 62.200 916.485 62.460 916.630 ;
        RECT 48.390 916.115 48.670 916.485 ;
        RECT 62.190 916.115 62.470 916.485 ;
        RECT 206.640 916.370 206.900 916.630 ;
        RECT 207.100 916.370 207.360 916.630 ;
        RECT 206.640 916.310 207.360 916.370 ;
        RECT 289.440 916.310 289.700 916.630 ;
        RECT 303.240 916.370 303.500 916.630 ;
        RECT 303.700 916.370 303.960 916.630 ;
        RECT 303.240 916.310 303.960 916.370 ;
        RECT 386.040 916.310 386.300 916.630 ;
        RECT 399.840 916.370 400.100 916.630 ;
        RECT 400.300 916.370 400.560 916.630 ;
        RECT 399.840 916.310 400.560 916.370 ;
        RECT 448.600 916.310 448.860 916.630 ;
        RECT 476.200 916.485 476.460 916.630 ;
        RECT 206.700 916.230 207.300 916.310 ;
        RECT 303.300 916.230 303.900 916.310 ;
        RECT 399.900 916.230 400.500 916.310 ;
        RECT 476.190 916.115 476.470 916.485 ;
        RECT 524.040 916.310 524.300 916.630 ;
        RECT 572.800 916.310 573.060 916.630 ;
        RECT 572.860 915.610 573.000 916.310 ;
        RECT 620.640 915.970 620.900 916.290 ;
        RECT 620.700 915.610 620.840 915.970 ;
        RECT 572.800 915.290 573.060 915.610 ;
        RECT 620.640 915.290 620.900 915.610 ;
        RECT 656.060 914.950 656.320 915.270 ;
        RECT 656.120 913.765 656.260 914.950 ;
        RECT 656.050 913.395 656.330 913.765 ;
      LAYER via2 ;
        RECT 40.570 2656.280 40.850 2656.560 ;
        RECT 41.950 2656.280 42.230 2656.560 ;
        RECT 40.570 2559.720 40.850 2560.000 ;
        RECT 41.950 2559.720 42.230 2560.000 ;
        RECT 39.650 2366.600 39.930 2366.880 ;
        RECT 40.570 2366.600 40.850 2366.880 ;
        RECT 39.190 1014.080 39.470 1014.360 ;
        RECT 40.110 1014.080 40.390 1014.360 ;
        RECT 40.570 931.800 40.850 932.080 ;
        RECT 40.110 931.120 40.390 931.400 ;
        RECT 241.590 916.840 241.870 917.120 ;
        RECT 289.430 916.840 289.710 917.120 ;
        RECT 338.190 916.840 338.470 917.120 ;
        RECT 386.030 916.840 386.310 917.120 ;
        RECT 524.030 916.840 524.310 917.120 ;
        RECT 48.390 916.160 48.670 916.440 ;
        RECT 62.190 916.160 62.470 916.440 ;
        RECT 476.190 916.160 476.470 916.440 ;
        RECT 656.050 913.440 656.330 913.720 ;
      LAYER met3 ;
        RECT 40.545 2656.570 40.875 2656.585 ;
        RECT 41.925 2656.570 42.255 2656.585 ;
        RECT 40.545 2656.270 42.255 2656.570 ;
        RECT 40.545 2656.255 40.875 2656.270 ;
        RECT 41.925 2656.255 42.255 2656.270 ;
        RECT 40.545 2560.010 40.875 2560.025 ;
        RECT 41.925 2560.010 42.255 2560.025 ;
        RECT 40.545 2559.710 42.255 2560.010 ;
        RECT 40.545 2559.695 40.875 2559.710 ;
        RECT 41.925 2559.695 42.255 2559.710 ;
        RECT 39.625 2366.890 39.955 2366.905 ;
        RECT 40.545 2366.890 40.875 2366.905 ;
        RECT 39.625 2366.590 40.875 2366.890 ;
        RECT 39.625 2366.575 39.955 2366.590 ;
        RECT 40.545 2366.575 40.875 2366.590 ;
        RECT 39.165 1014.370 39.495 1014.385 ;
        RECT 40.085 1014.370 40.415 1014.385 ;
        RECT 39.165 1014.070 40.415 1014.370 ;
        RECT 39.165 1014.055 39.495 1014.070 ;
        RECT 40.085 1014.055 40.415 1014.070 ;
        RECT 40.545 932.090 40.875 932.105 ;
        RECT 39.870 931.790 40.875 932.090 ;
        RECT 39.870 931.425 40.170 931.790 ;
        RECT 40.545 931.775 40.875 931.790 ;
        RECT 39.870 931.110 40.415 931.425 ;
        RECT 40.085 931.095 40.415 931.110 ;
        RECT 241.565 917.130 241.895 917.145 ;
        RECT 289.405 917.130 289.735 917.145 ;
        RECT 241.565 916.830 289.735 917.130 ;
        RECT 241.565 916.815 241.895 916.830 ;
        RECT 289.405 916.815 289.735 916.830 ;
        RECT 338.165 917.130 338.495 917.145 ;
        RECT 386.005 917.130 386.335 917.145 ;
        RECT 524.005 917.130 524.335 917.145 ;
        RECT 338.165 916.830 386.335 917.130 ;
        RECT 338.165 916.815 338.495 916.830 ;
        RECT 386.005 916.815 386.335 916.830 ;
        RECT 476.870 916.830 524.335 917.130 ;
        RECT 48.365 916.450 48.695 916.465 ;
        RECT 62.165 916.450 62.495 916.465 ;
        RECT 48.365 916.150 62.495 916.450 ;
        RECT 48.365 916.135 48.695 916.150 ;
        RECT 62.165 916.135 62.495 916.150 ;
        RECT 476.165 916.450 476.495 916.465 ;
        RECT 476.870 916.450 477.170 916.830 ;
        RECT 524.005 916.815 524.335 916.830 ;
        RECT 476.165 916.150 477.170 916.450 ;
        RECT 476.165 916.135 476.495 916.150 ;
        RECT 656.025 913.730 656.355 913.745 ;
        RECT 656.025 913.430 670.370 913.730 ;
        RECT 656.025 913.415 656.355 913.430 ;
        RECT 670.070 911.400 670.370 913.430 ;
        RECT 670.000 910.800 674.000 911.400 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 917.560 17.410 917.620 ;
        RECT 97.130 917.560 97.450 917.620 ;
        RECT 656.030 917.560 656.350 917.620 ;
        RECT 17.090 917.420 97.450 917.560 ;
        RECT 17.090 917.360 17.410 917.420 ;
        RECT 97.130 917.360 97.450 917.420 ;
        RECT 97.680 917.420 656.350 917.560 ;
        RECT 97.680 917.280 97.820 917.420 ;
        RECT 656.030 917.360 656.350 917.420 ;
        RECT 97.590 917.020 97.910 917.280 ;
      LAYER via ;
        RECT 17.120 917.360 17.380 917.620 ;
        RECT 97.160 917.360 97.420 917.620 ;
        RECT 656.060 917.360 656.320 917.620 ;
        RECT 97.620 917.020 97.880 917.280 ;
      LAYER met2 ;
        RECT 17.110 3267.555 17.390 3267.925 ;
        RECT 17.180 917.650 17.320 3267.555 ;
        RECT 17.120 917.330 17.380 917.650 ;
        RECT 97.160 917.330 97.420 917.650 ;
        RECT 656.060 917.330 656.320 917.650 ;
        RECT 97.220 917.050 97.360 917.330 ;
        RECT 97.620 917.050 97.880 917.310 ;
        RECT 97.220 916.990 97.880 917.050 ;
        RECT 97.220 916.910 97.820 916.990 ;
        RECT 656.120 915.805 656.260 917.330 ;
        RECT 656.050 915.435 656.330 915.805 ;
      LAYER via2 ;
        RECT 17.110 3267.600 17.390 3267.880 ;
        RECT 656.050 915.480 656.330 915.760 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 17.085 3267.890 17.415 3267.905 ;
        RECT -4.800 3267.590 17.415 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 17.085 3267.575 17.415 3267.590 ;
        RECT 656.025 915.770 656.355 915.785 ;
        RECT 670.000 915.770 674.000 916.160 ;
        RECT 656.025 915.560 674.000 915.770 ;
        RECT 656.025 915.470 670.220 915.560 ;
        RECT 656.025 915.455 656.355 915.470 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 924.360 18.330 924.420 ;
        RECT 656.030 924.360 656.350 924.420 ;
        RECT 18.010 924.220 656.350 924.360 ;
        RECT 18.010 924.160 18.330 924.220 ;
        RECT 656.030 924.160 656.350 924.220 ;
      LAYER via ;
        RECT 18.040 924.160 18.300 924.420 ;
        RECT 656.060 924.160 656.320 924.420 ;
      LAYER met2 ;
        RECT 18.030 2979.915 18.310 2980.285 ;
        RECT 18.100 924.450 18.240 2979.915 ;
        RECT 18.040 924.130 18.300 924.450 ;
        RECT 656.060 924.130 656.320 924.450 ;
        RECT 656.120 920.565 656.260 924.130 ;
        RECT 656.050 920.195 656.330 920.565 ;
      LAYER via2 ;
        RECT 18.030 2979.960 18.310 2980.240 ;
        RECT 656.050 920.240 656.330 920.520 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 18.005 2980.250 18.335 2980.265 ;
        RECT -4.800 2979.950 18.335 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 18.005 2979.935 18.335 2979.950 ;
        RECT 656.025 920.530 656.355 920.545 ;
        RECT 670.000 920.530 674.000 920.920 ;
        RECT 656.025 920.320 674.000 920.530 ;
        RECT 656.025 920.230 670.220 920.320 ;
        RECT 656.025 920.215 656.355 920.230 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2691.340 16.030 2691.400 ;
        RECT 24.450 2691.340 24.770 2691.400 ;
        RECT 15.710 2691.200 24.770 2691.340 ;
        RECT 15.710 2691.140 16.030 2691.200 ;
        RECT 24.450 2691.140 24.770 2691.200 ;
        RECT 24.450 931.500 24.770 931.560 ;
        RECT 24.450 931.360 656.720 931.500 ;
        RECT 24.450 931.300 24.770 931.360 ;
        RECT 656.030 930.140 656.350 930.200 ;
        RECT 656.580 930.140 656.720 931.360 ;
        RECT 656.030 930.000 656.720 930.140 ;
        RECT 656.030 929.940 656.350 930.000 ;
      LAYER via ;
        RECT 15.740 2691.140 16.000 2691.400 ;
        RECT 24.480 2691.140 24.740 2691.400 ;
        RECT 24.480 931.300 24.740 931.560 ;
        RECT 656.060 929.940 656.320 930.200 ;
      LAYER met2 ;
        RECT 15.730 2692.955 16.010 2693.325 ;
        RECT 15.800 2691.430 15.940 2692.955 ;
        RECT 15.740 2691.110 16.000 2691.430 ;
        RECT 24.480 2691.110 24.740 2691.430 ;
        RECT 24.540 931.590 24.680 2691.110 ;
        RECT 24.480 931.270 24.740 931.590 ;
        RECT 656.060 929.910 656.320 930.230 ;
        RECT 656.120 926.005 656.260 929.910 ;
        RECT 656.050 925.635 656.330 926.005 ;
      LAYER via2 ;
        RECT 15.730 2693.000 16.010 2693.280 ;
        RECT 656.050 925.680 656.330 925.960 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 15.705 2693.290 16.035 2693.305 ;
        RECT -4.800 2692.990 16.035 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 15.705 2692.975 16.035 2692.990 ;
        RECT 656.025 925.970 656.355 925.985 ;
        RECT 670.000 925.970 674.000 926.360 ;
        RECT 656.025 925.760 674.000 925.970 ;
        RECT 656.025 925.670 670.220 925.760 ;
        RECT 656.025 925.655 656.355 925.670 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2402.340 16.030 2402.400 ;
        RECT 24.910 2402.340 25.230 2402.400 ;
        RECT 15.710 2402.200 25.230 2402.340 ;
        RECT 15.710 2402.140 16.030 2402.200 ;
        RECT 24.910 2402.140 25.230 2402.200 ;
        RECT 24.910 931.160 25.230 931.220 ;
        RECT 656.030 931.160 656.350 931.220 ;
        RECT 24.910 931.020 656.350 931.160 ;
        RECT 24.910 930.960 25.230 931.020 ;
        RECT 656.030 930.960 656.350 931.020 ;
      LAYER via ;
        RECT 15.740 2402.140 16.000 2402.400 ;
        RECT 24.940 2402.140 25.200 2402.400 ;
        RECT 24.940 930.960 25.200 931.220 ;
        RECT 656.060 930.960 656.320 931.220 ;
      LAYER met2 ;
        RECT 15.730 2405.315 16.010 2405.685 ;
        RECT 15.800 2402.430 15.940 2405.315 ;
        RECT 15.740 2402.110 16.000 2402.430 ;
        RECT 24.940 2402.110 25.200 2402.430 ;
        RECT 25.000 931.250 25.140 2402.110 ;
        RECT 24.940 930.930 25.200 931.250 ;
        RECT 656.060 930.930 656.320 931.250 ;
        RECT 656.120 930.765 656.260 930.930 ;
        RECT 656.050 930.395 656.330 930.765 ;
      LAYER via2 ;
        RECT 15.730 2405.360 16.010 2405.640 ;
        RECT 656.050 930.440 656.330 930.720 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 15.705 2405.650 16.035 2405.665 ;
        RECT -4.800 2405.350 16.035 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 15.705 2405.335 16.035 2405.350 ;
        RECT 656.025 930.730 656.355 930.745 ;
        RECT 670.000 930.730 674.000 931.120 ;
        RECT 656.025 930.520 674.000 930.730 ;
        RECT 656.025 930.430 670.220 930.520 ;
        RECT 656.025 930.415 656.355 930.430 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 938.300 20.630 938.360 ;
        RECT 656.030 938.300 656.350 938.360 ;
        RECT 20.310 938.160 656.350 938.300 ;
        RECT 20.310 938.100 20.630 938.160 ;
        RECT 656.030 938.100 656.350 938.160 ;
      LAYER via ;
        RECT 20.340 938.100 20.600 938.360 ;
        RECT 656.060 938.100 656.320 938.360 ;
      LAYER met2 ;
        RECT 20.330 2118.355 20.610 2118.725 ;
        RECT 20.400 938.390 20.540 2118.355 ;
        RECT 20.340 938.070 20.600 938.390 ;
        RECT 656.060 938.070 656.320 938.390 ;
        RECT 656.120 936.205 656.260 938.070 ;
        RECT 656.050 935.835 656.330 936.205 ;
      LAYER via2 ;
        RECT 20.330 2118.400 20.610 2118.680 ;
        RECT 656.050 935.880 656.330 936.160 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 20.305 2118.690 20.635 2118.705 ;
        RECT -4.800 2118.390 20.635 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 20.305 2118.375 20.635 2118.390 ;
        RECT 656.025 936.170 656.355 936.185 ;
        RECT 670.000 936.170 674.000 936.560 ;
        RECT 656.025 935.960 674.000 936.170 ;
        RECT 656.025 935.870 670.220 935.960 ;
        RECT 656.025 935.855 656.355 935.870 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 1828.760 15.570 1828.820 ;
        RECT 25.370 1828.760 25.690 1828.820 ;
        RECT 15.250 1828.620 25.690 1828.760 ;
        RECT 15.250 1828.560 15.570 1828.620 ;
        RECT 25.370 1828.560 25.690 1828.620 ;
        RECT 25.370 945.100 25.690 945.160 ;
        RECT 656.030 945.100 656.350 945.160 ;
        RECT 25.370 944.960 656.350 945.100 ;
        RECT 25.370 944.900 25.690 944.960 ;
        RECT 656.030 944.900 656.350 944.960 ;
      LAYER via ;
        RECT 15.280 1828.560 15.540 1828.820 ;
        RECT 25.400 1828.560 25.660 1828.820 ;
        RECT 25.400 944.900 25.660 945.160 ;
        RECT 656.060 944.900 656.320 945.160 ;
      LAYER met2 ;
        RECT 15.270 1830.715 15.550 1831.085 ;
        RECT 15.340 1828.850 15.480 1830.715 ;
        RECT 15.280 1828.530 15.540 1828.850 ;
        RECT 25.400 1828.530 25.660 1828.850 ;
        RECT 25.460 945.190 25.600 1828.530 ;
        RECT 25.400 944.870 25.660 945.190 ;
        RECT 656.060 944.870 656.320 945.190 ;
        RECT 656.120 940.965 656.260 944.870 ;
        RECT 656.050 940.595 656.330 940.965 ;
      LAYER via2 ;
        RECT 15.270 1830.760 15.550 1831.040 ;
        RECT 656.050 940.640 656.330 940.920 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.245 1831.050 15.575 1831.065 ;
        RECT -4.800 1830.750 15.575 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.245 1830.735 15.575 1830.750 ;
        RECT 656.025 940.930 656.355 940.945 ;
        RECT 670.000 940.930 674.000 941.320 ;
        RECT 656.025 940.720 674.000 940.930 ;
        RECT 656.025 940.630 670.220 940.720 ;
        RECT 656.025 940.615 656.355 940.630 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2901.290 603.400 2901.610 603.460 ;
        RECT 694.760 603.260 2901.610 603.400 ;
        RECT 667.530 601.020 667.850 601.080 ;
        RECT 694.760 601.020 694.900 603.260 ;
        RECT 2901.290 603.200 2901.610 603.260 ;
        RECT 667.530 600.880 694.900 601.020 ;
        RECT 667.530 600.820 667.850 600.880 ;
      LAYER via ;
        RECT 667.560 600.820 667.820 601.080 ;
        RECT 2901.320 603.200 2901.580 603.460 ;
      LAYER met2 ;
        RECT 667.550 803.915 667.830 804.285 ;
        RECT 667.620 601.110 667.760 803.915 ;
        RECT 2901.310 674.035 2901.590 674.405 ;
        RECT 2901.380 603.490 2901.520 674.035 ;
        RECT 2901.320 603.170 2901.580 603.490 ;
        RECT 667.560 600.790 667.820 601.110 ;
      LAYER via2 ;
        RECT 667.550 803.960 667.830 804.240 ;
        RECT 2901.310 674.080 2901.590 674.360 ;
      LAYER met3 ;
        RECT 667.525 804.250 667.855 804.265 ;
        RECT 670.000 804.250 674.000 804.640 ;
        RECT 667.525 804.040 674.000 804.250 ;
        RECT 667.525 803.950 670.220 804.040 ;
        RECT 667.525 803.935 667.855 803.950 ;
        RECT 2901.285 674.370 2901.615 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2901.285 674.070 2924.800 674.370 ;
        RECT 2901.285 674.055 2901.615 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 1539.080 14.190 1539.140 ;
        RECT 25.830 1539.080 26.150 1539.140 ;
        RECT 13.870 1538.940 26.150 1539.080 ;
        RECT 13.870 1538.880 14.190 1538.940 ;
        RECT 25.830 1538.880 26.150 1538.940 ;
        RECT 25.830 952.240 26.150 952.300 ;
        RECT 25.830 952.100 656.720 952.240 ;
        RECT 25.830 952.040 26.150 952.100 ;
        RECT 656.030 950.540 656.350 950.600 ;
        RECT 656.580 950.540 656.720 952.100 ;
        RECT 656.030 950.400 656.720 950.540 ;
        RECT 656.030 950.340 656.350 950.400 ;
      LAYER via ;
        RECT 13.900 1538.880 14.160 1539.140 ;
        RECT 25.860 1538.880 26.120 1539.140 ;
        RECT 25.860 952.040 26.120 952.300 ;
        RECT 656.060 950.340 656.320 950.600 ;
      LAYER met2 ;
        RECT 13.890 1543.755 14.170 1544.125 ;
        RECT 13.960 1539.170 14.100 1543.755 ;
        RECT 13.900 1538.850 14.160 1539.170 ;
        RECT 25.860 1538.850 26.120 1539.170 ;
        RECT 25.920 952.330 26.060 1538.850 ;
        RECT 25.860 952.010 26.120 952.330 ;
        RECT 656.060 950.310 656.320 950.630 ;
        RECT 656.120 946.405 656.260 950.310 ;
        RECT 656.050 946.035 656.330 946.405 ;
      LAYER via2 ;
        RECT 13.890 1543.800 14.170 1544.080 ;
        RECT 656.050 946.080 656.330 946.360 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 13.865 1544.090 14.195 1544.105 ;
        RECT -4.800 1543.790 14.195 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 13.865 1543.775 14.195 1543.790 ;
        RECT 656.025 946.370 656.355 946.385 ;
        RECT 670.000 946.370 674.000 946.760 ;
        RECT 656.025 946.160 674.000 946.370 ;
        RECT 656.025 946.070 670.220 946.160 ;
        RECT 656.025 946.055 656.355 946.070 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 1324.880 15.110 1324.940 ;
        RECT 26.290 1324.880 26.610 1324.940 ;
        RECT 14.790 1324.740 26.610 1324.880 ;
        RECT 14.790 1324.680 15.110 1324.740 ;
        RECT 26.290 1324.680 26.610 1324.740 ;
        RECT 26.290 951.900 26.610 951.960 ;
        RECT 656.030 951.900 656.350 951.960 ;
        RECT 26.290 951.760 656.350 951.900 ;
        RECT 26.290 951.700 26.610 951.760 ;
        RECT 656.030 951.700 656.350 951.760 ;
      LAYER via ;
        RECT 14.820 1324.680 15.080 1324.940 ;
        RECT 26.320 1324.680 26.580 1324.940 ;
        RECT 26.320 951.700 26.580 951.960 ;
        RECT 656.060 951.700 656.320 951.960 ;
      LAYER met2 ;
        RECT 14.810 1328.195 15.090 1328.565 ;
        RECT 14.880 1324.970 15.020 1328.195 ;
        RECT 14.820 1324.650 15.080 1324.970 ;
        RECT 26.320 1324.650 26.580 1324.970 ;
        RECT 26.380 951.990 26.520 1324.650 ;
        RECT 26.320 951.670 26.580 951.990 ;
        RECT 656.060 951.670 656.320 951.990 ;
        RECT 656.120 951.165 656.260 951.670 ;
        RECT 656.050 950.795 656.330 951.165 ;
      LAYER via2 ;
        RECT 14.810 1328.240 15.090 1328.520 ;
        RECT 656.050 950.840 656.330 951.120 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 14.785 1328.530 15.115 1328.545 ;
        RECT -4.800 1328.230 15.115 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 14.785 1328.215 15.115 1328.230 ;
        RECT 656.025 951.130 656.355 951.145 ;
        RECT 670.000 951.130 674.000 951.520 ;
        RECT 656.025 950.920 674.000 951.130 ;
        RECT 656.025 950.830 670.220 950.920 ;
        RECT 656.025 950.815 656.355 950.830 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 1112.720 14.650 1112.780 ;
        RECT 27.210 1112.720 27.530 1112.780 ;
        RECT 14.330 1112.580 27.530 1112.720 ;
        RECT 14.330 1112.520 14.650 1112.580 ;
        RECT 27.210 1112.520 27.530 1112.580 ;
        RECT 27.210 958.700 27.530 958.760 ;
        RECT 656.030 958.700 656.350 958.760 ;
        RECT 27.210 958.560 656.350 958.700 ;
        RECT 27.210 958.500 27.530 958.560 ;
        RECT 656.030 958.500 656.350 958.560 ;
      LAYER via ;
        RECT 14.360 1112.520 14.620 1112.780 ;
        RECT 27.240 1112.520 27.500 1112.780 ;
        RECT 27.240 958.500 27.500 958.760 ;
        RECT 656.060 958.500 656.320 958.760 ;
      LAYER met2 ;
        RECT 14.350 1112.635 14.630 1113.005 ;
        RECT 14.360 1112.490 14.620 1112.635 ;
        RECT 27.240 1112.490 27.500 1112.810 ;
        RECT 27.300 958.790 27.440 1112.490 ;
        RECT 27.240 958.470 27.500 958.790 ;
        RECT 656.060 958.470 656.320 958.790 ;
        RECT 656.120 956.605 656.260 958.470 ;
        RECT 656.050 956.235 656.330 956.605 ;
      LAYER via2 ;
        RECT 14.350 1112.680 14.630 1112.960 ;
        RECT 656.050 956.280 656.330 956.560 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 14.325 1112.970 14.655 1112.985 ;
        RECT -4.800 1112.670 14.655 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 14.325 1112.655 14.655 1112.670 ;
        RECT 656.025 956.570 656.355 956.585 ;
        RECT 670.000 956.570 674.000 956.960 ;
        RECT 656.025 956.360 674.000 956.570 ;
        RECT 656.025 956.270 670.220 956.360 ;
        RECT 656.025 956.255 656.355 956.270 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 30.890 959.720 31.210 959.780 ;
        RECT 656.030 959.720 656.350 959.780 ;
        RECT 30.890 959.580 656.350 959.720 ;
        RECT 30.890 959.520 31.210 959.580 ;
        RECT 656.030 959.520 656.350 959.580 ;
        RECT 18.010 897.500 18.330 897.560 ;
        RECT 30.890 897.500 31.210 897.560 ;
        RECT 18.010 897.360 31.210 897.500 ;
        RECT 18.010 897.300 18.330 897.360 ;
        RECT 30.890 897.300 31.210 897.360 ;
      LAYER via ;
        RECT 30.920 959.520 31.180 959.780 ;
        RECT 656.060 959.520 656.320 959.780 ;
        RECT 18.040 897.300 18.300 897.560 ;
        RECT 30.920 897.300 31.180 897.560 ;
      LAYER met2 ;
        RECT 656.050 960.995 656.330 961.365 ;
        RECT 656.120 959.810 656.260 960.995 ;
        RECT 30.920 959.490 31.180 959.810 ;
        RECT 656.060 959.490 656.320 959.810 ;
        RECT 30.980 897.590 31.120 959.490 ;
        RECT 18.040 897.445 18.300 897.590 ;
        RECT 18.030 897.075 18.310 897.445 ;
        RECT 30.920 897.270 31.180 897.590 ;
      LAYER via2 ;
        RECT 656.050 961.040 656.330 961.320 ;
        RECT 18.030 897.120 18.310 897.400 ;
      LAYER met3 ;
        RECT 656.025 961.330 656.355 961.345 ;
        RECT 670.000 961.330 674.000 961.720 ;
        RECT 656.025 961.120 674.000 961.330 ;
        RECT 656.025 961.030 670.220 961.120 ;
        RECT 656.025 961.015 656.355 961.030 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 18.005 897.410 18.335 897.425 ;
        RECT -4.800 897.110 18.335 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 18.005 897.095 18.335 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.030 961.760 656.350 961.820 ;
        RECT 656.030 961.620 656.720 961.760 ;
        RECT 656.030 961.560 656.350 961.620 ;
        RECT 26.750 959.380 27.070 959.440 ;
        RECT 656.580 959.380 656.720 961.620 ;
        RECT 26.750 959.240 656.720 959.380 ;
        RECT 26.750 959.180 27.070 959.240 ;
        RECT 13.870 681.940 14.190 682.000 ;
        RECT 26.750 681.940 27.070 682.000 ;
        RECT 13.870 681.800 27.070 681.940 ;
        RECT 13.870 681.740 14.190 681.800 ;
        RECT 26.750 681.740 27.070 681.800 ;
      LAYER via ;
        RECT 656.060 961.560 656.320 961.820 ;
        RECT 26.780 959.180 27.040 959.440 ;
        RECT 13.900 681.740 14.160 682.000 ;
        RECT 26.780 681.740 27.040 682.000 ;
      LAYER met2 ;
        RECT 656.050 965.755 656.330 966.125 ;
        RECT 656.120 961.850 656.260 965.755 ;
        RECT 656.060 961.530 656.320 961.850 ;
        RECT 26.780 959.150 27.040 959.470 ;
        RECT 26.840 682.030 26.980 959.150 ;
        RECT 13.900 681.885 14.160 682.030 ;
        RECT 13.890 681.515 14.170 681.885 ;
        RECT 26.780 681.710 27.040 682.030 ;
      LAYER via2 ;
        RECT 656.050 965.800 656.330 966.080 ;
        RECT 13.890 681.560 14.170 681.840 ;
      LAYER met3 ;
        RECT 656.025 966.090 656.355 966.105 ;
        RECT 670.000 966.090 674.000 966.480 ;
        RECT 656.025 965.880 674.000 966.090 ;
        RECT 656.025 965.790 670.220 965.880 ;
        RECT 656.025 965.775 656.355 965.790 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 13.865 681.850 14.195 681.865 ;
        RECT -4.800 681.550 14.195 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 13.865 681.535 14.195 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.770 968.220 435.090 968.280 ;
        RECT 482.610 968.220 482.930 968.280 ;
        RECT 434.770 968.080 482.930 968.220 ;
        RECT 434.770 968.020 435.090 968.080 ;
        RECT 482.610 968.020 482.930 968.080 ;
        RECT 144.970 967.880 145.290 967.940 ;
        RECT 241.570 967.880 241.890 967.940 ;
        RECT 338.170 967.880 338.490 967.940 ;
        RECT 116.540 967.740 145.290 967.880 ;
        RECT 110.010 967.540 110.330 967.600 ;
        RECT 96.300 967.400 110.330 967.540 ;
        RECT 96.300 967.260 96.440 967.400 ;
        RECT 110.010 967.340 110.330 967.400 ;
        RECT 110.470 967.540 110.790 967.600 ;
        RECT 116.540 967.540 116.680 967.740 ;
        RECT 144.970 967.680 145.290 967.740 ;
        RECT 213.140 967.740 241.890 967.880 ;
        RECT 110.470 967.400 116.680 967.540 ;
        RECT 192.810 967.540 193.130 967.600 ;
        RECT 206.610 967.540 206.930 967.600 ;
        RECT 192.810 967.400 206.930 967.540 ;
        RECT 110.470 967.340 110.790 967.400 ;
        RECT 192.810 967.340 193.130 967.400 ;
        RECT 206.610 967.340 206.930 967.400 ;
        RECT 207.070 967.540 207.390 967.600 ;
        RECT 213.140 967.540 213.280 967.740 ;
        RECT 241.570 967.680 241.890 967.740 ;
        RECT 309.740 967.740 338.490 967.880 ;
        RECT 207.070 967.400 213.280 967.540 ;
        RECT 289.410 967.540 289.730 967.600 ;
        RECT 303.210 967.540 303.530 967.600 ;
        RECT 289.410 967.400 303.530 967.540 ;
        RECT 207.070 967.340 207.390 967.400 ;
        RECT 289.410 967.340 289.730 967.400 ;
        RECT 303.210 967.340 303.530 967.400 ;
        RECT 303.670 967.540 303.990 967.600 ;
        RECT 309.740 967.540 309.880 967.740 ;
        RECT 338.170 967.680 338.490 967.740 ;
        RECT 572.770 967.880 573.090 967.940 ;
        RECT 620.610 967.880 620.930 967.940 ;
        RECT 572.770 967.740 620.930 967.880 ;
        RECT 572.770 967.680 573.090 967.740 ;
        RECT 620.610 967.680 620.930 967.740 ;
        RECT 303.670 967.400 309.880 967.540 ;
        RECT 400.730 967.540 401.050 967.600 ;
        RECT 434.770 967.540 435.090 967.600 ;
        RECT 400.730 967.400 435.090 967.540 ;
        RECT 303.670 967.340 303.990 967.400 ;
        RECT 400.730 967.340 401.050 967.400 ;
        RECT 434.770 967.340 435.090 967.400 ;
        RECT 96.210 967.000 96.530 967.260 ;
        RECT 386.010 967.200 386.330 967.260 ;
        RECT 399.810 967.200 400.130 967.260 ;
        RECT 386.010 967.060 400.130 967.200 ;
        RECT 386.010 967.000 386.330 967.060 ;
        RECT 399.810 967.000 400.130 967.060 ;
        RECT 545.170 967.200 545.490 967.260 ;
        RECT 572.770 967.200 573.090 967.260 ;
        RECT 545.170 967.060 573.090 967.200 ;
        RECT 545.170 967.000 545.490 967.060 ;
        RECT 572.770 967.000 573.090 967.060 ;
        RECT 482.610 966.860 482.930 966.920 ;
        RECT 495.950 966.860 496.270 966.920 ;
        RECT 482.610 966.720 496.270 966.860 ;
        RECT 482.610 966.660 482.930 966.720 ;
        RECT 495.950 966.660 496.270 966.720 ;
        RECT 620.610 966.860 620.930 966.920 ;
        RECT 620.610 966.720 641.540 966.860 ;
        RECT 620.610 966.660 620.930 966.720 ;
        RECT 51.590 966.520 51.910 966.580 ;
        RECT 96.210 966.520 96.530 966.580 ;
        RECT 51.590 966.380 96.530 966.520 ;
        RECT 51.590 966.320 51.910 966.380 ;
        RECT 96.210 966.320 96.530 966.380 ;
        RECT 497.330 966.520 497.650 966.580 ;
        RECT 544.710 966.520 545.030 966.580 ;
        RECT 497.330 966.380 545.030 966.520 ;
        RECT 641.400 966.520 641.540 966.720 ;
        RECT 656.030 966.520 656.350 966.580 ;
        RECT 641.400 966.380 656.350 966.520 ;
        RECT 497.330 966.320 497.650 966.380 ;
        RECT 544.710 966.320 545.030 966.380 ;
        RECT 656.030 966.320 656.350 966.380 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 51.590 469.100 51.910 469.160 ;
        RECT 17.090 468.960 51.910 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 51.590 468.900 51.910 468.960 ;
      LAYER via ;
        RECT 434.800 968.020 435.060 968.280 ;
        RECT 482.640 968.020 482.900 968.280 ;
        RECT 110.040 967.340 110.300 967.600 ;
        RECT 110.500 967.340 110.760 967.600 ;
        RECT 145.000 967.680 145.260 967.940 ;
        RECT 192.840 967.340 193.100 967.600 ;
        RECT 206.640 967.340 206.900 967.600 ;
        RECT 207.100 967.340 207.360 967.600 ;
        RECT 241.600 967.680 241.860 967.940 ;
        RECT 289.440 967.340 289.700 967.600 ;
        RECT 303.240 967.340 303.500 967.600 ;
        RECT 303.700 967.340 303.960 967.600 ;
        RECT 338.200 967.680 338.460 967.940 ;
        RECT 572.800 967.680 573.060 967.940 ;
        RECT 620.640 967.680 620.900 967.940 ;
        RECT 400.760 967.340 401.020 967.600 ;
        RECT 434.800 967.340 435.060 967.600 ;
        RECT 96.240 967.000 96.500 967.260 ;
        RECT 386.040 967.000 386.300 967.260 ;
        RECT 399.840 967.000 400.100 967.260 ;
        RECT 545.200 967.000 545.460 967.260 ;
        RECT 572.800 967.000 573.060 967.260 ;
        RECT 482.640 966.660 482.900 966.920 ;
        RECT 495.980 966.660 496.240 966.920 ;
        RECT 620.640 966.660 620.900 966.920 ;
        RECT 51.620 966.320 51.880 966.580 ;
        RECT 96.240 966.320 96.500 966.580 ;
        RECT 497.360 966.320 497.620 966.580 ;
        RECT 544.740 966.320 545.000 966.580 ;
        RECT 656.060 966.320 656.320 966.580 ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 51.620 468.900 51.880 469.160 ;
      LAYER met2 ;
        RECT 656.050 971.195 656.330 971.565 ;
        RECT 144.990 967.795 145.270 968.165 ;
        RECT 192.830 967.795 193.110 968.165 ;
        RECT 241.590 967.795 241.870 968.165 ;
        RECT 289.430 967.795 289.710 968.165 ;
        RECT 338.190 967.795 338.470 968.165 ;
        RECT 385.110 967.795 385.390 968.165 ;
        RECT 434.800 967.990 435.060 968.310 ;
        RECT 482.640 967.990 482.900 968.310 ;
        RECT 145.000 967.650 145.260 967.795 ;
        RECT 192.900 967.630 193.040 967.795 ;
        RECT 241.600 967.650 241.860 967.795 ;
        RECT 289.500 967.630 289.640 967.795 ;
        RECT 338.200 967.650 338.460 967.795 ;
        RECT 110.040 967.370 110.300 967.630 ;
        RECT 110.500 967.370 110.760 967.630 ;
        RECT 110.040 967.310 110.760 967.370 ;
        RECT 192.840 967.310 193.100 967.630 ;
        RECT 206.640 967.370 206.900 967.630 ;
        RECT 207.100 967.370 207.360 967.630 ;
        RECT 206.640 967.310 207.360 967.370 ;
        RECT 289.440 967.310 289.700 967.630 ;
        RECT 303.240 967.370 303.500 967.630 ;
        RECT 303.700 967.370 303.960 967.630 ;
        RECT 303.240 967.310 303.960 967.370 ;
        RECT 96.240 966.970 96.500 967.290 ;
        RECT 110.100 967.230 110.700 967.310 ;
        RECT 206.700 967.230 207.300 967.310 ;
        RECT 303.300 967.230 303.900 967.310 ;
        RECT 96.300 966.610 96.440 966.970 ;
        RECT 385.180 966.690 385.320 967.795 ;
        RECT 434.860 967.630 435.000 967.990 ;
        RECT 400.760 967.370 401.020 967.630 ;
        RECT 399.900 967.310 401.020 967.370 ;
        RECT 434.800 967.310 435.060 967.630 ;
        RECT 399.900 967.290 400.960 967.310 ;
        RECT 386.040 966.970 386.300 967.290 ;
        RECT 399.840 967.230 400.960 967.290 ;
        RECT 399.840 966.970 400.100 967.230 ;
        RECT 386.100 966.690 386.240 966.970 ;
        RECT 482.700 966.950 482.840 967.990 ;
        RECT 572.800 967.650 573.060 967.970 ;
        RECT 620.640 967.650 620.900 967.970 ;
        RECT 572.860 967.290 573.000 967.650 ;
        RECT 545.200 966.970 545.460 967.290 ;
        RECT 572.800 966.970 573.060 967.290 ;
        RECT 51.620 966.290 51.880 966.610 ;
        RECT 96.240 966.290 96.500 966.610 ;
        RECT 385.180 966.550 386.240 966.690 ;
        RECT 482.640 966.630 482.900 966.950 ;
        RECT 495.980 966.805 496.240 966.950 ;
        RECT 495.970 966.435 496.250 966.805 ;
        RECT 497.350 966.435 497.630 966.805 ;
        RECT 545.260 966.690 545.400 966.970 ;
        RECT 620.700 966.950 620.840 967.650 ;
        RECT 544.800 966.610 545.400 966.690 ;
        RECT 620.640 966.630 620.900 966.950 ;
        RECT 656.120 966.610 656.260 971.195 ;
        RECT 544.740 966.550 545.400 966.610 ;
        RECT 497.360 966.290 497.620 966.435 ;
        RECT 544.740 966.290 545.000 966.550 ;
        RECT 656.060 966.290 656.320 966.610 ;
        RECT 51.680 469.190 51.820 966.290 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 51.620 468.870 51.880 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 656.050 971.240 656.330 971.520 ;
        RECT 144.990 967.840 145.270 968.120 ;
        RECT 192.830 967.840 193.110 968.120 ;
        RECT 241.590 967.840 241.870 968.120 ;
        RECT 289.430 967.840 289.710 968.120 ;
        RECT 338.190 967.840 338.470 968.120 ;
        RECT 385.110 967.840 385.390 968.120 ;
        RECT 495.970 966.480 496.250 966.760 ;
        RECT 497.350 966.480 497.630 966.760 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 656.025 971.530 656.355 971.545 ;
        RECT 670.000 971.530 674.000 971.920 ;
        RECT 656.025 971.320 674.000 971.530 ;
        RECT 656.025 971.230 670.220 971.320 ;
        RECT 656.025 971.215 656.355 971.230 ;
        RECT 144.965 968.130 145.295 968.145 ;
        RECT 192.805 968.130 193.135 968.145 ;
        RECT 144.965 967.830 193.135 968.130 ;
        RECT 144.965 967.815 145.295 967.830 ;
        RECT 192.805 967.815 193.135 967.830 ;
        RECT 241.565 968.130 241.895 968.145 ;
        RECT 289.405 968.130 289.735 968.145 ;
        RECT 241.565 967.830 289.735 968.130 ;
        RECT 241.565 967.815 241.895 967.830 ;
        RECT 289.405 967.815 289.735 967.830 ;
        RECT 338.165 968.130 338.495 968.145 ;
        RECT 385.085 968.130 385.415 968.145 ;
        RECT 338.165 967.830 385.415 968.130 ;
        RECT 338.165 967.815 338.495 967.830 ;
        RECT 385.085 967.815 385.415 967.830 ;
        RECT 495.945 966.770 496.275 966.785 ;
        RECT 497.325 966.770 497.655 966.785 ;
        RECT 495.945 966.470 497.655 966.770 ;
        RECT 495.945 966.455 496.275 966.470 ;
        RECT 497.325 966.455 497.655 966.470 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 972.980 16.490 973.040 ;
        RECT 656.030 972.980 656.350 973.040 ;
        RECT 16.170 972.840 656.350 972.980 ;
        RECT 16.170 972.780 16.490 972.840 ;
        RECT 656.030 972.780 656.350 972.840 ;
      LAYER via ;
        RECT 16.200 972.780 16.460 973.040 ;
        RECT 656.060 972.780 656.320 973.040 ;
      LAYER met2 ;
        RECT 656.050 975.955 656.330 976.325 ;
        RECT 656.120 973.070 656.260 975.955 ;
        RECT 16.200 972.750 16.460 973.070 ;
        RECT 656.060 972.750 656.320 973.070 ;
        RECT 16.260 250.765 16.400 972.750 ;
        RECT 16.190 250.395 16.470 250.765 ;
      LAYER via2 ;
        RECT 656.050 976.000 656.330 976.280 ;
        RECT 16.190 250.440 16.470 250.720 ;
      LAYER met3 ;
        RECT 656.025 976.290 656.355 976.305 ;
        RECT 670.000 976.290 674.000 976.680 ;
        RECT 656.025 976.080 674.000 976.290 ;
        RECT 656.025 975.990 670.220 976.080 ;
        RECT 656.025 975.975 656.355 975.990 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 16.165 250.730 16.495 250.745 ;
        RECT -4.800 250.430 16.495 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 16.165 250.415 16.495 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.390 980.120 19.710 980.180 ;
        RECT 656.030 980.120 656.350 980.180 ;
        RECT 19.390 979.980 656.350 980.120 ;
        RECT 19.390 979.920 19.710 979.980 ;
        RECT 656.030 979.920 656.350 979.980 ;
      LAYER via ;
        RECT 19.420 979.920 19.680 980.180 ;
        RECT 656.060 979.920 656.320 980.180 ;
      LAYER met2 ;
        RECT 656.050 981.395 656.330 981.765 ;
        RECT 656.120 980.210 656.260 981.395 ;
        RECT 19.420 979.890 19.680 980.210 ;
        RECT 656.060 979.890 656.320 980.210 ;
        RECT 19.480 35.885 19.620 979.890 ;
        RECT 19.410 35.515 19.690 35.885 ;
      LAYER via2 ;
        RECT 656.050 981.440 656.330 981.720 ;
        RECT 19.410 35.560 19.690 35.840 ;
      LAYER met3 ;
        RECT 656.025 981.730 656.355 981.745 ;
        RECT 670.000 981.730 674.000 982.120 ;
        RECT 656.025 981.520 674.000 981.730 ;
        RECT 656.025 981.430 670.220 981.520 ;
        RECT 656.025 981.415 656.355 981.430 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 19.385 35.850 19.715 35.865 ;
        RECT -4.800 35.550 19.715 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 19.385 35.535 19.715 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 958.250 1000.860 958.570 1000.920 ;
        RECT 933.960 1000.720 958.570 1000.860 ;
        RECT 933.960 1000.180 934.100 1000.720 ;
        RECT 958.250 1000.660 958.570 1000.720 ;
        RECT 2042.010 1000.520 2042.330 1000.580 ;
        RECT 883.820 1000.040 934.100 1000.180 ;
        RECT 1993.800 1000.380 2042.330 1000.520 ;
        RECT 863.030 999.840 863.350 999.900 ;
        RECT 883.820 999.840 883.960 1000.040 ;
        RECT 863.030 999.700 883.960 999.840 ;
        RECT 960.550 999.840 960.870 999.900 ;
        RECT 1464.710 999.840 1465.030 999.900 ;
        RECT 1837.770 999.840 1838.090 999.900 ;
        RECT 1883.770 999.840 1884.090 999.900 ;
        RECT 1993.800 999.840 1993.940 1000.380 ;
        RECT 2042.010 1000.320 2042.330 1000.380 ;
        RECT 2042.470 1000.520 2042.790 1000.580 ;
        RECT 2042.470 1000.380 2052.820 1000.520 ;
        RECT 2042.470 1000.320 2042.790 1000.380 ;
        RECT 2052.680 1000.180 2052.820 1000.380 ;
        RECT 2076.970 1000.180 2077.290 1000.240 ;
        RECT 2052.680 1000.040 2077.290 1000.180 ;
        RECT 2076.970 999.980 2077.290 1000.040 ;
        RECT 960.550 999.700 1072.100 999.840 ;
        RECT 863.030 999.640 863.350 999.700 ;
        RECT 960.550 999.640 960.870 999.700 ;
        RECT 668.450 999.500 668.770 999.560 ;
        RECT 668.450 999.360 835.200 999.500 ;
        RECT 668.450 999.300 668.770 999.360 ;
        RECT 835.060 998.820 835.200 999.360 ;
        RECT 863.030 998.960 863.350 999.220 ;
        RECT 863.120 998.820 863.260 998.960 ;
        RECT 835.060 998.680 863.260 998.820 ;
        RECT 1071.960 998.820 1072.100 999.700 ;
        RECT 1172.700 999.700 1252.880 999.840 ;
        RECT 1172.700 998.820 1172.840 999.700 ;
        RECT 1071.960 998.680 1172.840 998.820 ;
        RECT 1252.740 998.820 1252.880 999.700 ;
        RECT 1464.710 999.700 1564.300 999.840 ;
        RECT 1464.710 999.640 1465.030 999.700 ;
        RECT 1366.360 999.360 1371.100 999.500 ;
        RECT 1366.360 999.160 1366.500 999.360 ;
        RECT 1363.140 999.020 1366.500 999.160 ;
        RECT 1363.140 998.820 1363.280 999.020 ;
        RECT 1252.740 998.680 1363.280 998.820 ;
        RECT 1370.960 998.820 1371.100 999.360 ;
        RECT 1456.890 998.960 1457.210 999.220 ;
        RECT 1564.160 999.160 1564.300 999.700 ;
        RECT 1656.160 999.700 1763.940 999.840 ;
        RECT 1565.080 999.360 1570.740 999.500 ;
        RECT 1565.080 999.160 1565.220 999.360 ;
        RECT 1564.160 999.020 1565.220 999.160 ;
        RECT 1456.980 998.820 1457.120 998.960 ;
        RECT 1370.960 998.680 1457.120 998.820 ;
        RECT 1570.600 998.820 1570.740 999.360 ;
        RECT 1656.160 998.820 1656.300 999.700 ;
        RECT 1570.600 998.680 1656.300 998.820 ;
        RECT 1763.800 998.820 1763.940 999.700 ;
        RECT 1837.770 999.700 1884.090 999.840 ;
        RECT 1837.770 999.640 1838.090 999.700 ;
        RECT 1883.770 999.640 1884.090 999.700 ;
        RECT 1949.180 999.700 1993.940 999.840 ;
        RECT 1909.070 999.300 1909.390 999.560 ;
        RECT 1837.770 998.960 1838.090 999.220 ;
        RECT 1837.860 998.820 1838.000 998.960 ;
        RECT 1763.800 998.680 1838.000 998.820 ;
        RECT 1909.160 998.820 1909.300 999.300 ;
        RECT 1949.180 998.820 1949.320 999.700 ;
        RECT 2091.690 998.960 2092.010 999.220 ;
        RECT 2148.270 998.960 2148.590 999.220 ;
        RECT 1909.160 998.680 1949.320 998.820 ;
        RECT 2091.780 998.820 2091.920 998.960 ;
        RECT 2148.360 998.820 2148.500 998.960 ;
        RECT 2091.780 998.680 2148.500 998.820 ;
        RECT 2171.270 998.820 2171.590 998.880 ;
        RECT 2901.750 998.820 2902.070 998.880 ;
        RECT 2171.270 998.680 2902.070 998.820 ;
        RECT 2171.270 998.620 2171.590 998.680 ;
        RECT 2901.750 998.620 2902.070 998.680 ;
      LAYER via ;
        RECT 958.280 1000.660 958.540 1000.920 ;
        RECT 863.060 999.640 863.320 999.900 ;
        RECT 960.580 999.640 960.840 999.900 ;
        RECT 668.480 999.300 668.740 999.560 ;
        RECT 863.060 998.960 863.320 999.220 ;
        RECT 1464.740 999.640 1465.000 999.900 ;
        RECT 1456.920 998.960 1457.180 999.220 ;
        RECT 1837.800 999.640 1838.060 999.900 ;
        RECT 1883.800 999.640 1884.060 999.900 ;
        RECT 2042.040 1000.320 2042.300 1000.580 ;
        RECT 2042.500 1000.320 2042.760 1000.580 ;
        RECT 2077.000 999.980 2077.260 1000.240 ;
        RECT 1909.100 999.300 1909.360 999.560 ;
        RECT 1837.800 998.960 1838.060 999.220 ;
        RECT 2091.720 998.960 2091.980 999.220 ;
        RECT 2148.300 998.960 2148.560 999.220 ;
        RECT 2171.300 998.620 2171.560 998.880 ;
        RECT 2901.780 998.620 2902.040 998.880 ;
      LAYER met2 ;
        RECT 958.280 1000.635 958.540 1000.950 ;
        RECT 958.270 1000.265 958.550 1000.635 ;
        RECT 2042.100 1000.610 2042.700 1000.690 ;
        RECT 2042.040 1000.550 2042.760 1000.610 ;
        RECT 2042.040 1000.290 2042.300 1000.550 ;
        RECT 2042.500 1000.290 2042.760 1000.550 ;
        RECT 2077.000 1000.125 2077.260 1000.270 ;
        RECT 863.060 999.610 863.320 999.930 ;
        RECT 960.570 999.755 960.850 1000.125 ;
        RECT 1456.910 999.755 1457.190 1000.125 ;
        RECT 1464.730 999.755 1465.010 1000.125 ;
        RECT 960.580 999.610 960.840 999.755 ;
        RECT 668.480 999.270 668.740 999.590 ;
        RECT 668.540 809.725 668.680 999.270 ;
        RECT 863.120 999.250 863.260 999.610 ;
        RECT 1456.980 999.250 1457.120 999.755 ;
        RECT 1464.740 999.610 1465.000 999.755 ;
        RECT 1837.800 999.610 1838.060 999.930 ;
        RECT 1883.790 999.755 1884.070 1000.125 ;
        RECT 1909.090 999.755 1909.370 1000.125 ;
        RECT 2076.990 999.755 2077.270 1000.125 ;
        RECT 2091.710 999.755 2091.990 1000.125 ;
        RECT 1883.800 999.610 1884.060 999.755 ;
        RECT 1837.860 999.250 1838.000 999.610 ;
        RECT 1909.160 999.590 1909.300 999.755 ;
        RECT 1909.100 999.270 1909.360 999.590 ;
        RECT 2091.780 999.250 2091.920 999.755 ;
        RECT 863.060 998.930 863.320 999.250 ;
        RECT 1456.920 998.930 1457.180 999.250 ;
        RECT 1837.800 998.930 1838.060 999.250 ;
        RECT 2091.720 998.930 2091.980 999.250 ;
        RECT 2148.290 999.075 2148.570 999.445 ;
        RECT 2171.290 999.075 2171.570 999.445 ;
        RECT 2148.300 998.930 2148.560 999.075 ;
        RECT 2171.360 998.910 2171.500 999.075 ;
        RECT 2171.300 998.590 2171.560 998.910 ;
        RECT 2901.780 998.590 2902.040 998.910 ;
        RECT 2901.840 909.685 2901.980 998.590 ;
        RECT 2901.770 909.315 2902.050 909.685 ;
        RECT 668.470 809.355 668.750 809.725 ;
      LAYER via2 ;
        RECT 958.270 1000.310 958.550 1000.590 ;
        RECT 960.570 999.800 960.850 1000.080 ;
        RECT 1456.910 999.800 1457.190 1000.080 ;
        RECT 1464.730 999.800 1465.010 1000.080 ;
        RECT 1883.790 999.800 1884.070 1000.080 ;
        RECT 1909.090 999.800 1909.370 1000.080 ;
        RECT 2076.990 999.800 2077.270 1000.080 ;
        RECT 2091.710 999.800 2091.990 1000.080 ;
        RECT 2148.290 999.120 2148.570 999.400 ;
        RECT 2171.290 999.120 2171.570 999.400 ;
        RECT 2901.770 909.360 2902.050 909.640 ;
        RECT 668.470 809.400 668.750 809.680 ;
      LAYER met3 ;
        RECT 958.245 1000.600 958.575 1000.615 ;
        RECT 958.245 1000.300 959.250 1000.600 ;
        RECT 958.245 1000.285 958.575 1000.300 ;
        RECT 958.950 1000.090 959.250 1000.300 ;
        RECT 960.545 1000.090 960.875 1000.105 ;
        RECT 958.950 999.790 960.875 1000.090 ;
        RECT 960.545 999.775 960.875 999.790 ;
        RECT 1456.885 1000.090 1457.215 1000.105 ;
        RECT 1464.705 1000.090 1465.035 1000.105 ;
        RECT 1456.885 999.790 1465.035 1000.090 ;
        RECT 1456.885 999.775 1457.215 999.790 ;
        RECT 1464.705 999.775 1465.035 999.790 ;
        RECT 1883.765 1000.090 1884.095 1000.105 ;
        RECT 1909.065 1000.090 1909.395 1000.105 ;
        RECT 1883.765 999.790 1909.395 1000.090 ;
        RECT 1883.765 999.775 1884.095 999.790 ;
        RECT 1909.065 999.775 1909.395 999.790 ;
        RECT 2076.965 1000.090 2077.295 1000.105 ;
        RECT 2091.685 1000.090 2092.015 1000.105 ;
        RECT 2076.965 999.790 2092.015 1000.090 ;
        RECT 2076.965 999.775 2077.295 999.790 ;
        RECT 2091.685 999.775 2092.015 999.790 ;
        RECT 2148.265 999.410 2148.595 999.425 ;
        RECT 2171.265 999.410 2171.595 999.425 ;
        RECT 2148.265 999.110 2171.595 999.410 ;
        RECT 2148.265 999.095 2148.595 999.110 ;
        RECT 2171.265 999.095 2171.595 999.110 ;
        RECT 2901.745 909.650 2902.075 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2901.745 909.350 2924.800 909.650 ;
        RECT 2901.745 909.335 2902.075 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT 668.445 809.690 668.775 809.705 ;
        RECT 670.000 809.690 674.000 810.080 ;
        RECT 668.445 809.480 674.000 809.690 ;
        RECT 668.445 809.390 670.220 809.480 ;
        RECT 668.445 809.375 668.775 809.390 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 663.390 1138.900 663.710 1138.960 ;
        RECT 2898.990 1138.900 2899.310 1138.960 ;
        RECT 663.390 1138.760 2899.310 1138.900 ;
        RECT 663.390 1138.700 663.710 1138.760 ;
        RECT 2898.990 1138.700 2899.310 1138.760 ;
      LAYER via ;
        RECT 663.420 1138.700 663.680 1138.960 ;
        RECT 2899.020 1138.700 2899.280 1138.960 ;
      LAYER met2 ;
        RECT 2899.010 1143.915 2899.290 1144.285 ;
        RECT 2899.080 1138.990 2899.220 1143.915 ;
        RECT 663.420 1138.670 663.680 1138.990 ;
        RECT 2899.020 1138.670 2899.280 1138.990 ;
        RECT 663.480 814.485 663.620 1138.670 ;
        RECT 663.410 814.115 663.690 814.485 ;
      LAYER via2 ;
        RECT 2899.010 1143.960 2899.290 1144.240 ;
        RECT 663.410 814.160 663.690 814.440 ;
      LAYER met3 ;
        RECT 2898.985 1144.250 2899.315 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2898.985 1143.950 2924.800 1144.250 ;
        RECT 2898.985 1143.935 2899.315 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 663.385 814.450 663.715 814.465 ;
        RECT 670.000 814.450 674.000 814.840 ;
        RECT 663.385 814.240 674.000 814.450 ;
        RECT 663.385 814.150 670.220 814.240 ;
        RECT 663.385 814.135 663.715 814.150 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 650.050 1373.500 650.370 1373.560 ;
        RECT 2900.370 1373.500 2900.690 1373.560 ;
        RECT 650.050 1373.360 2900.690 1373.500 ;
        RECT 650.050 1373.300 650.370 1373.360 ;
        RECT 2900.370 1373.300 2900.690 1373.360 ;
        RECT 650.050 821.000 650.370 821.060 ;
        RECT 658.330 821.000 658.650 821.060 ;
        RECT 650.050 820.860 658.650 821.000 ;
        RECT 650.050 820.800 650.370 820.860 ;
        RECT 658.330 820.800 658.650 820.860 ;
      LAYER via ;
        RECT 650.080 1373.300 650.340 1373.560 ;
        RECT 2900.400 1373.300 2900.660 1373.560 ;
        RECT 650.080 820.800 650.340 821.060 ;
        RECT 658.360 820.800 658.620 821.060 ;
      LAYER met2 ;
        RECT 2900.390 1378.515 2900.670 1378.885 ;
        RECT 2900.460 1373.590 2900.600 1378.515 ;
        RECT 650.080 1373.270 650.340 1373.590 ;
        RECT 2900.400 1373.270 2900.660 1373.590 ;
        RECT 650.140 821.090 650.280 1373.270 ;
        RECT 650.080 820.770 650.340 821.090 ;
        RECT 658.360 820.770 658.620 821.090 ;
        RECT 658.420 819.925 658.560 820.770 ;
        RECT 658.350 819.555 658.630 819.925 ;
      LAYER via2 ;
        RECT 2900.390 1378.560 2900.670 1378.840 ;
        RECT 658.350 819.600 658.630 819.880 ;
      LAYER met3 ;
        RECT 2900.365 1378.850 2900.695 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.365 1378.550 2924.800 1378.850 ;
        RECT 2900.365 1378.535 2900.695 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 658.325 819.890 658.655 819.905 ;
        RECT 670.000 819.890 674.000 820.280 ;
        RECT 658.325 819.680 674.000 819.890 ;
        RECT 658.325 819.590 670.220 819.680 ;
        RECT 658.325 819.575 658.655 819.590 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 668.450 1608.100 668.770 1608.160 ;
        RECT 2900.370 1608.100 2900.690 1608.160 ;
        RECT 668.450 1607.960 2900.690 1608.100 ;
        RECT 668.450 1607.900 668.770 1607.960 ;
        RECT 2900.370 1607.900 2900.690 1607.960 ;
        RECT 664.310 1594.160 664.630 1594.220 ;
        RECT 668.450 1594.160 668.770 1594.220 ;
        RECT 664.310 1594.020 668.770 1594.160 ;
        RECT 664.310 1593.960 664.630 1594.020 ;
        RECT 668.450 1593.960 668.770 1594.020 ;
      LAYER via ;
        RECT 668.480 1607.900 668.740 1608.160 ;
        RECT 2900.400 1607.900 2900.660 1608.160 ;
        RECT 664.340 1593.960 664.600 1594.220 ;
        RECT 668.480 1593.960 668.740 1594.220 ;
      LAYER met2 ;
        RECT 2900.390 1613.115 2900.670 1613.485 ;
        RECT 2900.460 1608.190 2900.600 1613.115 ;
        RECT 668.480 1607.870 668.740 1608.190 ;
        RECT 2900.400 1607.870 2900.660 1608.190 ;
        RECT 668.540 1594.250 668.680 1607.870 ;
        RECT 664.340 1593.930 664.600 1594.250 ;
        RECT 668.480 1593.930 668.740 1594.250 ;
        RECT 664.400 824.685 664.540 1593.930 ;
        RECT 664.330 824.315 664.610 824.685 ;
      LAYER via2 ;
        RECT 2900.390 1613.160 2900.670 1613.440 ;
        RECT 664.330 824.360 664.610 824.640 ;
      LAYER met3 ;
        RECT 2900.365 1613.450 2900.695 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.365 1613.150 2924.800 1613.450 ;
        RECT 2900.365 1613.135 2900.695 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 664.305 824.650 664.635 824.665 ;
        RECT 670.000 824.650 674.000 825.040 ;
        RECT 664.305 824.440 674.000 824.650 ;
        RECT 664.305 824.350 670.220 824.440 ;
        RECT 664.305 824.335 664.635 824.350 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 655.570 1004.940 655.890 1005.000 ;
        RECT 2904.050 1004.940 2904.370 1005.000 ;
        RECT 655.570 1004.800 2904.370 1004.940 ;
        RECT 655.570 1004.740 655.890 1004.800 ;
        RECT 2904.050 1004.740 2904.370 1004.800 ;
      LAYER via ;
        RECT 655.600 1004.740 655.860 1005.000 ;
        RECT 2904.080 1004.740 2904.340 1005.000 ;
      LAYER met2 ;
        RECT 2904.070 1847.715 2904.350 1848.085 ;
        RECT 2904.140 1005.030 2904.280 1847.715 ;
        RECT 655.600 1004.710 655.860 1005.030 ;
        RECT 2904.080 1004.710 2904.340 1005.030 ;
        RECT 655.660 829.445 655.800 1004.710 ;
        RECT 655.590 829.075 655.870 829.445 ;
      LAYER via2 ;
        RECT 2904.070 1847.760 2904.350 1848.040 ;
        RECT 655.590 829.120 655.870 829.400 ;
      LAYER met3 ;
        RECT 2904.045 1848.050 2904.375 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2904.045 1847.750 2924.800 1848.050 ;
        RECT 2904.045 1847.735 2904.375 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 655.565 829.410 655.895 829.425 ;
        RECT 670.000 829.410 674.000 829.800 ;
        RECT 655.565 829.200 674.000 829.410 ;
        RECT 655.565 829.110 670.220 829.200 ;
        RECT 655.565 829.095 655.895 829.110 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 665.230 2077.300 665.550 2077.360 ;
        RECT 2898.990 2077.300 2899.310 2077.360 ;
        RECT 665.230 2077.160 2899.310 2077.300 ;
        RECT 665.230 2077.100 665.550 2077.160 ;
        RECT 2898.990 2077.100 2899.310 2077.160 ;
        RECT 665.230 839.160 665.550 839.420 ;
        RECT 665.320 838.400 665.460 839.160 ;
        RECT 665.230 838.140 665.550 838.400 ;
      LAYER via ;
        RECT 665.260 2077.100 665.520 2077.360 ;
        RECT 2899.020 2077.100 2899.280 2077.360 ;
        RECT 665.260 839.160 665.520 839.420 ;
        RECT 665.260 838.140 665.520 838.400 ;
      LAYER met2 ;
        RECT 2899.010 2082.315 2899.290 2082.685 ;
        RECT 2899.080 2077.390 2899.220 2082.315 ;
        RECT 665.260 2077.070 665.520 2077.390 ;
        RECT 2899.020 2077.070 2899.280 2077.390 ;
        RECT 665.320 839.450 665.460 2077.070 ;
        RECT 665.260 839.130 665.520 839.450 ;
        RECT 665.260 838.110 665.520 838.430 ;
        RECT 665.320 834.885 665.460 838.110 ;
        RECT 665.250 834.515 665.530 834.885 ;
      LAYER via2 ;
        RECT 2899.010 2082.360 2899.290 2082.640 ;
        RECT 665.250 834.560 665.530 834.840 ;
      LAYER met3 ;
        RECT 2898.985 2082.650 2899.315 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2898.985 2082.350 2924.800 2082.650 ;
        RECT 2898.985 2082.335 2899.315 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 665.225 834.850 665.555 834.865 ;
        RECT 670.000 834.850 674.000 835.240 ;
        RECT 665.225 834.640 674.000 834.850 ;
        RECT 665.225 834.550 670.220 834.640 ;
        RECT 665.225 834.535 665.555 834.550 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 665.690 2311.900 666.010 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 665.690 2311.760 2901.150 2311.900 ;
        RECT 665.690 2311.700 666.010 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
      LAYER via ;
        RECT 665.720 2311.700 665.980 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 665.720 2311.670 665.980 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 665.780 839.645 665.920 2311.670 ;
        RECT 665.710 839.275 665.990 839.645 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 665.710 839.320 665.990 839.600 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 665.685 839.610 666.015 839.625 ;
        RECT 670.000 839.610 674.000 840.000 ;
        RECT 665.685 839.400 674.000 839.610 ;
        RECT 665.685 839.310 670.220 839.400 ;
        RECT 665.685 839.295 666.015 839.310 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 151.540 662.330 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 662.010 151.400 2901.150 151.540 ;
        RECT 662.010 151.340 662.330 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 662.040 151.340 662.300 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 662.030 601.955 662.310 602.325 ;
        RECT 662.100 151.630 662.240 601.955 ;
        RECT 662.040 151.310 662.300 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 662.030 602.000 662.310 602.280 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 662.005 602.290 662.335 602.305 ;
        RECT 670.000 602.290 674.000 602.680 ;
        RECT 662.005 602.080 674.000 602.290 ;
        RECT 662.005 601.990 670.220 602.080 ;
        RECT 662.005 601.975 662.335 601.990 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 658.790 2491.080 659.110 2491.140 ;
        RECT 2899.450 2491.080 2899.770 2491.140 ;
        RECT 658.790 2490.940 2899.770 2491.080 ;
        RECT 658.790 2490.880 659.110 2490.940 ;
        RECT 2899.450 2490.880 2899.770 2490.940 ;
        RECT 658.790 822.160 659.110 822.420 ;
        RECT 658.880 821.400 659.020 822.160 ;
        RECT 658.790 821.140 659.110 821.400 ;
        RECT 658.790 784.760 659.110 785.020 ;
        RECT 658.880 784.000 659.020 784.760 ;
        RECT 658.790 783.740 659.110 784.000 ;
      LAYER via ;
        RECT 658.820 2490.880 659.080 2491.140 ;
        RECT 2899.480 2490.880 2899.740 2491.140 ;
        RECT 658.820 822.160 659.080 822.420 ;
        RECT 658.820 821.140 659.080 821.400 ;
        RECT 658.820 784.760 659.080 785.020 ;
        RECT 658.820 783.740 659.080 784.000 ;
      LAYER met2 ;
        RECT 2899.470 2493.035 2899.750 2493.405 ;
        RECT 2899.540 2491.170 2899.680 2493.035 ;
        RECT 658.820 2490.850 659.080 2491.170 ;
        RECT 2899.480 2490.850 2899.740 2491.170 ;
        RECT 658.880 822.450 659.020 2490.850 ;
        RECT 658.820 822.130 659.080 822.450 ;
        RECT 658.820 821.110 659.080 821.430 ;
        RECT 658.880 785.050 659.020 821.110 ;
        RECT 658.820 784.730 659.080 785.050 ;
        RECT 658.820 783.710 659.080 784.030 ;
        RECT 658.880 652.645 659.020 783.710 ;
        RECT 658.810 652.275 659.090 652.645 ;
      LAYER via2 ;
        RECT 2899.470 2493.080 2899.750 2493.360 ;
        RECT 658.810 652.320 659.090 652.600 ;
      LAYER met3 ;
        RECT 2899.445 2493.370 2899.775 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2899.445 2493.070 2924.800 2493.370 ;
        RECT 2899.445 2493.055 2899.775 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 658.785 652.610 659.115 652.625 ;
        RECT 670.000 652.610 674.000 653.000 ;
        RECT 658.785 652.400 674.000 652.610 ;
        RECT 658.785 652.310 670.220 652.400 ;
        RECT 658.785 652.295 659.115 652.310 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.030 1004.260 656.350 1004.320 ;
        RECT 2901.750 1004.260 2902.070 1004.320 ;
        RECT 656.030 1004.120 2902.070 1004.260 ;
        RECT 656.030 1004.060 656.350 1004.120 ;
        RECT 2901.750 1004.060 2902.070 1004.120 ;
        RECT 655.570 796.860 655.890 796.920 ;
        RECT 658.330 796.860 658.650 796.920 ;
        RECT 655.570 796.720 658.650 796.860 ;
        RECT 655.570 796.660 655.890 796.720 ;
        RECT 658.330 796.660 658.650 796.720 ;
        RECT 656.030 786.660 656.350 786.720 ;
        RECT 658.330 786.660 658.650 786.720 ;
        RECT 656.030 786.520 658.650 786.660 ;
        RECT 656.030 786.460 656.350 786.520 ;
        RECT 658.330 786.460 658.650 786.520 ;
      LAYER via ;
        RECT 656.060 1004.060 656.320 1004.320 ;
        RECT 2901.780 1004.060 2902.040 1004.320 ;
        RECT 655.600 796.660 655.860 796.920 ;
        RECT 658.360 796.660 658.620 796.920 ;
        RECT 656.060 786.460 656.320 786.720 ;
        RECT 658.360 786.460 658.620 786.720 ;
      LAYER met2 ;
        RECT 2901.770 2727.635 2902.050 2728.005 ;
        RECT 2901.840 1004.350 2901.980 2727.635 ;
        RECT 656.060 1004.030 656.320 1004.350 ;
        RECT 2901.780 1004.030 2902.040 1004.350 ;
        RECT 656.120 982.330 656.260 1004.030 ;
        RECT 656.120 982.190 656.720 982.330 ;
        RECT 656.580 932.125 656.720 982.190 ;
        RECT 656.510 931.755 656.790 932.125 ;
        RECT 656.050 904.555 656.330 904.925 ;
        RECT 656.120 821.000 656.260 904.555 ;
        RECT 655.660 820.860 656.260 821.000 ;
        RECT 655.660 796.950 655.800 820.860 ;
        RECT 655.600 796.630 655.860 796.950 ;
        RECT 658.360 796.630 658.620 796.950 ;
        RECT 658.420 786.750 658.560 796.630 ;
        RECT 656.060 786.430 656.320 786.750 ;
        RECT 658.360 786.430 658.620 786.750 ;
        RECT 656.120 737.530 656.260 786.430 ;
        RECT 655.660 737.390 656.260 737.530 ;
        RECT 655.660 732.090 655.800 737.390 ;
        RECT 655.660 731.950 656.260 732.090 ;
        RECT 656.120 725.290 656.260 731.950 ;
        RECT 655.200 725.150 656.260 725.290 ;
        RECT 655.200 722.570 655.340 725.150 ;
        RECT 655.200 722.430 655.800 722.570 ;
        RECT 655.660 657.405 655.800 722.430 ;
        RECT 655.590 657.035 655.870 657.405 ;
      LAYER via2 ;
        RECT 2901.770 2727.680 2902.050 2727.960 ;
        RECT 656.510 931.800 656.790 932.080 ;
        RECT 656.050 904.600 656.330 904.880 ;
        RECT 655.590 657.080 655.870 657.360 ;
      LAYER met3 ;
        RECT 2901.745 2727.970 2902.075 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2901.745 2727.670 2924.800 2727.970 ;
        RECT 2901.745 2727.655 2902.075 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 656.485 932.100 656.815 932.105 ;
        RECT 656.230 932.090 656.815 932.100 ;
        RECT 656.030 931.790 656.815 932.090 ;
        RECT 656.230 931.780 656.815 931.790 ;
        RECT 656.485 931.775 656.815 931.780 ;
        RECT 656.025 904.900 656.355 904.905 ;
        RECT 656.025 904.890 656.610 904.900 ;
        RECT 655.800 904.590 656.610 904.890 ;
        RECT 656.025 904.580 656.610 904.590 ;
        RECT 656.025 904.575 656.355 904.580 ;
        RECT 655.565 657.370 655.895 657.385 ;
        RECT 670.000 657.370 674.000 657.760 ;
        RECT 655.565 657.160 674.000 657.370 ;
        RECT 655.565 657.070 670.220 657.160 ;
        RECT 655.565 657.055 655.895 657.070 ;
      LAYER via3 ;
        RECT 656.260 931.780 656.580 932.100 ;
        RECT 656.260 904.580 656.580 904.900 ;
      LAYER met4 ;
        RECT 656.255 931.775 656.585 932.105 ;
        RECT 656.270 904.905 656.570 931.775 ;
        RECT 656.255 904.575 656.585 904.905 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 654.650 2960.280 654.970 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 654.650 2960.140 2901.150 2960.280 ;
        RECT 654.650 2960.080 654.970 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 654.680 2960.080 654.940 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 654.680 2960.050 654.940 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 654.740 662.845 654.880 2960.050 ;
        RECT 654.670 662.475 654.950 662.845 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
        RECT 654.670 662.520 654.950 662.800 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 654.645 662.810 654.975 662.825 ;
        RECT 670.000 662.810 674.000 663.200 ;
        RECT 654.645 662.600 674.000 662.810 ;
        RECT 654.645 662.510 670.220 662.600 ;
        RECT 654.645 662.495 654.975 662.510 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 659.710 3194.880 660.030 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 659.710 3194.740 2901.150 3194.880 ;
        RECT 659.710 3194.680 660.030 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 659.740 3194.680 660.000 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 659.740 3194.650 660.000 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 659.800 667.605 659.940 3194.650 ;
        RECT 659.730 667.235 660.010 667.605 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 659.730 667.280 660.010 667.560 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 659.705 667.570 660.035 667.585 ;
        RECT 670.000 667.570 674.000 667.960 ;
        RECT 659.705 667.360 674.000 667.570 ;
        RECT 659.705 667.270 670.220 667.360 ;
        RECT 659.705 667.255 660.035 667.270 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 660.170 3429.480 660.490 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 660.170 3429.340 2901.150 3429.480 ;
        RECT 660.170 3429.280 660.490 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 660.200 3429.280 660.460 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 660.200 3429.250 660.460 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 660.260 673.045 660.400 3429.250 ;
        RECT 660.190 672.675 660.470 673.045 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 660.190 672.720 660.470 673.000 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 660.165 673.010 660.495 673.025 ;
        RECT 670.000 673.010 674.000 673.400 ;
        RECT 660.165 672.800 674.000 673.010 ;
        RECT 660.165 672.710 670.220 672.800 ;
        RECT 660.165 672.695 660.495 672.710 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 3501.560 662.330 3501.620 ;
        RECT 2717.290 3501.560 2717.610 3501.620 ;
        RECT 662.010 3501.420 2717.610 3501.560 ;
        RECT 662.010 3501.360 662.330 3501.420 ;
        RECT 2717.290 3501.360 2717.610 3501.420 ;
      LAYER via ;
        RECT 662.040 3501.360 662.300 3501.620 ;
        RECT 2717.320 3501.360 2717.580 3501.620 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.650 2717.520 3517.600 ;
        RECT 662.040 3501.330 662.300 3501.650 ;
        RECT 2717.320 3501.330 2717.580 3501.650 ;
        RECT 662.100 677.805 662.240 3501.330 ;
        RECT 662.030 677.435 662.310 677.805 ;
      LAYER via2 ;
        RECT 662.030 677.480 662.310 677.760 ;
      LAYER met3 ;
        RECT 662.005 677.770 662.335 677.785 ;
        RECT 670.000 677.770 674.000 678.160 ;
        RECT 662.005 677.560 674.000 677.770 ;
        RECT 662.005 677.470 670.220 677.560 ;
        RECT 662.005 677.455 662.335 677.470 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 661.550 3502.580 661.870 3502.640 ;
        RECT 2392.530 3502.580 2392.850 3502.640 ;
        RECT 661.550 3502.440 2392.850 3502.580 ;
        RECT 661.550 3502.380 661.870 3502.440 ;
        RECT 2392.530 3502.380 2392.850 3502.440 ;
      LAYER via ;
        RECT 661.580 3502.380 661.840 3502.640 ;
        RECT 2392.560 3502.380 2392.820 3502.640 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3502.670 2392.760 3517.600 ;
        RECT 661.580 3502.350 661.840 3502.670 ;
        RECT 2392.560 3502.350 2392.820 3502.670 ;
        RECT 661.640 683.245 661.780 3502.350 ;
        RECT 661.570 682.875 661.850 683.245 ;
      LAYER via2 ;
        RECT 661.570 682.920 661.850 683.200 ;
      LAYER met3 ;
        RECT 661.545 683.210 661.875 683.225 ;
        RECT 670.000 683.210 674.000 683.600 ;
        RECT 661.545 683.000 674.000 683.210 ;
        RECT 661.545 682.910 670.220 683.000 ;
        RECT 661.545 682.895 661.875 682.910 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 661.090 3503.600 661.410 3503.660 ;
        RECT 2068.230 3503.600 2068.550 3503.660 ;
        RECT 661.090 3503.460 2068.550 3503.600 ;
        RECT 661.090 3503.400 661.410 3503.460 ;
        RECT 2068.230 3503.400 2068.550 3503.460 ;
      LAYER via ;
        RECT 661.120 3503.400 661.380 3503.660 ;
        RECT 2068.260 3503.400 2068.520 3503.660 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3503.690 2068.460 3517.600 ;
        RECT 661.120 3503.370 661.380 3503.690 ;
        RECT 2068.260 3503.370 2068.520 3503.690 ;
        RECT 661.180 688.005 661.320 3503.370 ;
        RECT 661.110 687.635 661.390 688.005 ;
      LAYER via2 ;
        RECT 661.110 687.680 661.390 687.960 ;
      LAYER met3 ;
        RECT 661.085 687.970 661.415 687.985 ;
        RECT 670.000 687.970 674.000 688.360 ;
        RECT 661.085 687.760 674.000 687.970 ;
        RECT 661.085 687.670 670.220 687.760 ;
        RECT 661.085 687.655 661.415 687.670 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 668.910 3504.620 669.230 3504.680 ;
        RECT 1743.930 3504.620 1744.250 3504.680 ;
        RECT 668.910 3504.480 1744.250 3504.620 ;
        RECT 668.910 3504.420 669.230 3504.480 ;
        RECT 1743.930 3504.420 1744.250 3504.480 ;
      LAYER via ;
        RECT 668.940 3504.420 669.200 3504.680 ;
        RECT 1743.960 3504.420 1744.220 3504.680 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3504.710 1744.160 3517.600 ;
        RECT 668.940 3504.390 669.200 3504.710 ;
        RECT 1743.960 3504.390 1744.220 3504.710 ;
        RECT 669.000 692.765 669.140 3504.390 ;
        RECT 668.930 692.395 669.210 692.765 ;
      LAYER via2 ;
        RECT 668.930 692.440 669.210 692.720 ;
      LAYER met3 ;
        RECT 668.905 692.730 669.235 692.745 ;
        RECT 670.000 692.730 674.000 693.120 ;
        RECT 668.905 692.520 674.000 692.730 ;
        RECT 668.905 692.430 670.220 692.520 ;
        RECT 668.905 692.415 669.235 692.430 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 648.210 3500.880 648.530 3500.940 ;
        RECT 1419.170 3500.880 1419.490 3500.940 ;
        RECT 648.210 3500.740 1419.490 3500.880 ;
        RECT 648.210 3500.680 648.530 3500.740 ;
        RECT 1419.170 3500.680 1419.490 3500.740 ;
        RECT 648.210 703.360 648.530 703.420 ;
        RECT 658.330 703.360 658.650 703.420 ;
        RECT 648.210 703.220 658.650 703.360 ;
        RECT 648.210 703.160 648.530 703.220 ;
        RECT 658.330 703.160 658.650 703.220 ;
      LAYER via ;
        RECT 648.240 3500.680 648.500 3500.940 ;
        RECT 1419.200 3500.680 1419.460 3500.940 ;
        RECT 648.240 703.160 648.500 703.420 ;
        RECT 658.360 703.160 658.620 703.420 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3500.970 1419.400 3517.600 ;
        RECT 648.240 3500.650 648.500 3500.970 ;
        RECT 1419.200 3500.650 1419.460 3500.970 ;
        RECT 648.300 703.450 648.440 3500.650 ;
        RECT 648.240 703.130 648.500 703.450 ;
        RECT 658.360 703.130 658.620 703.450 ;
        RECT 658.420 698.205 658.560 703.130 ;
        RECT 658.350 697.835 658.630 698.205 ;
      LAYER via2 ;
        RECT 658.350 697.880 658.630 698.160 ;
      LAYER met3 ;
        RECT 658.325 698.170 658.655 698.185 ;
        RECT 670.000 698.170 674.000 698.560 ;
        RECT 658.325 697.960 674.000 698.170 ;
        RECT 658.325 697.870 670.220 697.960 ;
        RECT 658.325 697.855 658.655 697.870 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 661.090 386.140 661.410 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 661.090 386.000 1176.520 386.140 ;
        RECT 661.090 385.940 661.410 386.000 ;
        RECT 1176.380 385.800 1176.520 386.000 ;
        RECT 1188.340 386.000 2901.150 386.140 ;
        RECT 1188.340 385.800 1188.480 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
        RECT 1176.380 385.660 1188.480 385.800 ;
      LAYER via ;
        RECT 661.120 385.940 661.380 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 661.110 606.715 661.390 607.085 ;
        RECT 661.180 386.230 661.320 606.715 ;
        RECT 661.120 385.910 661.380 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 661.110 606.760 661.390 607.040 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 661.085 607.050 661.415 607.065 ;
        RECT 670.000 607.050 674.000 607.440 ;
        RECT 661.085 606.840 674.000 607.050 ;
        RECT 661.085 606.750 670.220 606.840 ;
        RECT 661.085 606.735 661.415 606.750 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 3498.500 1069.430 3498.560 ;
        RECT 1094.870 3498.500 1095.190 3498.560 ;
        RECT 1069.110 3498.360 1095.190 3498.500 ;
        RECT 1069.110 3498.300 1069.430 3498.360 ;
        RECT 1094.870 3498.300 1095.190 3498.360 ;
        RECT 986.770 3487.960 987.090 3488.020 ;
        RECT 1069.110 3487.960 1069.430 3488.020 ;
        RECT 986.770 3487.820 1069.430 3487.960 ;
        RECT 986.770 3487.760 987.090 3487.820 ;
        RECT 1069.110 3487.760 1069.430 3487.820 ;
        RECT 935.710 3474.020 936.030 3474.080 ;
        RECT 986.770 3474.020 987.090 3474.080 ;
        RECT 935.710 3473.880 987.090 3474.020 ;
        RECT 935.710 3473.820 936.030 3473.880 ;
        RECT 986.770 3473.820 987.090 3473.880 ;
        RECT 869.010 3432.540 869.330 3432.600 ;
        RECT 935.710 3432.540 936.030 3432.600 ;
        RECT 869.010 3432.400 936.030 3432.540 ;
        RECT 869.010 3432.340 869.330 3432.400 ;
        RECT 935.710 3432.340 936.030 3432.400 ;
        RECT 851.990 3415.880 852.310 3415.940 ;
        RECT 869.010 3415.880 869.330 3415.940 ;
        RECT 851.990 3415.740 869.330 3415.880 ;
        RECT 851.990 3415.680 852.310 3415.740 ;
        RECT 869.010 3415.680 869.330 3415.740 ;
        RECT 830.830 3370.320 831.150 3370.380 ;
        RECT 851.990 3370.320 852.310 3370.380 ;
        RECT 830.830 3370.180 852.310 3370.320 ;
        RECT 830.830 3370.120 831.150 3370.180 ;
        RECT 851.990 3370.120 852.310 3370.180 ;
        RECT 819.330 3346.860 819.650 3346.920 ;
        RECT 830.830 3346.860 831.150 3346.920 ;
        RECT 819.330 3346.720 831.150 3346.860 ;
        RECT 819.330 3346.660 819.650 3346.720 ;
        RECT 830.830 3346.660 831.150 3346.720 ;
        RECT 803.690 3318.980 804.010 3319.040 ;
        RECT 819.330 3318.980 819.650 3319.040 ;
        RECT 803.690 3318.840 819.650 3318.980 ;
        RECT 803.690 3318.780 804.010 3318.840 ;
        RECT 819.330 3318.780 819.650 3318.840 ;
        RECT 755.390 3253.360 755.710 3253.420 ;
        RECT 803.690 3253.360 804.010 3253.420 ;
        RECT 755.390 3253.220 804.010 3253.360 ;
        RECT 755.390 3253.160 755.710 3253.220 ;
        RECT 803.690 3253.160 804.010 3253.220 ;
        RECT 727.790 3180.940 728.110 3181.000 ;
        RECT 755.390 3180.940 755.710 3181.000 ;
        RECT 727.790 3180.800 755.710 3180.940 ;
        RECT 727.790 3180.740 728.110 3180.800 ;
        RECT 755.390 3180.740 755.710 3180.800 ;
        RECT 703.870 3004.820 704.190 3004.880 ;
        RECT 727.790 3004.820 728.110 3004.880 ;
        RECT 703.870 3004.680 728.110 3004.820 ;
        RECT 703.870 3004.620 704.190 3004.680 ;
        RECT 727.790 3004.620 728.110 3004.680 ;
        RECT 664.770 2991.560 665.090 2991.620 ;
        RECT 703.870 2991.560 704.190 2991.620 ;
        RECT 664.770 2991.420 704.190 2991.560 ;
        RECT 664.770 2991.360 665.090 2991.420 ;
        RECT 703.870 2991.360 704.190 2991.420 ;
        RECT 658.330 2070.160 658.650 2070.220 ;
        RECT 664.770 2070.160 665.090 2070.220 ;
        RECT 658.330 2070.020 665.090 2070.160 ;
        RECT 658.330 2069.960 658.650 2070.020 ;
        RECT 664.770 2069.960 665.090 2070.020 ;
        RECT 650.510 1002.560 650.830 1002.620 ;
        RECT 658.330 1002.560 658.650 1002.620 ;
        RECT 650.510 1002.420 658.650 1002.560 ;
        RECT 650.510 1002.360 650.830 1002.420 ;
        RECT 658.330 1002.360 658.650 1002.420 ;
        RECT 650.510 703.700 650.830 703.760 ;
        RECT 656.030 703.700 656.350 703.760 ;
        RECT 650.510 703.560 656.350 703.700 ;
        RECT 650.510 703.500 650.830 703.560 ;
        RECT 656.030 703.500 656.350 703.560 ;
      LAYER via ;
        RECT 1069.140 3498.300 1069.400 3498.560 ;
        RECT 1094.900 3498.300 1095.160 3498.560 ;
        RECT 986.800 3487.760 987.060 3488.020 ;
        RECT 1069.140 3487.760 1069.400 3488.020 ;
        RECT 935.740 3473.820 936.000 3474.080 ;
        RECT 986.800 3473.820 987.060 3474.080 ;
        RECT 869.040 3432.340 869.300 3432.600 ;
        RECT 935.740 3432.340 936.000 3432.600 ;
        RECT 852.020 3415.680 852.280 3415.940 ;
        RECT 869.040 3415.680 869.300 3415.940 ;
        RECT 830.860 3370.120 831.120 3370.380 ;
        RECT 852.020 3370.120 852.280 3370.380 ;
        RECT 819.360 3346.660 819.620 3346.920 ;
        RECT 830.860 3346.660 831.120 3346.920 ;
        RECT 803.720 3318.780 803.980 3319.040 ;
        RECT 819.360 3318.780 819.620 3319.040 ;
        RECT 755.420 3253.160 755.680 3253.420 ;
        RECT 803.720 3253.160 803.980 3253.420 ;
        RECT 727.820 3180.740 728.080 3181.000 ;
        RECT 755.420 3180.740 755.680 3181.000 ;
        RECT 703.900 3004.620 704.160 3004.880 ;
        RECT 727.820 3004.620 728.080 3004.880 ;
        RECT 664.800 2991.360 665.060 2991.620 ;
        RECT 703.900 2991.360 704.160 2991.620 ;
        RECT 658.360 2069.960 658.620 2070.220 ;
        RECT 664.800 2069.960 665.060 2070.220 ;
        RECT 650.540 1002.360 650.800 1002.620 ;
        RECT 658.360 1002.360 658.620 1002.620 ;
        RECT 650.540 703.500 650.800 703.760 ;
        RECT 656.060 703.500 656.320 703.760 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3498.590 1095.100 3517.600 ;
        RECT 1069.140 3498.270 1069.400 3498.590 ;
        RECT 1094.900 3498.270 1095.160 3498.590 ;
        RECT 1069.200 3488.050 1069.340 3498.270 ;
        RECT 986.800 3487.730 987.060 3488.050 ;
        RECT 1069.140 3487.730 1069.400 3488.050 ;
        RECT 986.860 3474.110 987.000 3487.730 ;
        RECT 935.740 3473.790 936.000 3474.110 ;
        RECT 986.800 3473.790 987.060 3474.110 ;
        RECT 935.800 3432.630 935.940 3473.790 ;
        RECT 869.040 3432.310 869.300 3432.630 ;
        RECT 935.740 3432.310 936.000 3432.630 ;
        RECT 869.100 3415.970 869.240 3432.310 ;
        RECT 852.020 3415.650 852.280 3415.970 ;
        RECT 869.040 3415.650 869.300 3415.970 ;
        RECT 852.080 3370.410 852.220 3415.650 ;
        RECT 830.860 3370.090 831.120 3370.410 ;
        RECT 852.020 3370.090 852.280 3370.410 ;
        RECT 830.920 3346.950 831.060 3370.090 ;
        RECT 819.360 3346.630 819.620 3346.950 ;
        RECT 830.860 3346.630 831.120 3346.950 ;
        RECT 819.420 3319.070 819.560 3346.630 ;
        RECT 803.720 3318.750 803.980 3319.070 ;
        RECT 819.360 3318.750 819.620 3319.070 ;
        RECT 803.780 3253.450 803.920 3318.750 ;
        RECT 755.420 3253.130 755.680 3253.450 ;
        RECT 803.720 3253.130 803.980 3253.450 ;
        RECT 755.480 3181.030 755.620 3253.130 ;
        RECT 727.820 3180.710 728.080 3181.030 ;
        RECT 755.420 3180.710 755.680 3181.030 ;
        RECT 727.880 3004.910 728.020 3180.710 ;
        RECT 703.900 3004.590 704.160 3004.910 ;
        RECT 727.820 3004.590 728.080 3004.910 ;
        RECT 703.960 2991.650 704.100 3004.590 ;
        RECT 664.800 2991.330 665.060 2991.650 ;
        RECT 703.900 2991.330 704.160 2991.650 ;
        RECT 664.860 2070.250 665.000 2991.330 ;
        RECT 658.360 2069.930 658.620 2070.250 ;
        RECT 664.800 2069.930 665.060 2070.250 ;
        RECT 658.420 1002.650 658.560 2069.930 ;
        RECT 650.540 1002.330 650.800 1002.650 ;
        RECT 658.360 1002.330 658.620 1002.650 ;
        RECT 650.600 703.790 650.740 1002.330 ;
        RECT 650.540 703.470 650.800 703.790 ;
        RECT 656.060 703.470 656.320 703.790 ;
        RECT 656.120 702.965 656.260 703.470 ;
        RECT 656.050 702.595 656.330 702.965 ;
      LAYER via2 ;
        RECT 656.050 702.640 656.330 702.920 ;
      LAYER met3 ;
        RECT 656.025 702.930 656.355 702.945 ;
        RECT 670.000 702.930 674.000 703.320 ;
        RECT 656.025 702.720 674.000 702.930 ;
        RECT 656.025 702.630 670.220 702.720 ;
        RECT 656.025 702.615 656.355 702.630 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 660.630 3504.280 660.950 3504.340 ;
        RECT 770.570 3504.280 770.890 3504.340 ;
        RECT 660.630 3504.140 770.890 3504.280 ;
        RECT 660.630 3504.080 660.950 3504.140 ;
        RECT 770.570 3504.080 770.890 3504.140 ;
        RECT 660.630 737.700 660.950 737.760 ;
        RECT 660.630 737.560 661.320 737.700 ;
        RECT 660.630 737.500 660.950 737.560 ;
        RECT 658.330 736.340 658.650 736.400 ;
        RECT 661.180 736.340 661.320 737.560 ;
        RECT 658.330 736.200 661.320 736.340 ;
        RECT 658.330 736.140 658.650 736.200 ;
      LAYER via ;
        RECT 660.660 3504.080 660.920 3504.340 ;
        RECT 770.600 3504.080 770.860 3504.340 ;
        RECT 660.660 737.500 660.920 737.760 ;
        RECT 658.360 736.140 658.620 736.400 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3504.370 770.800 3517.600 ;
        RECT 660.660 3504.050 660.920 3504.370 ;
        RECT 770.600 3504.050 770.860 3504.370 ;
        RECT 660.720 737.790 660.860 3504.050 ;
        RECT 660.660 737.470 660.920 737.790 ;
        RECT 658.360 736.110 658.620 736.430 ;
        RECT 658.420 708.405 658.560 736.110 ;
        RECT 658.350 708.035 658.630 708.405 ;
      LAYER via2 ;
        RECT 658.350 708.080 658.630 708.360 ;
      LAYER met3 ;
        RECT 658.325 708.370 658.655 708.385 ;
        RECT 670.000 708.370 674.000 708.760 ;
        RECT 658.325 708.160 674.000 708.370 ;
        RECT 658.325 708.070 670.220 708.160 ;
        RECT 658.325 708.055 658.655 708.070 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 2763.420 448.430 2763.480 ;
        RECT 644.990 2763.420 645.310 2763.480 ;
        RECT 448.110 2763.280 645.310 2763.420 ;
        RECT 448.110 2763.220 448.430 2763.280 ;
        RECT 644.990 2763.220 645.310 2763.280 ;
        RECT 644.990 713.900 645.310 713.960 ;
        RECT 656.030 713.900 656.350 713.960 ;
        RECT 644.990 713.760 656.350 713.900 ;
        RECT 644.990 713.700 645.310 713.760 ;
        RECT 656.030 713.700 656.350 713.760 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 2763.220 448.400 2763.480 ;
        RECT 645.020 2763.220 645.280 2763.480 ;
        RECT 645.020 713.700 645.280 713.960 ;
        RECT 656.060 713.700 656.320 713.960 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 2763.510 448.340 3498.270 ;
        RECT 448.140 2763.190 448.400 2763.510 ;
        RECT 645.020 2763.190 645.280 2763.510 ;
        RECT 645.080 713.990 645.220 2763.190 ;
        RECT 645.020 713.670 645.280 713.990 ;
        RECT 656.060 713.670 656.320 713.990 ;
        RECT 656.120 713.165 656.260 713.670 ;
        RECT 656.050 712.795 656.330 713.165 ;
      LAYER via2 ;
        RECT 656.050 712.840 656.330 713.120 ;
      LAYER met3 ;
        RECT 656.025 713.130 656.355 713.145 ;
        RECT 670.000 713.130 674.000 713.520 ;
        RECT 656.025 712.920 674.000 713.130 ;
        RECT 656.025 712.830 670.220 712.920 ;
        RECT 656.025 712.815 656.355 712.830 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 724.100 124.130 724.160 ;
        RECT 656.030 724.100 656.350 724.160 ;
        RECT 123.810 723.960 579.900 724.100 ;
        RECT 123.810 723.900 124.130 723.960 ;
        RECT 579.760 723.760 579.900 723.960 ;
        RECT 613.340 723.960 656.350 724.100 ;
        RECT 613.340 723.760 613.480 723.960 ;
        RECT 656.030 723.900 656.350 723.960 ;
        RECT 579.760 723.620 613.480 723.760 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 723.900 124.100 724.160 ;
        RECT 656.060 723.900 656.320 724.160 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 724.190 124.040 3498.270 ;
        RECT 123.840 723.870 124.100 724.190 ;
        RECT 656.060 723.870 656.320 724.190 ;
        RECT 656.120 718.605 656.260 723.870 ;
        RECT 656.050 718.235 656.330 718.605 ;
      LAYER via2 ;
        RECT 656.050 718.280 656.330 718.560 ;
      LAYER met3 ;
        RECT 656.025 718.570 656.355 718.585 ;
        RECT 670.000 718.570 674.000 718.960 ;
        RECT 656.025 718.360 674.000 718.570 ;
        RECT 656.025 718.270 670.220 718.360 ;
        RECT 656.025 718.255 656.355 718.270 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 23.990 724.440 24.310 724.500 ;
        RECT 603.590 724.440 603.910 724.500 ;
        RECT 23.990 724.300 603.910 724.440 ;
        RECT 23.990 724.240 24.310 724.300 ;
        RECT 603.590 724.240 603.910 724.300 ;
        RECT 614.630 724.440 614.950 724.500 ;
        RECT 655.570 724.440 655.890 724.500 ;
        RECT 614.630 724.300 655.890 724.440 ;
        RECT 614.630 724.240 614.950 724.300 ;
        RECT 655.570 724.240 655.890 724.300 ;
        RECT 603.590 723.080 603.910 723.140 ;
        RECT 614.630 723.080 614.950 723.140 ;
        RECT 603.590 722.940 614.950 723.080 ;
        RECT 603.590 722.880 603.910 722.940 ;
        RECT 614.630 722.880 614.950 722.940 ;
      LAYER via ;
        RECT 24.020 724.240 24.280 724.500 ;
        RECT 603.620 724.240 603.880 724.500 ;
        RECT 614.660 724.240 614.920 724.500 ;
        RECT 655.600 724.240 655.860 724.500 ;
        RECT 603.620 722.880 603.880 723.140 ;
        RECT 614.660 722.880 614.920 723.140 ;
      LAYER met2 ;
        RECT 24.010 3339.635 24.290 3340.005 ;
        RECT 24.080 724.530 24.220 3339.635 ;
        RECT 24.020 724.210 24.280 724.530 ;
        RECT 603.620 724.210 603.880 724.530 ;
        RECT 614.660 724.210 614.920 724.530 ;
        RECT 655.600 724.210 655.860 724.530 ;
        RECT 603.680 723.170 603.820 724.210 ;
        RECT 614.720 723.170 614.860 724.210 ;
        RECT 655.660 723.365 655.800 724.210 ;
        RECT 603.620 722.850 603.880 723.170 ;
        RECT 614.660 722.850 614.920 723.170 ;
        RECT 655.590 722.995 655.870 723.365 ;
      LAYER via2 ;
        RECT 24.010 3339.680 24.290 3339.960 ;
        RECT 655.590 723.040 655.870 723.320 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 23.985 3339.970 24.315 3339.985 ;
        RECT -4.800 3339.670 24.315 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 23.985 3339.655 24.315 3339.670 ;
        RECT 655.565 723.330 655.895 723.345 ;
        RECT 670.000 723.330 674.000 723.720 ;
        RECT 655.565 723.120 674.000 723.330 ;
        RECT 655.565 723.030 670.220 723.120 ;
        RECT 655.565 723.015 655.895 723.030 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 731.240 17.870 731.300 ;
        RECT 655.570 731.240 655.890 731.300 ;
        RECT 17.550 731.100 655.890 731.240 ;
        RECT 17.550 731.040 17.870 731.100 ;
        RECT 655.570 731.040 655.890 731.100 ;
      LAYER via ;
        RECT 17.580 731.040 17.840 731.300 ;
        RECT 655.600 731.040 655.860 731.300 ;
      LAYER met2 ;
        RECT 17.570 3051.995 17.850 3052.365 ;
        RECT 17.640 731.330 17.780 3051.995 ;
        RECT 17.580 731.010 17.840 731.330 ;
        RECT 655.600 731.010 655.860 731.330 ;
        RECT 655.660 728.805 655.800 731.010 ;
        RECT 655.590 728.435 655.870 728.805 ;
      LAYER via2 ;
        RECT 17.570 3052.040 17.850 3052.320 ;
        RECT 655.590 728.480 655.870 728.760 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.545 3052.330 17.875 3052.345 ;
        RECT -4.800 3052.030 17.875 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.545 3052.015 17.875 3052.030 ;
        RECT 655.565 728.770 655.895 728.785 ;
        RECT 670.000 728.770 674.000 729.160 ;
        RECT 655.565 728.560 674.000 728.770 ;
        RECT 655.565 728.470 670.220 728.560 ;
        RECT 655.565 728.455 655.895 728.470 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 737.700 18.790 737.760 ;
        RECT 18.470 737.560 653.040 737.700 ;
        RECT 18.470 737.500 18.790 737.560 ;
        RECT 652.900 736.680 653.040 737.560 ;
        RECT 656.030 736.680 656.350 736.740 ;
        RECT 652.900 736.540 656.350 736.680 ;
        RECT 656.030 736.480 656.350 736.540 ;
      LAYER via ;
        RECT 18.500 737.500 18.760 737.760 ;
        RECT 656.060 736.480 656.320 736.740 ;
      LAYER met2 ;
        RECT 18.490 2765.035 18.770 2765.405 ;
        RECT 18.560 737.790 18.700 2765.035 ;
        RECT 18.500 737.470 18.760 737.790 ;
        RECT 656.060 736.450 656.320 736.770 ;
        RECT 656.120 733.565 656.260 736.450 ;
        RECT 656.050 733.195 656.330 733.565 ;
      LAYER via2 ;
        RECT 18.490 2765.080 18.770 2765.360 ;
        RECT 656.050 733.240 656.330 733.520 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 18.465 2765.370 18.795 2765.385 ;
        RECT -4.800 2765.070 18.795 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 18.465 2765.055 18.795 2765.070 ;
        RECT 656.025 733.530 656.355 733.545 ;
        RECT 670.000 733.530 674.000 733.920 ;
        RECT 656.025 733.320 674.000 733.530 ;
        RECT 656.025 733.230 670.220 733.320 ;
        RECT 656.025 733.215 656.355 733.230 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 738.040 19.250 738.100 ;
        RECT 655.570 738.040 655.890 738.100 ;
        RECT 18.930 737.900 655.890 738.040 ;
        RECT 18.930 737.840 19.250 737.900 ;
        RECT 655.570 737.840 655.890 737.900 ;
      LAYER via ;
        RECT 18.960 737.840 19.220 738.100 ;
        RECT 655.600 737.840 655.860 738.100 ;
      LAYER met2 ;
        RECT 18.950 2477.395 19.230 2477.765 ;
        RECT 19.020 738.130 19.160 2477.395 ;
        RECT 18.960 737.810 19.220 738.130 ;
        RECT 655.590 737.955 655.870 738.325 ;
        RECT 655.600 737.810 655.860 737.955 ;
      LAYER via2 ;
        RECT 18.950 2477.440 19.230 2477.720 ;
        RECT 655.590 738.000 655.870 738.280 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 18.925 2477.730 19.255 2477.745 ;
        RECT -4.800 2477.430 19.255 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 18.925 2477.415 19.255 2477.430 ;
        RECT 655.565 738.290 655.895 738.305 ;
        RECT 670.000 738.290 674.000 738.680 ;
        RECT 655.565 738.080 674.000 738.290 ;
        RECT 655.565 737.990 670.220 738.080 ;
        RECT 655.565 737.975 655.895 737.990 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 745.180 20.170 745.240 ;
        RECT 655.570 745.180 655.890 745.240 ;
        RECT 19.850 745.040 655.890 745.180 ;
        RECT 19.850 744.980 20.170 745.040 ;
        RECT 655.570 744.980 655.890 745.040 ;
      LAYER via ;
        RECT 19.880 744.980 20.140 745.240 ;
        RECT 655.600 744.980 655.860 745.240 ;
      LAYER met2 ;
        RECT 19.870 2189.755 20.150 2190.125 ;
        RECT 19.940 745.270 20.080 2189.755 ;
        RECT 19.880 744.950 20.140 745.270 ;
        RECT 655.600 744.950 655.860 745.270 ;
        RECT 655.660 743.765 655.800 744.950 ;
        RECT 655.590 743.395 655.870 743.765 ;
      LAYER via2 ;
        RECT 19.870 2189.800 20.150 2190.080 ;
        RECT 655.590 743.440 655.870 743.720 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 19.845 2190.090 20.175 2190.105 ;
        RECT -4.800 2189.790 20.175 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 19.845 2189.775 20.175 2189.790 ;
        RECT 655.565 743.730 655.895 743.745 ;
        RECT 670.000 743.730 674.000 744.120 ;
        RECT 655.565 743.520 674.000 743.730 ;
        RECT 655.565 743.430 670.220 743.520 ;
        RECT 655.565 743.415 655.895 743.430 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 751.980 16.950 752.040 ;
        RECT 655.570 751.980 655.890 752.040 ;
        RECT 16.630 751.840 655.890 751.980 ;
        RECT 16.630 751.780 16.950 751.840 ;
        RECT 655.570 751.780 655.890 751.840 ;
      LAYER via ;
        RECT 16.660 751.780 16.920 752.040 ;
        RECT 655.600 751.780 655.860 752.040 ;
      LAYER met2 ;
        RECT 16.650 1902.795 16.930 1903.165 ;
        RECT 16.720 752.070 16.860 1902.795 ;
        RECT 16.660 751.750 16.920 752.070 ;
        RECT 655.600 751.750 655.860 752.070 ;
        RECT 655.660 748.525 655.800 751.750 ;
        RECT 655.590 748.155 655.870 748.525 ;
      LAYER via2 ;
        RECT 16.650 1902.840 16.930 1903.120 ;
        RECT 655.590 748.200 655.870 748.480 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.625 1903.130 16.955 1903.145 ;
        RECT -4.800 1902.830 16.955 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.625 1902.815 16.955 1902.830 ;
        RECT 655.565 748.490 655.895 748.505 ;
        RECT 670.000 748.490 674.000 748.880 ;
        RECT 655.565 748.280 674.000 748.490 ;
        RECT 655.565 748.190 670.220 748.280 ;
        RECT 655.565 748.175 655.895 748.190 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2904.510 604.080 2904.830 604.140 ;
        RECT 693.380 603.940 2904.830 604.080 ;
        RECT 669.370 603.740 669.690 603.800 ;
        RECT 669.370 603.600 670.060 603.740 ;
        RECT 669.370 603.540 669.690 603.600 ;
        RECT 669.920 603.060 670.060 603.600 ;
        RECT 693.380 603.400 693.520 603.940 ;
        RECT 2904.510 603.880 2904.830 603.940 ;
        RECT 692.920 603.260 693.520 603.400 ;
        RECT 692.920 603.060 693.060 603.260 ;
        RECT 669.920 602.920 693.060 603.060 ;
      LAYER via ;
        RECT 669.400 603.540 669.660 603.800 ;
        RECT 2904.540 603.880 2904.800 604.140 ;
      LAYER met2 ;
        RECT 2904.530 615.555 2904.810 615.925 ;
        RECT 669.390 608.755 669.670 609.125 ;
        RECT 669.460 603.830 669.600 608.755 ;
        RECT 2904.600 604.170 2904.740 615.555 ;
        RECT 2904.540 603.850 2904.800 604.170 ;
        RECT 669.400 603.510 669.660 603.830 ;
      LAYER via2 ;
        RECT 2904.530 615.600 2904.810 615.880 ;
        RECT 669.390 608.800 669.670 609.080 ;
      LAYER met3 ;
        RECT 2904.505 615.890 2904.835 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2904.505 615.590 2924.800 615.890 ;
        RECT 2904.505 615.575 2904.835 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
        RECT 670.000 611.600 674.000 612.200 ;
        RECT 669.365 609.090 669.695 609.105 ;
        RECT 670.070 609.090 670.370 611.600 ;
        RECT 669.365 608.790 670.370 609.090 ;
        RECT 669.365 608.775 669.695 608.790 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 758.440 16.030 758.500 ;
        RECT 656.490 758.440 656.810 758.500 ;
        RECT 15.710 758.300 656.810 758.440 ;
        RECT 15.710 758.240 16.030 758.300 ;
        RECT 656.490 758.240 656.810 758.300 ;
      LAYER via ;
        RECT 15.740 758.240 16.000 758.500 ;
        RECT 656.520 758.240 656.780 758.500 ;
      LAYER met2 ;
        RECT 15.730 1615.155 16.010 1615.525 ;
        RECT 15.800 758.530 15.940 1615.155 ;
        RECT 15.740 758.210 16.000 758.530 ;
        RECT 656.520 758.210 656.780 758.530 ;
        RECT 656.580 753.965 656.720 758.210 ;
        RECT 656.510 753.595 656.790 753.965 ;
      LAYER via2 ;
        RECT 15.730 1615.200 16.010 1615.480 ;
        RECT 656.510 753.640 656.790 753.920 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 15.705 1615.490 16.035 1615.505 ;
        RECT -4.800 1615.190 16.035 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 15.705 1615.175 16.035 1615.190 ;
        RECT 656.485 753.930 656.815 753.945 ;
        RECT 670.000 753.930 674.000 754.320 ;
        RECT 656.485 753.720 674.000 753.930 ;
        RECT 656.485 753.630 670.220 753.720 ;
        RECT 656.485 753.615 656.815 753.630 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 758.100 15.570 758.160 ;
        RECT 655.570 758.100 655.890 758.160 ;
        RECT 15.250 757.960 655.890 758.100 ;
        RECT 15.250 757.900 15.570 757.960 ;
        RECT 655.570 757.900 655.890 757.960 ;
      LAYER via ;
        RECT 15.280 757.900 15.540 758.160 ;
        RECT 655.600 757.900 655.860 758.160 ;
      LAYER met2 ;
        RECT 15.270 1400.275 15.550 1400.645 ;
        RECT 15.340 758.190 15.480 1400.275 ;
        RECT 655.590 758.355 655.870 758.725 ;
        RECT 655.660 758.190 655.800 758.355 ;
        RECT 15.280 757.870 15.540 758.190 ;
        RECT 655.600 757.870 655.860 758.190 ;
      LAYER via2 ;
        RECT 15.270 1400.320 15.550 1400.600 ;
        RECT 655.590 758.400 655.870 758.680 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 15.245 1400.610 15.575 1400.625 ;
        RECT -4.800 1400.310 15.575 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 15.245 1400.295 15.575 1400.310 ;
        RECT 655.565 758.690 655.895 758.705 ;
        RECT 670.000 758.690 674.000 759.080 ;
        RECT 655.565 758.480 674.000 758.690 ;
        RECT 655.565 758.390 670.220 758.480 ;
        RECT 655.565 758.375 655.895 758.390 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 765.920 15.110 765.980 ;
        RECT 655.570 765.920 655.890 765.980 ;
        RECT 14.790 765.780 655.890 765.920 ;
        RECT 14.790 765.720 15.110 765.780 ;
        RECT 655.570 765.720 655.890 765.780 ;
      LAYER via ;
        RECT 14.820 765.720 15.080 765.980 ;
        RECT 655.600 765.720 655.860 765.980 ;
      LAYER met2 ;
        RECT 14.810 1184.715 15.090 1185.085 ;
        RECT 14.880 766.010 15.020 1184.715 ;
        RECT 14.820 765.690 15.080 766.010 ;
        RECT 655.600 765.690 655.860 766.010 ;
        RECT 655.660 764.165 655.800 765.690 ;
        RECT 655.590 763.795 655.870 764.165 ;
      LAYER via2 ;
        RECT 14.810 1184.760 15.090 1185.040 ;
        RECT 655.590 763.840 655.870 764.120 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 14.785 1185.050 15.115 1185.065 ;
        RECT -4.800 1184.750 15.115 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 14.785 1184.735 15.115 1184.750 ;
        RECT 655.565 764.130 655.895 764.145 ;
        RECT 670.000 764.130 674.000 764.520 ;
        RECT 655.565 763.920 674.000 764.130 ;
        RECT 655.565 763.830 670.220 763.920 ;
        RECT 655.565 763.815 655.895 763.830 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 772.720 14.650 772.780 ;
        RECT 655.570 772.720 655.890 772.780 ;
        RECT 14.330 772.580 655.890 772.720 ;
        RECT 14.330 772.520 14.650 772.580 ;
        RECT 655.570 772.520 655.890 772.580 ;
      LAYER via ;
        RECT 14.360 772.520 14.620 772.780 ;
        RECT 655.600 772.520 655.860 772.780 ;
      LAYER met2 ;
        RECT 14.350 969.155 14.630 969.525 ;
        RECT 14.420 772.810 14.560 969.155 ;
        RECT 14.360 772.490 14.620 772.810 ;
        RECT 655.600 772.490 655.860 772.810 ;
        RECT 655.660 768.925 655.800 772.490 ;
        RECT 655.590 768.555 655.870 768.925 ;
      LAYER via2 ;
        RECT 14.350 969.200 14.630 969.480 ;
        RECT 655.590 768.600 655.870 768.880 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 14.325 969.490 14.655 969.505 ;
        RECT -4.800 969.190 14.655 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 14.325 969.175 14.655 969.190 ;
        RECT 655.565 768.890 655.895 768.905 ;
        RECT 670.000 768.890 674.000 769.280 ;
        RECT 655.565 768.680 674.000 768.890 ;
        RECT 655.565 768.590 670.220 768.680 ;
        RECT 655.565 768.575 655.895 768.590 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 24.910 773.400 25.230 773.460 ;
        RECT 655.570 773.400 655.890 773.460 ;
        RECT 24.910 773.260 655.890 773.400 ;
        RECT 24.910 773.200 25.230 773.260 ;
        RECT 655.570 773.200 655.890 773.260 ;
        RECT 13.870 755.720 14.190 755.780 ;
        RECT 24.910 755.720 25.230 755.780 ;
        RECT 13.870 755.580 25.230 755.720 ;
        RECT 13.870 755.520 14.190 755.580 ;
        RECT 24.910 755.520 25.230 755.580 ;
      LAYER via ;
        RECT 24.940 773.200 25.200 773.460 ;
        RECT 655.600 773.200 655.860 773.460 ;
        RECT 13.900 755.520 14.160 755.780 ;
        RECT 24.940 755.520 25.200 755.780 ;
      LAYER met2 ;
        RECT 655.590 773.995 655.870 774.365 ;
        RECT 655.660 773.490 655.800 773.995 ;
        RECT 24.940 773.170 25.200 773.490 ;
        RECT 655.600 773.170 655.860 773.490 ;
        RECT 25.000 755.810 25.140 773.170 ;
        RECT 13.900 755.490 14.160 755.810 ;
        RECT 24.940 755.490 25.200 755.810 ;
        RECT 13.960 753.965 14.100 755.490 ;
        RECT 13.890 753.595 14.170 753.965 ;
      LAYER via2 ;
        RECT 655.590 774.040 655.870 774.320 ;
        RECT 13.890 753.640 14.170 753.920 ;
      LAYER met3 ;
        RECT 655.565 774.330 655.895 774.345 ;
        RECT 670.000 774.330 674.000 774.720 ;
        RECT 655.565 774.120 674.000 774.330 ;
        RECT 655.565 774.030 670.220 774.120 ;
        RECT 655.565 774.015 655.895 774.030 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 13.865 753.930 14.195 753.945 ;
        RECT -4.800 753.630 14.195 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 13.865 753.615 14.195 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 773.060 17.410 773.120 ;
        RECT 656.490 773.060 656.810 773.120 ;
        RECT 17.090 772.920 656.810 773.060 ;
        RECT 17.090 772.860 17.410 772.920 ;
        RECT 656.490 772.860 656.810 772.920 ;
      LAYER via ;
        RECT 17.120 772.860 17.380 773.120 ;
        RECT 656.520 772.860 656.780 773.120 ;
      LAYER met2 ;
        RECT 656.510 778.755 656.790 779.125 ;
        RECT 656.580 773.150 656.720 778.755 ;
        RECT 17.120 772.830 17.380 773.150 ;
        RECT 656.520 772.830 656.780 773.150 ;
        RECT 17.180 538.405 17.320 772.830 ;
        RECT 17.110 538.035 17.390 538.405 ;
      LAYER via2 ;
        RECT 656.510 778.800 656.790 779.080 ;
        RECT 17.110 538.080 17.390 538.360 ;
      LAYER met3 ;
        RECT 656.485 779.090 656.815 779.105 ;
        RECT 670.000 779.090 674.000 779.480 ;
        RECT 656.485 778.880 674.000 779.090 ;
        RECT 656.485 778.790 670.220 778.880 ;
        RECT 656.485 778.775 656.815 778.790 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 17.085 538.370 17.415 538.385 ;
        RECT -4.800 538.070 17.415 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 17.085 538.055 17.415 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 659.250 324.260 659.570 324.320 ;
        RECT 16.630 324.120 659.570 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 659.250 324.060 659.570 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 659.280 324.060 659.540 324.320 ;
      LAYER met2 ;
        RECT 659.270 783.515 659.550 783.885 ;
        RECT 659.340 324.350 659.480 783.515 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 659.280 324.030 659.540 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 659.270 783.560 659.550 783.840 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 659.245 783.850 659.575 783.865 ;
        RECT 670.000 783.850 674.000 784.240 ;
        RECT 659.245 783.640 674.000 783.850 ;
        RECT 659.245 783.550 670.220 783.640 ;
        RECT 659.245 783.535 659.575 783.550 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 24.450 787.000 24.770 787.060 ;
        RECT 655.570 787.000 655.890 787.060 ;
        RECT 24.450 786.860 655.890 787.000 ;
        RECT 24.450 786.800 24.770 786.860 ;
        RECT 655.570 786.800 655.890 786.860 ;
        RECT 13.870 107.340 14.190 107.400 ;
        RECT 24.450 107.340 24.770 107.400 ;
        RECT 13.870 107.200 24.770 107.340 ;
        RECT 13.870 107.140 14.190 107.200 ;
        RECT 24.450 107.140 24.770 107.200 ;
      LAYER via ;
        RECT 24.480 786.800 24.740 787.060 ;
        RECT 655.600 786.800 655.860 787.060 ;
        RECT 13.900 107.140 14.160 107.400 ;
        RECT 24.480 107.140 24.740 107.400 ;
      LAYER met2 ;
        RECT 655.590 788.955 655.870 789.325 ;
        RECT 655.660 787.090 655.800 788.955 ;
        RECT 24.480 786.770 24.740 787.090 ;
        RECT 655.600 786.770 655.860 787.090 ;
        RECT 24.540 107.430 24.680 786.770 ;
        RECT 13.900 107.285 14.160 107.430 ;
        RECT 13.890 106.915 14.170 107.285 ;
        RECT 24.480 107.110 24.740 107.430 ;
      LAYER via2 ;
        RECT 655.590 789.000 655.870 789.280 ;
        RECT 13.890 106.960 14.170 107.240 ;
      LAYER met3 ;
        RECT 655.565 789.290 655.895 789.305 ;
        RECT 670.000 789.290 674.000 789.680 ;
        RECT 655.565 789.080 674.000 789.290 ;
        RECT 655.565 788.990 670.220 789.080 ;
        RECT 655.565 788.975 655.895 788.990 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 13.865 107.250 14.195 107.265 ;
        RECT -4.800 106.950 14.195 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 13.865 106.935 14.195 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2901.750 603.740 2902.070 603.800 ;
        RECT 694.300 603.600 2902.070 603.740 ;
        RECT 668.910 602.040 669.230 602.100 ;
        RECT 694.300 602.040 694.440 603.600 ;
        RECT 2901.750 603.540 2902.070 603.600 ;
        RECT 668.910 601.900 694.440 602.040 ;
        RECT 668.910 601.840 669.230 601.900 ;
      LAYER via ;
        RECT 668.940 601.840 669.200 602.100 ;
        RECT 2901.780 603.540 2902.040 603.800 ;
      LAYER met2 ;
        RECT 2901.770 850.155 2902.050 850.525 ;
        RECT 668.930 614.195 669.210 614.565 ;
        RECT 669.000 602.130 669.140 614.195 ;
        RECT 2901.840 603.830 2901.980 850.155 ;
        RECT 2901.780 603.510 2902.040 603.830 ;
        RECT 668.940 601.810 669.200 602.130 ;
      LAYER via2 ;
        RECT 2901.770 850.200 2902.050 850.480 ;
        RECT 668.930 614.240 669.210 614.520 ;
      LAYER met3 ;
        RECT 2901.745 850.490 2902.075 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2901.745 850.190 2924.800 850.490 ;
        RECT 2901.745 850.175 2902.075 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT 670.000 617.040 674.000 617.640 ;
        RECT 668.905 614.530 669.235 614.545 ;
        RECT 670.070 614.530 670.370 617.040 ;
        RECT 668.905 614.230 670.370 614.530 ;
        RECT 668.905 614.215 669.235 614.230 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 663.850 1083.480 664.170 1083.540 ;
        RECT 2899.910 1083.480 2900.230 1083.540 ;
        RECT 663.850 1083.340 2900.230 1083.480 ;
        RECT 663.850 1083.280 664.170 1083.340 ;
        RECT 2899.910 1083.280 2900.230 1083.340 ;
      LAYER via ;
        RECT 663.880 1083.280 664.140 1083.540 ;
        RECT 2899.940 1083.280 2900.200 1083.540 ;
      LAYER met2 ;
        RECT 2899.930 1084.755 2900.210 1085.125 ;
        RECT 2900.000 1083.570 2900.140 1084.755 ;
        RECT 663.880 1083.250 664.140 1083.570 ;
        RECT 2899.940 1083.250 2900.200 1083.570 ;
        RECT 663.940 622.045 664.080 1083.250 ;
        RECT 663.870 621.675 664.150 622.045 ;
      LAYER via2 ;
        RECT 2899.930 1084.800 2900.210 1085.080 ;
        RECT 663.870 621.720 664.150 622.000 ;
      LAYER met3 ;
        RECT 2899.905 1085.090 2900.235 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2899.905 1084.790 2924.800 1085.090 ;
        RECT 2899.905 1084.775 2900.235 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
        RECT 663.845 622.010 664.175 622.025 ;
        RECT 670.000 622.010 674.000 622.400 ;
        RECT 663.845 621.800 674.000 622.010 ;
        RECT 663.845 621.710 670.220 621.800 ;
        RECT 663.845 621.695 664.175 621.710 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 657.410 1318.080 657.730 1318.140 ;
        RECT 2898.990 1318.080 2899.310 1318.140 ;
        RECT 657.410 1317.940 2899.310 1318.080 ;
        RECT 657.410 1317.880 657.730 1317.940 ;
        RECT 2898.990 1317.880 2899.310 1317.940 ;
      LAYER via ;
        RECT 657.440 1317.880 657.700 1318.140 ;
        RECT 2899.020 1317.880 2899.280 1318.140 ;
      LAYER met2 ;
        RECT 2899.010 1319.355 2899.290 1319.725 ;
        RECT 2899.080 1318.170 2899.220 1319.355 ;
        RECT 657.440 1317.850 657.700 1318.170 ;
        RECT 2899.020 1317.850 2899.280 1318.170 ;
        RECT 657.500 627.485 657.640 1317.850 ;
        RECT 657.430 627.115 657.710 627.485 ;
      LAYER via2 ;
        RECT 2899.010 1319.400 2899.290 1319.680 ;
        RECT 657.430 627.160 657.710 627.440 ;
      LAYER met3 ;
        RECT 2898.985 1319.690 2899.315 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2898.985 1319.390 2924.800 1319.690 ;
        RECT 2898.985 1319.375 2899.315 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 657.405 627.450 657.735 627.465 ;
        RECT 670.000 627.450 674.000 627.840 ;
        RECT 657.405 627.240 674.000 627.450 ;
        RECT 657.405 627.150 670.220 627.240 ;
        RECT 657.405 627.135 657.735 627.150 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 657.870 1552.680 658.190 1552.740 ;
        RECT 2900.370 1552.680 2900.690 1552.740 ;
        RECT 657.870 1552.540 2900.690 1552.680 ;
        RECT 657.870 1552.480 658.190 1552.540 ;
        RECT 2900.370 1552.480 2900.690 1552.540 ;
      LAYER via ;
        RECT 657.900 1552.480 658.160 1552.740 ;
        RECT 2900.400 1552.480 2900.660 1552.740 ;
      LAYER met2 ;
        RECT 2900.390 1553.955 2900.670 1554.325 ;
        RECT 2900.460 1552.770 2900.600 1553.955 ;
        RECT 657.900 1552.450 658.160 1552.770 ;
        RECT 2900.400 1552.450 2900.660 1552.770 ;
        RECT 657.960 632.245 658.100 1552.450 ;
        RECT 657.890 631.875 658.170 632.245 ;
      LAYER via2 ;
        RECT 2900.390 1554.000 2900.670 1554.280 ;
        RECT 657.890 631.920 658.170 632.200 ;
      LAYER met3 ;
        RECT 2900.365 1554.290 2900.695 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.365 1553.990 2924.800 1554.290 ;
        RECT 2900.365 1553.975 2900.695 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 657.865 632.210 658.195 632.225 ;
        RECT 670.000 632.210 674.000 632.600 ;
        RECT 657.865 632.000 674.000 632.210 ;
        RECT 657.865 631.910 670.220 632.000 ;
        RECT 657.865 631.895 658.195 631.910 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 1004.600 657.270 1004.660 ;
        RECT 2900.830 1004.600 2901.150 1004.660 ;
        RECT 656.950 1004.460 2901.150 1004.600 ;
        RECT 656.950 1004.400 657.270 1004.460 ;
        RECT 2900.830 1004.400 2901.150 1004.460 ;
        RECT 658.330 737.020 658.650 737.080 ;
        RECT 660.630 737.020 660.950 737.080 ;
        RECT 658.330 736.880 660.950 737.020 ;
        RECT 658.330 736.820 658.650 736.880 ;
        RECT 660.630 736.820 660.950 736.880 ;
        RECT 658.330 665.960 658.650 666.020 ;
        RECT 660.630 665.960 660.950 666.020 ;
        RECT 658.330 665.820 660.950 665.960 ;
        RECT 658.330 665.760 658.650 665.820 ;
        RECT 660.630 665.760 660.950 665.820 ;
      LAYER via ;
        RECT 656.980 1004.400 657.240 1004.660 ;
        RECT 2900.860 1004.400 2901.120 1004.660 ;
        RECT 658.360 736.820 658.620 737.080 ;
        RECT 660.660 736.820 660.920 737.080 ;
        RECT 658.360 665.760 658.620 666.020 ;
        RECT 660.660 665.760 660.920 666.020 ;
      LAYER met2 ;
        RECT 2900.850 1789.235 2901.130 1789.605 ;
        RECT 2900.920 1004.690 2901.060 1789.235 ;
        RECT 656.980 1004.370 657.240 1004.690 ;
        RECT 2900.860 1004.370 2901.120 1004.690 ;
        RECT 657.040 983.805 657.180 1004.370 ;
        RECT 656.970 983.435 657.250 983.805 ;
        RECT 658.350 978.675 658.630 979.045 ;
        RECT 658.420 903.565 658.560 978.675 ;
        RECT 658.350 903.195 658.630 903.565 ;
        RECT 658.350 882.795 658.630 883.165 ;
        RECT 658.420 821.850 658.560 882.795 ;
        RECT 658.420 821.710 659.480 821.850 ;
        RECT 659.340 784.450 659.480 821.710 ;
        RECT 658.420 784.310 659.480 784.450 ;
        RECT 658.420 737.110 658.560 784.310 ;
        RECT 658.360 736.790 658.620 737.110 ;
        RECT 660.660 736.790 660.920 737.110 ;
        RECT 660.720 666.050 660.860 736.790 ;
        RECT 658.360 665.730 658.620 666.050 ;
        RECT 660.660 665.730 660.920 666.050 ;
        RECT 658.420 637.685 658.560 665.730 ;
        RECT 658.350 637.315 658.630 637.685 ;
      LAYER via2 ;
        RECT 2900.850 1789.280 2901.130 1789.560 ;
        RECT 656.970 983.480 657.250 983.760 ;
        RECT 658.350 978.720 658.630 979.000 ;
        RECT 658.350 903.240 658.630 903.520 ;
        RECT 658.350 882.840 658.630 883.120 ;
        RECT 658.350 637.360 658.630 637.640 ;
      LAYER met3 ;
        RECT 2900.825 1789.570 2901.155 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.825 1789.270 2924.800 1789.570 ;
        RECT 2900.825 1789.255 2901.155 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 656.945 983.770 657.275 983.785 ;
        RECT 658.070 983.770 658.450 983.780 ;
        RECT 656.945 983.470 658.450 983.770 ;
        RECT 656.945 983.455 657.275 983.470 ;
        RECT 658.070 983.460 658.450 983.470 ;
        RECT 658.325 979.020 658.655 979.025 ;
        RECT 658.070 979.010 658.655 979.020 ;
        RECT 657.870 978.710 658.655 979.010 ;
        RECT 658.070 978.700 658.655 978.710 ;
        RECT 658.325 978.695 658.655 978.700 ;
        RECT 658.325 903.540 658.655 903.545 ;
        RECT 658.070 903.530 658.655 903.540 ;
        RECT 657.870 903.230 658.655 903.530 ;
        RECT 658.070 903.220 658.655 903.230 ;
        RECT 658.325 903.215 658.655 903.220 ;
        RECT 658.325 883.140 658.655 883.145 ;
        RECT 658.070 883.130 658.655 883.140 ;
        RECT 657.870 882.830 658.655 883.130 ;
        RECT 658.070 882.820 658.655 882.830 ;
        RECT 658.325 882.815 658.655 882.820 ;
        RECT 658.325 637.650 658.655 637.665 ;
        RECT 670.000 637.650 674.000 638.040 ;
        RECT 658.325 637.440 674.000 637.650 ;
        RECT 658.325 637.350 670.220 637.440 ;
        RECT 658.325 637.335 658.655 637.350 ;
      LAYER via3 ;
        RECT 658.100 983.460 658.420 983.780 ;
        RECT 658.100 978.700 658.420 979.020 ;
        RECT 658.100 903.220 658.420 903.540 ;
        RECT 658.100 882.820 658.420 883.140 ;
      LAYER met4 ;
        RECT 658.095 983.455 658.425 983.785 ;
        RECT 658.110 979.025 658.410 983.455 ;
        RECT 658.095 978.695 658.425 979.025 ;
        RECT 658.095 903.215 658.425 903.545 ;
        RECT 658.110 883.145 658.410 903.215 ;
        RECT 658.095 882.815 658.425 883.145 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.490 1003.920 656.810 1003.980 ;
        RECT 2903.590 1003.920 2903.910 1003.980 ;
        RECT 656.490 1003.780 2903.910 1003.920 ;
        RECT 656.490 1003.720 656.810 1003.780 ;
        RECT 2903.590 1003.720 2903.910 1003.780 ;
        RECT 655.110 787.340 655.430 787.400 ;
        RECT 656.950 787.340 657.270 787.400 ;
        RECT 655.110 787.200 657.270 787.340 ;
        RECT 655.110 787.140 655.430 787.200 ;
        RECT 656.950 787.140 657.270 787.200 ;
        RECT 655.570 774.760 655.890 774.820 ;
        RECT 656.950 774.760 657.270 774.820 ;
        RECT 655.570 774.620 657.270 774.760 ;
        RECT 655.570 774.560 655.890 774.620 ;
        RECT 656.950 774.560 657.270 774.620 ;
        RECT 656.950 738.040 657.270 738.100 ;
        RECT 656.580 737.900 657.270 738.040 ;
        RECT 653.270 737.360 653.590 737.420 ;
        RECT 656.580 737.360 656.720 737.900 ;
        RECT 656.950 737.840 657.270 737.900 ;
        RECT 653.270 737.220 656.720 737.360 ;
        RECT 653.270 737.160 653.590 737.220 ;
        RECT 653.270 714.240 653.590 714.300 ;
        RECT 656.490 714.240 656.810 714.300 ;
        RECT 653.270 714.100 656.810 714.240 ;
        RECT 653.270 714.040 653.590 714.100 ;
        RECT 656.490 714.040 656.810 714.100 ;
      LAYER via ;
        RECT 656.520 1003.720 656.780 1003.980 ;
        RECT 2903.620 1003.720 2903.880 1003.980 ;
        RECT 655.140 787.140 655.400 787.400 ;
        RECT 656.980 787.140 657.240 787.400 ;
        RECT 655.600 774.560 655.860 774.820 ;
        RECT 656.980 774.560 657.240 774.820 ;
        RECT 653.300 737.160 653.560 737.420 ;
        RECT 656.980 737.840 657.240 738.100 ;
        RECT 653.300 714.040 653.560 714.300 ;
        RECT 656.520 714.040 656.780 714.300 ;
      LAYER met2 ;
        RECT 2903.610 2023.835 2903.890 2024.205 ;
        RECT 2903.680 1004.010 2903.820 2023.835 ;
        RECT 656.520 1003.690 656.780 1004.010 ;
        RECT 2903.620 1003.690 2903.880 1004.010 ;
        RECT 656.580 983.010 656.720 1003.690 ;
        RECT 656.580 982.870 657.180 983.010 ;
        RECT 657.040 903.565 657.180 982.870 ;
        RECT 656.970 903.195 657.250 903.565 ;
        RECT 656.970 882.795 657.250 883.165 ;
        RECT 657.040 787.430 657.180 882.795 ;
        RECT 655.140 787.110 655.400 787.430 ;
        RECT 656.980 787.110 657.240 787.430 ;
        RECT 655.200 786.490 655.340 787.110 ;
        RECT 655.200 786.350 655.800 786.490 ;
        RECT 655.660 774.850 655.800 786.350 ;
        RECT 655.600 774.530 655.860 774.850 ;
        RECT 656.980 774.530 657.240 774.850 ;
        RECT 657.040 738.130 657.180 774.530 ;
        RECT 656.980 737.810 657.240 738.130 ;
        RECT 653.300 737.130 653.560 737.450 ;
        RECT 653.360 714.330 653.500 737.130 ;
        RECT 653.300 714.010 653.560 714.330 ;
        RECT 656.520 714.010 656.780 714.330 ;
        RECT 656.580 702.170 656.720 714.010 ;
        RECT 656.120 702.030 656.720 702.170 ;
        RECT 656.120 642.445 656.260 702.030 ;
        RECT 656.050 642.075 656.330 642.445 ;
      LAYER via2 ;
        RECT 2903.610 2023.880 2903.890 2024.160 ;
        RECT 656.970 903.240 657.250 903.520 ;
        RECT 656.970 882.840 657.250 883.120 ;
        RECT 656.050 642.120 656.330 642.400 ;
      LAYER met3 ;
        RECT 2903.585 2024.170 2903.915 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2903.585 2023.870 2924.800 2024.170 ;
        RECT 2903.585 2023.855 2903.915 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 656.945 903.540 657.275 903.545 ;
        RECT 656.945 903.530 657.530 903.540 ;
        RECT 656.720 903.230 657.530 903.530 ;
        RECT 656.945 903.220 657.530 903.230 ;
        RECT 656.945 903.215 657.275 903.220 ;
        RECT 656.945 883.140 657.275 883.145 ;
        RECT 656.945 883.130 657.530 883.140 ;
        RECT 656.720 882.830 657.530 883.130 ;
        RECT 656.945 882.820 657.530 882.830 ;
        RECT 656.945 882.815 657.275 882.820 ;
        RECT 656.025 642.410 656.355 642.425 ;
        RECT 670.000 642.410 674.000 642.800 ;
        RECT 656.025 642.200 674.000 642.410 ;
        RECT 656.025 642.110 670.220 642.200 ;
        RECT 656.025 642.095 656.355 642.110 ;
      LAYER via3 ;
        RECT 657.180 903.220 657.500 903.540 ;
        RECT 657.180 882.820 657.500 883.140 ;
      LAYER met4 ;
        RECT 657.175 903.215 657.505 903.545 ;
        RECT 657.190 883.145 657.490 903.215 ;
        RECT 657.175 882.815 657.505 883.145 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 669.370 2256.480 669.690 2256.540 ;
        RECT 2899.450 2256.480 2899.770 2256.540 ;
        RECT 669.370 2256.340 2899.770 2256.480 ;
        RECT 669.370 2256.280 669.690 2256.340 ;
        RECT 2899.450 2256.280 2899.770 2256.340 ;
        RECT 666.150 738.040 666.470 738.100 ;
        RECT 669.370 738.040 669.690 738.100 ;
        RECT 666.150 737.900 669.690 738.040 ;
        RECT 666.150 737.840 666.470 737.900 ;
        RECT 669.370 737.840 669.690 737.900 ;
      LAYER via ;
        RECT 669.400 2256.280 669.660 2256.540 ;
        RECT 2899.480 2256.280 2899.740 2256.540 ;
        RECT 666.180 737.840 666.440 738.100 ;
        RECT 669.400 737.840 669.660 738.100 ;
      LAYER met2 ;
        RECT 2899.470 2258.435 2899.750 2258.805 ;
        RECT 2899.540 2256.570 2899.680 2258.435 ;
        RECT 669.400 2256.250 669.660 2256.570 ;
        RECT 2899.480 2256.250 2899.740 2256.570 ;
        RECT 669.460 738.130 669.600 2256.250 ;
        RECT 666.180 737.810 666.440 738.130 ;
        RECT 669.400 737.810 669.660 738.130 ;
        RECT 666.240 648.565 666.380 737.810 ;
        RECT 666.170 648.195 666.450 648.565 ;
      LAYER via2 ;
        RECT 2899.470 2258.480 2899.750 2258.760 ;
        RECT 666.170 648.240 666.450 648.520 ;
      LAYER met3 ;
        RECT 2899.445 2258.770 2899.775 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2899.445 2258.470 2924.800 2258.770 ;
        RECT 2899.445 2258.455 2899.775 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 666.145 648.530 666.475 648.545 ;
        RECT 666.145 648.230 670.370 648.530 ;
        RECT 666.145 648.215 666.475 648.230 ;
        RECT 670.070 647.560 670.370 648.230 ;
        RECT 670.000 646.960 674.000 647.560 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 993.670 367.920 993.990 368.180 ;
        RECT 993.760 366.140 993.900 367.920 ;
        RECT 993.670 365.880 993.990 366.140 ;
        RECT 633.030 36.960 633.350 37.020 ;
        RECT 993.670 36.960 993.990 37.020 ;
        RECT 633.030 36.820 993.990 36.960 ;
        RECT 633.030 36.760 633.350 36.820 ;
        RECT 993.670 36.760 993.990 36.820 ;
      LAYER via ;
        RECT 993.700 367.920 993.960 368.180 ;
        RECT 993.700 365.880 993.960 366.140 ;
        RECT 633.060 36.760 633.320 37.020 ;
        RECT 993.700 36.760 993.960 37.020 ;
      LAYER met2 ;
        RECT 995.310 600.170 995.590 604.000 ;
        RECT 993.760 600.030 995.590 600.170 ;
        RECT 993.760 368.210 993.900 600.030 ;
        RECT 995.310 600.000 995.590 600.030 ;
        RECT 993.700 367.890 993.960 368.210 ;
        RECT 993.700 365.850 993.960 366.170 ;
        RECT 993.760 37.050 993.900 365.850 ;
        RECT 633.060 36.730 633.320 37.050 ;
        RECT 993.700 36.730 993.960 37.050 ;
        RECT 633.120 2.400 633.260 36.730 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1913.210 587.080 1913.530 587.140 ;
        RECT 1917.350 587.080 1917.670 587.140 ;
        RECT 1913.210 586.940 1917.670 587.080 ;
        RECT 1913.210 586.880 1913.530 586.940 ;
        RECT 1917.350 586.880 1917.670 586.940 ;
        RECT 1917.350 36.620 1917.670 36.680 ;
        RECT 2417.370 36.620 2417.690 36.680 ;
        RECT 1917.350 36.480 2417.690 36.620 ;
        RECT 1917.350 36.420 1917.670 36.480 ;
        RECT 2417.370 36.420 2417.690 36.480 ;
      LAYER via ;
        RECT 1913.240 586.880 1913.500 587.140 ;
        RECT 1917.380 586.880 1917.640 587.140 ;
        RECT 1917.380 36.420 1917.640 36.680 ;
        RECT 2417.400 36.420 2417.660 36.680 ;
      LAYER met2 ;
        RECT 1911.630 600.170 1911.910 604.000 ;
        RECT 1911.630 600.030 1913.440 600.170 ;
        RECT 1911.630 600.000 1911.910 600.030 ;
        RECT 1913.300 587.170 1913.440 600.030 ;
        RECT 1913.240 586.850 1913.500 587.170 ;
        RECT 1917.380 586.850 1917.640 587.170 ;
        RECT 1917.440 36.710 1917.580 586.850 ;
        RECT 1917.380 36.390 1917.640 36.710 ;
        RECT 2417.400 36.390 2417.660 36.710 ;
        RECT 2417.460 2.400 2417.600 36.390 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1923.330 462.640 1923.650 462.700 ;
        RECT 1923.790 462.640 1924.110 462.700 ;
        RECT 1923.330 462.500 1924.110 462.640 ;
        RECT 1923.330 462.440 1923.650 462.500 ;
        RECT 1923.790 462.440 1924.110 462.500 ;
        RECT 1922.410 414.020 1922.730 414.080 ;
        RECT 1923.330 414.020 1923.650 414.080 ;
        RECT 1922.410 413.880 1923.650 414.020 ;
        RECT 1922.410 413.820 1922.730 413.880 ;
        RECT 1923.330 413.820 1923.650 413.880 ;
        RECT 1921.950 366.080 1922.270 366.140 ;
        RECT 1922.410 366.080 1922.730 366.140 ;
        RECT 1921.950 365.940 1922.730 366.080 ;
        RECT 1921.950 365.880 1922.270 365.940 ;
        RECT 1922.410 365.880 1922.730 365.940 ;
        RECT 1921.950 324.260 1922.270 324.320 ;
        RECT 1922.870 324.260 1923.190 324.320 ;
        RECT 1921.950 324.120 1923.190 324.260 ;
        RECT 1921.950 324.060 1922.270 324.120 ;
        RECT 1922.870 324.060 1923.190 324.120 ;
        RECT 1921.950 276.320 1922.270 276.380 ;
        RECT 1924.250 276.320 1924.570 276.380 ;
        RECT 1921.950 276.180 1924.570 276.320 ;
        RECT 1921.950 276.120 1922.270 276.180 ;
        RECT 1924.250 276.120 1924.570 276.180 ;
        RECT 1921.950 227.700 1922.270 227.760 ;
        RECT 1922.870 227.700 1923.190 227.760 ;
        RECT 1921.950 227.560 1923.190 227.700 ;
        RECT 1921.950 227.500 1922.270 227.560 ;
        RECT 1922.870 227.500 1923.190 227.560 ;
        RECT 1921.950 179.760 1922.270 179.820 ;
        RECT 1923.330 179.760 1923.650 179.820 ;
        RECT 1921.950 179.620 1923.650 179.760 ;
        RECT 1921.950 179.560 1922.270 179.620 ;
        RECT 1923.330 179.560 1923.650 179.620 ;
        RECT 1923.330 158.680 1923.650 158.740 ;
        RECT 1924.250 158.680 1924.570 158.740 ;
        RECT 1923.330 158.540 1924.570 158.680 ;
        RECT 1923.330 158.480 1923.650 158.540 ;
        RECT 1924.250 158.480 1924.570 158.540 ;
        RECT 1923.330 96.800 1923.650 96.860 ;
        RECT 1923.790 96.800 1924.110 96.860 ;
        RECT 1923.330 96.660 1924.110 96.800 ;
        RECT 1923.330 96.600 1923.650 96.660 ;
        RECT 1923.790 96.600 1924.110 96.660 ;
        RECT 1922.410 96.120 1922.730 96.180 ;
        RECT 1923.790 96.120 1924.110 96.180 ;
        RECT 1922.410 95.980 1924.110 96.120 ;
        RECT 1922.410 95.920 1922.730 95.980 ;
        RECT 1923.790 95.920 1924.110 95.980 ;
        RECT 1922.410 48.520 1922.730 48.580 ;
        RECT 1924.250 48.520 1924.570 48.580 ;
        RECT 1922.410 48.380 1924.570 48.520 ;
        RECT 1922.410 48.320 1922.730 48.380 ;
        RECT 1924.250 48.320 1924.570 48.380 ;
        RECT 1924.250 36.960 1924.570 37.020 ;
        RECT 2434.850 36.960 2435.170 37.020 ;
        RECT 1924.250 36.820 2435.170 36.960 ;
        RECT 1924.250 36.760 1924.570 36.820 ;
        RECT 2434.850 36.760 2435.170 36.820 ;
      LAYER via ;
        RECT 1923.360 462.440 1923.620 462.700 ;
        RECT 1923.820 462.440 1924.080 462.700 ;
        RECT 1922.440 413.820 1922.700 414.080 ;
        RECT 1923.360 413.820 1923.620 414.080 ;
        RECT 1921.980 365.880 1922.240 366.140 ;
        RECT 1922.440 365.880 1922.700 366.140 ;
        RECT 1921.980 324.060 1922.240 324.320 ;
        RECT 1922.900 324.060 1923.160 324.320 ;
        RECT 1921.980 276.120 1922.240 276.380 ;
        RECT 1924.280 276.120 1924.540 276.380 ;
        RECT 1921.980 227.500 1922.240 227.760 ;
        RECT 1922.900 227.500 1923.160 227.760 ;
        RECT 1921.980 179.560 1922.240 179.820 ;
        RECT 1923.360 179.560 1923.620 179.820 ;
        RECT 1923.360 158.480 1923.620 158.740 ;
        RECT 1924.280 158.480 1924.540 158.740 ;
        RECT 1923.360 96.600 1923.620 96.860 ;
        RECT 1923.820 96.600 1924.080 96.860 ;
        RECT 1922.440 95.920 1922.700 96.180 ;
        RECT 1923.820 95.920 1924.080 96.180 ;
        RECT 1922.440 48.320 1922.700 48.580 ;
        RECT 1924.280 48.320 1924.540 48.580 ;
        RECT 1924.280 36.760 1924.540 37.020 ;
        RECT 2434.880 36.760 2435.140 37.020 ;
      LAYER met2 ;
        RECT 1920.830 600.170 1921.110 604.000 ;
        RECT 1920.830 600.030 1923.100 600.170 ;
        RECT 1920.830 600.000 1921.110 600.030 ;
        RECT 1922.960 555.970 1923.100 600.030 ;
        RECT 1922.960 555.830 1924.020 555.970 ;
        RECT 1923.880 462.730 1924.020 555.830 ;
        RECT 1923.360 462.410 1923.620 462.730 ;
        RECT 1923.820 462.410 1924.080 462.730 ;
        RECT 1923.420 414.110 1923.560 462.410 ;
        RECT 1922.440 413.790 1922.700 414.110 ;
        RECT 1923.360 413.790 1923.620 414.110 ;
        RECT 1922.500 366.170 1922.640 413.790 ;
        RECT 1921.980 365.850 1922.240 366.170 ;
        RECT 1922.440 365.850 1922.700 366.170 ;
        RECT 1922.040 324.885 1922.180 365.850 ;
        RECT 1921.970 324.515 1922.250 324.885 ;
        RECT 1922.890 324.515 1923.170 324.885 ;
        RECT 1922.960 324.350 1923.100 324.515 ;
        RECT 1921.980 324.030 1922.240 324.350 ;
        RECT 1922.900 324.030 1923.160 324.350 ;
        RECT 1922.040 276.410 1922.180 324.030 ;
        RECT 1921.980 276.090 1922.240 276.410 ;
        RECT 1924.280 276.090 1924.540 276.410 ;
        RECT 1924.340 235.010 1924.480 276.090 ;
        RECT 1922.960 234.870 1924.480 235.010 ;
        RECT 1922.960 227.790 1923.100 234.870 ;
        RECT 1921.980 227.470 1922.240 227.790 ;
        RECT 1922.900 227.470 1923.160 227.790 ;
        RECT 1922.040 179.850 1922.180 227.470 ;
        RECT 1921.980 179.530 1922.240 179.850 ;
        RECT 1923.360 179.530 1923.620 179.850 ;
        RECT 1923.420 158.770 1923.560 179.530 ;
        RECT 1923.360 158.450 1923.620 158.770 ;
        RECT 1924.280 158.450 1924.540 158.770 ;
        RECT 1924.340 120.770 1924.480 158.450 ;
        RECT 1923.420 120.630 1924.480 120.770 ;
        RECT 1923.420 96.890 1923.560 120.630 ;
        RECT 1923.360 96.570 1923.620 96.890 ;
        RECT 1923.820 96.570 1924.080 96.890 ;
        RECT 1923.880 96.210 1924.020 96.570 ;
        RECT 1922.440 95.890 1922.700 96.210 ;
        RECT 1923.820 95.890 1924.080 96.210 ;
        RECT 1922.500 48.610 1922.640 95.890 ;
        RECT 1922.440 48.290 1922.700 48.610 ;
        RECT 1924.280 48.290 1924.540 48.610 ;
        RECT 1924.340 37.050 1924.480 48.290 ;
        RECT 1924.280 36.730 1924.540 37.050 ;
        RECT 2434.880 36.730 2435.140 37.050 ;
        RECT 2434.940 2.400 2435.080 36.730 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
      LAYER via2 ;
        RECT 1921.970 324.560 1922.250 324.840 ;
        RECT 1922.890 324.560 1923.170 324.840 ;
      LAYER met3 ;
        RECT 1921.945 324.850 1922.275 324.865 ;
        RECT 1922.865 324.850 1923.195 324.865 ;
        RECT 1921.945 324.550 1923.195 324.850 ;
        RECT 1921.945 324.535 1922.275 324.550 ;
        RECT 1922.865 324.535 1923.195 324.550 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1931.610 37.300 1931.930 37.360 ;
        RECT 2452.790 37.300 2453.110 37.360 ;
        RECT 1931.610 37.160 2453.110 37.300 ;
        RECT 1931.610 37.100 1931.930 37.160 ;
        RECT 2452.790 37.100 2453.110 37.160 ;
      LAYER via ;
        RECT 1931.640 37.100 1931.900 37.360 ;
        RECT 2452.820 37.100 2453.080 37.360 ;
      LAYER met2 ;
        RECT 1930.030 600.170 1930.310 604.000 ;
        RECT 1930.030 600.030 1931.840 600.170 ;
        RECT 1930.030 600.000 1930.310 600.030 ;
        RECT 1931.700 37.390 1931.840 600.030 ;
        RECT 1931.640 37.070 1931.900 37.390 ;
        RECT 2452.820 37.070 2453.080 37.390 ;
        RECT 2452.880 2.400 2453.020 37.070 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1940.810 587.080 1941.130 587.140 ;
        RECT 1944.950 587.080 1945.270 587.140 ;
        RECT 1940.810 586.940 1945.270 587.080 ;
        RECT 1940.810 586.880 1941.130 586.940 ;
        RECT 1944.950 586.880 1945.270 586.940 ;
        RECT 1944.950 37.640 1945.270 37.700 ;
        RECT 2470.730 37.640 2471.050 37.700 ;
        RECT 1944.950 37.500 2471.050 37.640 ;
        RECT 1944.950 37.440 1945.270 37.500 ;
        RECT 2470.730 37.440 2471.050 37.500 ;
      LAYER via ;
        RECT 1940.840 586.880 1941.100 587.140 ;
        RECT 1944.980 586.880 1945.240 587.140 ;
        RECT 1944.980 37.440 1945.240 37.700 ;
        RECT 2470.760 37.440 2471.020 37.700 ;
      LAYER met2 ;
        RECT 1939.230 600.170 1939.510 604.000 ;
        RECT 1939.230 600.030 1941.040 600.170 ;
        RECT 1939.230 600.000 1939.510 600.030 ;
        RECT 1940.900 587.170 1941.040 600.030 ;
        RECT 1940.840 586.850 1941.100 587.170 ;
        RECT 1944.980 586.850 1945.240 587.170 ;
        RECT 1945.040 37.730 1945.180 586.850 ;
        RECT 1944.980 37.410 1945.240 37.730 ;
        RECT 2470.760 37.410 2471.020 37.730 ;
        RECT 2470.820 2.400 2470.960 37.410 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1948.630 579.940 1948.950 580.000 ;
        RECT 1949.550 579.940 1949.870 580.000 ;
        RECT 1948.630 579.800 1949.870 579.940 ;
        RECT 1948.630 579.740 1948.950 579.800 ;
        RECT 1949.550 579.740 1949.870 579.800 ;
        RECT 1949.550 579.260 1949.870 579.320 ;
        RECT 1950.930 579.260 1951.250 579.320 ;
        RECT 1949.550 579.120 1951.250 579.260 ;
        RECT 1949.550 579.060 1949.870 579.120 ;
        RECT 1950.930 579.060 1951.250 579.120 ;
        RECT 1950.470 524.180 1950.790 524.240 ;
        RECT 1951.390 524.180 1951.710 524.240 ;
        RECT 1950.470 524.040 1951.710 524.180 ;
        RECT 1950.470 523.980 1950.790 524.040 ;
        RECT 1951.390 523.980 1951.710 524.040 ;
        RECT 1950.470 476.240 1950.790 476.300 ;
        RECT 1951.390 476.240 1951.710 476.300 ;
        RECT 1950.470 476.100 1951.710 476.240 ;
        RECT 1950.470 476.040 1950.790 476.100 ;
        RECT 1951.390 476.040 1951.710 476.100 ;
        RECT 1951.390 448.700 1951.710 448.760 ;
        RECT 1951.390 448.560 1952.080 448.700 ;
        RECT 1951.390 448.500 1951.710 448.560 ;
        RECT 1951.940 448.420 1952.080 448.560 ;
        RECT 1951.850 448.160 1952.170 448.420 ;
        RECT 1950.470 434.760 1950.790 434.820 ;
        RECT 1951.390 434.760 1951.710 434.820 ;
        RECT 1950.470 434.620 1951.710 434.760 ;
        RECT 1950.470 434.560 1950.790 434.620 ;
        RECT 1951.390 434.560 1951.710 434.620 ;
        RECT 1950.470 386.480 1950.790 386.540 ;
        RECT 1950.930 386.480 1951.250 386.540 ;
        RECT 1950.470 386.340 1951.250 386.480 ;
        RECT 1950.470 386.280 1950.790 386.340 ;
        RECT 1950.930 386.280 1951.250 386.340 ;
        RECT 1950.930 338.340 1951.250 338.600 ;
        RECT 1951.020 337.580 1951.160 338.340 ;
        RECT 1950.930 337.320 1951.250 337.580 ;
        RECT 1950.930 303.660 1951.250 303.920 ;
        RECT 1951.020 303.240 1951.160 303.660 ;
        RECT 1950.930 302.980 1951.250 303.240 ;
        RECT 1950.930 255.380 1951.250 255.640 ;
        RECT 1951.020 254.620 1951.160 255.380 ;
        RECT 1950.930 254.360 1951.250 254.620 ;
        RECT 1950.930 158.680 1951.250 158.740 ;
        RECT 1951.850 158.680 1952.170 158.740 ;
        RECT 1950.930 158.540 1952.170 158.680 ;
        RECT 1950.930 158.480 1951.250 158.540 ;
        RECT 1951.850 158.480 1952.170 158.540 ;
        RECT 1950.470 144.740 1950.790 144.800 ;
        RECT 1951.850 144.740 1952.170 144.800 ;
        RECT 1950.470 144.600 1952.170 144.740 ;
        RECT 1950.470 144.540 1950.790 144.600 ;
        RECT 1951.850 144.540 1952.170 144.600 ;
        RECT 1950.470 96.800 1950.790 96.860 ;
        RECT 1951.390 96.800 1951.710 96.860 ;
        RECT 1950.470 96.660 1951.710 96.800 ;
        RECT 1950.470 96.600 1950.790 96.660 ;
        RECT 1951.390 96.600 1951.710 96.660 ;
        RECT 1951.390 47.160 1951.710 47.220 ;
        RECT 2488.670 47.160 2488.990 47.220 ;
        RECT 1951.390 47.020 2488.990 47.160 ;
        RECT 1951.390 46.960 1951.710 47.020 ;
        RECT 2488.670 46.960 2488.990 47.020 ;
      LAYER via ;
        RECT 1948.660 579.740 1948.920 580.000 ;
        RECT 1949.580 579.740 1949.840 580.000 ;
        RECT 1949.580 579.060 1949.840 579.320 ;
        RECT 1950.960 579.060 1951.220 579.320 ;
        RECT 1950.500 523.980 1950.760 524.240 ;
        RECT 1951.420 523.980 1951.680 524.240 ;
        RECT 1950.500 476.040 1950.760 476.300 ;
        RECT 1951.420 476.040 1951.680 476.300 ;
        RECT 1951.420 448.500 1951.680 448.760 ;
        RECT 1951.880 448.160 1952.140 448.420 ;
        RECT 1950.500 434.560 1950.760 434.820 ;
        RECT 1951.420 434.560 1951.680 434.820 ;
        RECT 1950.500 386.280 1950.760 386.540 ;
        RECT 1950.960 386.280 1951.220 386.540 ;
        RECT 1950.960 338.340 1951.220 338.600 ;
        RECT 1950.960 337.320 1951.220 337.580 ;
        RECT 1950.960 303.660 1951.220 303.920 ;
        RECT 1950.960 302.980 1951.220 303.240 ;
        RECT 1950.960 255.380 1951.220 255.640 ;
        RECT 1950.960 254.360 1951.220 254.620 ;
        RECT 1950.960 158.480 1951.220 158.740 ;
        RECT 1951.880 158.480 1952.140 158.740 ;
        RECT 1950.500 144.540 1950.760 144.800 ;
        RECT 1951.880 144.540 1952.140 144.800 ;
        RECT 1950.500 96.600 1950.760 96.860 ;
        RECT 1951.420 96.600 1951.680 96.860 ;
        RECT 1951.420 46.960 1951.680 47.220 ;
        RECT 2488.700 46.960 2488.960 47.220 ;
      LAYER met2 ;
        RECT 1948.430 600.000 1948.710 604.000 ;
        RECT 1948.490 598.810 1948.630 600.000 ;
        RECT 1948.490 598.670 1948.860 598.810 ;
        RECT 1948.720 580.030 1948.860 598.670 ;
        RECT 1948.660 579.710 1948.920 580.030 ;
        RECT 1949.580 579.710 1949.840 580.030 ;
        RECT 1949.640 579.350 1949.780 579.710 ;
        RECT 1949.580 579.030 1949.840 579.350 ;
        RECT 1950.960 579.030 1951.220 579.350 ;
        RECT 1951.020 543.730 1951.160 579.030 ;
        RECT 1951.020 543.590 1951.620 543.730 ;
        RECT 1951.480 524.270 1951.620 543.590 ;
        RECT 1950.500 523.950 1950.760 524.270 ;
        RECT 1951.420 523.950 1951.680 524.270 ;
        RECT 1950.560 476.330 1950.700 523.950 ;
        RECT 1950.500 476.010 1950.760 476.330 ;
        RECT 1951.420 476.010 1951.680 476.330 ;
        RECT 1951.480 448.790 1951.620 476.010 ;
        RECT 1951.420 448.470 1951.680 448.790 ;
        RECT 1951.880 448.130 1952.140 448.450 ;
        RECT 1951.940 434.930 1952.080 448.130 ;
        RECT 1951.480 434.850 1952.080 434.930 ;
        RECT 1950.500 434.530 1950.760 434.850 ;
        RECT 1951.420 434.790 1952.080 434.850 ;
        RECT 1951.420 434.530 1951.680 434.790 ;
        RECT 1950.560 386.570 1950.700 434.530 ;
        RECT 1950.500 386.250 1950.760 386.570 ;
        RECT 1950.960 386.250 1951.220 386.570 ;
        RECT 1951.020 338.630 1951.160 386.250 ;
        RECT 1950.960 338.310 1951.220 338.630 ;
        RECT 1950.960 337.290 1951.220 337.610 ;
        RECT 1951.020 303.950 1951.160 337.290 ;
        RECT 1950.960 303.630 1951.220 303.950 ;
        RECT 1950.960 302.950 1951.220 303.270 ;
        RECT 1951.020 255.670 1951.160 302.950 ;
        RECT 1950.960 255.350 1951.220 255.670 ;
        RECT 1950.960 254.330 1951.220 254.650 ;
        RECT 1951.020 207.245 1951.160 254.330 ;
        RECT 1950.950 206.875 1951.230 207.245 ;
        RECT 1950.950 206.195 1951.230 206.565 ;
        RECT 1951.020 158.770 1951.160 206.195 ;
        RECT 1950.960 158.450 1951.220 158.770 ;
        RECT 1951.880 158.450 1952.140 158.770 ;
        RECT 1951.940 144.830 1952.080 158.450 ;
        RECT 1950.500 144.510 1950.760 144.830 ;
        RECT 1951.880 144.510 1952.140 144.830 ;
        RECT 1950.560 96.890 1950.700 144.510 ;
        RECT 1950.500 96.570 1950.760 96.890 ;
        RECT 1951.420 96.570 1951.680 96.890 ;
        RECT 1951.480 47.250 1951.620 96.570 ;
        RECT 1951.420 46.930 1951.680 47.250 ;
        RECT 2488.700 46.930 2488.960 47.250 ;
        RECT 2488.760 2.400 2488.900 46.930 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
      LAYER via2 ;
        RECT 1950.950 206.920 1951.230 207.200 ;
        RECT 1950.950 206.240 1951.230 206.520 ;
      LAYER met3 ;
        RECT 1950.925 207.210 1951.255 207.225 ;
        RECT 1950.710 206.895 1951.255 207.210 ;
        RECT 1950.710 206.545 1951.010 206.895 ;
        RECT 1950.710 206.230 1951.255 206.545 ;
        RECT 1950.925 206.215 1951.255 206.230 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1959.210 46.820 1959.530 46.880 ;
        RECT 2506.150 46.820 2506.470 46.880 ;
        RECT 1959.210 46.680 2506.470 46.820 ;
        RECT 1959.210 46.620 1959.530 46.680 ;
        RECT 2506.150 46.620 2506.470 46.680 ;
      LAYER via ;
        RECT 1959.240 46.620 1959.500 46.880 ;
        RECT 2506.180 46.620 2506.440 46.880 ;
      LAYER met2 ;
        RECT 1957.630 600.170 1957.910 604.000 ;
        RECT 1957.630 600.030 1959.440 600.170 ;
        RECT 1957.630 600.000 1957.910 600.030 ;
        RECT 1959.300 46.910 1959.440 600.030 ;
        RECT 1959.240 46.590 1959.500 46.910 ;
        RECT 2506.180 46.590 2506.440 46.910 ;
        RECT 2506.240 2.400 2506.380 46.590 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1968.410 587.080 1968.730 587.140 ;
        RECT 1972.550 587.080 1972.870 587.140 ;
        RECT 1968.410 586.940 1972.870 587.080 ;
        RECT 1968.410 586.880 1968.730 586.940 ;
        RECT 1972.550 586.880 1972.870 586.940 ;
        RECT 1972.550 46.480 1972.870 46.540 ;
        RECT 2524.090 46.480 2524.410 46.540 ;
        RECT 1972.550 46.340 2524.410 46.480 ;
        RECT 1972.550 46.280 1972.870 46.340 ;
        RECT 2524.090 46.280 2524.410 46.340 ;
      LAYER via ;
        RECT 1968.440 586.880 1968.700 587.140 ;
        RECT 1972.580 586.880 1972.840 587.140 ;
        RECT 1972.580 46.280 1972.840 46.540 ;
        RECT 2524.120 46.280 2524.380 46.540 ;
      LAYER met2 ;
        RECT 1966.830 600.170 1967.110 604.000 ;
        RECT 1966.830 600.030 1968.640 600.170 ;
        RECT 1966.830 600.000 1967.110 600.030 ;
        RECT 1968.500 587.170 1968.640 600.030 ;
        RECT 1968.440 586.850 1968.700 587.170 ;
        RECT 1972.580 586.850 1972.840 587.170 ;
        RECT 1972.640 46.570 1972.780 586.850 ;
        RECT 1972.580 46.250 1972.840 46.570 ;
        RECT 2524.120 46.250 2524.380 46.570 ;
        RECT 2524.180 2.400 2524.320 46.250 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1977.150 586.740 1977.470 586.800 ;
        RECT 1979.450 586.740 1979.770 586.800 ;
        RECT 1977.150 586.600 1979.770 586.740 ;
        RECT 1977.150 586.540 1977.470 586.600 ;
        RECT 1979.450 586.540 1979.770 586.600 ;
        RECT 1979.450 46.140 1979.770 46.200 ;
        RECT 2542.030 46.140 2542.350 46.200 ;
        RECT 1979.450 46.000 2542.350 46.140 ;
        RECT 1979.450 45.940 1979.770 46.000 ;
        RECT 2542.030 45.940 2542.350 46.000 ;
      LAYER via ;
        RECT 1977.180 586.540 1977.440 586.800 ;
        RECT 1979.480 586.540 1979.740 586.800 ;
        RECT 1979.480 45.940 1979.740 46.200 ;
        RECT 2542.060 45.940 2542.320 46.200 ;
      LAYER met2 ;
        RECT 1975.570 600.170 1975.850 604.000 ;
        RECT 1975.570 600.030 1977.380 600.170 ;
        RECT 1975.570 600.000 1975.850 600.030 ;
        RECT 1977.240 586.830 1977.380 600.030 ;
        RECT 1977.180 586.510 1977.440 586.830 ;
        RECT 1979.480 586.510 1979.740 586.830 ;
        RECT 1979.540 46.230 1979.680 586.510 ;
        RECT 1979.480 45.910 1979.740 46.230 ;
        RECT 2542.060 45.910 2542.320 46.230 ;
        RECT 2542.120 2.400 2542.260 45.910 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1986.810 45.800 1987.130 45.860 ;
        RECT 2559.970 45.800 2560.290 45.860 ;
        RECT 1986.810 45.660 2560.290 45.800 ;
        RECT 1986.810 45.600 1987.130 45.660 ;
        RECT 2559.970 45.600 2560.290 45.660 ;
      LAYER via ;
        RECT 1986.840 45.600 1987.100 45.860 ;
        RECT 2560.000 45.600 2560.260 45.860 ;
      LAYER met2 ;
        RECT 1984.770 600.170 1985.050 604.000 ;
        RECT 1984.770 600.030 1987.040 600.170 ;
        RECT 1984.770 600.000 1985.050 600.030 ;
        RECT 1986.900 45.890 1987.040 600.030 ;
        RECT 1986.840 45.570 1987.100 45.890 ;
        RECT 2560.000 45.570 2560.260 45.890 ;
        RECT 2560.060 2.400 2560.200 45.570 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1995.550 586.740 1995.870 586.800 ;
        RECT 2000.610 586.740 2000.930 586.800 ;
        RECT 1995.550 586.600 2000.930 586.740 ;
        RECT 1995.550 586.540 1995.870 586.600 ;
        RECT 2000.610 586.540 2000.930 586.600 ;
        RECT 2000.610 21.320 2000.930 21.380 ;
        RECT 2577.910 21.320 2578.230 21.380 ;
        RECT 2000.610 21.180 2578.230 21.320 ;
        RECT 2000.610 21.120 2000.930 21.180 ;
        RECT 2577.910 21.120 2578.230 21.180 ;
      LAYER via ;
        RECT 1995.580 586.540 1995.840 586.800 ;
        RECT 2000.640 586.540 2000.900 586.800 ;
        RECT 2000.640 21.120 2000.900 21.380 ;
        RECT 2577.940 21.120 2578.200 21.380 ;
      LAYER met2 ;
        RECT 1993.970 600.170 1994.250 604.000 ;
        RECT 1993.970 600.030 1995.780 600.170 ;
        RECT 1993.970 600.000 1994.250 600.030 ;
        RECT 1995.640 586.830 1995.780 600.030 ;
        RECT 1995.580 586.510 1995.840 586.830 ;
        RECT 2000.640 586.510 2000.900 586.830 ;
        RECT 2000.700 21.410 2000.840 586.510 ;
        RECT 2000.640 21.090 2000.900 21.410 ;
        RECT 2577.940 21.090 2578.200 21.410 ;
        RECT 2578.000 2.400 2578.140 21.090 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 811.510 17.240 811.830 17.300 ;
        RECT 1084.750 17.240 1085.070 17.300 ;
        RECT 811.510 17.100 1085.070 17.240 ;
        RECT 811.510 17.040 811.830 17.100 ;
        RECT 1084.750 17.040 1085.070 17.100 ;
      LAYER via ;
        RECT 811.540 17.040 811.800 17.300 ;
        RECT 1084.780 17.040 1085.040 17.300 ;
      LAYER met2 ;
        RECT 1086.850 600.170 1087.130 604.000 ;
        RECT 1084.840 600.030 1087.130 600.170 ;
        RECT 1084.840 17.330 1084.980 600.030 ;
        RECT 1086.850 600.000 1087.130 600.030 ;
        RECT 811.540 17.010 811.800 17.330 ;
        RECT 1084.780 17.010 1085.040 17.330 ;
        RECT 811.600 2.400 811.740 17.010 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2004.750 586.740 2005.070 586.800 ;
        RECT 2007.510 586.740 2007.830 586.800 ;
        RECT 2004.750 586.600 2007.830 586.740 ;
        RECT 2004.750 586.540 2005.070 586.600 ;
        RECT 2007.510 586.540 2007.830 586.600 ;
        RECT 2007.510 21.660 2007.830 21.720 ;
        RECT 2595.390 21.660 2595.710 21.720 ;
        RECT 2007.510 21.520 2595.710 21.660 ;
        RECT 2007.510 21.460 2007.830 21.520 ;
        RECT 2595.390 21.460 2595.710 21.520 ;
      LAYER via ;
        RECT 2004.780 586.540 2005.040 586.800 ;
        RECT 2007.540 586.540 2007.800 586.800 ;
        RECT 2007.540 21.460 2007.800 21.720 ;
        RECT 2595.420 21.460 2595.680 21.720 ;
      LAYER met2 ;
        RECT 2003.170 600.170 2003.450 604.000 ;
        RECT 2003.170 600.030 2004.980 600.170 ;
        RECT 2003.170 600.000 2003.450 600.030 ;
        RECT 2004.840 586.830 2004.980 600.030 ;
        RECT 2004.780 586.510 2005.040 586.830 ;
        RECT 2007.540 586.510 2007.800 586.830 ;
        RECT 2007.600 21.750 2007.740 586.510 ;
        RECT 2007.540 21.430 2007.800 21.750 ;
        RECT 2595.420 21.430 2595.680 21.750 ;
        RECT 2595.480 2.400 2595.620 21.430 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2014.410 22.000 2014.730 22.060 ;
        RECT 2613.330 22.000 2613.650 22.060 ;
        RECT 2014.410 21.860 2613.650 22.000 ;
        RECT 2014.410 21.800 2014.730 21.860 ;
        RECT 2613.330 21.800 2613.650 21.860 ;
      LAYER via ;
        RECT 2014.440 21.800 2014.700 22.060 ;
        RECT 2613.360 21.800 2613.620 22.060 ;
      LAYER met2 ;
        RECT 2012.370 600.170 2012.650 604.000 ;
        RECT 2012.370 600.030 2014.640 600.170 ;
        RECT 2012.370 600.000 2012.650 600.030 ;
        RECT 2014.500 22.090 2014.640 600.030 ;
        RECT 2014.440 21.770 2014.700 22.090 ;
        RECT 2613.360 21.770 2613.620 22.090 ;
        RECT 2613.420 2.400 2613.560 21.770 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2023.150 586.740 2023.470 586.800 ;
        RECT 2028.210 586.740 2028.530 586.800 ;
        RECT 2023.150 586.600 2028.530 586.740 ;
        RECT 2023.150 586.540 2023.470 586.600 ;
        RECT 2028.210 586.540 2028.530 586.600 ;
        RECT 2028.210 22.340 2028.530 22.400 ;
        RECT 2631.270 22.340 2631.590 22.400 ;
        RECT 2028.210 22.200 2631.590 22.340 ;
        RECT 2028.210 22.140 2028.530 22.200 ;
        RECT 2631.270 22.140 2631.590 22.200 ;
      LAYER via ;
        RECT 2023.180 586.540 2023.440 586.800 ;
        RECT 2028.240 586.540 2028.500 586.800 ;
        RECT 2028.240 22.140 2028.500 22.400 ;
        RECT 2631.300 22.140 2631.560 22.400 ;
      LAYER met2 ;
        RECT 2021.570 600.170 2021.850 604.000 ;
        RECT 2021.570 600.030 2023.380 600.170 ;
        RECT 2021.570 600.000 2021.850 600.030 ;
        RECT 2023.240 586.830 2023.380 600.030 ;
        RECT 2023.180 586.510 2023.440 586.830 ;
        RECT 2028.240 586.510 2028.500 586.830 ;
        RECT 2028.300 22.430 2028.440 586.510 ;
        RECT 2028.240 22.110 2028.500 22.430 ;
        RECT 2631.300 22.110 2631.560 22.430 ;
        RECT 2631.360 2.400 2631.500 22.110 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2032.350 586.740 2032.670 586.800 ;
        RECT 2035.110 586.740 2035.430 586.800 ;
        RECT 2032.350 586.600 2035.430 586.740 ;
        RECT 2032.350 586.540 2032.670 586.600 ;
        RECT 2035.110 586.540 2035.430 586.600 ;
        RECT 2035.110 22.680 2035.430 22.740 ;
        RECT 2649.210 22.680 2649.530 22.740 ;
        RECT 2035.110 22.540 2649.530 22.680 ;
        RECT 2035.110 22.480 2035.430 22.540 ;
        RECT 2649.210 22.480 2649.530 22.540 ;
      LAYER via ;
        RECT 2032.380 586.540 2032.640 586.800 ;
        RECT 2035.140 586.540 2035.400 586.800 ;
        RECT 2035.140 22.480 2035.400 22.740 ;
        RECT 2649.240 22.480 2649.500 22.740 ;
      LAYER met2 ;
        RECT 2030.770 600.170 2031.050 604.000 ;
        RECT 2030.770 600.030 2032.580 600.170 ;
        RECT 2030.770 600.000 2031.050 600.030 ;
        RECT 2032.440 586.830 2032.580 600.030 ;
        RECT 2032.380 586.510 2032.640 586.830 ;
        RECT 2035.140 586.510 2035.400 586.830 ;
        RECT 2035.200 22.770 2035.340 586.510 ;
        RECT 2035.140 22.450 2035.400 22.770 ;
        RECT 2649.240 22.450 2649.500 22.770 ;
        RECT 2649.300 2.400 2649.440 22.450 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2041.550 23.020 2041.870 23.080 ;
        RECT 2667.150 23.020 2667.470 23.080 ;
        RECT 2041.550 22.880 2667.470 23.020 ;
        RECT 2041.550 22.820 2041.870 22.880 ;
        RECT 2667.150 22.820 2667.470 22.880 ;
      LAYER via ;
        RECT 2041.580 22.820 2041.840 23.080 ;
        RECT 2667.180 22.820 2667.440 23.080 ;
      LAYER met2 ;
        RECT 2039.970 600.170 2040.250 604.000 ;
        RECT 2039.970 600.030 2041.780 600.170 ;
        RECT 2039.970 600.000 2040.250 600.030 ;
        RECT 2041.640 23.110 2041.780 600.030 ;
        RECT 2041.580 22.790 2041.840 23.110 ;
        RECT 2667.180 22.790 2667.440 23.110 ;
        RECT 2667.240 2.400 2667.380 22.790 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2050.750 586.740 2051.070 586.800 ;
        RECT 2055.350 586.740 2055.670 586.800 ;
        RECT 2050.750 586.600 2055.670 586.740 ;
        RECT 2050.750 586.540 2051.070 586.600 ;
        RECT 2055.350 586.540 2055.670 586.600 ;
        RECT 2055.350 23.360 2055.670 23.420 ;
        RECT 2684.630 23.360 2684.950 23.420 ;
        RECT 2055.350 23.220 2684.950 23.360 ;
        RECT 2055.350 23.160 2055.670 23.220 ;
        RECT 2684.630 23.160 2684.950 23.220 ;
      LAYER via ;
        RECT 2050.780 586.540 2051.040 586.800 ;
        RECT 2055.380 586.540 2055.640 586.800 ;
        RECT 2055.380 23.160 2055.640 23.420 ;
        RECT 2684.660 23.160 2684.920 23.420 ;
      LAYER met2 ;
        RECT 2049.170 600.170 2049.450 604.000 ;
        RECT 2049.170 600.030 2050.980 600.170 ;
        RECT 2049.170 600.000 2049.450 600.030 ;
        RECT 2050.840 586.830 2050.980 600.030 ;
        RECT 2050.780 586.510 2051.040 586.830 ;
        RECT 2055.380 586.510 2055.640 586.830 ;
        RECT 2055.440 23.450 2055.580 586.510 ;
        RECT 2055.380 23.130 2055.640 23.450 ;
        RECT 2684.660 23.130 2684.920 23.450 ;
        RECT 2684.720 2.400 2684.860 23.130 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2059.950 586.740 2060.270 586.800 ;
        RECT 2062.710 586.740 2063.030 586.800 ;
        RECT 2059.950 586.600 2063.030 586.740 ;
        RECT 2059.950 586.540 2060.270 586.600 ;
        RECT 2062.710 586.540 2063.030 586.600 ;
        RECT 2062.710 23.700 2063.030 23.760 ;
        RECT 2702.570 23.700 2702.890 23.760 ;
        RECT 2062.710 23.560 2702.890 23.700 ;
        RECT 2062.710 23.500 2063.030 23.560 ;
        RECT 2702.570 23.500 2702.890 23.560 ;
      LAYER via ;
        RECT 2059.980 586.540 2060.240 586.800 ;
        RECT 2062.740 586.540 2063.000 586.800 ;
        RECT 2062.740 23.500 2063.000 23.760 ;
        RECT 2702.600 23.500 2702.860 23.760 ;
      LAYER met2 ;
        RECT 2058.370 600.170 2058.650 604.000 ;
        RECT 2058.370 600.030 2060.180 600.170 ;
        RECT 2058.370 600.000 2058.650 600.030 ;
        RECT 2060.040 586.830 2060.180 600.030 ;
        RECT 2059.980 586.510 2060.240 586.830 ;
        RECT 2062.740 586.510 2063.000 586.830 ;
        RECT 2062.800 23.790 2062.940 586.510 ;
        RECT 2062.740 23.470 2063.000 23.790 ;
        RECT 2702.600 23.470 2702.860 23.790 ;
        RECT 2702.660 2.400 2702.800 23.470 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2069.610 27.440 2069.930 27.500 ;
        RECT 2720.510 27.440 2720.830 27.500 ;
        RECT 2069.610 27.300 2720.830 27.440 ;
        RECT 2069.610 27.240 2069.930 27.300 ;
        RECT 2720.510 27.240 2720.830 27.300 ;
      LAYER via ;
        RECT 2069.640 27.240 2069.900 27.500 ;
        RECT 2720.540 27.240 2720.800 27.500 ;
      LAYER met2 ;
        RECT 2067.570 600.170 2067.850 604.000 ;
        RECT 2067.570 600.030 2069.840 600.170 ;
        RECT 2067.570 600.000 2067.850 600.030 ;
        RECT 2069.700 27.530 2069.840 600.030 ;
        RECT 2069.640 27.210 2069.900 27.530 ;
        RECT 2720.540 27.210 2720.800 27.530 ;
        RECT 2720.600 2.400 2720.740 27.210 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2078.350 586.740 2078.670 586.800 ;
        RECT 2083.410 586.740 2083.730 586.800 ;
        RECT 2078.350 586.600 2083.730 586.740 ;
        RECT 2078.350 586.540 2078.670 586.600 ;
        RECT 2083.410 586.540 2083.730 586.600 ;
        RECT 2083.410 27.100 2083.730 27.160 ;
        RECT 2738.450 27.100 2738.770 27.160 ;
        RECT 2083.410 26.960 2738.770 27.100 ;
        RECT 2083.410 26.900 2083.730 26.960 ;
        RECT 2738.450 26.900 2738.770 26.960 ;
      LAYER via ;
        RECT 2078.380 586.540 2078.640 586.800 ;
        RECT 2083.440 586.540 2083.700 586.800 ;
        RECT 2083.440 26.900 2083.700 27.160 ;
        RECT 2738.480 26.900 2738.740 27.160 ;
      LAYER met2 ;
        RECT 2076.770 600.170 2077.050 604.000 ;
        RECT 2076.770 600.030 2078.580 600.170 ;
        RECT 2076.770 600.000 2077.050 600.030 ;
        RECT 2078.440 586.830 2078.580 600.030 ;
        RECT 2078.380 586.510 2078.640 586.830 ;
        RECT 2083.440 586.510 2083.700 586.830 ;
        RECT 2083.500 27.190 2083.640 586.510 ;
        RECT 2083.440 26.870 2083.700 27.190 ;
        RECT 2738.480 26.870 2738.740 27.190 ;
        RECT 2738.540 2.400 2738.680 26.870 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2087.550 586.740 2087.870 586.800 ;
        RECT 2090.310 586.740 2090.630 586.800 ;
        RECT 2087.550 586.600 2090.630 586.740 ;
        RECT 2087.550 586.540 2087.870 586.600 ;
        RECT 2090.310 586.540 2090.630 586.600 ;
        RECT 2090.310 26.760 2090.630 26.820 ;
        RECT 2755.930 26.760 2756.250 26.820 ;
        RECT 2090.310 26.620 2756.250 26.760 ;
        RECT 2090.310 26.560 2090.630 26.620 ;
        RECT 2755.930 26.560 2756.250 26.620 ;
      LAYER via ;
        RECT 2087.580 586.540 2087.840 586.800 ;
        RECT 2090.340 586.540 2090.600 586.800 ;
        RECT 2090.340 26.560 2090.600 26.820 ;
        RECT 2755.960 26.560 2756.220 26.820 ;
      LAYER met2 ;
        RECT 2085.970 600.170 2086.250 604.000 ;
        RECT 2085.970 600.030 2087.780 600.170 ;
        RECT 2085.970 600.000 2086.250 600.030 ;
        RECT 2087.640 586.830 2087.780 600.030 ;
        RECT 2087.580 586.510 2087.840 586.830 ;
        RECT 2090.340 586.510 2090.600 586.830 ;
        RECT 2090.400 26.850 2090.540 586.510 ;
        RECT 2090.340 26.530 2090.600 26.850 ;
        RECT 2755.960 26.530 2756.220 26.850 ;
        RECT 2756.020 2.400 2756.160 26.530 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1091.650 476.240 1091.970 476.300 ;
        RECT 1093.950 476.240 1094.270 476.300 ;
        RECT 1091.650 476.100 1094.270 476.240 ;
        RECT 1091.650 476.040 1091.970 476.100 ;
        RECT 1093.950 476.040 1094.270 476.100 ;
        RECT 1091.650 324.260 1091.970 324.320 ;
        RECT 1092.110 324.260 1092.430 324.320 ;
        RECT 1091.650 324.120 1092.430 324.260 ;
        RECT 1091.650 324.060 1091.970 324.120 ;
        RECT 1092.110 324.060 1092.430 324.120 ;
        RECT 1091.190 234.840 1091.510 234.900 ;
        RECT 1092.110 234.840 1092.430 234.900 ;
        RECT 1091.190 234.700 1092.430 234.840 ;
        RECT 1091.190 234.640 1091.510 234.700 ;
        RECT 1092.110 234.640 1092.430 234.700 ;
        RECT 1091.190 186.700 1091.510 186.960 ;
        RECT 1091.280 186.560 1091.420 186.700 ;
        RECT 1091.650 186.560 1091.970 186.620 ;
        RECT 1091.280 186.420 1091.970 186.560 ;
        RECT 1091.650 186.360 1091.970 186.420 ;
        RECT 1091.650 159.020 1091.970 159.080 ;
        RECT 1091.280 158.880 1091.970 159.020 ;
        RECT 1091.280 158.740 1091.420 158.880 ;
        RECT 1091.650 158.820 1091.970 158.880 ;
        RECT 1091.190 158.480 1091.510 158.740 ;
        RECT 1091.190 41.720 1091.510 41.780 ;
        RECT 1091.650 41.720 1091.970 41.780 ;
        RECT 1091.190 41.580 1091.970 41.720 ;
        RECT 1091.190 41.520 1091.510 41.580 ;
        RECT 1091.650 41.520 1091.970 41.580 ;
        RECT 829.450 17.580 829.770 17.640 ;
        RECT 1039.210 17.580 1039.530 17.640 ;
        RECT 829.450 17.440 1039.530 17.580 ;
        RECT 829.450 17.380 829.770 17.440 ;
        RECT 1039.210 17.380 1039.530 17.440 ;
        RECT 1039.210 15.200 1039.530 15.260 ;
        RECT 1091.190 15.200 1091.510 15.260 ;
        RECT 1039.210 15.060 1091.510 15.200 ;
        RECT 1039.210 15.000 1039.530 15.060 ;
        RECT 1091.190 15.000 1091.510 15.060 ;
      LAYER via ;
        RECT 1091.680 476.040 1091.940 476.300 ;
        RECT 1093.980 476.040 1094.240 476.300 ;
        RECT 1091.680 324.060 1091.940 324.320 ;
        RECT 1092.140 324.060 1092.400 324.320 ;
        RECT 1091.220 234.640 1091.480 234.900 ;
        RECT 1092.140 234.640 1092.400 234.900 ;
        RECT 1091.220 186.700 1091.480 186.960 ;
        RECT 1091.680 186.360 1091.940 186.620 ;
        RECT 1091.680 158.820 1091.940 159.080 ;
        RECT 1091.220 158.480 1091.480 158.740 ;
        RECT 1091.220 41.520 1091.480 41.780 ;
        RECT 1091.680 41.520 1091.940 41.780 ;
        RECT 829.480 17.380 829.740 17.640 ;
        RECT 1039.240 17.380 1039.500 17.640 ;
        RECT 1039.240 15.000 1039.500 15.260 ;
        RECT 1091.220 15.000 1091.480 15.260 ;
      LAYER met2 ;
        RECT 1096.050 600.170 1096.330 604.000 ;
        RECT 1095.420 600.030 1096.330 600.170 ;
        RECT 1095.420 579.885 1095.560 600.030 ;
        RECT 1096.050 600.000 1096.330 600.030 ;
        RECT 1093.970 579.515 1094.250 579.885 ;
        RECT 1095.350 579.515 1095.630 579.885 ;
        RECT 1094.040 476.330 1094.180 579.515 ;
        RECT 1091.680 476.010 1091.940 476.330 ;
        RECT 1093.980 476.010 1094.240 476.330 ;
        RECT 1091.740 458.730 1091.880 476.010 ;
        RECT 1091.740 458.590 1092.340 458.730 ;
        RECT 1092.200 331.570 1092.340 458.590 ;
        RECT 1091.740 331.430 1092.340 331.570 ;
        RECT 1091.740 324.350 1091.880 331.430 ;
        RECT 1091.680 324.030 1091.940 324.350 ;
        RECT 1092.140 324.030 1092.400 324.350 ;
        RECT 1092.200 234.930 1092.340 324.030 ;
        RECT 1091.220 234.610 1091.480 234.930 ;
        RECT 1092.140 234.610 1092.400 234.930 ;
        RECT 1091.280 186.990 1091.420 234.610 ;
        RECT 1091.220 186.670 1091.480 186.990 ;
        RECT 1091.680 186.330 1091.940 186.650 ;
        RECT 1091.740 159.110 1091.880 186.330 ;
        RECT 1091.680 158.790 1091.940 159.110 ;
        RECT 1091.220 158.450 1091.480 158.770 ;
        RECT 1091.280 130.970 1091.420 158.450 ;
        RECT 1091.280 130.830 1091.880 130.970 ;
        RECT 1091.740 41.810 1091.880 130.830 ;
        RECT 1091.220 41.490 1091.480 41.810 ;
        RECT 1091.680 41.490 1091.940 41.810 ;
        RECT 829.480 17.350 829.740 17.670 ;
        RECT 1039.240 17.350 1039.500 17.670 ;
        RECT 829.540 2.400 829.680 17.350 ;
        RECT 1039.300 15.290 1039.440 17.350 ;
        RECT 1091.280 15.290 1091.420 41.490 ;
        RECT 1039.240 14.970 1039.500 15.290 ;
        RECT 1091.220 14.970 1091.480 15.290 ;
        RECT 829.330 -4.800 829.890 2.400 ;
      LAYER via2 ;
        RECT 1093.970 579.560 1094.250 579.840 ;
        RECT 1095.350 579.560 1095.630 579.840 ;
      LAYER met3 ;
        RECT 1093.945 579.850 1094.275 579.865 ;
        RECT 1095.325 579.850 1095.655 579.865 ;
        RECT 1093.945 579.550 1095.655 579.850 ;
        RECT 1093.945 579.535 1094.275 579.550 ;
        RECT 1095.325 579.535 1095.655 579.550 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2096.750 26.420 2097.070 26.480 ;
        RECT 2773.870 26.420 2774.190 26.480 ;
        RECT 2096.750 26.280 2774.190 26.420 ;
        RECT 2096.750 26.220 2097.070 26.280 ;
        RECT 2773.870 26.220 2774.190 26.280 ;
      LAYER via ;
        RECT 2096.780 26.220 2097.040 26.480 ;
        RECT 2773.900 26.220 2774.160 26.480 ;
      LAYER met2 ;
        RECT 2094.710 600.170 2094.990 604.000 ;
        RECT 2094.710 600.030 2096.980 600.170 ;
        RECT 2094.710 600.000 2094.990 600.030 ;
        RECT 2096.840 26.510 2096.980 600.030 ;
        RECT 2096.780 26.190 2097.040 26.510 ;
        RECT 2773.900 26.190 2774.160 26.510 ;
        RECT 2773.960 2.400 2774.100 26.190 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2104.110 26.080 2104.430 26.140 ;
        RECT 2791.810 26.080 2792.130 26.140 ;
        RECT 2104.110 25.940 2792.130 26.080 ;
        RECT 2104.110 25.880 2104.430 25.940 ;
        RECT 2791.810 25.880 2792.130 25.940 ;
      LAYER via ;
        RECT 2104.140 25.880 2104.400 26.140 ;
        RECT 2791.840 25.880 2792.100 26.140 ;
      LAYER met2 ;
        RECT 2103.910 600.000 2104.190 604.000 ;
        RECT 2103.970 598.810 2104.110 600.000 ;
        RECT 2103.970 598.670 2104.340 598.810 ;
        RECT 2104.200 26.170 2104.340 598.670 ;
        RECT 2104.140 25.850 2104.400 26.170 ;
        RECT 2791.840 25.850 2792.100 26.170 ;
        RECT 2791.900 2.400 2792.040 25.850 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2114.690 586.740 2115.010 586.800 ;
        RECT 2117.910 586.740 2118.230 586.800 ;
        RECT 2114.690 586.600 2118.230 586.740 ;
        RECT 2114.690 586.540 2115.010 586.600 ;
        RECT 2117.910 586.540 2118.230 586.600 ;
        RECT 2117.910 25.740 2118.230 25.800 ;
        RECT 2809.750 25.740 2810.070 25.800 ;
        RECT 2117.910 25.600 2810.070 25.740 ;
        RECT 2117.910 25.540 2118.230 25.600 ;
        RECT 2809.750 25.540 2810.070 25.600 ;
      LAYER via ;
        RECT 2114.720 586.540 2114.980 586.800 ;
        RECT 2117.940 586.540 2118.200 586.800 ;
        RECT 2117.940 25.540 2118.200 25.800 ;
        RECT 2809.780 25.540 2810.040 25.800 ;
      LAYER met2 ;
        RECT 2113.110 600.170 2113.390 604.000 ;
        RECT 2113.110 600.030 2114.920 600.170 ;
        RECT 2113.110 600.000 2113.390 600.030 ;
        RECT 2114.780 586.830 2114.920 600.030 ;
        RECT 2114.720 586.510 2114.980 586.830 ;
        RECT 2117.940 586.510 2118.200 586.830 ;
        RECT 2118.000 25.830 2118.140 586.510 ;
        RECT 2117.940 25.510 2118.200 25.830 ;
        RECT 2809.780 25.510 2810.040 25.830 ;
        RECT 2809.840 2.400 2809.980 25.510 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2124.810 25.400 2125.130 25.460 ;
        RECT 2827.690 25.400 2828.010 25.460 ;
        RECT 2124.810 25.260 2828.010 25.400 ;
        RECT 2124.810 25.200 2125.130 25.260 ;
        RECT 2827.690 25.200 2828.010 25.260 ;
      LAYER via ;
        RECT 2124.840 25.200 2125.100 25.460 ;
        RECT 2827.720 25.200 2827.980 25.460 ;
      LAYER met2 ;
        RECT 2122.310 600.170 2122.590 604.000 ;
        RECT 2122.310 600.030 2125.040 600.170 ;
        RECT 2122.310 600.000 2122.590 600.030 ;
        RECT 2124.900 25.490 2125.040 600.030 ;
        RECT 2124.840 25.170 2125.100 25.490 ;
        RECT 2827.720 25.170 2827.980 25.490 ;
        RECT 2827.780 2.400 2827.920 25.170 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2129.870 592.520 2130.190 592.580 ;
        RECT 2130.790 592.520 2131.110 592.580 ;
        RECT 2129.870 592.380 2131.110 592.520 ;
        RECT 2129.870 592.320 2130.190 592.380 ;
        RECT 2130.790 592.320 2131.110 592.380 ;
        RECT 2129.870 545.260 2130.190 545.320 ;
        RECT 2131.250 545.260 2131.570 545.320 ;
        RECT 2129.870 545.120 2131.570 545.260 ;
        RECT 2129.870 545.060 2130.190 545.120 ;
        RECT 2131.250 545.060 2131.570 545.120 ;
        RECT 2131.250 497.320 2131.570 497.380 ;
        RECT 2130.420 497.180 2131.570 497.320 ;
        RECT 2130.420 497.040 2130.560 497.180 ;
        RECT 2131.250 497.120 2131.570 497.180 ;
        RECT 2130.330 496.780 2130.650 497.040 ;
        RECT 2130.330 448.700 2130.650 448.760 ;
        RECT 2131.250 448.700 2131.570 448.760 ;
        RECT 2130.330 448.560 2131.570 448.700 ;
        RECT 2130.330 448.500 2130.650 448.560 ;
        RECT 2131.250 448.500 2131.570 448.560 ;
        RECT 2131.250 400.760 2131.570 400.820 ;
        RECT 2130.420 400.620 2131.570 400.760 ;
        RECT 2130.420 400.480 2130.560 400.620 ;
        RECT 2131.250 400.560 2131.570 400.620 ;
        RECT 2130.330 400.220 2130.650 400.480 ;
        RECT 2130.330 352.140 2130.650 352.200 ;
        RECT 2131.250 352.140 2131.570 352.200 ;
        RECT 2130.330 352.000 2131.570 352.140 ;
        RECT 2130.330 351.940 2130.650 352.000 ;
        RECT 2131.250 351.940 2131.570 352.000 ;
        RECT 2131.250 304.200 2131.570 304.260 ;
        RECT 2130.420 304.060 2131.570 304.200 ;
        RECT 2130.420 303.920 2130.560 304.060 ;
        RECT 2131.250 304.000 2131.570 304.060 ;
        RECT 2130.330 303.660 2130.650 303.920 ;
        RECT 2130.330 255.580 2130.650 255.640 ;
        RECT 2131.250 255.580 2131.570 255.640 ;
        RECT 2130.330 255.440 2131.570 255.580 ;
        RECT 2130.330 255.380 2130.650 255.440 ;
        RECT 2131.250 255.380 2131.570 255.440 ;
        RECT 2130.330 207.300 2130.650 207.360 ;
        RECT 2131.250 207.300 2131.570 207.360 ;
        RECT 2130.330 207.160 2131.570 207.300 ;
        RECT 2130.330 207.100 2130.650 207.160 ;
        RECT 2131.250 207.100 2131.570 207.160 ;
        RECT 2130.330 159.020 2130.650 159.080 ;
        RECT 2131.250 159.020 2131.570 159.080 ;
        RECT 2130.330 158.880 2131.570 159.020 ;
        RECT 2130.330 158.820 2130.650 158.880 ;
        RECT 2131.250 158.820 2131.570 158.880 ;
        RECT 2130.330 62.460 2130.650 62.520 ;
        RECT 2131.250 62.460 2131.570 62.520 ;
        RECT 2130.330 62.320 2131.570 62.460 ;
        RECT 2130.330 62.260 2130.650 62.320 ;
        RECT 2131.250 62.260 2131.570 62.320 ;
        RECT 2130.330 24.720 2130.650 24.780 ;
        RECT 2845.170 24.720 2845.490 24.780 ;
        RECT 2130.330 24.580 2845.490 24.720 ;
        RECT 2130.330 24.520 2130.650 24.580 ;
        RECT 2845.170 24.520 2845.490 24.580 ;
      LAYER via ;
        RECT 2129.900 592.320 2130.160 592.580 ;
        RECT 2130.820 592.320 2131.080 592.580 ;
        RECT 2129.900 545.060 2130.160 545.320 ;
        RECT 2131.280 545.060 2131.540 545.320 ;
        RECT 2131.280 497.120 2131.540 497.380 ;
        RECT 2130.360 496.780 2130.620 497.040 ;
        RECT 2130.360 448.500 2130.620 448.760 ;
        RECT 2131.280 448.500 2131.540 448.760 ;
        RECT 2131.280 400.560 2131.540 400.820 ;
        RECT 2130.360 400.220 2130.620 400.480 ;
        RECT 2130.360 351.940 2130.620 352.200 ;
        RECT 2131.280 351.940 2131.540 352.200 ;
        RECT 2131.280 304.000 2131.540 304.260 ;
        RECT 2130.360 303.660 2130.620 303.920 ;
        RECT 2130.360 255.380 2130.620 255.640 ;
        RECT 2131.280 255.380 2131.540 255.640 ;
        RECT 2130.360 207.100 2130.620 207.360 ;
        RECT 2131.280 207.100 2131.540 207.360 ;
        RECT 2130.360 158.820 2130.620 159.080 ;
        RECT 2131.280 158.820 2131.540 159.080 ;
        RECT 2130.360 62.260 2130.620 62.520 ;
        RECT 2131.280 62.260 2131.540 62.520 ;
        RECT 2130.360 24.520 2130.620 24.780 ;
        RECT 2845.200 24.520 2845.460 24.780 ;
      LAYER met2 ;
        RECT 2131.510 600.170 2131.790 604.000 ;
        RECT 2130.880 600.030 2131.790 600.170 ;
        RECT 2130.880 592.610 2131.020 600.030 ;
        RECT 2131.510 600.000 2131.790 600.030 ;
        RECT 2129.900 592.290 2130.160 592.610 ;
        RECT 2130.820 592.290 2131.080 592.610 ;
        RECT 2129.960 545.350 2130.100 592.290 ;
        RECT 2129.900 545.030 2130.160 545.350 ;
        RECT 2131.280 545.030 2131.540 545.350 ;
        RECT 2131.340 497.410 2131.480 545.030 ;
        RECT 2131.280 497.090 2131.540 497.410 ;
        RECT 2130.360 496.750 2130.620 497.070 ;
        RECT 2130.420 448.790 2130.560 496.750 ;
        RECT 2130.360 448.470 2130.620 448.790 ;
        RECT 2131.280 448.470 2131.540 448.790 ;
        RECT 2131.340 400.850 2131.480 448.470 ;
        RECT 2131.280 400.530 2131.540 400.850 ;
        RECT 2130.360 400.190 2130.620 400.510 ;
        RECT 2130.420 352.230 2130.560 400.190 ;
        RECT 2130.360 351.910 2130.620 352.230 ;
        RECT 2131.280 351.910 2131.540 352.230 ;
        RECT 2131.340 304.290 2131.480 351.910 ;
        RECT 2131.280 303.970 2131.540 304.290 ;
        RECT 2130.360 303.630 2130.620 303.950 ;
        RECT 2130.420 255.670 2130.560 303.630 ;
        RECT 2130.360 255.350 2130.620 255.670 ;
        RECT 2131.280 255.350 2131.540 255.670 ;
        RECT 2131.340 207.390 2131.480 255.350 ;
        RECT 2130.360 207.070 2130.620 207.390 ;
        RECT 2131.280 207.070 2131.540 207.390 ;
        RECT 2130.420 159.110 2130.560 207.070 ;
        RECT 2130.360 158.790 2130.620 159.110 ;
        RECT 2131.280 158.790 2131.540 159.110 ;
        RECT 2131.340 62.550 2131.480 158.790 ;
        RECT 2130.360 62.230 2130.620 62.550 ;
        RECT 2131.280 62.230 2131.540 62.550 ;
        RECT 2130.420 24.810 2130.560 62.230 ;
        RECT 2130.360 24.490 2130.620 24.810 ;
        RECT 2845.200 24.490 2845.460 24.810 ;
        RECT 2845.260 2.400 2845.400 24.490 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2140.680 598.980 2141.000 599.040 ;
        RECT 2145.510 598.980 2145.830 599.040 ;
        RECT 2140.680 598.840 2145.830 598.980 ;
        RECT 2140.680 598.780 2141.000 598.840 ;
        RECT 2145.510 598.780 2145.830 598.840 ;
        RECT 2145.510 25.060 2145.830 25.120 ;
        RECT 2863.110 25.060 2863.430 25.120 ;
        RECT 2145.510 24.920 2863.430 25.060 ;
        RECT 2145.510 24.860 2145.830 24.920 ;
        RECT 2863.110 24.860 2863.430 24.920 ;
      LAYER via ;
        RECT 2140.710 598.780 2140.970 599.040 ;
        RECT 2145.540 598.780 2145.800 599.040 ;
        RECT 2145.540 24.860 2145.800 25.120 ;
        RECT 2863.140 24.860 2863.400 25.120 ;
      LAYER met2 ;
        RECT 2140.710 600.000 2140.990 604.000 ;
        RECT 2140.770 599.070 2140.910 600.000 ;
        RECT 2140.710 598.750 2140.970 599.070 ;
        RECT 2145.540 598.750 2145.800 599.070 ;
        RECT 2145.600 25.150 2145.740 598.750 ;
        RECT 2145.540 24.830 2145.800 25.150 ;
        RECT 2863.140 24.830 2863.400 25.150 ;
        RECT 2863.200 2.400 2863.340 24.830 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2152.410 24.380 2152.730 24.440 ;
        RECT 2881.050 24.380 2881.370 24.440 ;
        RECT 2152.410 24.240 2881.370 24.380 ;
        RECT 2152.410 24.180 2152.730 24.240 ;
        RECT 2881.050 24.180 2881.370 24.240 ;
      LAYER via ;
        RECT 2152.440 24.180 2152.700 24.440 ;
        RECT 2881.080 24.180 2881.340 24.440 ;
      LAYER met2 ;
        RECT 2149.910 600.170 2150.190 604.000 ;
        RECT 2149.910 600.030 2152.640 600.170 ;
        RECT 2149.910 600.000 2150.190 600.030 ;
        RECT 2152.500 24.470 2152.640 600.030 ;
        RECT 2152.440 24.150 2152.700 24.470 ;
        RECT 2881.080 24.150 2881.340 24.470 ;
        RECT 2881.140 2.400 2881.280 24.150 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2159.310 24.040 2159.630 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 2159.310 23.900 2899.310 24.040 ;
        RECT 2159.310 23.840 2159.630 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 2159.340 23.840 2159.600 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 2159.110 600.000 2159.390 604.000 ;
        RECT 2159.170 598.810 2159.310 600.000 ;
        RECT 2159.170 598.670 2159.540 598.810 ;
        RECT 2159.400 24.130 2159.540 598.670 ;
        RECT 2159.340 23.810 2159.600 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.400 2899.220 23.810 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 846.930 17.920 847.250 17.980 ;
        RECT 1104.070 17.920 1104.390 17.980 ;
        RECT 846.930 17.780 1104.390 17.920 ;
        RECT 846.930 17.720 847.250 17.780 ;
        RECT 1104.070 17.720 1104.390 17.780 ;
      LAYER via ;
        RECT 846.960 17.720 847.220 17.980 ;
        RECT 1104.100 17.720 1104.360 17.980 ;
      LAYER met2 ;
        RECT 1105.250 600.170 1105.530 604.000 ;
        RECT 1104.160 600.030 1105.530 600.170 ;
        RECT 1104.160 18.010 1104.300 600.030 ;
        RECT 1105.250 600.000 1105.530 600.030 ;
        RECT 846.960 17.690 847.220 18.010 ;
        RECT 1104.100 17.690 1104.360 18.010 ;
        RECT 847.020 2.400 847.160 17.690 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 900.290 18.260 900.610 18.320 ;
        RECT 1111.890 18.260 1112.210 18.320 ;
        RECT 900.290 18.120 1112.210 18.260 ;
        RECT 900.290 18.060 900.610 18.120 ;
        RECT 1111.890 18.060 1112.210 18.120 ;
        RECT 864.870 15.880 865.190 15.940 ;
        RECT 900.290 15.880 900.610 15.940 ;
        RECT 864.870 15.740 900.610 15.880 ;
        RECT 864.870 15.680 865.190 15.740 ;
        RECT 900.290 15.680 900.610 15.740 ;
      LAYER via ;
        RECT 900.320 18.060 900.580 18.320 ;
        RECT 1111.920 18.060 1112.180 18.320 ;
        RECT 864.900 15.680 865.160 15.940 ;
        RECT 900.320 15.680 900.580 15.940 ;
      LAYER met2 ;
        RECT 1114.450 600.170 1114.730 604.000 ;
        RECT 1111.980 600.030 1114.730 600.170 ;
        RECT 1111.980 18.350 1112.120 600.030 ;
        RECT 1114.450 600.000 1114.730 600.030 ;
        RECT 900.320 18.030 900.580 18.350 ;
        RECT 1111.920 18.030 1112.180 18.350 ;
        RECT 900.380 15.970 900.520 18.030 ;
        RECT 864.900 15.650 865.160 15.970 ;
        RECT 900.320 15.650 900.580 15.970 ;
        RECT 864.960 2.400 865.100 15.650 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1117.870 483.040 1118.190 483.100 ;
        RECT 1118.330 483.040 1118.650 483.100 ;
        RECT 1117.870 482.900 1118.650 483.040 ;
        RECT 1117.870 482.840 1118.190 482.900 ;
        RECT 1118.330 482.840 1118.650 482.900 ;
        RECT 1117.410 410.620 1117.730 410.680 ;
        RECT 1118.790 410.620 1119.110 410.680 ;
        RECT 1117.410 410.480 1119.110 410.620 ;
        RECT 1117.410 410.420 1117.730 410.480 ;
        RECT 1118.790 410.420 1119.110 410.480 ;
        RECT 1117.410 386.480 1117.730 386.540 ;
        RECT 1118.330 386.480 1118.650 386.540 ;
        RECT 1117.410 386.340 1118.650 386.480 ;
        RECT 1117.410 386.280 1117.730 386.340 ;
        RECT 1118.330 386.280 1118.650 386.340 ;
        RECT 1118.330 351.940 1118.650 352.200 ;
        RECT 1118.420 351.520 1118.560 351.940 ;
        RECT 1118.330 351.260 1118.650 351.520 ;
        RECT 1117.870 331.060 1118.190 331.120 ;
        RECT 1118.330 331.060 1118.650 331.120 ;
        RECT 1117.870 330.920 1118.650 331.060 ;
        RECT 1117.870 330.860 1118.190 330.920 ;
        RECT 1118.330 330.860 1118.650 330.920 ;
        RECT 1117.410 193.020 1117.730 193.080 ;
        RECT 1118.330 193.020 1118.650 193.080 ;
        RECT 1117.410 192.880 1118.650 193.020 ;
        RECT 1117.410 192.820 1117.730 192.880 ;
        RECT 1118.330 192.820 1118.650 192.880 ;
        RECT 1117.410 145.080 1117.730 145.140 ;
        RECT 1118.330 145.080 1118.650 145.140 ;
        RECT 1117.410 144.940 1118.650 145.080 ;
        RECT 1117.410 144.880 1117.730 144.940 ;
        RECT 1118.330 144.880 1118.650 144.940 ;
        RECT 1117.870 22.000 1118.190 22.060 ;
        RECT 1021.820 21.860 1118.190 22.000 ;
        RECT 979.410 21.320 979.730 21.380 ;
        RECT 1000.570 21.320 1000.890 21.380 ;
        RECT 979.410 21.180 1000.890 21.320 ;
        RECT 979.410 21.120 979.730 21.180 ;
        RECT 1000.570 21.120 1000.890 21.180 ;
        RECT 1000.570 20.640 1000.890 20.700 ;
        RECT 1021.820 20.640 1021.960 21.860 ;
        RECT 1117.870 21.800 1118.190 21.860 ;
        RECT 1000.570 20.500 1021.960 20.640 ;
        RECT 1000.570 20.440 1000.890 20.500 ;
        RECT 882.350 20.300 882.670 20.360 ;
        RECT 979.410 20.300 979.730 20.360 ;
        RECT 882.350 20.160 979.730 20.300 ;
        RECT 882.350 20.100 882.670 20.160 ;
        RECT 979.410 20.100 979.730 20.160 ;
      LAYER via ;
        RECT 1117.900 482.840 1118.160 483.100 ;
        RECT 1118.360 482.840 1118.620 483.100 ;
        RECT 1117.440 410.420 1117.700 410.680 ;
        RECT 1118.820 410.420 1119.080 410.680 ;
        RECT 1117.440 386.280 1117.700 386.540 ;
        RECT 1118.360 386.280 1118.620 386.540 ;
        RECT 1118.360 351.940 1118.620 352.200 ;
        RECT 1118.360 351.260 1118.620 351.520 ;
        RECT 1117.900 330.860 1118.160 331.120 ;
        RECT 1118.360 330.860 1118.620 331.120 ;
        RECT 1117.440 192.820 1117.700 193.080 ;
        RECT 1118.360 192.820 1118.620 193.080 ;
        RECT 1117.440 144.880 1117.700 145.140 ;
        RECT 1118.360 144.880 1118.620 145.140 ;
        RECT 979.440 21.120 979.700 21.380 ;
        RECT 1000.600 21.120 1000.860 21.380 ;
        RECT 1000.600 20.440 1000.860 20.700 ;
        RECT 1117.900 21.800 1118.160 22.060 ;
        RECT 882.380 20.100 882.640 20.360 ;
        RECT 979.440 20.100 979.700 20.360 ;
      LAYER met2 ;
        RECT 1123.190 600.170 1123.470 604.000 ;
        RECT 1121.180 600.030 1123.470 600.170 ;
        RECT 1121.180 569.570 1121.320 600.030 ;
        RECT 1123.190 600.000 1123.470 600.030 ;
        RECT 1118.420 569.430 1121.320 569.570 ;
        RECT 1118.420 507.010 1118.560 569.430 ;
        RECT 1117.960 506.870 1118.560 507.010 ;
        RECT 1117.960 483.130 1118.100 506.870 ;
        RECT 1117.900 482.810 1118.160 483.130 ;
        RECT 1118.360 482.810 1118.620 483.130 ;
        RECT 1118.420 434.930 1118.560 482.810 ;
        RECT 1118.420 434.790 1119.020 434.930 ;
        RECT 1118.880 410.710 1119.020 434.790 ;
        RECT 1117.440 410.390 1117.700 410.710 ;
        RECT 1118.820 410.390 1119.080 410.710 ;
        RECT 1117.500 386.570 1117.640 410.390 ;
        RECT 1117.440 386.250 1117.700 386.570 ;
        RECT 1118.360 386.250 1118.620 386.570 ;
        RECT 1118.420 352.230 1118.560 386.250 ;
        RECT 1118.360 351.910 1118.620 352.230 ;
        RECT 1118.360 351.230 1118.620 351.550 ;
        RECT 1118.420 331.150 1118.560 351.230 ;
        RECT 1117.900 330.830 1118.160 331.150 ;
        RECT 1118.360 330.830 1118.620 331.150 ;
        RECT 1117.960 264.930 1118.100 330.830 ;
        RECT 1117.960 264.790 1118.560 264.930 ;
        RECT 1118.420 193.110 1118.560 264.790 ;
        RECT 1117.440 192.790 1117.700 193.110 ;
        RECT 1118.360 192.790 1118.620 193.110 ;
        RECT 1117.500 145.170 1117.640 192.790 ;
        RECT 1117.440 144.850 1117.700 145.170 ;
        RECT 1118.360 144.850 1118.620 145.170 ;
        RECT 1118.420 62.290 1118.560 144.850 ;
        RECT 1117.960 62.150 1118.560 62.290 ;
        RECT 1117.960 22.090 1118.100 62.150 ;
        RECT 1117.900 21.770 1118.160 22.090 ;
        RECT 979.440 21.090 979.700 21.410 ;
        RECT 1000.600 21.090 1000.860 21.410 ;
        RECT 979.500 20.390 979.640 21.090 ;
        RECT 1000.660 20.730 1000.800 21.090 ;
        RECT 1000.600 20.410 1000.860 20.730 ;
        RECT 882.380 20.070 882.640 20.390 ;
        RECT 979.440 20.070 979.700 20.390 ;
        RECT 882.440 10.610 882.580 20.070 ;
        RECT 882.440 10.470 883.040 10.610 ;
        RECT 882.900 2.400 883.040 10.470 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1021.270 23.020 1021.590 23.080 ;
        RECT 1132.130 23.020 1132.450 23.080 ;
        RECT 1021.270 22.880 1132.450 23.020 ;
        RECT 1021.270 22.820 1021.590 22.880 ;
        RECT 1132.130 22.820 1132.450 22.880 ;
        RECT 900.750 15.880 901.070 15.940 ;
        RECT 1021.270 15.880 1021.590 15.940 ;
        RECT 900.750 15.740 1021.590 15.880 ;
        RECT 900.750 15.680 901.070 15.740 ;
        RECT 1021.270 15.680 1021.590 15.740 ;
      LAYER via ;
        RECT 1021.300 22.820 1021.560 23.080 ;
        RECT 1132.160 22.820 1132.420 23.080 ;
        RECT 900.780 15.680 901.040 15.940 ;
        RECT 1021.300 15.680 1021.560 15.940 ;
      LAYER met2 ;
        RECT 1132.390 600.000 1132.670 604.000 ;
        RECT 1132.450 598.810 1132.590 600.000 ;
        RECT 1132.220 598.670 1132.590 598.810 ;
        RECT 1132.220 23.110 1132.360 598.670 ;
        RECT 1021.300 22.790 1021.560 23.110 ;
        RECT 1132.160 22.790 1132.420 23.110 ;
        RECT 1021.360 15.970 1021.500 22.790 ;
        RECT 900.780 15.650 901.040 15.970 ;
        RECT 1021.300 15.650 1021.560 15.970 ;
        RECT 900.840 2.400 900.980 15.650 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.570 386.480 1138.890 386.540 ;
        RECT 1139.490 386.480 1139.810 386.540 ;
        RECT 1138.570 386.340 1139.810 386.480 ;
        RECT 1138.570 386.280 1138.890 386.340 ;
        RECT 1139.490 386.280 1139.810 386.340 ;
        RECT 1139.030 303.520 1139.350 303.580 ;
        RECT 1139.950 303.520 1140.270 303.580 ;
        RECT 1139.030 303.380 1140.270 303.520 ;
        RECT 1139.030 303.320 1139.350 303.380 ;
        RECT 1139.950 303.320 1140.270 303.380 ;
        RECT 1139.950 252.660 1140.270 252.920 ;
        RECT 1140.040 252.240 1140.180 252.660 ;
        RECT 1139.950 251.980 1140.270 252.240 ;
        RECT 1138.570 193.360 1138.890 193.420 ;
        RECT 1139.950 193.360 1140.270 193.420 ;
        RECT 1138.570 193.220 1140.270 193.360 ;
        RECT 1138.570 193.160 1138.890 193.220 ;
        RECT 1139.950 193.160 1140.270 193.220 ;
        RECT 1139.030 110.400 1139.350 110.460 ;
        RECT 1139.950 110.400 1140.270 110.460 ;
        RECT 1139.030 110.260 1140.270 110.400 ;
        RECT 1139.030 110.200 1139.350 110.260 ;
        RECT 1139.950 110.200 1140.270 110.260 ;
        RECT 1139.030 96.460 1139.350 96.520 ;
        RECT 1139.950 96.460 1140.270 96.520 ;
        RECT 1139.030 96.320 1140.270 96.460 ;
        RECT 1139.030 96.260 1139.350 96.320 ;
        RECT 1139.950 96.260 1140.270 96.320 ;
        RECT 1014.370 23.360 1014.690 23.420 ;
        RECT 1139.950 23.360 1140.270 23.420 ;
        RECT 1014.370 23.220 1140.270 23.360 ;
        RECT 1014.370 23.160 1014.690 23.220 ;
        RECT 1139.950 23.160 1140.270 23.220 ;
        RECT 918.690 20.640 919.010 20.700 ;
        RECT 918.690 20.500 989.760 20.640 ;
        RECT 918.690 20.440 919.010 20.500 ;
        RECT 989.620 19.960 989.760 20.500 ;
        RECT 1014.370 19.960 1014.690 20.020 ;
        RECT 989.620 19.820 1014.690 19.960 ;
        RECT 1014.370 19.760 1014.690 19.820 ;
      LAYER via ;
        RECT 1138.600 386.280 1138.860 386.540 ;
        RECT 1139.520 386.280 1139.780 386.540 ;
        RECT 1139.060 303.320 1139.320 303.580 ;
        RECT 1139.980 303.320 1140.240 303.580 ;
        RECT 1139.980 252.660 1140.240 252.920 ;
        RECT 1139.980 251.980 1140.240 252.240 ;
        RECT 1138.600 193.160 1138.860 193.420 ;
        RECT 1139.980 193.160 1140.240 193.420 ;
        RECT 1139.060 110.200 1139.320 110.460 ;
        RECT 1139.980 110.200 1140.240 110.460 ;
        RECT 1139.060 96.260 1139.320 96.520 ;
        RECT 1139.980 96.260 1140.240 96.520 ;
        RECT 1014.400 23.160 1014.660 23.420 ;
        RECT 1139.980 23.160 1140.240 23.420 ;
        RECT 918.720 20.440 918.980 20.700 ;
        RECT 1014.400 19.760 1014.660 20.020 ;
      LAYER met2 ;
        RECT 1141.590 600.170 1141.870 604.000 ;
        RECT 1139.580 600.030 1141.870 600.170 ;
        RECT 1139.580 386.570 1139.720 600.030 ;
        RECT 1141.590 600.000 1141.870 600.030 ;
        RECT 1138.600 386.250 1138.860 386.570 ;
        RECT 1139.520 386.250 1139.780 386.570 ;
        RECT 1138.660 351.290 1138.800 386.250 ;
        RECT 1138.660 351.150 1139.260 351.290 ;
        RECT 1139.120 303.610 1139.260 351.150 ;
        RECT 1139.060 303.290 1139.320 303.610 ;
        RECT 1139.980 303.290 1140.240 303.610 ;
        RECT 1140.040 252.950 1140.180 303.290 ;
        RECT 1139.980 252.630 1140.240 252.950 ;
        RECT 1139.980 251.950 1140.240 252.270 ;
        RECT 1140.040 193.450 1140.180 251.950 ;
        RECT 1138.600 193.130 1138.860 193.450 ;
        RECT 1139.980 193.130 1140.240 193.450 ;
        RECT 1138.660 158.170 1138.800 193.130 ;
        RECT 1138.660 158.030 1139.260 158.170 ;
        RECT 1139.120 110.490 1139.260 158.030 ;
        RECT 1139.060 110.170 1139.320 110.490 ;
        RECT 1139.980 110.170 1140.240 110.490 ;
        RECT 1140.040 96.550 1140.180 110.170 ;
        RECT 1139.060 96.230 1139.320 96.550 ;
        RECT 1139.980 96.230 1140.240 96.550 ;
        RECT 1139.120 58.890 1139.260 96.230 ;
        RECT 1139.120 58.750 1140.180 58.890 ;
        RECT 1140.040 23.450 1140.180 58.750 ;
        RECT 1014.400 23.130 1014.660 23.450 ;
        RECT 1139.980 23.130 1140.240 23.450 ;
        RECT 918.720 20.410 918.980 20.730 ;
        RECT 918.780 2.400 918.920 20.410 ;
        RECT 1014.460 20.050 1014.600 23.130 ;
        RECT 1014.400 19.730 1014.660 20.050 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 936.170 19.280 936.490 19.340 ;
        RECT 936.170 19.140 1081.760 19.280 ;
        RECT 936.170 19.080 936.490 19.140 ;
        RECT 1081.620 18.940 1081.760 19.140 ;
        RECT 1146.390 18.940 1146.710 19.000 ;
        RECT 1081.620 18.800 1146.710 18.940 ;
        RECT 1146.390 18.740 1146.710 18.800 ;
      LAYER via ;
        RECT 936.200 19.080 936.460 19.340 ;
        RECT 1146.420 18.740 1146.680 19.000 ;
      LAYER met2 ;
        RECT 1150.790 600.170 1151.070 604.000 ;
        RECT 1148.780 600.030 1151.070 600.170 ;
        RECT 1148.780 592.010 1148.920 600.030 ;
        RECT 1150.790 600.000 1151.070 600.030 ;
        RECT 1146.940 591.870 1148.920 592.010 ;
        RECT 1146.940 569.570 1147.080 591.870 ;
        RECT 1146.480 569.430 1147.080 569.570 ;
        RECT 936.200 19.050 936.460 19.370 ;
        RECT 936.260 2.400 936.400 19.050 ;
        RECT 1146.480 19.030 1146.620 569.430 ;
        RECT 1146.420 18.710 1146.680 19.030 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1033.690 27.440 1034.010 27.500 ;
        RECT 1159.730 27.440 1160.050 27.500 ;
        RECT 1033.690 27.300 1160.050 27.440 ;
        RECT 1033.690 27.240 1034.010 27.300 ;
        RECT 1159.730 27.240 1160.050 27.300 ;
        RECT 954.110 16.900 954.430 16.960 ;
        RECT 1003.790 16.900 1004.110 16.960 ;
        RECT 954.110 16.760 1004.110 16.900 ;
        RECT 954.110 16.700 954.430 16.760 ;
        RECT 1003.790 16.700 1004.110 16.760 ;
        RECT 1003.790 14.860 1004.110 14.920 ;
        RECT 1033.690 14.860 1034.010 14.920 ;
        RECT 1003.790 14.720 1034.010 14.860 ;
        RECT 1003.790 14.660 1004.110 14.720 ;
        RECT 1033.690 14.660 1034.010 14.720 ;
      LAYER via ;
        RECT 1033.720 27.240 1033.980 27.500 ;
        RECT 1159.760 27.240 1160.020 27.500 ;
        RECT 954.140 16.700 954.400 16.960 ;
        RECT 1003.820 16.700 1004.080 16.960 ;
        RECT 1003.820 14.660 1004.080 14.920 ;
        RECT 1033.720 14.660 1033.980 14.920 ;
      LAYER met2 ;
        RECT 1159.990 600.000 1160.270 604.000 ;
        RECT 1160.050 598.810 1160.190 600.000 ;
        RECT 1159.820 598.670 1160.190 598.810 ;
        RECT 1159.820 27.530 1159.960 598.670 ;
        RECT 1033.720 27.210 1033.980 27.530 ;
        RECT 1159.760 27.210 1160.020 27.530 ;
        RECT 954.140 16.670 954.400 16.990 ;
        RECT 1003.820 16.670 1004.080 16.990 ;
        RECT 954.200 2.400 954.340 16.670 ;
        RECT 1003.880 14.950 1004.020 16.670 ;
        RECT 1033.780 14.950 1033.920 27.210 ;
        RECT 1003.820 14.630 1004.080 14.950 ;
        RECT 1033.720 14.630 1033.980 14.950 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1036.910 23.700 1037.230 23.760 ;
        RECT 1166.630 23.700 1166.950 23.760 ;
        RECT 1036.910 23.560 1166.950 23.700 ;
        RECT 1036.910 23.500 1037.230 23.560 ;
        RECT 1166.630 23.500 1166.950 23.560 ;
        RECT 972.050 15.200 972.370 15.260 ;
        RECT 1036.910 15.200 1037.230 15.260 ;
        RECT 972.050 15.060 1037.230 15.200 ;
        RECT 972.050 15.000 972.370 15.060 ;
        RECT 1036.910 15.000 1037.230 15.060 ;
      LAYER via ;
        RECT 1036.940 23.500 1037.200 23.760 ;
        RECT 1166.660 23.500 1166.920 23.760 ;
        RECT 972.080 15.000 972.340 15.260 ;
        RECT 1036.940 15.000 1037.200 15.260 ;
      LAYER met2 ;
        RECT 1169.190 600.170 1169.470 604.000 ;
        RECT 1166.720 600.030 1169.470 600.170 ;
        RECT 1166.720 23.790 1166.860 600.030 ;
        RECT 1169.190 600.000 1169.470 600.030 ;
        RECT 1036.940 23.470 1037.200 23.790 ;
        RECT 1166.660 23.470 1166.920 23.790 ;
        RECT 1037.000 15.290 1037.140 23.470 ;
        RECT 972.080 14.970 972.340 15.290 ;
        RECT 1036.940 14.970 1037.200 15.290 ;
        RECT 972.140 2.400 972.280 14.970 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1002.410 497.320 1002.730 497.380 ;
        RECT 1001.580 497.180 1002.730 497.320 ;
        RECT 1001.580 497.040 1001.720 497.180 ;
        RECT 1002.410 497.120 1002.730 497.180 ;
        RECT 1001.490 496.780 1001.810 497.040 ;
        RECT 1000.570 451.760 1000.890 451.820 ;
        RECT 1001.490 451.760 1001.810 451.820 ;
        RECT 1000.570 451.620 1001.810 451.760 ;
        RECT 1000.570 451.560 1000.890 451.620 ;
        RECT 1001.490 451.560 1001.810 451.620 ;
        RECT 650.970 36.280 651.290 36.340 ;
        RECT 1000.570 36.280 1000.890 36.340 ;
        RECT 650.970 36.140 1000.890 36.280 ;
        RECT 650.970 36.080 651.290 36.140 ;
        RECT 1000.570 36.080 1000.890 36.140 ;
      LAYER via ;
        RECT 1002.440 497.120 1002.700 497.380 ;
        RECT 1001.520 496.780 1001.780 497.040 ;
        RECT 1000.600 451.560 1000.860 451.820 ;
        RECT 1001.520 451.560 1001.780 451.820 ;
        RECT 651.000 36.080 651.260 36.340 ;
        RECT 1000.600 36.080 1000.860 36.340 ;
      LAYER met2 ;
        RECT 1004.050 600.170 1004.330 604.000 ;
        RECT 1002.500 600.030 1004.330 600.170 ;
        RECT 1002.500 497.410 1002.640 600.030 ;
        RECT 1004.050 600.000 1004.330 600.030 ;
        RECT 1002.440 497.090 1002.700 497.410 ;
        RECT 1001.520 496.750 1001.780 497.070 ;
        RECT 1001.580 451.850 1001.720 496.750 ;
        RECT 1000.600 451.530 1000.860 451.850 ;
        RECT 1001.520 451.530 1001.780 451.850 ;
        RECT 1000.660 36.370 1000.800 451.530 ;
        RECT 651.000 36.050 651.260 36.370 ;
        RECT 1000.600 36.050 1000.860 36.370 ;
        RECT 651.060 2.400 651.200 36.050 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1173.530 496.780 1173.850 497.040 ;
        RECT 1173.070 496.640 1173.390 496.700 ;
        RECT 1173.620 496.640 1173.760 496.780 ;
        RECT 1173.070 496.500 1173.760 496.640 ;
        RECT 1173.070 496.440 1173.390 496.500 ;
        RECT 1173.530 427.620 1173.850 427.680 ;
        RECT 1173.990 427.620 1174.310 427.680 ;
        RECT 1173.530 427.480 1174.310 427.620 ;
        RECT 1173.530 427.420 1173.850 427.480 ;
        RECT 1173.990 427.420 1174.310 427.480 ;
        RECT 1173.530 338.200 1173.850 338.260 ;
        RECT 1173.990 338.200 1174.310 338.260 ;
        RECT 1173.530 338.060 1174.310 338.200 ;
        RECT 1173.530 338.000 1173.850 338.060 ;
        RECT 1173.990 338.000 1174.310 338.060 ;
        RECT 1173.070 282.780 1173.390 282.840 ;
        RECT 1173.990 282.780 1174.310 282.840 ;
        RECT 1173.070 282.640 1174.310 282.780 ;
        RECT 1173.070 282.580 1173.390 282.640 ;
        RECT 1173.990 282.580 1174.310 282.640 ;
        RECT 1173.990 186.220 1174.310 186.280 ;
        RECT 1174.910 186.220 1175.230 186.280 ;
        RECT 1173.990 186.080 1175.230 186.220 ;
        RECT 1173.990 186.020 1174.310 186.080 ;
        RECT 1174.910 186.020 1175.230 186.080 ;
        RECT 1173.530 138.280 1173.850 138.340 ;
        RECT 1174.910 138.280 1175.230 138.340 ;
        RECT 1173.530 138.140 1175.230 138.280 ;
        RECT 1173.530 138.080 1173.850 138.140 ;
        RECT 1174.910 138.080 1175.230 138.140 ;
        RECT 1173.070 89.660 1173.390 89.720 ;
        RECT 1173.530 89.660 1173.850 89.720 ;
        RECT 1173.070 89.520 1173.850 89.660 ;
        RECT 1173.070 89.460 1173.390 89.520 ;
        RECT 1173.530 89.460 1173.850 89.520 ;
        RECT 1173.070 41.720 1173.390 41.780 ;
        RECT 1173.990 41.720 1174.310 41.780 ;
        RECT 1173.070 41.580 1174.310 41.720 ;
        RECT 1173.070 41.520 1173.390 41.580 ;
        RECT 1173.990 41.520 1174.310 41.580 ;
        RECT 989.990 31.860 990.310 31.920 ;
        RECT 1173.990 31.860 1174.310 31.920 ;
        RECT 989.990 31.720 1174.310 31.860 ;
        RECT 989.990 31.660 990.310 31.720 ;
        RECT 1173.990 31.660 1174.310 31.720 ;
      LAYER via ;
        RECT 1173.560 496.780 1173.820 497.040 ;
        RECT 1173.100 496.440 1173.360 496.700 ;
        RECT 1173.560 427.420 1173.820 427.680 ;
        RECT 1174.020 427.420 1174.280 427.680 ;
        RECT 1173.560 338.000 1173.820 338.260 ;
        RECT 1174.020 338.000 1174.280 338.260 ;
        RECT 1173.100 282.580 1173.360 282.840 ;
        RECT 1174.020 282.580 1174.280 282.840 ;
        RECT 1174.020 186.020 1174.280 186.280 ;
        RECT 1174.940 186.020 1175.200 186.280 ;
        RECT 1173.560 138.080 1173.820 138.340 ;
        RECT 1174.940 138.080 1175.200 138.340 ;
        RECT 1173.100 89.460 1173.360 89.720 ;
        RECT 1173.560 89.460 1173.820 89.720 ;
        RECT 1173.100 41.520 1173.360 41.780 ;
        RECT 1174.020 41.520 1174.280 41.780 ;
        RECT 990.020 31.660 990.280 31.920 ;
        RECT 1174.020 31.660 1174.280 31.920 ;
      LAYER met2 ;
        RECT 1178.390 600.850 1178.670 604.000 ;
        RECT 1175.920 600.710 1178.670 600.850 ;
        RECT 1175.920 596.770 1176.060 600.710 ;
        RECT 1178.390 600.000 1178.670 600.710 ;
        RECT 1174.080 596.630 1176.060 596.770 ;
        RECT 1174.080 545.090 1174.220 596.630 ;
        RECT 1173.620 544.950 1174.220 545.090 ;
        RECT 1173.620 497.070 1173.760 544.950 ;
        RECT 1173.560 496.750 1173.820 497.070 ;
        RECT 1173.100 496.410 1173.360 496.730 ;
        RECT 1173.160 483.325 1173.300 496.410 ;
        RECT 1173.090 482.955 1173.370 483.325 ;
        RECT 1174.010 482.955 1174.290 483.325 ;
        RECT 1174.080 448.530 1174.220 482.955 ;
        RECT 1173.620 448.390 1174.220 448.530 ;
        RECT 1173.620 427.710 1173.760 448.390 ;
        RECT 1173.560 427.390 1173.820 427.710 ;
        RECT 1174.020 427.390 1174.280 427.710 ;
        RECT 1174.080 338.290 1174.220 427.390 ;
        RECT 1173.560 337.970 1173.820 338.290 ;
        RECT 1174.020 337.970 1174.280 338.290 ;
        RECT 1173.620 307.090 1173.760 337.970 ;
        RECT 1173.620 306.950 1174.220 307.090 ;
        RECT 1174.080 282.870 1174.220 306.950 ;
        RECT 1173.100 282.550 1173.360 282.870 ;
        RECT 1174.020 282.550 1174.280 282.870 ;
        RECT 1173.160 254.050 1173.300 282.550 ;
        RECT 1173.160 253.910 1174.220 254.050 ;
        RECT 1174.080 234.330 1174.220 253.910 ;
        RECT 1173.160 234.190 1174.220 234.330 ;
        RECT 1173.160 186.845 1173.300 234.190 ;
        RECT 1173.090 186.475 1173.370 186.845 ;
        RECT 1174.010 186.475 1174.290 186.845 ;
        RECT 1174.080 186.310 1174.220 186.475 ;
        RECT 1174.020 185.990 1174.280 186.310 ;
        RECT 1174.940 185.990 1175.200 186.310 ;
        RECT 1175.000 138.370 1175.140 185.990 ;
        RECT 1173.560 138.050 1173.820 138.370 ;
        RECT 1174.940 138.050 1175.200 138.370 ;
        RECT 1173.620 137.770 1173.760 138.050 ;
        RECT 1173.160 137.630 1173.760 137.770 ;
        RECT 1173.160 113.290 1173.300 137.630 ;
        RECT 1173.160 113.150 1173.760 113.290 ;
        RECT 1173.620 89.750 1173.760 113.150 ;
        RECT 1173.100 89.430 1173.360 89.750 ;
        RECT 1173.560 89.430 1173.820 89.750 ;
        RECT 1173.160 41.810 1173.300 89.430 ;
        RECT 1173.100 41.490 1173.360 41.810 ;
        RECT 1174.020 41.490 1174.280 41.810 ;
        RECT 1174.080 31.950 1174.220 41.490 ;
        RECT 990.020 31.630 990.280 31.950 ;
        RECT 1174.020 31.630 1174.280 31.950 ;
        RECT 990.080 2.400 990.220 31.630 ;
        RECT 989.870 -4.800 990.430 2.400 ;
      LAYER via2 ;
        RECT 1173.090 483.000 1173.370 483.280 ;
        RECT 1174.010 483.000 1174.290 483.280 ;
        RECT 1173.090 186.520 1173.370 186.800 ;
        RECT 1174.010 186.520 1174.290 186.800 ;
      LAYER met3 ;
        RECT 1173.065 483.290 1173.395 483.305 ;
        RECT 1173.985 483.290 1174.315 483.305 ;
        RECT 1173.065 482.990 1174.315 483.290 ;
        RECT 1173.065 482.975 1173.395 482.990 ;
        RECT 1173.985 482.975 1174.315 482.990 ;
        RECT 1173.065 186.810 1173.395 186.825 ;
        RECT 1173.985 186.810 1174.315 186.825 ;
        RECT 1173.065 186.510 1174.315 186.810 ;
        RECT 1173.065 186.495 1173.395 186.510 ;
        RECT 1173.985 186.495 1174.315 186.510 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.470 32.200 1007.790 32.260 ;
        RECT 1187.330 32.200 1187.650 32.260 ;
        RECT 1007.470 32.060 1187.650 32.200 ;
        RECT 1007.470 32.000 1007.790 32.060 ;
        RECT 1187.330 32.000 1187.650 32.060 ;
      LAYER via ;
        RECT 1007.500 32.000 1007.760 32.260 ;
        RECT 1187.360 32.000 1187.620 32.260 ;
      LAYER met2 ;
        RECT 1187.590 600.000 1187.870 604.000 ;
        RECT 1187.650 598.810 1187.790 600.000 ;
        RECT 1187.420 598.670 1187.790 598.810 ;
        RECT 1187.420 387.445 1187.560 598.670 ;
        RECT 1187.350 387.075 1187.630 387.445 ;
        RECT 1187.350 385.715 1187.630 386.085 ;
        RECT 1187.420 32.290 1187.560 385.715 ;
        RECT 1007.500 31.970 1007.760 32.290 ;
        RECT 1187.360 31.970 1187.620 32.290 ;
        RECT 1007.560 2.400 1007.700 31.970 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
      LAYER via2 ;
        RECT 1187.350 387.120 1187.630 387.400 ;
        RECT 1187.350 385.760 1187.630 386.040 ;
      LAYER met3 ;
        RECT 1187.325 387.410 1187.655 387.425 ;
        RECT 1187.110 387.095 1187.655 387.410 ;
        RECT 1187.110 386.065 1187.410 387.095 ;
        RECT 1187.110 385.750 1187.655 386.065 ;
        RECT 1187.325 385.735 1187.655 385.750 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.510 24.040 1041.830 24.100 ;
        RECT 1194.230 24.040 1194.550 24.100 ;
        RECT 1041.510 23.900 1194.550 24.040 ;
        RECT 1041.510 23.840 1041.830 23.900 ;
        RECT 1194.230 23.840 1194.550 23.900 ;
        RECT 1025.410 14.180 1025.730 14.240 ;
        RECT 1041.510 14.180 1041.830 14.240 ;
        RECT 1025.410 14.040 1041.830 14.180 ;
        RECT 1025.410 13.980 1025.730 14.040 ;
        RECT 1041.510 13.980 1041.830 14.040 ;
      LAYER via ;
        RECT 1041.540 23.840 1041.800 24.100 ;
        RECT 1194.260 23.840 1194.520 24.100 ;
        RECT 1025.440 13.980 1025.700 14.240 ;
        RECT 1041.540 13.980 1041.800 14.240 ;
      LAYER met2 ;
        RECT 1196.790 600.170 1197.070 604.000 ;
        RECT 1194.320 600.030 1197.070 600.170 ;
        RECT 1194.320 24.130 1194.460 600.030 ;
        RECT 1196.790 600.000 1197.070 600.030 ;
        RECT 1041.540 23.810 1041.800 24.130 ;
        RECT 1194.260 23.810 1194.520 24.130 ;
        RECT 1041.600 14.270 1041.740 23.810 ;
        RECT 1025.440 13.950 1025.700 14.270 ;
        RECT 1041.540 13.950 1041.800 14.270 ;
        RECT 1025.500 2.400 1025.640 13.950 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1201.130 496.780 1201.450 497.040 ;
        RECT 1200.670 496.640 1200.990 496.700 ;
        RECT 1201.220 496.640 1201.360 496.780 ;
        RECT 1200.670 496.500 1201.360 496.640 ;
        RECT 1200.670 496.440 1200.990 496.500 ;
        RECT 1201.130 427.620 1201.450 427.680 ;
        RECT 1202.510 427.620 1202.830 427.680 ;
        RECT 1201.130 427.480 1202.830 427.620 ;
        RECT 1201.130 427.420 1201.450 427.480 ;
        RECT 1202.510 427.420 1202.830 427.480 ;
        RECT 1201.590 379.680 1201.910 379.740 ;
        RECT 1202.510 379.680 1202.830 379.740 ;
        RECT 1201.590 379.540 1202.830 379.680 ;
        RECT 1201.590 379.480 1201.910 379.540 ;
        RECT 1202.510 379.480 1202.830 379.540 ;
        RECT 1201.130 331.740 1201.450 331.800 ;
        RECT 1202.510 331.740 1202.830 331.800 ;
        RECT 1201.130 331.600 1202.830 331.740 ;
        RECT 1201.130 331.540 1201.450 331.600 ;
        RECT 1202.510 331.540 1202.830 331.600 ;
        RECT 1201.130 331.060 1201.450 331.120 ;
        RECT 1201.590 331.060 1201.910 331.120 ;
        RECT 1201.130 330.920 1201.910 331.060 ;
        RECT 1201.130 330.860 1201.450 330.920 ;
        RECT 1201.590 330.860 1201.910 330.920 ;
        RECT 1201.590 324.260 1201.910 324.320 ;
        RECT 1202.510 324.260 1202.830 324.320 ;
        RECT 1201.590 324.120 1202.830 324.260 ;
        RECT 1201.590 324.060 1201.910 324.120 ;
        RECT 1202.510 324.060 1202.830 324.120 ;
        RECT 1201.590 276.320 1201.910 276.380 ;
        RECT 1202.510 276.320 1202.830 276.380 ;
        RECT 1201.590 276.180 1202.830 276.320 ;
        RECT 1201.590 276.120 1201.910 276.180 ;
        RECT 1202.510 276.120 1202.830 276.180 ;
        RECT 1201.590 255.380 1201.910 255.640 ;
        RECT 1201.680 254.900 1201.820 255.380 ;
        RECT 1202.050 254.900 1202.370 254.960 ;
        RECT 1201.680 254.760 1202.370 254.900 ;
        RECT 1202.050 254.700 1202.370 254.760 ;
        RECT 1201.130 227.700 1201.450 227.760 ;
        RECT 1202.050 227.700 1202.370 227.760 ;
        RECT 1201.130 227.560 1202.370 227.700 ;
        RECT 1201.130 227.500 1201.450 227.560 ;
        RECT 1202.050 227.500 1202.370 227.560 ;
        RECT 1201.130 179.760 1201.450 179.820 ;
        RECT 1201.590 179.760 1201.910 179.820 ;
        RECT 1201.130 179.620 1201.910 179.760 ;
        RECT 1201.130 179.560 1201.450 179.620 ;
        RECT 1201.590 179.560 1201.910 179.620 ;
        RECT 1201.590 159.020 1201.910 159.080 ;
        RECT 1201.220 158.880 1201.910 159.020 ;
        RECT 1201.220 158.740 1201.360 158.880 ;
        RECT 1201.590 158.820 1201.910 158.880 ;
        RECT 1201.130 158.480 1201.450 158.740 ;
        RECT 1200.670 110.400 1200.990 110.460 ;
        RECT 1201.590 110.400 1201.910 110.460 ;
        RECT 1200.670 110.260 1201.910 110.400 ;
        RECT 1200.670 110.200 1200.990 110.260 ;
        RECT 1201.590 110.200 1201.910 110.260 ;
        RECT 1043.350 24.720 1043.670 24.780 ;
        RECT 1201.590 24.720 1201.910 24.780 ;
        RECT 1043.350 24.580 1201.910 24.720 ;
        RECT 1043.350 24.520 1043.670 24.580 ;
        RECT 1201.590 24.520 1201.910 24.580 ;
      LAYER via ;
        RECT 1201.160 496.780 1201.420 497.040 ;
        RECT 1200.700 496.440 1200.960 496.700 ;
        RECT 1201.160 427.420 1201.420 427.680 ;
        RECT 1202.540 427.420 1202.800 427.680 ;
        RECT 1201.620 379.480 1201.880 379.740 ;
        RECT 1202.540 379.480 1202.800 379.740 ;
        RECT 1201.160 331.540 1201.420 331.800 ;
        RECT 1202.540 331.540 1202.800 331.800 ;
        RECT 1201.160 330.860 1201.420 331.120 ;
        RECT 1201.620 330.860 1201.880 331.120 ;
        RECT 1201.620 324.060 1201.880 324.320 ;
        RECT 1202.540 324.060 1202.800 324.320 ;
        RECT 1201.620 276.120 1201.880 276.380 ;
        RECT 1202.540 276.120 1202.800 276.380 ;
        RECT 1201.620 255.380 1201.880 255.640 ;
        RECT 1202.080 254.700 1202.340 254.960 ;
        RECT 1201.160 227.500 1201.420 227.760 ;
        RECT 1202.080 227.500 1202.340 227.760 ;
        RECT 1201.160 179.560 1201.420 179.820 ;
        RECT 1201.620 179.560 1201.880 179.820 ;
        RECT 1201.620 158.820 1201.880 159.080 ;
        RECT 1201.160 158.480 1201.420 158.740 ;
        RECT 1200.700 110.200 1200.960 110.460 ;
        RECT 1201.620 110.200 1201.880 110.460 ;
        RECT 1043.380 24.520 1043.640 24.780 ;
        RECT 1201.620 24.520 1201.880 24.780 ;
      LAYER met2 ;
        RECT 1205.990 600.850 1206.270 604.000 ;
        RECT 1203.520 600.710 1206.270 600.850 ;
        RECT 1203.520 596.770 1203.660 600.710 ;
        RECT 1205.990 600.000 1206.270 600.710 ;
        RECT 1201.680 596.630 1203.660 596.770 ;
        RECT 1201.680 545.090 1201.820 596.630 ;
        RECT 1201.220 544.950 1201.820 545.090 ;
        RECT 1201.220 497.070 1201.360 544.950 ;
        RECT 1201.160 496.750 1201.420 497.070 ;
        RECT 1200.700 496.410 1200.960 496.730 ;
        RECT 1200.760 483.325 1200.900 496.410 ;
        RECT 1200.690 482.955 1200.970 483.325 ;
        RECT 1201.610 482.955 1201.890 483.325 ;
        RECT 1201.680 448.530 1201.820 482.955 ;
        RECT 1201.220 448.390 1201.820 448.530 ;
        RECT 1201.220 427.710 1201.360 448.390 ;
        RECT 1201.160 427.390 1201.420 427.710 ;
        RECT 1202.540 427.390 1202.800 427.710 ;
        RECT 1202.600 379.770 1202.740 427.390 ;
        RECT 1201.620 379.450 1201.880 379.770 ;
        RECT 1202.540 379.450 1202.800 379.770 ;
        RECT 1201.680 379.285 1201.820 379.450 ;
        RECT 1201.610 378.915 1201.890 379.285 ;
        RECT 1202.530 378.235 1202.810 378.605 ;
        RECT 1202.600 331.830 1202.740 378.235 ;
        RECT 1201.160 331.510 1201.420 331.830 ;
        RECT 1202.540 331.510 1202.800 331.830 ;
        RECT 1201.220 331.150 1201.360 331.510 ;
        RECT 1201.160 330.830 1201.420 331.150 ;
        RECT 1201.620 330.830 1201.880 331.150 ;
        RECT 1201.680 324.350 1201.820 330.830 ;
        RECT 1201.620 324.030 1201.880 324.350 ;
        RECT 1202.540 324.030 1202.800 324.350 ;
        RECT 1202.600 276.410 1202.740 324.030 ;
        RECT 1201.620 276.090 1201.880 276.410 ;
        RECT 1202.540 276.090 1202.800 276.410 ;
        RECT 1201.680 255.670 1201.820 276.090 ;
        RECT 1201.620 255.350 1201.880 255.670 ;
        RECT 1202.080 254.670 1202.340 254.990 ;
        RECT 1202.140 227.790 1202.280 254.670 ;
        RECT 1201.160 227.470 1201.420 227.790 ;
        RECT 1202.080 227.470 1202.340 227.790 ;
        RECT 1201.220 179.850 1201.360 227.470 ;
        RECT 1201.160 179.530 1201.420 179.850 ;
        RECT 1201.620 179.530 1201.880 179.850 ;
        RECT 1201.680 159.110 1201.820 179.530 ;
        RECT 1201.620 158.790 1201.880 159.110 ;
        RECT 1201.160 158.450 1201.420 158.770 ;
        RECT 1201.220 110.570 1201.360 158.450 ;
        RECT 1200.760 110.490 1201.360 110.570 ;
        RECT 1200.700 110.430 1201.360 110.490 ;
        RECT 1200.700 110.170 1200.960 110.430 ;
        RECT 1201.620 110.170 1201.880 110.490 ;
        RECT 1201.680 60.250 1201.820 110.170 ;
        RECT 1201.680 60.110 1202.280 60.250 ;
        RECT 1202.140 58.890 1202.280 60.110 ;
        RECT 1201.680 58.750 1202.280 58.890 ;
        RECT 1201.680 24.810 1201.820 58.750 ;
        RECT 1043.380 24.490 1043.640 24.810 ;
        RECT 1201.620 24.490 1201.880 24.810 ;
        RECT 1043.440 2.400 1043.580 24.490 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
      LAYER via2 ;
        RECT 1200.690 483.000 1200.970 483.280 ;
        RECT 1201.610 483.000 1201.890 483.280 ;
        RECT 1201.610 378.960 1201.890 379.240 ;
        RECT 1202.530 378.280 1202.810 378.560 ;
      LAYER met3 ;
        RECT 1200.665 483.290 1200.995 483.305 ;
        RECT 1201.585 483.290 1201.915 483.305 ;
        RECT 1200.665 482.990 1201.915 483.290 ;
        RECT 1200.665 482.975 1200.995 482.990 ;
        RECT 1201.585 482.975 1201.915 482.990 ;
        RECT 1201.585 379.250 1201.915 379.265 ;
        RECT 1200.910 378.950 1201.915 379.250 ;
        RECT 1200.910 378.570 1201.210 378.950 ;
        RECT 1201.585 378.935 1201.915 378.950 ;
        RECT 1202.505 378.570 1202.835 378.585 ;
        RECT 1200.910 378.270 1202.835 378.570 ;
        RECT 1202.505 378.255 1202.835 378.270 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1061.290 24.380 1061.610 24.440 ;
        RECT 1214.930 24.380 1215.250 24.440 ;
        RECT 1061.290 24.240 1215.250 24.380 ;
        RECT 1061.290 24.180 1061.610 24.240 ;
        RECT 1214.930 24.180 1215.250 24.240 ;
      LAYER via ;
        RECT 1061.320 24.180 1061.580 24.440 ;
        RECT 1214.960 24.180 1215.220 24.440 ;
      LAYER met2 ;
        RECT 1215.190 600.000 1215.470 604.000 ;
        RECT 1215.250 598.810 1215.390 600.000 ;
        RECT 1215.020 598.670 1215.390 598.810 ;
        RECT 1215.020 24.470 1215.160 598.670 ;
        RECT 1061.320 24.150 1061.580 24.470 ;
        RECT 1214.960 24.150 1215.220 24.470 ;
        RECT 1061.380 2.400 1061.520 24.150 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1079.230 25.060 1079.550 25.120 ;
        RECT 1221.830 25.060 1222.150 25.120 ;
        RECT 1079.230 24.920 1222.150 25.060 ;
        RECT 1079.230 24.860 1079.550 24.920 ;
        RECT 1221.830 24.860 1222.150 24.920 ;
      LAYER via ;
        RECT 1079.260 24.860 1079.520 25.120 ;
        RECT 1221.860 24.860 1222.120 25.120 ;
      LAYER met2 ;
        RECT 1224.390 600.170 1224.670 604.000 ;
        RECT 1221.920 600.030 1224.670 600.170 ;
        RECT 1221.920 25.150 1222.060 600.030 ;
        RECT 1224.390 600.000 1224.670 600.030 ;
        RECT 1079.260 24.830 1079.520 25.150 ;
        RECT 1221.860 24.830 1222.120 25.150 ;
        RECT 1079.320 2.400 1079.460 24.830 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1228.730 569.400 1229.050 569.460 ;
        RECT 1231.950 569.400 1232.270 569.460 ;
        RECT 1228.730 569.260 1232.270 569.400 ;
        RECT 1228.730 569.200 1229.050 569.260 ;
        RECT 1231.950 569.200 1232.270 569.260 ;
        RECT 1096.710 25.400 1097.030 25.460 ;
        RECT 1228.730 25.400 1229.050 25.460 ;
        RECT 1096.710 25.260 1229.050 25.400 ;
        RECT 1096.710 25.200 1097.030 25.260 ;
        RECT 1228.730 25.200 1229.050 25.260 ;
      LAYER via ;
        RECT 1228.760 569.200 1229.020 569.460 ;
        RECT 1231.980 569.200 1232.240 569.460 ;
        RECT 1096.740 25.200 1097.000 25.460 ;
        RECT 1228.760 25.200 1229.020 25.460 ;
      LAYER met2 ;
        RECT 1233.590 600.170 1233.870 604.000 ;
        RECT 1232.040 600.030 1233.870 600.170 ;
        RECT 1232.040 569.490 1232.180 600.030 ;
        RECT 1233.590 600.000 1233.870 600.030 ;
        RECT 1228.760 569.170 1229.020 569.490 ;
        RECT 1231.980 569.170 1232.240 569.490 ;
        RECT 1228.820 25.490 1228.960 569.170 ;
        RECT 1096.740 25.170 1097.000 25.490 ;
        RECT 1228.760 25.170 1229.020 25.490 ;
        RECT 1096.800 2.400 1096.940 25.170 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1114.650 17.580 1114.970 17.640 ;
        RECT 1242.530 17.580 1242.850 17.640 ;
        RECT 1114.650 17.440 1242.850 17.580 ;
        RECT 1114.650 17.380 1114.970 17.440 ;
        RECT 1242.530 17.380 1242.850 17.440 ;
      LAYER via ;
        RECT 1114.680 17.380 1114.940 17.640 ;
        RECT 1242.560 17.380 1242.820 17.640 ;
      LAYER met2 ;
        RECT 1242.330 600.000 1242.610 604.000 ;
        RECT 1242.390 598.810 1242.530 600.000 ;
        RECT 1242.390 598.670 1242.760 598.810 ;
        RECT 1242.620 17.670 1242.760 598.670 ;
        RECT 1114.680 17.350 1114.940 17.670 ;
        RECT 1242.560 17.350 1242.820 17.670 ;
        RECT 1114.740 2.400 1114.880 17.350 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1249.430 569.400 1249.750 569.460 ;
        RECT 1250.350 569.400 1250.670 569.460 ;
        RECT 1249.430 569.260 1250.670 569.400 ;
        RECT 1249.430 569.200 1249.750 569.260 ;
        RECT 1250.350 569.200 1250.670 569.260 ;
        RECT 1132.590 18.260 1132.910 18.320 ;
        RECT 1249.430 18.260 1249.750 18.320 ;
        RECT 1132.590 18.120 1249.750 18.260 ;
        RECT 1132.590 18.060 1132.910 18.120 ;
        RECT 1249.430 18.060 1249.750 18.120 ;
      LAYER via ;
        RECT 1249.460 569.200 1249.720 569.460 ;
        RECT 1250.380 569.200 1250.640 569.460 ;
        RECT 1132.620 18.060 1132.880 18.320 ;
        RECT 1249.460 18.060 1249.720 18.320 ;
      LAYER met2 ;
        RECT 1251.530 600.170 1251.810 604.000 ;
        RECT 1250.440 600.030 1251.810 600.170 ;
        RECT 1250.440 569.490 1250.580 600.030 ;
        RECT 1251.530 600.000 1251.810 600.030 ;
        RECT 1249.460 569.170 1249.720 569.490 ;
        RECT 1250.380 569.170 1250.640 569.490 ;
        RECT 1249.520 18.350 1249.660 569.170 ;
        RECT 1132.620 18.030 1132.880 18.350 ;
        RECT 1249.460 18.030 1249.720 18.350 ;
        RECT 1132.680 2.400 1132.820 18.030 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1256.330 496.780 1256.650 497.040 ;
        RECT 1255.870 496.640 1256.190 496.700 ;
        RECT 1256.420 496.640 1256.560 496.780 ;
        RECT 1255.870 496.500 1256.560 496.640 ;
        RECT 1255.870 496.440 1256.190 496.500 ;
        RECT 1256.790 385.800 1257.110 385.860 ;
        RECT 1258.170 385.800 1258.490 385.860 ;
        RECT 1256.790 385.660 1258.490 385.800 ;
        RECT 1256.790 385.600 1257.110 385.660 ;
        RECT 1258.170 385.600 1258.490 385.660 ;
        RECT 1256.330 338.200 1256.650 338.260 ;
        RECT 1258.170 338.200 1258.490 338.260 ;
        RECT 1256.330 338.060 1258.490 338.200 ;
        RECT 1256.330 338.000 1256.650 338.060 ;
        RECT 1258.170 338.000 1258.490 338.060 ;
        RECT 1255.870 289.580 1256.190 289.640 ;
        RECT 1256.790 289.580 1257.110 289.640 ;
        RECT 1255.870 289.440 1257.110 289.580 ;
        RECT 1255.870 289.380 1256.190 289.440 ;
        RECT 1256.790 289.380 1257.110 289.440 ;
        RECT 1255.870 241.640 1256.190 241.700 ;
        RECT 1257.250 241.640 1257.570 241.700 ;
        RECT 1255.870 241.500 1257.570 241.640 ;
        RECT 1255.870 241.440 1256.190 241.500 ;
        RECT 1257.250 241.440 1257.570 241.500 ;
        RECT 1256.790 193.020 1257.110 193.080 ;
        RECT 1257.710 193.020 1258.030 193.080 ;
        RECT 1256.790 192.880 1258.030 193.020 ;
        RECT 1256.790 192.820 1257.110 192.880 ;
        RECT 1257.710 192.820 1258.030 192.880 ;
        RECT 1256.330 145.080 1256.650 145.140 ;
        RECT 1257.710 145.080 1258.030 145.140 ;
        RECT 1256.330 144.940 1258.030 145.080 ;
        RECT 1256.330 144.880 1256.650 144.940 ;
        RECT 1257.710 144.880 1258.030 144.940 ;
        RECT 1255.870 110.400 1256.190 110.460 ;
        RECT 1256.790 110.400 1257.110 110.460 ;
        RECT 1255.870 110.260 1257.110 110.400 ;
        RECT 1255.870 110.200 1256.190 110.260 ;
        RECT 1256.790 110.200 1257.110 110.260 ;
        RECT 1255.870 96.460 1256.190 96.520 ;
        RECT 1256.790 96.460 1257.110 96.520 ;
        RECT 1255.870 96.320 1257.110 96.460 ;
        RECT 1255.870 96.260 1256.190 96.320 ;
        RECT 1256.790 96.260 1257.110 96.320 ;
        RECT 1150.530 19.620 1150.850 19.680 ;
        RECT 1159.270 19.620 1159.590 19.680 ;
        RECT 1256.790 19.620 1257.110 19.680 ;
        RECT 1150.530 19.480 1159.590 19.620 ;
        RECT 1150.530 19.420 1150.850 19.480 ;
        RECT 1159.270 19.420 1159.590 19.480 ;
        RECT 1255.500 19.480 1257.110 19.620 ;
        RECT 1207.570 19.280 1207.890 19.340 ;
        RECT 1187.420 19.140 1207.890 19.280 ;
        RECT 1159.270 18.600 1159.590 18.660 ;
        RECT 1187.420 18.600 1187.560 19.140 ;
        RECT 1207.570 19.080 1207.890 19.140 ;
        RECT 1226.430 19.280 1226.750 19.340 ;
        RECT 1255.500 19.280 1255.640 19.480 ;
        RECT 1256.790 19.420 1257.110 19.480 ;
        RECT 1226.430 19.140 1255.640 19.280 ;
        RECT 1226.430 19.080 1226.750 19.140 ;
        RECT 1159.270 18.460 1187.560 18.600 ;
        RECT 1159.270 18.400 1159.590 18.460 ;
      LAYER via ;
        RECT 1256.360 496.780 1256.620 497.040 ;
        RECT 1255.900 496.440 1256.160 496.700 ;
        RECT 1256.820 385.600 1257.080 385.860 ;
        RECT 1258.200 385.600 1258.460 385.860 ;
        RECT 1256.360 338.000 1256.620 338.260 ;
        RECT 1258.200 338.000 1258.460 338.260 ;
        RECT 1255.900 289.380 1256.160 289.640 ;
        RECT 1256.820 289.380 1257.080 289.640 ;
        RECT 1255.900 241.440 1256.160 241.700 ;
        RECT 1257.280 241.440 1257.540 241.700 ;
        RECT 1256.820 192.820 1257.080 193.080 ;
        RECT 1257.740 192.820 1258.000 193.080 ;
        RECT 1256.360 144.880 1256.620 145.140 ;
        RECT 1257.740 144.880 1258.000 145.140 ;
        RECT 1255.900 110.200 1256.160 110.460 ;
        RECT 1256.820 110.200 1257.080 110.460 ;
        RECT 1255.900 96.260 1256.160 96.520 ;
        RECT 1256.820 96.260 1257.080 96.520 ;
        RECT 1150.560 19.420 1150.820 19.680 ;
        RECT 1159.300 19.420 1159.560 19.680 ;
        RECT 1159.300 18.400 1159.560 18.660 ;
        RECT 1207.600 19.080 1207.860 19.340 ;
        RECT 1226.460 19.080 1226.720 19.340 ;
        RECT 1256.820 19.420 1257.080 19.680 ;
      LAYER met2 ;
        RECT 1260.730 600.850 1261.010 604.000 ;
        RECT 1258.720 600.710 1261.010 600.850 ;
        RECT 1258.720 596.770 1258.860 600.710 ;
        RECT 1260.730 600.000 1261.010 600.710 ;
        RECT 1256.880 596.630 1258.860 596.770 ;
        RECT 1256.880 545.090 1257.020 596.630 ;
        RECT 1256.420 544.950 1257.020 545.090 ;
        RECT 1256.420 497.070 1256.560 544.950 ;
        RECT 1256.360 496.750 1256.620 497.070 ;
        RECT 1255.900 496.410 1256.160 496.730 ;
        RECT 1255.960 483.325 1256.100 496.410 ;
        RECT 1255.890 482.955 1256.170 483.325 ;
        RECT 1256.810 482.955 1257.090 483.325 ;
        RECT 1256.880 448.530 1257.020 482.955 ;
        RECT 1256.420 448.390 1257.020 448.530 ;
        RECT 1256.420 410.450 1256.560 448.390 ;
        RECT 1256.420 410.310 1257.020 410.450 ;
        RECT 1256.880 385.890 1257.020 410.310 ;
        RECT 1256.820 385.570 1257.080 385.890 ;
        RECT 1258.200 385.570 1258.460 385.890 ;
        RECT 1258.260 338.290 1258.400 385.570 ;
        RECT 1256.360 337.970 1256.620 338.290 ;
        RECT 1258.200 337.970 1258.460 338.290 ;
        RECT 1256.420 337.805 1256.560 337.970 ;
        RECT 1256.350 337.435 1256.630 337.805 ;
        RECT 1256.810 303.435 1257.090 303.805 ;
        RECT 1256.880 289.670 1257.020 303.435 ;
        RECT 1255.900 289.350 1256.160 289.670 ;
        RECT 1256.820 289.350 1257.080 289.670 ;
        RECT 1255.960 241.730 1256.100 289.350 ;
        RECT 1255.900 241.410 1256.160 241.730 ;
        RECT 1257.280 241.410 1257.540 241.730 ;
        RECT 1257.340 207.925 1257.480 241.410 ;
        RECT 1257.270 207.555 1257.550 207.925 ;
        RECT 1256.810 193.275 1257.090 193.645 ;
        RECT 1256.880 193.110 1257.020 193.275 ;
        RECT 1256.820 192.790 1257.080 193.110 ;
        RECT 1257.740 192.790 1258.000 193.110 ;
        RECT 1257.800 145.170 1257.940 192.790 ;
        RECT 1256.360 144.850 1256.620 145.170 ;
        RECT 1257.740 144.850 1258.000 145.170 ;
        RECT 1256.420 110.570 1256.560 144.850 ;
        RECT 1255.960 110.490 1256.560 110.570 ;
        RECT 1255.900 110.430 1256.560 110.490 ;
        RECT 1255.900 110.170 1256.160 110.430 ;
        RECT 1256.820 110.170 1257.080 110.490 ;
        RECT 1256.880 96.550 1257.020 110.170 ;
        RECT 1255.900 96.230 1256.160 96.550 ;
        RECT 1256.820 96.230 1257.080 96.550 ;
        RECT 1255.960 60.930 1256.100 96.230 ;
        RECT 1255.960 60.790 1257.020 60.930 ;
        RECT 1256.880 19.710 1257.020 60.790 ;
        RECT 1150.560 19.390 1150.820 19.710 ;
        RECT 1159.300 19.390 1159.560 19.710 ;
        RECT 1150.620 2.400 1150.760 19.390 ;
        RECT 1159.360 18.690 1159.500 19.390 ;
        RECT 1207.590 19.195 1207.870 19.565 ;
        RECT 1226.450 19.195 1226.730 19.565 ;
        RECT 1256.820 19.390 1257.080 19.710 ;
        RECT 1207.600 19.050 1207.860 19.195 ;
        RECT 1226.460 19.050 1226.720 19.195 ;
        RECT 1159.300 18.370 1159.560 18.690 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
      LAYER via2 ;
        RECT 1255.890 483.000 1256.170 483.280 ;
        RECT 1256.810 483.000 1257.090 483.280 ;
        RECT 1256.350 337.480 1256.630 337.760 ;
        RECT 1256.810 303.480 1257.090 303.760 ;
        RECT 1257.270 207.600 1257.550 207.880 ;
        RECT 1256.810 193.320 1257.090 193.600 ;
        RECT 1207.590 19.240 1207.870 19.520 ;
        RECT 1226.450 19.240 1226.730 19.520 ;
      LAYER met3 ;
        RECT 1255.865 483.290 1256.195 483.305 ;
        RECT 1256.785 483.290 1257.115 483.305 ;
        RECT 1255.865 482.990 1257.115 483.290 ;
        RECT 1255.865 482.975 1256.195 482.990 ;
        RECT 1256.785 482.975 1257.115 482.990 ;
        RECT 1256.325 337.780 1256.655 337.785 ;
        RECT 1256.070 337.770 1256.655 337.780 ;
        RECT 1256.070 337.470 1256.880 337.770 ;
        RECT 1256.070 337.460 1256.655 337.470 ;
        RECT 1256.325 337.455 1256.655 337.460 ;
        RECT 1256.070 303.770 1256.450 303.780 ;
        RECT 1256.785 303.770 1257.115 303.785 ;
        RECT 1256.070 303.470 1257.115 303.770 ;
        RECT 1256.070 303.460 1256.450 303.470 ;
        RECT 1256.785 303.455 1257.115 303.470 ;
        RECT 1257.245 207.900 1257.575 207.905 ;
        RECT 1256.990 207.890 1257.575 207.900 ;
        RECT 1256.790 207.590 1257.575 207.890 ;
        RECT 1256.990 207.580 1257.575 207.590 ;
        RECT 1257.245 207.575 1257.575 207.580 ;
        RECT 1256.785 193.620 1257.115 193.625 ;
        RECT 1256.785 193.610 1257.370 193.620 ;
        RECT 1256.785 193.310 1257.570 193.610 ;
        RECT 1256.785 193.300 1257.370 193.310 ;
        RECT 1256.785 193.295 1257.115 193.300 ;
        RECT 1207.565 19.530 1207.895 19.545 ;
        RECT 1226.425 19.530 1226.755 19.545 ;
        RECT 1207.565 19.230 1226.755 19.530 ;
        RECT 1207.565 19.215 1207.895 19.230 ;
        RECT 1226.425 19.215 1226.755 19.230 ;
      LAYER via3 ;
        RECT 1256.100 337.460 1256.420 337.780 ;
        RECT 1256.100 303.460 1256.420 303.780 ;
        RECT 1257.020 207.580 1257.340 207.900 ;
        RECT 1257.020 193.300 1257.340 193.620 ;
      LAYER met4 ;
        RECT 1256.095 337.455 1256.425 337.785 ;
        RECT 1256.110 303.785 1256.410 337.455 ;
        RECT 1256.095 303.455 1256.425 303.785 ;
        RECT 1257.015 207.575 1257.345 207.905 ;
        RECT 1257.030 193.625 1257.330 207.575 ;
        RECT 1257.015 193.295 1257.345 193.625 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.470 569.400 1007.790 569.460 ;
        RECT 1011.610 569.400 1011.930 569.460 ;
        RECT 1007.470 569.260 1011.930 569.400 ;
        RECT 1007.470 569.200 1007.790 569.260 ;
        RECT 1011.610 569.200 1011.930 569.260 ;
        RECT 668.910 35.940 669.230 36.000 ;
        RECT 1007.470 35.940 1007.790 36.000 ;
        RECT 668.910 35.800 1007.790 35.940 ;
        RECT 668.910 35.740 669.230 35.800 ;
        RECT 1007.470 35.740 1007.790 35.800 ;
      LAYER via ;
        RECT 1007.500 569.200 1007.760 569.460 ;
        RECT 1011.640 569.200 1011.900 569.460 ;
        RECT 668.940 35.740 669.200 36.000 ;
        RECT 1007.500 35.740 1007.760 36.000 ;
      LAYER met2 ;
        RECT 1013.250 600.170 1013.530 604.000 ;
        RECT 1011.700 600.030 1013.530 600.170 ;
        RECT 1011.700 569.490 1011.840 600.030 ;
        RECT 1013.250 600.000 1013.530 600.030 ;
        RECT 1007.500 569.170 1007.760 569.490 ;
        RECT 1011.640 569.170 1011.900 569.490 ;
        RECT 1007.560 36.030 1007.700 569.170 ;
        RECT 668.940 35.710 669.200 36.030 ;
        RECT 1007.500 35.710 1007.760 36.030 ;
        RECT 669.000 2.400 669.140 35.710 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1172.610 591.500 1172.930 591.560 ;
        RECT 1172.610 591.360 1197.220 591.500 ;
        RECT 1172.610 591.300 1172.930 591.360 ;
        RECT 1197.080 591.160 1197.220 591.360 ;
        RECT 1269.670 591.160 1269.990 591.220 ;
        RECT 1197.080 591.020 1269.990 591.160 ;
        RECT 1269.670 590.960 1269.990 591.020 ;
        RECT 1168.470 19.960 1168.790 20.020 ;
        RECT 1172.610 19.960 1172.930 20.020 ;
        RECT 1168.470 19.820 1172.930 19.960 ;
        RECT 1168.470 19.760 1168.790 19.820 ;
        RECT 1172.610 19.760 1172.930 19.820 ;
      LAYER via ;
        RECT 1172.640 591.300 1172.900 591.560 ;
        RECT 1269.700 590.960 1269.960 591.220 ;
        RECT 1168.500 19.760 1168.760 20.020 ;
        RECT 1172.640 19.760 1172.900 20.020 ;
      LAYER met2 ;
        RECT 1269.930 600.000 1270.210 604.000 ;
        RECT 1269.990 598.810 1270.130 600.000 ;
        RECT 1269.760 598.670 1270.130 598.810 ;
        RECT 1172.640 591.270 1172.900 591.590 ;
        RECT 1172.700 20.050 1172.840 591.270 ;
        RECT 1269.760 591.250 1269.900 598.670 ;
        RECT 1269.700 590.930 1269.960 591.250 ;
        RECT 1168.500 19.730 1168.760 20.050 ;
        RECT 1172.640 19.730 1172.900 20.050 ;
        RECT 1168.560 2.400 1168.700 19.730 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1277.490 592.520 1277.810 592.580 ;
        RECT 1201.680 592.380 1277.810 592.520 ;
        RECT 1186.410 592.180 1186.730 592.240 ;
        RECT 1201.680 592.180 1201.820 592.380 ;
        RECT 1277.490 592.320 1277.810 592.380 ;
        RECT 1186.410 592.040 1201.820 592.180 ;
        RECT 1186.410 591.980 1186.730 592.040 ;
        RECT 1186.410 572.460 1186.730 572.520 ;
        RECT 1187.790 572.460 1188.110 572.520 ;
        RECT 1186.410 572.320 1188.110 572.460 ;
        RECT 1186.410 572.260 1186.730 572.320 ;
        RECT 1187.790 572.260 1188.110 572.320 ;
        RECT 1186.410 524.520 1186.730 524.580 ;
        RECT 1187.790 524.520 1188.110 524.580 ;
        RECT 1186.410 524.380 1188.110 524.520 ;
        RECT 1186.410 524.320 1186.730 524.380 ;
        RECT 1187.790 524.320 1188.110 524.380 ;
        RECT 1185.030 475.900 1185.350 475.960 ;
        RECT 1186.410 475.900 1186.730 475.960 ;
        RECT 1185.030 475.760 1186.730 475.900 ;
        RECT 1185.030 475.700 1185.350 475.760 ;
        RECT 1186.410 475.700 1186.730 475.760 ;
        RECT 1185.030 427.960 1185.350 428.020 ;
        RECT 1186.410 427.960 1186.730 428.020 ;
        RECT 1185.030 427.820 1186.730 427.960 ;
        RECT 1185.030 427.760 1185.350 427.820 ;
        RECT 1186.410 427.760 1186.730 427.820 ;
        RECT 1186.410 426.260 1186.730 426.320 ;
        RECT 1187.790 426.260 1188.110 426.320 ;
        RECT 1186.410 426.120 1188.110 426.260 ;
        RECT 1186.410 426.060 1186.730 426.120 ;
        RECT 1187.790 426.060 1188.110 426.120 ;
        RECT 1186.410 338.200 1186.730 338.260 ;
        RECT 1187.790 338.200 1188.110 338.260 ;
        RECT 1186.410 338.060 1188.110 338.200 ;
        RECT 1186.410 338.000 1186.730 338.060 ;
        RECT 1187.790 338.000 1188.110 338.060 ;
        RECT 1186.410 234.500 1186.730 234.560 ;
        RECT 1187.790 234.500 1188.110 234.560 ;
        RECT 1186.410 234.360 1188.110 234.500 ;
        RECT 1186.410 234.300 1186.730 234.360 ;
        RECT 1187.790 234.300 1188.110 234.360 ;
        RECT 1186.410 186.560 1186.730 186.620 ;
        RECT 1187.790 186.560 1188.110 186.620 ;
        RECT 1186.410 186.420 1188.110 186.560 ;
        RECT 1186.410 186.360 1186.730 186.420 ;
        RECT 1187.790 186.360 1188.110 186.420 ;
        RECT 1186.410 137.940 1186.730 138.000 ;
        RECT 1187.790 137.940 1188.110 138.000 ;
        RECT 1186.410 137.800 1188.110 137.940 ;
        RECT 1186.410 137.740 1186.730 137.800 ;
        RECT 1187.790 137.740 1188.110 137.800 ;
        RECT 1186.410 90.000 1186.730 90.060 ;
        RECT 1187.790 90.000 1188.110 90.060 ;
        RECT 1186.410 89.860 1188.110 90.000 ;
        RECT 1186.410 89.800 1186.730 89.860 ;
        RECT 1187.790 89.800 1188.110 89.860 ;
        RECT 1186.410 62.800 1186.730 62.860 ;
        RECT 1185.580 62.660 1186.730 62.800 ;
        RECT 1185.580 62.180 1185.720 62.660 ;
        RECT 1186.410 62.600 1186.730 62.660 ;
        RECT 1185.490 61.920 1185.810 62.180 ;
        RECT 1185.490 23.700 1185.810 23.760 ;
        RECT 1186.410 23.700 1186.730 23.760 ;
        RECT 1185.490 23.560 1186.730 23.700 ;
        RECT 1185.490 23.500 1185.810 23.560 ;
        RECT 1186.410 23.500 1186.730 23.560 ;
      LAYER via ;
        RECT 1186.440 591.980 1186.700 592.240 ;
        RECT 1277.520 592.320 1277.780 592.580 ;
        RECT 1186.440 572.260 1186.700 572.520 ;
        RECT 1187.820 572.260 1188.080 572.520 ;
        RECT 1186.440 524.320 1186.700 524.580 ;
        RECT 1187.820 524.320 1188.080 524.580 ;
        RECT 1185.060 475.700 1185.320 475.960 ;
        RECT 1186.440 475.700 1186.700 475.960 ;
        RECT 1185.060 427.760 1185.320 428.020 ;
        RECT 1186.440 427.760 1186.700 428.020 ;
        RECT 1186.440 426.060 1186.700 426.320 ;
        RECT 1187.820 426.060 1188.080 426.320 ;
        RECT 1186.440 338.000 1186.700 338.260 ;
        RECT 1187.820 338.000 1188.080 338.260 ;
        RECT 1186.440 234.300 1186.700 234.560 ;
        RECT 1187.820 234.300 1188.080 234.560 ;
        RECT 1186.440 186.360 1186.700 186.620 ;
        RECT 1187.820 186.360 1188.080 186.620 ;
        RECT 1186.440 137.740 1186.700 138.000 ;
        RECT 1187.820 137.740 1188.080 138.000 ;
        RECT 1186.440 89.800 1186.700 90.060 ;
        RECT 1187.820 89.800 1188.080 90.060 ;
        RECT 1186.440 62.600 1186.700 62.860 ;
        RECT 1185.520 61.920 1185.780 62.180 ;
        RECT 1185.520 23.500 1185.780 23.760 ;
        RECT 1186.440 23.500 1186.700 23.760 ;
      LAYER met2 ;
        RECT 1279.130 600.170 1279.410 604.000 ;
        RECT 1277.580 600.030 1279.410 600.170 ;
        RECT 1277.580 592.610 1277.720 600.030 ;
        RECT 1279.130 600.000 1279.410 600.030 ;
        RECT 1277.520 592.290 1277.780 592.610 ;
        RECT 1186.440 591.950 1186.700 592.270 ;
        RECT 1186.500 572.550 1186.640 591.950 ;
        RECT 1186.440 572.230 1186.700 572.550 ;
        RECT 1187.820 572.230 1188.080 572.550 ;
        RECT 1187.880 524.610 1188.020 572.230 ;
        RECT 1186.440 524.290 1186.700 524.610 ;
        RECT 1187.820 524.290 1188.080 524.610 ;
        RECT 1186.500 475.990 1186.640 524.290 ;
        RECT 1185.060 475.670 1185.320 475.990 ;
        RECT 1186.440 475.670 1186.700 475.990 ;
        RECT 1185.120 428.050 1185.260 475.670 ;
        RECT 1185.060 427.730 1185.320 428.050 ;
        RECT 1186.440 427.730 1186.700 428.050 ;
        RECT 1186.500 426.350 1186.640 427.730 ;
        RECT 1186.440 426.030 1186.700 426.350 ;
        RECT 1187.820 426.030 1188.080 426.350 ;
        RECT 1187.880 338.290 1188.020 426.030 ;
        RECT 1186.440 337.970 1186.700 338.290 ;
        RECT 1187.820 337.970 1188.080 338.290 ;
        RECT 1186.500 234.590 1186.640 337.970 ;
        RECT 1186.440 234.270 1186.700 234.590 ;
        RECT 1187.820 234.270 1188.080 234.590 ;
        RECT 1187.880 186.650 1188.020 234.270 ;
        RECT 1186.440 186.330 1186.700 186.650 ;
        RECT 1187.820 186.330 1188.080 186.650 ;
        RECT 1186.500 138.030 1186.640 186.330 ;
        RECT 1186.440 137.710 1186.700 138.030 ;
        RECT 1187.820 137.710 1188.080 138.030 ;
        RECT 1187.880 90.090 1188.020 137.710 ;
        RECT 1186.440 89.770 1186.700 90.090 ;
        RECT 1187.820 89.770 1188.080 90.090 ;
        RECT 1186.500 62.890 1186.640 89.770 ;
        RECT 1186.440 62.570 1186.700 62.890 ;
        RECT 1185.520 61.890 1185.780 62.210 ;
        RECT 1185.580 23.790 1185.720 61.890 ;
        RECT 1185.520 23.470 1185.780 23.790 ;
        RECT 1186.440 23.470 1186.700 23.790 ;
        RECT 1186.500 22.850 1186.640 23.470 ;
        RECT 1186.040 22.710 1186.640 22.850 ;
        RECT 1186.040 2.400 1186.180 22.710 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.110 589.460 1207.430 589.520 ;
        RECT 1286.690 589.460 1287.010 589.520 ;
        RECT 1207.110 589.320 1287.010 589.460 ;
        RECT 1207.110 589.260 1207.430 589.320 ;
        RECT 1286.690 589.260 1287.010 589.320 ;
        RECT 1203.890 20.640 1204.210 20.700 ;
        RECT 1207.110 20.640 1207.430 20.700 ;
        RECT 1203.890 20.500 1207.430 20.640 ;
        RECT 1203.890 20.440 1204.210 20.500 ;
        RECT 1207.110 20.440 1207.430 20.500 ;
      LAYER via ;
        RECT 1207.140 589.260 1207.400 589.520 ;
        RECT 1286.720 589.260 1286.980 589.520 ;
        RECT 1203.920 20.440 1204.180 20.700 ;
        RECT 1207.140 20.440 1207.400 20.700 ;
      LAYER met2 ;
        RECT 1288.330 600.170 1288.610 604.000 ;
        RECT 1286.780 600.030 1288.610 600.170 ;
        RECT 1286.780 589.550 1286.920 600.030 ;
        RECT 1288.330 600.000 1288.610 600.030 ;
        RECT 1207.140 589.230 1207.400 589.550 ;
        RECT 1286.720 589.230 1286.980 589.550 ;
        RECT 1207.200 20.730 1207.340 589.230 ;
        RECT 1203.920 20.410 1204.180 20.730 ;
        RECT 1207.140 20.410 1207.400 20.730 ;
        RECT 1203.980 2.400 1204.120 20.410 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1227.350 589.120 1227.670 589.180 ;
        RECT 1297.730 589.120 1298.050 589.180 ;
        RECT 1227.350 588.980 1298.050 589.120 ;
        RECT 1227.350 588.920 1227.670 588.980 ;
        RECT 1297.730 588.920 1298.050 588.980 ;
        RECT 1221.830 16.560 1222.150 16.620 ;
        RECT 1227.350 16.560 1227.670 16.620 ;
        RECT 1221.830 16.420 1227.670 16.560 ;
        RECT 1221.830 16.360 1222.150 16.420 ;
        RECT 1227.350 16.360 1227.670 16.420 ;
      LAYER via ;
        RECT 1227.380 588.920 1227.640 589.180 ;
        RECT 1297.760 588.920 1298.020 589.180 ;
        RECT 1221.860 16.360 1222.120 16.620 ;
        RECT 1227.380 16.360 1227.640 16.620 ;
      LAYER met2 ;
        RECT 1297.530 600.000 1297.810 604.000 ;
        RECT 1297.590 598.810 1297.730 600.000 ;
        RECT 1297.590 598.670 1297.960 598.810 ;
        RECT 1297.820 589.210 1297.960 598.670 ;
        RECT 1227.380 588.890 1227.640 589.210 ;
        RECT 1297.760 588.890 1298.020 589.210 ;
        RECT 1227.440 16.650 1227.580 588.890 ;
        RECT 1221.860 16.330 1222.120 16.650 ;
        RECT 1227.380 16.330 1227.640 16.650 ;
        RECT 1221.920 2.400 1222.060 16.330 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.610 588.780 1241.930 588.840 ;
        RECT 1305.090 588.780 1305.410 588.840 ;
        RECT 1241.610 588.640 1305.410 588.780 ;
        RECT 1241.610 588.580 1241.930 588.640 ;
        RECT 1305.090 588.580 1305.410 588.640 ;
        RECT 1239.770 2.960 1240.090 3.020 ;
        RECT 1241.610 2.960 1241.930 3.020 ;
        RECT 1239.770 2.820 1241.930 2.960 ;
        RECT 1239.770 2.760 1240.090 2.820 ;
        RECT 1241.610 2.760 1241.930 2.820 ;
      LAYER via ;
        RECT 1241.640 588.580 1241.900 588.840 ;
        RECT 1305.120 588.580 1305.380 588.840 ;
        RECT 1239.800 2.760 1240.060 3.020 ;
        RECT 1241.640 2.760 1241.900 3.020 ;
      LAYER met2 ;
        RECT 1306.730 600.170 1307.010 604.000 ;
        RECT 1305.180 600.030 1307.010 600.170 ;
        RECT 1305.180 588.870 1305.320 600.030 ;
        RECT 1306.730 600.000 1307.010 600.030 ;
        RECT 1241.640 588.550 1241.900 588.870 ;
        RECT 1305.120 588.550 1305.380 588.870 ;
        RECT 1241.700 3.050 1241.840 588.550 ;
        RECT 1239.800 2.730 1240.060 3.050 ;
        RECT 1241.640 2.730 1241.900 3.050 ;
        RECT 1239.860 2.400 1240.000 2.730 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 587.760 1262.630 587.820 ;
        RECT 1314.290 587.760 1314.610 587.820 ;
        RECT 1262.310 587.620 1314.610 587.760 ;
        RECT 1262.310 587.560 1262.630 587.620 ;
        RECT 1314.290 587.560 1314.610 587.620 ;
        RECT 1257.250 20.640 1257.570 20.700 ;
        RECT 1262.310 20.640 1262.630 20.700 ;
        RECT 1257.250 20.500 1262.630 20.640 ;
        RECT 1257.250 20.440 1257.570 20.500 ;
        RECT 1262.310 20.440 1262.630 20.500 ;
      LAYER via ;
        RECT 1262.340 587.560 1262.600 587.820 ;
        RECT 1314.320 587.560 1314.580 587.820 ;
        RECT 1257.280 20.440 1257.540 20.700 ;
        RECT 1262.340 20.440 1262.600 20.700 ;
      LAYER met2 ;
        RECT 1315.930 600.170 1316.210 604.000 ;
        RECT 1314.380 600.030 1316.210 600.170 ;
        RECT 1314.380 587.850 1314.520 600.030 ;
        RECT 1315.930 600.000 1316.210 600.030 ;
        RECT 1262.340 587.530 1262.600 587.850 ;
        RECT 1314.320 587.530 1314.580 587.850 ;
        RECT 1262.400 20.730 1262.540 587.530 ;
        RECT 1257.280 20.410 1257.540 20.730 ;
        RECT 1262.340 20.410 1262.600 20.730 ;
        RECT 1257.340 2.400 1257.480 20.410 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.110 590.820 1276.430 590.880 ;
        RECT 1324.870 590.820 1325.190 590.880 ;
        RECT 1276.110 590.680 1325.190 590.820 ;
        RECT 1276.110 590.620 1276.430 590.680 ;
        RECT 1324.870 590.620 1325.190 590.680 ;
      LAYER via ;
        RECT 1276.140 590.620 1276.400 590.880 ;
        RECT 1324.900 590.620 1325.160 590.880 ;
      LAYER met2 ;
        RECT 1325.130 600.000 1325.410 604.000 ;
        RECT 1325.190 598.810 1325.330 600.000 ;
        RECT 1324.960 598.670 1325.330 598.810 ;
        RECT 1324.960 590.910 1325.100 598.670 ;
        RECT 1276.140 590.590 1276.400 590.910 ;
        RECT 1324.900 590.590 1325.160 590.910 ;
        RECT 1276.200 16.730 1276.340 590.590 ;
        RECT 1275.280 16.590 1276.340 16.730 ;
        RECT 1275.280 2.400 1275.420 16.590 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 587.420 1297.130 587.480 ;
        RECT 1332.690 587.420 1333.010 587.480 ;
        RECT 1296.810 587.280 1333.010 587.420 ;
        RECT 1296.810 587.220 1297.130 587.280 ;
        RECT 1332.690 587.220 1333.010 587.280 ;
        RECT 1293.130 15.540 1293.450 15.600 ;
        RECT 1296.810 15.540 1297.130 15.600 ;
        RECT 1293.130 15.400 1297.130 15.540 ;
        RECT 1293.130 15.340 1293.450 15.400 ;
        RECT 1296.810 15.340 1297.130 15.400 ;
      LAYER via ;
        RECT 1296.840 587.220 1297.100 587.480 ;
        RECT 1332.720 587.220 1332.980 587.480 ;
        RECT 1293.160 15.340 1293.420 15.600 ;
        RECT 1296.840 15.340 1297.100 15.600 ;
      LAYER met2 ;
        RECT 1334.330 600.170 1334.610 604.000 ;
        RECT 1332.780 600.030 1334.610 600.170 ;
        RECT 1332.780 587.510 1332.920 600.030 ;
        RECT 1334.330 600.000 1334.610 600.030 ;
        RECT 1296.840 587.190 1297.100 587.510 ;
        RECT 1332.720 587.190 1332.980 587.510 ;
        RECT 1296.900 15.630 1297.040 587.190 ;
        RECT 1293.160 15.310 1293.420 15.630 ;
        RECT 1296.840 15.310 1297.100 15.630 ;
        RECT 1293.220 2.400 1293.360 15.310 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1317.510 589.460 1317.830 589.520 ;
        RECT 1341.890 589.460 1342.210 589.520 ;
        RECT 1317.510 589.320 1342.210 589.460 ;
        RECT 1317.510 589.260 1317.830 589.320 ;
        RECT 1341.890 589.260 1342.210 589.320 ;
        RECT 1311.070 17.580 1311.390 17.640 ;
        RECT 1317.510 17.580 1317.830 17.640 ;
        RECT 1311.070 17.440 1317.830 17.580 ;
        RECT 1311.070 17.380 1311.390 17.440 ;
        RECT 1317.510 17.380 1317.830 17.440 ;
      LAYER via ;
        RECT 1317.540 589.260 1317.800 589.520 ;
        RECT 1341.920 589.260 1342.180 589.520 ;
        RECT 1311.100 17.380 1311.360 17.640 ;
        RECT 1317.540 17.380 1317.800 17.640 ;
      LAYER met2 ;
        RECT 1343.530 600.170 1343.810 604.000 ;
        RECT 1341.980 600.030 1343.810 600.170 ;
        RECT 1341.980 589.550 1342.120 600.030 ;
        RECT 1343.530 600.000 1343.810 600.030 ;
        RECT 1317.540 589.230 1317.800 589.550 ;
        RECT 1341.920 589.230 1342.180 589.550 ;
        RECT 1317.600 17.670 1317.740 589.230 ;
        RECT 1311.100 17.350 1311.360 17.670 ;
        RECT 1317.540 17.350 1317.800 17.670 ;
        RECT 1311.160 2.400 1311.300 17.350 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.310 589.800 1331.630 589.860 ;
        RECT 1352.470 589.800 1352.790 589.860 ;
        RECT 1331.310 589.660 1352.790 589.800 ;
        RECT 1331.310 589.600 1331.630 589.660 ;
        RECT 1352.470 589.600 1352.790 589.660 ;
        RECT 1329.010 17.580 1329.330 17.640 ;
        RECT 1331.310 17.580 1331.630 17.640 ;
        RECT 1329.010 17.440 1331.630 17.580 ;
        RECT 1329.010 17.380 1329.330 17.440 ;
        RECT 1331.310 17.380 1331.630 17.440 ;
      LAYER via ;
        RECT 1331.340 589.600 1331.600 589.860 ;
        RECT 1352.500 589.600 1352.760 589.860 ;
        RECT 1329.040 17.380 1329.300 17.640 ;
        RECT 1331.340 17.380 1331.600 17.640 ;
      LAYER met2 ;
        RECT 1352.730 600.000 1353.010 604.000 ;
        RECT 1352.790 598.810 1352.930 600.000 ;
        RECT 1352.560 598.670 1352.930 598.810 ;
        RECT 1352.560 589.890 1352.700 598.670 ;
        RECT 1331.340 589.570 1331.600 589.890 ;
        RECT 1352.500 589.570 1352.760 589.890 ;
        RECT 1331.400 17.670 1331.540 589.570 ;
        RECT 1329.040 17.350 1329.300 17.670 ;
        RECT 1331.340 17.350 1331.600 17.670 ;
        RECT 1329.100 2.400 1329.240 17.350 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 37.980 686.710 38.040 ;
        RECT 1021.730 37.980 1022.050 38.040 ;
        RECT 686.390 37.840 1022.050 37.980 ;
        RECT 686.390 37.780 686.710 37.840 ;
        RECT 1021.730 37.780 1022.050 37.840 ;
      LAYER via ;
        RECT 686.420 37.780 686.680 38.040 ;
        RECT 1021.760 37.780 1022.020 38.040 ;
      LAYER met2 ;
        RECT 1022.450 600.170 1022.730 604.000 ;
        RECT 1021.820 600.030 1022.730 600.170 ;
        RECT 1021.820 38.070 1021.960 600.030 ;
        RECT 1022.450 600.000 1022.730 600.030 ;
        RECT 686.420 37.750 686.680 38.070 ;
        RECT 1021.760 37.750 1022.020 38.070 ;
        RECT 686.480 2.400 686.620 37.750 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.490 17.240 1346.810 17.300 ;
        RECT 1360.290 17.240 1360.610 17.300 ;
        RECT 1346.490 17.100 1360.610 17.240 ;
        RECT 1346.490 17.040 1346.810 17.100 ;
        RECT 1360.290 17.040 1360.610 17.100 ;
      LAYER via ;
        RECT 1346.520 17.040 1346.780 17.300 ;
        RECT 1360.320 17.040 1360.580 17.300 ;
      LAYER met2 ;
        RECT 1361.470 600.170 1361.750 604.000 ;
        RECT 1360.380 600.030 1361.750 600.170 ;
        RECT 1360.380 17.330 1360.520 600.030 ;
        RECT 1361.470 600.000 1361.750 600.030 ;
        RECT 1346.520 17.010 1346.780 17.330 ;
        RECT 1360.320 17.010 1360.580 17.330 ;
        RECT 1346.580 2.400 1346.720 17.010 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1367.650 497.320 1367.970 497.380 ;
        RECT 1367.280 497.180 1367.970 497.320 ;
        RECT 1367.280 496.700 1367.420 497.180 ;
        RECT 1367.650 497.120 1367.970 497.180 ;
        RECT 1367.190 496.440 1367.510 496.700 ;
        RECT 1365.810 427.620 1366.130 427.680 ;
        RECT 1367.650 427.620 1367.970 427.680 ;
        RECT 1365.810 427.480 1367.970 427.620 ;
        RECT 1365.810 427.420 1366.130 427.480 ;
        RECT 1367.650 427.420 1367.970 427.480 ;
        RECT 1365.810 379.680 1366.130 379.740 ;
        RECT 1366.730 379.680 1367.050 379.740 ;
        RECT 1365.810 379.540 1367.050 379.680 ;
        RECT 1365.810 379.480 1366.130 379.540 ;
        RECT 1366.730 379.480 1367.050 379.540 ;
        RECT 1365.810 379.000 1366.130 379.060 ;
        RECT 1366.730 379.000 1367.050 379.060 ;
        RECT 1365.810 378.860 1367.050 379.000 ;
        RECT 1365.810 378.800 1366.130 378.860 ;
        RECT 1366.730 378.800 1367.050 378.860 ;
        RECT 1365.810 351.460 1366.130 351.520 ;
        RECT 1367.190 351.460 1367.510 351.520 ;
        RECT 1365.810 351.320 1367.510 351.460 ;
        RECT 1365.810 351.260 1366.130 351.320 ;
        RECT 1367.190 351.260 1367.510 351.320 ;
        RECT 1367.190 303.520 1367.510 303.580 ;
        RECT 1368.110 303.520 1368.430 303.580 ;
        RECT 1367.190 303.380 1368.430 303.520 ;
        RECT 1367.190 303.320 1367.510 303.380 ;
        RECT 1368.110 303.320 1368.430 303.380 ;
        RECT 1366.730 289.580 1367.050 289.640 ;
        RECT 1368.110 289.580 1368.430 289.640 ;
        RECT 1366.730 289.440 1368.430 289.580 ;
        RECT 1366.730 289.380 1367.050 289.440 ;
        RECT 1368.110 289.380 1368.430 289.440 ;
        RECT 1366.730 241.640 1367.050 241.700 ;
        RECT 1367.650 241.640 1367.970 241.700 ;
        RECT 1366.730 241.500 1367.970 241.640 ;
        RECT 1366.730 241.440 1367.050 241.500 ;
        RECT 1367.650 241.440 1367.970 241.500 ;
        RECT 1367.650 210.360 1367.970 210.420 ;
        RECT 1368.570 210.360 1368.890 210.420 ;
        RECT 1367.650 210.220 1368.890 210.360 ;
        RECT 1367.650 210.160 1367.970 210.220 ;
        RECT 1368.570 210.160 1368.890 210.220 ;
        RECT 1367.650 186.560 1367.970 186.620 ;
        RECT 1368.570 186.560 1368.890 186.620 ;
        RECT 1367.650 186.420 1368.890 186.560 ;
        RECT 1367.650 186.360 1367.970 186.420 ;
        RECT 1368.570 186.360 1368.890 186.420 ;
        RECT 1367.190 110.400 1367.510 110.460 ;
        RECT 1368.110 110.400 1368.430 110.460 ;
        RECT 1367.190 110.260 1368.430 110.400 ;
        RECT 1367.190 110.200 1367.510 110.260 ;
        RECT 1368.110 110.200 1368.430 110.260 ;
        RECT 1367.190 96.460 1367.510 96.520 ;
        RECT 1368.110 96.460 1368.430 96.520 ;
        RECT 1367.190 96.320 1368.430 96.460 ;
        RECT 1367.190 96.260 1367.510 96.320 ;
        RECT 1368.110 96.260 1368.430 96.320 ;
        RECT 1364.430 20.640 1364.750 20.700 ;
        RECT 1368.110 20.640 1368.430 20.700 ;
        RECT 1364.430 20.500 1368.430 20.640 ;
        RECT 1364.430 20.440 1364.750 20.500 ;
        RECT 1368.110 20.440 1368.430 20.500 ;
      LAYER via ;
        RECT 1367.680 497.120 1367.940 497.380 ;
        RECT 1367.220 496.440 1367.480 496.700 ;
        RECT 1365.840 427.420 1366.100 427.680 ;
        RECT 1367.680 427.420 1367.940 427.680 ;
        RECT 1365.840 379.480 1366.100 379.740 ;
        RECT 1366.760 379.480 1367.020 379.740 ;
        RECT 1365.840 378.800 1366.100 379.060 ;
        RECT 1366.760 378.800 1367.020 379.060 ;
        RECT 1365.840 351.260 1366.100 351.520 ;
        RECT 1367.220 351.260 1367.480 351.520 ;
        RECT 1367.220 303.320 1367.480 303.580 ;
        RECT 1368.140 303.320 1368.400 303.580 ;
        RECT 1366.760 289.380 1367.020 289.640 ;
        RECT 1368.140 289.380 1368.400 289.640 ;
        RECT 1366.760 241.440 1367.020 241.700 ;
        RECT 1367.680 241.440 1367.940 241.700 ;
        RECT 1367.680 210.160 1367.940 210.420 ;
        RECT 1368.600 210.160 1368.860 210.420 ;
        RECT 1367.680 186.360 1367.940 186.620 ;
        RECT 1368.600 186.360 1368.860 186.620 ;
        RECT 1367.220 110.200 1367.480 110.460 ;
        RECT 1368.140 110.200 1368.400 110.460 ;
        RECT 1367.220 96.260 1367.480 96.520 ;
        RECT 1368.140 96.260 1368.400 96.520 ;
        RECT 1364.460 20.440 1364.720 20.700 ;
        RECT 1368.140 20.440 1368.400 20.700 ;
      LAYER met2 ;
        RECT 1370.670 600.170 1370.950 604.000 ;
        RECT 1369.580 600.030 1370.950 600.170 ;
        RECT 1369.580 579.885 1369.720 600.030 ;
        RECT 1370.670 600.000 1370.950 600.030 ;
        RECT 1368.590 579.515 1368.870 579.885 ;
        RECT 1369.510 579.515 1369.790 579.885 ;
        RECT 1368.660 545.090 1368.800 579.515 ;
        RECT 1367.740 544.950 1368.800 545.090 ;
        RECT 1367.740 497.410 1367.880 544.950 ;
        RECT 1367.680 497.090 1367.940 497.410 ;
        RECT 1367.220 496.410 1367.480 496.730 ;
        RECT 1367.280 434.930 1367.420 496.410 ;
        RECT 1367.280 434.790 1367.880 434.930 ;
        RECT 1367.740 427.710 1367.880 434.790 ;
        RECT 1365.840 427.390 1366.100 427.710 ;
        RECT 1367.680 427.390 1367.940 427.710 ;
        RECT 1365.900 379.770 1366.040 427.390 ;
        RECT 1365.840 379.450 1366.100 379.770 ;
        RECT 1366.760 379.450 1367.020 379.770 ;
        RECT 1366.820 379.090 1366.960 379.450 ;
        RECT 1365.840 378.770 1366.100 379.090 ;
        RECT 1366.760 378.770 1367.020 379.090 ;
        RECT 1365.900 351.550 1366.040 378.770 ;
        RECT 1365.840 351.230 1366.100 351.550 ;
        RECT 1367.220 351.230 1367.480 351.550 ;
        RECT 1367.280 303.610 1367.420 351.230 ;
        RECT 1367.220 303.290 1367.480 303.610 ;
        RECT 1368.140 303.290 1368.400 303.610 ;
        RECT 1368.200 289.670 1368.340 303.290 ;
        RECT 1366.760 289.350 1367.020 289.670 ;
        RECT 1368.140 289.350 1368.400 289.670 ;
        RECT 1366.820 241.730 1366.960 289.350 ;
        RECT 1366.760 241.410 1367.020 241.730 ;
        RECT 1367.680 241.410 1367.940 241.730 ;
        RECT 1367.740 210.450 1367.880 241.410 ;
        RECT 1367.680 210.130 1367.940 210.450 ;
        RECT 1368.600 210.130 1368.860 210.450 ;
        RECT 1368.660 186.650 1368.800 210.130 ;
        RECT 1367.680 186.330 1367.940 186.650 ;
        RECT 1368.600 186.330 1368.860 186.650 ;
        RECT 1367.740 157.490 1367.880 186.330 ;
        RECT 1367.280 157.350 1367.880 157.490 ;
        RECT 1367.280 110.490 1367.420 157.350 ;
        RECT 1367.220 110.170 1367.480 110.490 ;
        RECT 1368.140 110.170 1368.400 110.490 ;
        RECT 1368.200 96.550 1368.340 110.170 ;
        RECT 1367.220 96.230 1367.480 96.550 ;
        RECT 1368.140 96.230 1368.400 96.550 ;
        RECT 1367.280 60.930 1367.420 96.230 ;
        RECT 1367.280 60.790 1368.340 60.930 ;
        RECT 1368.200 20.730 1368.340 60.790 ;
        RECT 1364.460 20.410 1364.720 20.730 ;
        RECT 1368.140 20.410 1368.400 20.730 ;
        RECT 1364.520 2.400 1364.660 20.410 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
      LAYER via2 ;
        RECT 1368.590 579.560 1368.870 579.840 ;
        RECT 1369.510 579.560 1369.790 579.840 ;
      LAYER met3 ;
        RECT 1368.565 579.850 1368.895 579.865 ;
        RECT 1369.485 579.850 1369.815 579.865 ;
        RECT 1368.565 579.550 1369.815 579.850 ;
        RECT 1368.565 579.535 1368.895 579.550 ;
        RECT 1369.485 579.535 1369.815 579.550 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.990 579.600 1381.310 579.660 ;
        RECT 1381.910 579.600 1382.230 579.660 ;
        RECT 1380.990 579.460 1382.230 579.600 ;
        RECT 1380.990 579.400 1381.310 579.460 ;
        RECT 1381.910 579.400 1382.230 579.460 ;
        RECT 1380.990 531.660 1381.310 531.720 ;
        RECT 1381.910 531.660 1382.230 531.720 ;
        RECT 1380.990 531.520 1382.230 531.660 ;
        RECT 1380.990 531.460 1381.310 531.520 ;
        RECT 1381.910 531.460 1382.230 531.520 ;
        RECT 1380.990 483.040 1381.310 483.100 ;
        RECT 1381.910 483.040 1382.230 483.100 ;
        RECT 1380.990 482.900 1382.230 483.040 ;
        RECT 1380.990 482.840 1381.310 482.900 ;
        RECT 1381.910 482.840 1382.230 482.900 ;
        RECT 1380.990 435.100 1381.310 435.160 ;
        RECT 1381.910 435.100 1382.230 435.160 ;
        RECT 1380.990 434.960 1382.230 435.100 ;
        RECT 1380.990 434.900 1381.310 434.960 ;
        RECT 1381.910 434.900 1382.230 434.960 ;
        RECT 1380.990 289.580 1381.310 289.640 ;
        RECT 1381.910 289.580 1382.230 289.640 ;
        RECT 1380.990 289.440 1382.230 289.580 ;
        RECT 1380.990 289.380 1381.310 289.440 ;
        RECT 1381.910 289.380 1382.230 289.440 ;
        RECT 1380.990 241.640 1381.310 241.700 ;
        RECT 1381.910 241.640 1382.230 241.700 ;
        RECT 1380.990 241.500 1382.230 241.640 ;
        RECT 1380.990 241.440 1381.310 241.500 ;
        RECT 1381.910 241.440 1382.230 241.500 ;
        RECT 1380.990 193.020 1381.310 193.080 ;
        RECT 1381.910 193.020 1382.230 193.080 ;
        RECT 1380.990 192.880 1382.230 193.020 ;
        RECT 1380.990 192.820 1381.310 192.880 ;
        RECT 1381.910 192.820 1382.230 192.880 ;
        RECT 1380.990 145.080 1381.310 145.140 ;
        RECT 1381.910 145.080 1382.230 145.140 ;
        RECT 1380.990 144.940 1382.230 145.080 ;
        RECT 1380.990 144.880 1381.310 144.940 ;
        RECT 1381.910 144.880 1382.230 144.940 ;
        RECT 1380.990 96.460 1381.310 96.520 ;
        RECT 1381.910 96.460 1382.230 96.520 ;
        RECT 1380.990 96.320 1382.230 96.460 ;
        RECT 1380.990 96.260 1381.310 96.320 ;
        RECT 1381.910 96.260 1382.230 96.320 ;
        RECT 1380.990 48.520 1381.310 48.580 ;
        RECT 1381.910 48.520 1382.230 48.580 ;
        RECT 1380.990 48.380 1382.230 48.520 ;
        RECT 1380.990 48.320 1381.310 48.380 ;
        RECT 1381.910 48.320 1382.230 48.380 ;
        RECT 1380.990 13.980 1381.310 14.240 ;
        RECT 1381.080 13.840 1381.220 13.980 ;
        RECT 1381.910 13.840 1382.230 13.900 ;
        RECT 1381.080 13.700 1382.230 13.840 ;
        RECT 1381.910 13.640 1382.230 13.700 ;
        RECT 1381.910 2.960 1382.230 3.020 ;
        RECT 1382.370 2.960 1382.690 3.020 ;
        RECT 1381.910 2.820 1382.690 2.960 ;
        RECT 1381.910 2.760 1382.230 2.820 ;
        RECT 1382.370 2.760 1382.690 2.820 ;
      LAYER via ;
        RECT 1381.020 579.400 1381.280 579.660 ;
        RECT 1381.940 579.400 1382.200 579.660 ;
        RECT 1381.020 531.460 1381.280 531.720 ;
        RECT 1381.940 531.460 1382.200 531.720 ;
        RECT 1381.020 482.840 1381.280 483.100 ;
        RECT 1381.940 482.840 1382.200 483.100 ;
        RECT 1381.020 434.900 1381.280 435.160 ;
        RECT 1381.940 434.900 1382.200 435.160 ;
        RECT 1381.020 289.380 1381.280 289.640 ;
        RECT 1381.940 289.380 1382.200 289.640 ;
        RECT 1381.020 241.440 1381.280 241.700 ;
        RECT 1381.940 241.440 1382.200 241.700 ;
        RECT 1381.020 192.820 1381.280 193.080 ;
        RECT 1381.940 192.820 1382.200 193.080 ;
        RECT 1381.020 144.880 1381.280 145.140 ;
        RECT 1381.940 144.880 1382.200 145.140 ;
        RECT 1381.020 96.260 1381.280 96.520 ;
        RECT 1381.940 96.260 1382.200 96.520 ;
        RECT 1381.020 48.320 1381.280 48.580 ;
        RECT 1381.940 48.320 1382.200 48.580 ;
        RECT 1381.020 13.980 1381.280 14.240 ;
        RECT 1381.940 13.640 1382.200 13.900 ;
        RECT 1381.940 2.760 1382.200 3.020 ;
        RECT 1382.400 2.760 1382.660 3.020 ;
      LAYER met2 ;
        RECT 1379.870 600.170 1380.150 604.000 ;
        RECT 1379.870 600.030 1381.220 600.170 ;
        RECT 1379.870 600.000 1380.150 600.030 ;
        RECT 1381.080 579.690 1381.220 600.030 ;
        RECT 1381.020 579.370 1381.280 579.690 ;
        RECT 1381.940 579.370 1382.200 579.690 ;
        RECT 1382.000 531.750 1382.140 579.370 ;
        RECT 1381.020 531.430 1381.280 531.750 ;
        RECT 1381.940 531.430 1382.200 531.750 ;
        RECT 1381.080 483.130 1381.220 531.430 ;
        RECT 1381.020 482.810 1381.280 483.130 ;
        RECT 1381.940 482.810 1382.200 483.130 ;
        RECT 1382.000 435.190 1382.140 482.810 ;
        RECT 1381.020 434.870 1381.280 435.190 ;
        RECT 1381.940 434.870 1382.200 435.190 ;
        RECT 1381.080 289.670 1381.220 434.870 ;
        RECT 1381.020 289.350 1381.280 289.670 ;
        RECT 1381.940 289.350 1382.200 289.670 ;
        RECT 1382.000 241.730 1382.140 289.350 ;
        RECT 1381.020 241.410 1381.280 241.730 ;
        RECT 1381.940 241.410 1382.200 241.730 ;
        RECT 1381.080 193.110 1381.220 241.410 ;
        RECT 1381.020 192.790 1381.280 193.110 ;
        RECT 1381.940 192.790 1382.200 193.110 ;
        RECT 1382.000 145.170 1382.140 192.790 ;
        RECT 1381.020 144.850 1381.280 145.170 ;
        RECT 1381.940 144.850 1382.200 145.170 ;
        RECT 1381.080 96.550 1381.220 144.850 ;
        RECT 1381.020 96.230 1381.280 96.550 ;
        RECT 1381.940 96.230 1382.200 96.550 ;
        RECT 1382.000 48.610 1382.140 96.230 ;
        RECT 1381.020 48.290 1381.280 48.610 ;
        RECT 1381.940 48.290 1382.200 48.610 ;
        RECT 1381.080 14.270 1381.220 48.290 ;
        RECT 1381.020 13.950 1381.280 14.270 ;
        RECT 1381.940 13.610 1382.200 13.930 ;
        RECT 1382.000 3.050 1382.140 13.610 ;
        RECT 1381.940 2.730 1382.200 3.050 ;
        RECT 1382.400 2.730 1382.660 3.050 ;
        RECT 1382.460 2.400 1382.600 2.730 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1390.650 586.740 1390.970 586.800 ;
        RECT 1393.410 586.740 1393.730 586.800 ;
        RECT 1390.650 586.600 1393.730 586.740 ;
        RECT 1390.650 586.540 1390.970 586.600 ;
        RECT 1393.410 586.540 1393.730 586.600 ;
        RECT 1393.410 20.300 1393.730 20.360 ;
        RECT 1400.310 20.300 1400.630 20.360 ;
        RECT 1393.410 20.160 1400.630 20.300 ;
        RECT 1393.410 20.100 1393.730 20.160 ;
        RECT 1400.310 20.100 1400.630 20.160 ;
      LAYER via ;
        RECT 1390.680 586.540 1390.940 586.800 ;
        RECT 1393.440 586.540 1393.700 586.800 ;
        RECT 1393.440 20.100 1393.700 20.360 ;
        RECT 1400.340 20.100 1400.600 20.360 ;
      LAYER met2 ;
        RECT 1389.070 600.170 1389.350 604.000 ;
        RECT 1389.070 600.030 1390.880 600.170 ;
        RECT 1389.070 600.000 1389.350 600.030 ;
        RECT 1390.740 586.830 1390.880 600.030 ;
        RECT 1390.680 586.510 1390.940 586.830 ;
        RECT 1393.440 586.510 1393.700 586.830 ;
        RECT 1393.500 20.390 1393.640 586.510 ;
        RECT 1393.440 20.070 1393.700 20.390 ;
        RECT 1400.340 20.070 1400.600 20.390 ;
        RECT 1400.400 2.400 1400.540 20.070 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1399.850 17.580 1400.170 17.640 ;
        RECT 1418.250 17.580 1418.570 17.640 ;
        RECT 1399.850 17.440 1418.570 17.580 ;
        RECT 1399.850 17.380 1400.170 17.440 ;
        RECT 1418.250 17.380 1418.570 17.440 ;
      LAYER via ;
        RECT 1399.880 17.380 1400.140 17.640 ;
        RECT 1418.280 17.380 1418.540 17.640 ;
      LAYER met2 ;
        RECT 1398.270 600.170 1398.550 604.000 ;
        RECT 1398.270 600.030 1400.080 600.170 ;
        RECT 1398.270 600.000 1398.550 600.030 ;
        RECT 1399.940 17.670 1400.080 600.030 ;
        RECT 1399.880 17.350 1400.140 17.670 ;
        RECT 1418.280 17.350 1418.540 17.670 ;
        RECT 1418.340 2.400 1418.480 17.350 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1409.050 586.740 1409.370 586.800 ;
        RECT 1413.190 586.740 1413.510 586.800 ;
        RECT 1409.050 586.600 1413.510 586.740 ;
        RECT 1409.050 586.540 1409.370 586.600 ;
        RECT 1413.190 586.540 1413.510 586.600 ;
        RECT 1413.190 19.620 1413.510 19.680 ;
        RECT 1435.730 19.620 1436.050 19.680 ;
        RECT 1413.190 19.480 1436.050 19.620 ;
        RECT 1413.190 19.420 1413.510 19.480 ;
        RECT 1435.730 19.420 1436.050 19.480 ;
      LAYER via ;
        RECT 1409.080 586.540 1409.340 586.800 ;
        RECT 1413.220 586.540 1413.480 586.800 ;
        RECT 1413.220 19.420 1413.480 19.680 ;
        RECT 1435.760 19.420 1436.020 19.680 ;
      LAYER met2 ;
        RECT 1407.470 600.170 1407.750 604.000 ;
        RECT 1407.470 600.030 1409.280 600.170 ;
        RECT 1407.470 600.000 1407.750 600.030 ;
        RECT 1409.140 586.830 1409.280 600.030 ;
        RECT 1409.080 586.510 1409.340 586.830 ;
        RECT 1413.220 586.510 1413.480 586.830 ;
        RECT 1413.280 19.710 1413.420 586.510 ;
        RECT 1413.220 19.390 1413.480 19.710 ;
        RECT 1435.760 19.390 1436.020 19.710 ;
        RECT 1435.820 2.400 1435.960 19.390 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1418.250 586.740 1418.570 586.800 ;
        RECT 1421.010 586.740 1421.330 586.800 ;
        RECT 1418.250 586.600 1421.330 586.740 ;
        RECT 1418.250 586.540 1418.570 586.600 ;
        RECT 1421.010 586.540 1421.330 586.600 ;
        RECT 1421.010 18.600 1421.330 18.660 ;
        RECT 1453.670 18.600 1453.990 18.660 ;
        RECT 1421.010 18.460 1453.990 18.600 ;
        RECT 1421.010 18.400 1421.330 18.460 ;
        RECT 1453.670 18.400 1453.990 18.460 ;
      LAYER via ;
        RECT 1418.280 586.540 1418.540 586.800 ;
        RECT 1421.040 586.540 1421.300 586.800 ;
        RECT 1421.040 18.400 1421.300 18.660 ;
        RECT 1453.700 18.400 1453.960 18.660 ;
      LAYER met2 ;
        RECT 1416.670 600.170 1416.950 604.000 ;
        RECT 1416.670 600.030 1418.480 600.170 ;
        RECT 1416.670 600.000 1416.950 600.030 ;
        RECT 1418.340 586.830 1418.480 600.030 ;
        RECT 1418.280 586.510 1418.540 586.830 ;
        RECT 1421.040 586.510 1421.300 586.830 ;
        RECT 1421.100 18.690 1421.240 586.510 ;
        RECT 1421.040 18.370 1421.300 18.690 ;
        RECT 1453.700 18.370 1453.960 18.690 ;
        RECT 1453.760 2.400 1453.900 18.370 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1427.450 17.580 1427.770 17.640 ;
        RECT 1427.450 17.440 1430.440 17.580 ;
        RECT 1427.450 17.380 1427.770 17.440 ;
        RECT 1430.300 17.240 1430.440 17.440 ;
        RECT 1471.610 17.240 1471.930 17.300 ;
        RECT 1430.300 17.100 1471.930 17.240 ;
        RECT 1471.610 17.040 1471.930 17.100 ;
      LAYER via ;
        RECT 1427.480 17.380 1427.740 17.640 ;
        RECT 1471.640 17.040 1471.900 17.300 ;
      LAYER met2 ;
        RECT 1425.870 600.170 1426.150 604.000 ;
        RECT 1425.870 600.030 1427.680 600.170 ;
        RECT 1425.870 600.000 1426.150 600.030 ;
        RECT 1427.540 17.670 1427.680 600.030 ;
        RECT 1427.480 17.350 1427.740 17.670 ;
        RECT 1471.640 17.010 1471.900 17.330 ;
        RECT 1471.700 2.400 1471.840 17.010 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1436.650 586.740 1436.970 586.800 ;
        RECT 1440.790 586.740 1441.110 586.800 ;
        RECT 1436.650 586.600 1441.110 586.740 ;
        RECT 1436.650 586.540 1436.970 586.600 ;
        RECT 1440.790 586.540 1441.110 586.600 ;
        RECT 1440.790 16.900 1441.110 16.960 ;
        RECT 1489.550 16.900 1489.870 16.960 ;
        RECT 1440.790 16.760 1489.870 16.900 ;
        RECT 1440.790 16.700 1441.110 16.760 ;
        RECT 1489.550 16.700 1489.870 16.760 ;
      LAYER via ;
        RECT 1436.680 586.540 1436.940 586.800 ;
        RECT 1440.820 586.540 1441.080 586.800 ;
        RECT 1440.820 16.700 1441.080 16.960 ;
        RECT 1489.580 16.700 1489.840 16.960 ;
      LAYER met2 ;
        RECT 1435.070 600.170 1435.350 604.000 ;
        RECT 1435.070 600.030 1436.880 600.170 ;
        RECT 1435.070 600.000 1435.350 600.030 ;
        RECT 1436.740 586.830 1436.880 600.030 ;
        RECT 1436.680 586.510 1436.940 586.830 ;
        RECT 1440.820 586.510 1441.080 586.830 ;
        RECT 1440.880 16.990 1441.020 586.510 ;
        RECT 1440.820 16.670 1441.080 16.990 ;
        RECT 1489.580 16.670 1489.840 16.990 ;
        RECT 1489.640 2.400 1489.780 16.670 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1445.850 590.820 1446.170 590.880 ;
        RECT 1504.730 590.820 1505.050 590.880 ;
        RECT 1445.850 590.680 1505.050 590.820 ;
        RECT 1445.850 590.620 1446.170 590.680 ;
        RECT 1504.730 590.620 1505.050 590.680 ;
        RECT 1504.730 2.960 1505.050 3.020 ;
        RECT 1507.030 2.960 1507.350 3.020 ;
        RECT 1504.730 2.820 1507.350 2.960 ;
        RECT 1504.730 2.760 1505.050 2.820 ;
        RECT 1507.030 2.760 1507.350 2.820 ;
      LAYER via ;
        RECT 1445.880 590.620 1446.140 590.880 ;
        RECT 1504.760 590.620 1505.020 590.880 ;
        RECT 1504.760 2.760 1505.020 3.020 ;
        RECT 1507.060 2.760 1507.320 3.020 ;
      LAYER met2 ;
        RECT 1444.270 600.170 1444.550 604.000 ;
        RECT 1444.270 600.030 1446.080 600.170 ;
        RECT 1444.270 600.000 1444.550 600.030 ;
        RECT 1445.940 590.910 1446.080 600.030 ;
        RECT 1445.880 590.590 1446.140 590.910 ;
        RECT 1504.760 590.590 1505.020 590.910 ;
        RECT 1504.820 3.050 1504.960 590.590 ;
        RECT 1504.760 2.730 1505.020 3.050 ;
        RECT 1507.060 2.730 1507.320 3.050 ;
        RECT 1507.120 2.400 1507.260 2.730 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1029.090 496.980 1029.410 497.040 ;
        RECT 1030.010 496.980 1030.330 497.040 ;
        RECT 1029.090 496.840 1030.330 496.980 ;
        RECT 1029.090 496.780 1029.410 496.840 ;
        RECT 1030.010 496.780 1030.330 496.840 ;
        RECT 1028.170 449.380 1028.490 449.440 ;
        RECT 1029.090 449.380 1029.410 449.440 ;
        RECT 1028.170 449.240 1029.410 449.380 ;
        RECT 1028.170 449.180 1028.490 449.240 ;
        RECT 1029.090 449.180 1029.410 449.240 ;
        RECT 704.330 38.320 704.650 38.380 ;
        RECT 1028.170 38.320 1028.490 38.380 ;
        RECT 704.330 38.180 1028.490 38.320 ;
        RECT 704.330 38.120 704.650 38.180 ;
        RECT 1028.170 38.120 1028.490 38.180 ;
      LAYER via ;
        RECT 1029.120 496.780 1029.380 497.040 ;
        RECT 1030.040 496.780 1030.300 497.040 ;
        RECT 1028.200 449.180 1028.460 449.440 ;
        RECT 1029.120 449.180 1029.380 449.440 ;
        RECT 704.360 38.120 704.620 38.380 ;
        RECT 1028.200 38.120 1028.460 38.380 ;
      LAYER met2 ;
        RECT 1031.650 600.170 1031.930 604.000 ;
        RECT 1030.100 600.030 1031.930 600.170 ;
        RECT 1030.100 497.070 1030.240 600.030 ;
        RECT 1031.650 600.000 1031.930 600.030 ;
        RECT 1029.120 496.750 1029.380 497.070 ;
        RECT 1030.040 496.750 1030.300 497.070 ;
        RECT 1029.180 449.470 1029.320 496.750 ;
        RECT 1028.200 449.150 1028.460 449.470 ;
        RECT 1029.120 449.150 1029.380 449.470 ;
        RECT 1028.260 38.410 1028.400 449.150 ;
        RECT 704.360 38.090 704.620 38.410 ;
        RECT 1028.200 38.090 1028.460 38.410 ;
        RECT 704.420 2.400 704.560 38.090 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.050 590.140 1455.370 590.200 ;
        RECT 1525.430 590.140 1525.750 590.200 ;
        RECT 1455.050 590.000 1525.750 590.140 ;
        RECT 1455.050 589.940 1455.370 590.000 ;
        RECT 1525.430 589.940 1525.750 590.000 ;
      LAYER via ;
        RECT 1455.080 589.940 1455.340 590.200 ;
        RECT 1525.460 589.940 1525.720 590.200 ;
      LAYER met2 ;
        RECT 1453.470 600.170 1453.750 604.000 ;
        RECT 1453.470 600.030 1455.280 600.170 ;
        RECT 1453.470 600.000 1453.750 600.030 ;
        RECT 1455.140 590.230 1455.280 600.030 ;
        RECT 1455.080 589.910 1455.340 590.230 ;
        RECT 1525.460 589.910 1525.720 590.230 ;
        RECT 1525.520 3.130 1525.660 589.910 ;
        RECT 1525.060 2.990 1525.660 3.130 ;
        RECT 1525.060 2.400 1525.200 2.990 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1464.250 588.440 1464.570 588.500 ;
        RECT 1540.150 588.440 1540.470 588.500 ;
        RECT 1464.250 588.300 1540.470 588.440 ;
        RECT 1464.250 588.240 1464.570 588.300 ;
        RECT 1540.150 588.240 1540.470 588.300 ;
        RECT 1540.150 2.960 1540.470 3.020 ;
        RECT 1542.910 2.960 1543.230 3.020 ;
        RECT 1540.150 2.820 1543.230 2.960 ;
        RECT 1540.150 2.760 1540.470 2.820 ;
        RECT 1542.910 2.760 1543.230 2.820 ;
      LAYER via ;
        RECT 1464.280 588.240 1464.540 588.500 ;
        RECT 1540.180 588.240 1540.440 588.500 ;
        RECT 1540.180 2.760 1540.440 3.020 ;
        RECT 1542.940 2.760 1543.200 3.020 ;
      LAYER met2 ;
        RECT 1462.670 600.170 1462.950 604.000 ;
        RECT 1462.670 600.030 1464.480 600.170 ;
        RECT 1462.670 600.000 1462.950 600.030 ;
        RECT 1464.340 588.530 1464.480 600.030 ;
        RECT 1464.280 588.210 1464.540 588.530 ;
        RECT 1540.180 588.210 1540.440 588.530 ;
        RECT 1540.240 3.050 1540.380 588.210 ;
        RECT 1540.180 2.730 1540.440 3.050 ;
        RECT 1542.940 2.730 1543.200 3.050 ;
        RECT 1543.000 2.400 1543.140 2.730 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1473.450 592.860 1473.770 592.920 ;
        RECT 1560.390 592.860 1560.710 592.920 ;
        RECT 1473.450 592.720 1560.710 592.860 ;
        RECT 1473.450 592.660 1473.770 592.720 ;
        RECT 1560.390 592.660 1560.710 592.720 ;
      LAYER via ;
        RECT 1473.480 592.660 1473.740 592.920 ;
        RECT 1560.420 592.660 1560.680 592.920 ;
      LAYER met2 ;
        RECT 1471.870 600.170 1472.150 604.000 ;
        RECT 1471.870 600.030 1473.680 600.170 ;
        RECT 1471.870 600.000 1472.150 600.030 ;
        RECT 1473.540 592.950 1473.680 600.030 ;
        RECT 1473.480 592.630 1473.740 592.950 ;
        RECT 1560.420 592.630 1560.680 592.950 ;
        RECT 1560.480 3.130 1560.620 592.630 ;
        RECT 1560.480 2.990 1561.080 3.130 ;
        RECT 1560.940 2.400 1561.080 2.990 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1482.190 589.460 1482.510 589.520 ;
        RECT 1573.270 589.460 1573.590 589.520 ;
        RECT 1482.190 589.320 1573.590 589.460 ;
        RECT 1482.190 589.260 1482.510 589.320 ;
        RECT 1573.270 589.260 1573.590 589.320 ;
        RECT 1573.270 2.960 1573.590 3.020 ;
        RECT 1578.790 2.960 1579.110 3.020 ;
        RECT 1573.270 2.820 1579.110 2.960 ;
        RECT 1573.270 2.760 1573.590 2.820 ;
        RECT 1578.790 2.760 1579.110 2.820 ;
      LAYER via ;
        RECT 1482.220 589.260 1482.480 589.520 ;
        RECT 1573.300 589.260 1573.560 589.520 ;
        RECT 1573.300 2.760 1573.560 3.020 ;
        RECT 1578.820 2.760 1579.080 3.020 ;
      LAYER met2 ;
        RECT 1481.070 600.170 1481.350 604.000 ;
        RECT 1481.070 600.030 1482.420 600.170 ;
        RECT 1481.070 600.000 1481.350 600.030 ;
        RECT 1482.280 589.550 1482.420 600.030 ;
        RECT 1482.220 589.230 1482.480 589.550 ;
        RECT 1573.300 589.230 1573.560 589.550 ;
        RECT 1573.360 3.050 1573.500 589.230 ;
        RECT 1573.300 2.730 1573.560 3.050 ;
        RECT 1578.820 2.730 1579.080 3.050 ;
        RECT 1578.880 2.400 1579.020 2.730 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 588.100 1490.330 588.160 ;
        RECT 1595.350 588.100 1595.670 588.160 ;
        RECT 1490.010 587.960 1595.670 588.100 ;
        RECT 1490.010 587.900 1490.330 587.960 ;
        RECT 1595.350 587.900 1595.670 587.960 ;
        RECT 1595.350 579.600 1595.670 579.660 ;
        RECT 1596.270 579.600 1596.590 579.660 ;
        RECT 1595.350 579.460 1596.590 579.600 ;
        RECT 1595.350 579.400 1595.670 579.460 ;
        RECT 1596.270 579.400 1596.590 579.460 ;
        RECT 1595.350 531.660 1595.670 531.720 ;
        RECT 1596.270 531.660 1596.590 531.720 ;
        RECT 1595.350 531.520 1596.590 531.660 ;
        RECT 1595.350 531.460 1595.670 531.520 ;
        RECT 1596.270 531.460 1596.590 531.520 ;
        RECT 1595.350 289.580 1595.670 289.640 ;
        RECT 1596.270 289.580 1596.590 289.640 ;
        RECT 1595.350 289.440 1596.590 289.580 ;
        RECT 1595.350 289.380 1595.670 289.440 ;
        RECT 1596.270 289.380 1596.590 289.440 ;
        RECT 1595.350 241.640 1595.670 241.700 ;
        RECT 1596.270 241.640 1596.590 241.700 ;
        RECT 1595.350 241.500 1596.590 241.640 ;
        RECT 1595.350 241.440 1595.670 241.500 ;
        RECT 1596.270 241.440 1596.590 241.500 ;
        RECT 1595.350 193.020 1595.670 193.080 ;
        RECT 1596.270 193.020 1596.590 193.080 ;
        RECT 1595.350 192.880 1596.590 193.020 ;
        RECT 1595.350 192.820 1595.670 192.880 ;
        RECT 1596.270 192.820 1596.590 192.880 ;
        RECT 1595.350 145.080 1595.670 145.140 ;
        RECT 1596.270 145.080 1596.590 145.140 ;
        RECT 1595.350 144.940 1596.590 145.080 ;
        RECT 1595.350 144.880 1595.670 144.940 ;
        RECT 1596.270 144.880 1596.590 144.940 ;
        RECT 1595.350 96.460 1595.670 96.520 ;
        RECT 1596.270 96.460 1596.590 96.520 ;
        RECT 1595.350 96.320 1596.590 96.460 ;
        RECT 1595.350 96.260 1595.670 96.320 ;
        RECT 1596.270 96.260 1596.590 96.320 ;
        RECT 1595.350 48.520 1595.670 48.580 ;
        RECT 1596.270 48.520 1596.590 48.580 ;
        RECT 1595.350 48.380 1596.590 48.520 ;
        RECT 1595.350 48.320 1595.670 48.380 ;
        RECT 1596.270 48.320 1596.590 48.380 ;
        RECT 1595.350 14.180 1595.670 14.240 ;
        RECT 1595.350 14.040 1596.040 14.180 ;
        RECT 1595.350 13.980 1595.670 14.040 ;
        RECT 1595.900 13.900 1596.040 14.040 ;
        RECT 1595.810 13.640 1596.130 13.900 ;
        RECT 1595.810 2.960 1596.130 3.020 ;
        RECT 1596.270 2.960 1596.590 3.020 ;
        RECT 1595.810 2.820 1596.590 2.960 ;
        RECT 1595.810 2.760 1596.130 2.820 ;
        RECT 1596.270 2.760 1596.590 2.820 ;
      LAYER via ;
        RECT 1490.040 587.900 1490.300 588.160 ;
        RECT 1595.380 587.900 1595.640 588.160 ;
        RECT 1595.380 579.400 1595.640 579.660 ;
        RECT 1596.300 579.400 1596.560 579.660 ;
        RECT 1595.380 531.460 1595.640 531.720 ;
        RECT 1596.300 531.460 1596.560 531.720 ;
        RECT 1595.380 289.380 1595.640 289.640 ;
        RECT 1596.300 289.380 1596.560 289.640 ;
        RECT 1595.380 241.440 1595.640 241.700 ;
        RECT 1596.300 241.440 1596.560 241.700 ;
        RECT 1595.380 192.820 1595.640 193.080 ;
        RECT 1596.300 192.820 1596.560 193.080 ;
        RECT 1595.380 144.880 1595.640 145.140 ;
        RECT 1596.300 144.880 1596.560 145.140 ;
        RECT 1595.380 96.260 1595.640 96.520 ;
        RECT 1596.300 96.260 1596.560 96.520 ;
        RECT 1595.380 48.320 1595.640 48.580 ;
        RECT 1596.300 48.320 1596.560 48.580 ;
        RECT 1595.380 13.980 1595.640 14.240 ;
        RECT 1595.840 13.640 1596.100 13.900 ;
        RECT 1595.840 2.760 1596.100 3.020 ;
        RECT 1596.300 2.760 1596.560 3.020 ;
      LAYER met2 ;
        RECT 1489.810 600.000 1490.090 604.000 ;
        RECT 1489.870 598.810 1490.010 600.000 ;
        RECT 1489.870 598.670 1490.240 598.810 ;
        RECT 1490.100 588.190 1490.240 598.670 ;
        RECT 1490.040 587.870 1490.300 588.190 ;
        RECT 1595.380 587.870 1595.640 588.190 ;
        RECT 1595.440 579.690 1595.580 587.870 ;
        RECT 1595.380 579.370 1595.640 579.690 ;
        RECT 1596.300 579.370 1596.560 579.690 ;
        RECT 1596.360 531.750 1596.500 579.370 ;
        RECT 1595.380 531.430 1595.640 531.750 ;
        RECT 1596.300 531.430 1596.560 531.750 ;
        RECT 1595.440 289.670 1595.580 531.430 ;
        RECT 1595.380 289.350 1595.640 289.670 ;
        RECT 1596.300 289.350 1596.560 289.670 ;
        RECT 1596.360 241.730 1596.500 289.350 ;
        RECT 1595.380 241.410 1595.640 241.730 ;
        RECT 1596.300 241.410 1596.560 241.730 ;
        RECT 1595.440 193.110 1595.580 241.410 ;
        RECT 1595.380 192.790 1595.640 193.110 ;
        RECT 1596.300 192.790 1596.560 193.110 ;
        RECT 1596.360 145.170 1596.500 192.790 ;
        RECT 1595.380 144.850 1595.640 145.170 ;
        RECT 1596.300 144.850 1596.560 145.170 ;
        RECT 1595.440 96.550 1595.580 144.850 ;
        RECT 1595.380 96.230 1595.640 96.550 ;
        RECT 1596.300 96.230 1596.560 96.550 ;
        RECT 1596.360 48.610 1596.500 96.230 ;
        RECT 1595.380 48.290 1595.640 48.610 ;
        RECT 1596.300 48.290 1596.560 48.610 ;
        RECT 1595.440 14.270 1595.580 48.290 ;
        RECT 1595.380 13.950 1595.640 14.270 ;
        RECT 1595.840 13.610 1596.100 13.930 ;
        RECT 1595.900 3.050 1596.040 13.610 ;
        RECT 1595.840 2.730 1596.100 3.050 ;
        RECT 1596.300 2.730 1596.560 3.050 ;
        RECT 1596.360 2.400 1596.500 2.730 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 592.520 1500.910 592.580 ;
        RECT 1608.230 592.520 1608.550 592.580 ;
        RECT 1500.590 592.380 1608.550 592.520 ;
        RECT 1500.590 592.320 1500.910 592.380 ;
        RECT 1608.230 592.320 1608.550 592.380 ;
        RECT 1608.230 37.980 1608.550 38.040 ;
        RECT 1614.210 37.980 1614.530 38.040 ;
        RECT 1608.230 37.840 1614.530 37.980 ;
        RECT 1608.230 37.780 1608.550 37.840 ;
        RECT 1614.210 37.780 1614.530 37.840 ;
      LAYER via ;
        RECT 1500.620 592.320 1500.880 592.580 ;
        RECT 1608.260 592.320 1608.520 592.580 ;
        RECT 1608.260 37.780 1608.520 38.040 ;
        RECT 1614.240 37.780 1614.500 38.040 ;
      LAYER met2 ;
        RECT 1499.010 600.170 1499.290 604.000 ;
        RECT 1499.010 600.030 1500.820 600.170 ;
        RECT 1499.010 600.000 1499.290 600.030 ;
        RECT 1500.680 592.610 1500.820 600.030 ;
        RECT 1500.620 592.290 1500.880 592.610 ;
        RECT 1608.260 592.290 1608.520 592.610 ;
        RECT 1608.320 38.070 1608.460 592.290 ;
        RECT 1608.260 37.750 1608.520 38.070 ;
        RECT 1614.240 37.750 1614.500 38.070 ;
        RECT 1614.300 2.400 1614.440 37.750 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 587.420 1545.530 587.480 ;
        RECT 1545.210 587.280 1593.970 587.420 ;
        RECT 1545.210 587.220 1545.530 587.280 ;
        RECT 1593.830 587.080 1593.970 587.280 ;
        RECT 1606.390 587.080 1606.710 587.140 ;
        RECT 1593.830 586.940 1606.710 587.080 ;
        RECT 1606.390 586.880 1606.710 586.940 ;
        RECT 1606.390 583.340 1606.710 583.400 ;
        RECT 1629.390 583.340 1629.710 583.400 ;
        RECT 1606.390 583.200 1629.710 583.340 ;
        RECT 1606.390 583.140 1606.710 583.200 ;
        RECT 1629.390 583.140 1629.710 583.200 ;
        RECT 1629.390 2.960 1629.710 3.020 ;
        RECT 1632.150 2.960 1632.470 3.020 ;
        RECT 1629.390 2.820 1632.470 2.960 ;
        RECT 1629.390 2.760 1629.710 2.820 ;
        RECT 1632.150 2.760 1632.470 2.820 ;
      LAYER via ;
        RECT 1545.240 587.220 1545.500 587.480 ;
        RECT 1606.420 586.880 1606.680 587.140 ;
        RECT 1606.420 583.140 1606.680 583.400 ;
        RECT 1629.420 583.140 1629.680 583.400 ;
        RECT 1629.420 2.760 1629.680 3.020 ;
        RECT 1632.180 2.760 1632.440 3.020 ;
      LAYER met2 ;
        RECT 1508.210 600.170 1508.490 604.000 ;
        RECT 1508.210 600.030 1510.020 600.170 ;
        RECT 1508.210 600.000 1508.490 600.030 ;
        RECT 1509.880 587.365 1510.020 600.030 ;
        RECT 1545.240 587.365 1545.500 587.510 ;
        RECT 1509.810 586.995 1510.090 587.365 ;
        RECT 1545.230 586.995 1545.510 587.365 ;
        RECT 1606.420 586.850 1606.680 587.170 ;
        RECT 1606.480 583.430 1606.620 586.850 ;
        RECT 1606.420 583.110 1606.680 583.430 ;
        RECT 1629.420 583.110 1629.680 583.430 ;
        RECT 1629.480 3.050 1629.620 583.110 ;
        RECT 1629.420 2.730 1629.680 3.050 ;
        RECT 1632.180 2.730 1632.440 3.050 ;
        RECT 1632.240 2.400 1632.380 2.730 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
      LAYER via2 ;
        RECT 1509.810 587.040 1510.090 587.320 ;
        RECT 1545.230 587.040 1545.510 587.320 ;
      LAYER met3 ;
        RECT 1509.785 587.330 1510.115 587.345 ;
        RECT 1545.205 587.330 1545.535 587.345 ;
        RECT 1509.785 587.030 1545.535 587.330 ;
        RECT 1509.785 587.015 1510.115 587.030 ;
        RECT 1545.205 587.015 1545.535 587.030 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.150 591.160 1517.470 591.220 ;
        RECT 1651.010 591.160 1651.330 591.220 ;
        RECT 1517.150 591.020 1651.330 591.160 ;
        RECT 1517.150 590.960 1517.470 591.020 ;
        RECT 1651.010 590.960 1651.330 591.020 ;
        RECT 1651.010 531.120 1651.330 531.380 ;
        RECT 1651.100 530.980 1651.240 531.120 ;
        RECT 1651.930 530.980 1652.250 531.040 ;
        RECT 1651.100 530.840 1652.250 530.980 ;
        RECT 1651.930 530.780 1652.250 530.840 ;
        RECT 1649.170 434.760 1649.490 434.820 ;
        RECT 1650.550 434.760 1650.870 434.820 ;
        RECT 1649.170 434.620 1650.870 434.760 ;
        RECT 1649.170 434.560 1649.490 434.620 ;
        RECT 1650.550 434.560 1650.870 434.620 ;
        RECT 1649.170 386.480 1649.490 386.540 ;
        RECT 1650.090 386.480 1650.410 386.540 ;
        RECT 1649.170 386.340 1650.410 386.480 ;
        RECT 1649.170 386.280 1649.490 386.340 ;
        RECT 1650.090 386.280 1650.410 386.340 ;
        RECT 1650.090 331.060 1650.410 331.120 ;
        RECT 1650.550 331.060 1650.870 331.120 ;
        RECT 1650.090 330.920 1650.870 331.060 ;
        RECT 1650.090 330.860 1650.410 330.920 ;
        RECT 1650.550 330.860 1650.870 330.920 ;
        RECT 1650.090 283.120 1650.410 283.180 ;
        RECT 1651.010 283.120 1651.330 283.180 ;
        RECT 1650.090 282.980 1651.330 283.120 ;
        RECT 1650.090 282.920 1650.410 282.980 ;
        RECT 1651.010 282.920 1651.330 282.980 ;
        RECT 1649.170 234.500 1649.490 234.560 ;
        RECT 1651.010 234.500 1651.330 234.560 ;
        RECT 1649.170 234.360 1651.330 234.500 ;
        RECT 1649.170 234.300 1649.490 234.360 ;
        RECT 1651.010 234.300 1651.330 234.360 ;
        RECT 1649.170 186.560 1649.490 186.620 ;
        RECT 1650.090 186.560 1650.410 186.620 ;
        RECT 1649.170 186.420 1650.410 186.560 ;
        RECT 1649.170 186.360 1649.490 186.420 ;
        RECT 1650.090 186.360 1650.410 186.420 ;
        RECT 1650.550 138.280 1650.870 138.340 ;
        RECT 1651.930 138.280 1652.250 138.340 ;
        RECT 1650.550 138.140 1652.250 138.280 ;
        RECT 1650.550 138.080 1650.870 138.140 ;
        RECT 1651.930 138.080 1652.250 138.140 ;
        RECT 1650.550 110.400 1650.870 110.460 ;
        RECT 1651.470 110.400 1651.790 110.460 ;
        RECT 1650.550 110.260 1651.790 110.400 ;
        RECT 1650.550 110.200 1650.870 110.260 ;
        RECT 1651.470 110.200 1651.790 110.260 ;
        RECT 1650.090 96.460 1650.410 96.520 ;
        RECT 1651.470 96.460 1651.790 96.520 ;
        RECT 1650.090 96.320 1651.790 96.460 ;
        RECT 1650.090 96.260 1650.410 96.320 ;
        RECT 1651.470 96.260 1651.790 96.320 ;
        RECT 1650.090 48.520 1650.410 48.580 ;
        RECT 1651.010 48.520 1651.330 48.580 ;
        RECT 1650.090 48.380 1651.330 48.520 ;
        RECT 1650.090 48.320 1650.410 48.380 ;
        RECT 1651.010 48.320 1651.330 48.380 ;
        RECT 1650.090 2.960 1650.410 3.020 ;
        RECT 1651.010 2.960 1651.330 3.020 ;
        RECT 1650.090 2.820 1651.330 2.960 ;
        RECT 1650.090 2.760 1650.410 2.820 ;
        RECT 1651.010 2.760 1651.330 2.820 ;
      LAYER via ;
        RECT 1517.180 590.960 1517.440 591.220 ;
        RECT 1651.040 590.960 1651.300 591.220 ;
        RECT 1651.040 531.120 1651.300 531.380 ;
        RECT 1651.960 530.780 1652.220 531.040 ;
        RECT 1649.200 434.560 1649.460 434.820 ;
        RECT 1650.580 434.560 1650.840 434.820 ;
        RECT 1649.200 386.280 1649.460 386.540 ;
        RECT 1650.120 386.280 1650.380 386.540 ;
        RECT 1650.120 330.860 1650.380 331.120 ;
        RECT 1650.580 330.860 1650.840 331.120 ;
        RECT 1650.120 282.920 1650.380 283.180 ;
        RECT 1651.040 282.920 1651.300 283.180 ;
        RECT 1649.200 234.300 1649.460 234.560 ;
        RECT 1651.040 234.300 1651.300 234.560 ;
        RECT 1649.200 186.360 1649.460 186.620 ;
        RECT 1650.120 186.360 1650.380 186.620 ;
        RECT 1650.580 138.080 1650.840 138.340 ;
        RECT 1651.960 138.080 1652.220 138.340 ;
        RECT 1650.580 110.200 1650.840 110.460 ;
        RECT 1651.500 110.200 1651.760 110.460 ;
        RECT 1650.120 96.260 1650.380 96.520 ;
        RECT 1651.500 96.260 1651.760 96.520 ;
        RECT 1650.120 48.320 1650.380 48.580 ;
        RECT 1651.040 48.320 1651.300 48.580 ;
        RECT 1650.120 2.760 1650.380 3.020 ;
        RECT 1651.040 2.760 1651.300 3.020 ;
      LAYER met2 ;
        RECT 1517.410 600.000 1517.690 604.000 ;
        RECT 1517.470 598.810 1517.610 600.000 ;
        RECT 1517.240 598.670 1517.610 598.810 ;
        RECT 1517.240 591.250 1517.380 598.670 ;
        RECT 1517.180 590.930 1517.440 591.250 ;
        RECT 1651.040 590.930 1651.300 591.250 ;
        RECT 1651.100 531.410 1651.240 590.930 ;
        RECT 1651.040 531.090 1651.300 531.410 ;
        RECT 1651.960 530.750 1652.220 531.070 ;
        RECT 1652.020 448.530 1652.160 530.750 ;
        RECT 1650.640 448.390 1652.160 448.530 ;
        RECT 1650.640 434.850 1650.780 448.390 ;
        RECT 1649.200 434.530 1649.460 434.850 ;
        RECT 1650.580 434.530 1650.840 434.850 ;
        RECT 1649.260 386.570 1649.400 434.530 ;
        RECT 1649.200 386.250 1649.460 386.570 ;
        RECT 1650.120 386.250 1650.380 386.570 ;
        RECT 1650.180 351.290 1650.320 386.250 ;
        RECT 1650.180 351.150 1650.780 351.290 ;
        RECT 1650.640 331.150 1650.780 351.150 ;
        RECT 1650.120 330.830 1650.380 331.150 ;
        RECT 1650.580 330.830 1650.840 331.150 ;
        RECT 1650.180 283.210 1650.320 330.830 ;
        RECT 1650.120 282.890 1650.380 283.210 ;
        RECT 1651.040 282.890 1651.300 283.210 ;
        RECT 1651.100 255.410 1651.240 282.890 ;
        RECT 1650.640 255.270 1651.240 255.410 ;
        RECT 1650.640 254.730 1650.780 255.270 ;
        RECT 1650.640 254.590 1651.240 254.730 ;
        RECT 1651.100 234.590 1651.240 254.590 ;
        RECT 1649.200 234.270 1649.460 234.590 ;
        RECT 1651.040 234.270 1651.300 234.590 ;
        RECT 1649.260 186.650 1649.400 234.270 ;
        RECT 1649.200 186.330 1649.460 186.650 ;
        RECT 1650.120 186.330 1650.380 186.650 ;
        RECT 1650.180 186.165 1650.320 186.330 ;
        RECT 1650.110 185.795 1650.390 186.165 ;
        RECT 1651.950 185.795 1652.230 186.165 ;
        RECT 1652.020 138.370 1652.160 185.795 ;
        RECT 1650.580 138.050 1650.840 138.370 ;
        RECT 1651.960 138.050 1652.220 138.370 ;
        RECT 1650.640 110.490 1650.780 138.050 ;
        RECT 1650.580 110.170 1650.840 110.490 ;
        RECT 1651.500 110.170 1651.760 110.490 ;
        RECT 1651.560 96.550 1651.700 110.170 ;
        RECT 1650.120 96.230 1650.380 96.550 ;
        RECT 1651.500 96.230 1651.760 96.550 ;
        RECT 1650.180 48.610 1650.320 96.230 ;
        RECT 1650.120 48.290 1650.380 48.610 ;
        RECT 1651.040 48.290 1651.300 48.610 ;
        RECT 1651.100 3.050 1651.240 48.290 ;
        RECT 1650.120 2.730 1650.380 3.050 ;
        RECT 1651.040 2.730 1651.300 3.050 ;
        RECT 1650.180 2.400 1650.320 2.730 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
      LAYER via2 ;
        RECT 1650.110 185.840 1650.390 186.120 ;
        RECT 1651.950 185.840 1652.230 186.120 ;
      LAYER met3 ;
        RECT 1650.085 186.130 1650.415 186.145 ;
        RECT 1651.925 186.130 1652.255 186.145 ;
        RECT 1650.085 185.830 1652.255 186.130 ;
        RECT 1650.085 185.815 1650.415 185.830 ;
        RECT 1651.925 185.815 1652.255 185.830 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1528.190 591.840 1528.510 591.900 ;
        RECT 1528.190 591.700 1546.360 591.840 ;
        RECT 1528.190 591.640 1528.510 591.700 ;
        RECT 1546.220 591.500 1546.360 591.700 ;
        RECT 1663.890 591.500 1664.210 591.560 ;
        RECT 1546.220 591.360 1664.210 591.500 ;
        RECT 1663.890 591.300 1664.210 591.360 ;
        RECT 1663.890 62.120 1664.210 62.180 ;
        RECT 1668.030 62.120 1668.350 62.180 ;
        RECT 1663.890 61.980 1668.350 62.120 ;
        RECT 1663.890 61.920 1664.210 61.980 ;
        RECT 1668.030 61.920 1668.350 61.980 ;
      LAYER via ;
        RECT 1528.220 591.640 1528.480 591.900 ;
        RECT 1663.920 591.300 1664.180 591.560 ;
        RECT 1663.920 61.920 1664.180 62.180 ;
        RECT 1668.060 61.920 1668.320 62.180 ;
      LAYER met2 ;
        RECT 1526.610 600.170 1526.890 604.000 ;
        RECT 1526.610 600.030 1528.420 600.170 ;
        RECT 1526.610 600.000 1526.890 600.030 ;
        RECT 1528.280 591.930 1528.420 600.030 ;
        RECT 1528.220 591.610 1528.480 591.930 ;
        RECT 1663.920 591.270 1664.180 591.590 ;
        RECT 1663.980 62.210 1664.120 591.270 ;
        RECT 1663.920 61.890 1664.180 62.210 ;
        RECT 1668.060 61.890 1668.320 62.210 ;
        RECT 1668.120 2.400 1668.260 61.890 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1537.390 590.820 1537.710 590.880 ;
        RECT 1683.670 590.820 1683.990 590.880 ;
        RECT 1537.390 590.680 1683.990 590.820 ;
        RECT 1537.390 590.620 1537.710 590.680 ;
        RECT 1683.670 590.620 1683.990 590.680 ;
        RECT 1683.670 2.960 1683.990 3.020 ;
        RECT 1685.510 2.960 1685.830 3.020 ;
        RECT 1683.670 2.820 1685.830 2.960 ;
        RECT 1683.670 2.760 1683.990 2.820 ;
        RECT 1685.510 2.760 1685.830 2.820 ;
      LAYER via ;
        RECT 1537.420 590.620 1537.680 590.880 ;
        RECT 1683.700 590.620 1683.960 590.880 ;
        RECT 1683.700 2.760 1683.960 3.020 ;
        RECT 1685.540 2.760 1685.800 3.020 ;
      LAYER met2 ;
        RECT 1535.810 600.170 1536.090 604.000 ;
        RECT 1535.810 600.030 1537.620 600.170 ;
        RECT 1535.810 600.000 1536.090 600.030 ;
        RECT 1537.480 590.910 1537.620 600.030 ;
        RECT 1537.420 590.590 1537.680 590.910 ;
        RECT 1683.700 590.590 1683.960 590.910 ;
        RECT 1683.760 3.050 1683.900 590.590 ;
        RECT 1683.700 2.730 1683.960 3.050 ;
        RECT 1685.540 2.730 1685.800 3.050 ;
        RECT 1685.600 2.400 1685.740 2.730 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1035.530 569.400 1035.850 569.460 ;
        RECT 1039.210 569.400 1039.530 569.460 ;
        RECT 1035.530 569.260 1039.530 569.400 ;
        RECT 1035.530 569.200 1035.850 569.260 ;
        RECT 1039.210 569.200 1039.530 569.260 ;
        RECT 722.270 38.660 722.590 38.720 ;
        RECT 1035.530 38.660 1035.850 38.720 ;
        RECT 722.270 38.520 1035.850 38.660 ;
        RECT 722.270 38.460 722.590 38.520 ;
        RECT 1035.530 38.460 1035.850 38.520 ;
      LAYER via ;
        RECT 1035.560 569.200 1035.820 569.460 ;
        RECT 1039.240 569.200 1039.500 569.460 ;
        RECT 722.300 38.460 722.560 38.720 ;
        RECT 1035.560 38.460 1035.820 38.720 ;
      LAYER met2 ;
        RECT 1040.850 600.170 1041.130 604.000 ;
        RECT 1039.300 600.030 1041.130 600.170 ;
        RECT 1039.300 569.490 1039.440 600.030 ;
        RECT 1040.850 600.000 1041.130 600.030 ;
        RECT 1035.560 569.170 1035.820 569.490 ;
        RECT 1039.240 569.170 1039.500 569.490 ;
        RECT 1035.620 38.750 1035.760 569.170 ;
        RECT 722.300 38.430 722.560 38.750 ;
        RECT 1035.560 38.430 1035.820 38.750 ;
        RECT 722.360 2.400 722.500 38.430 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.670 590.480 1545.990 590.540 ;
        RECT 1697.930 590.480 1698.250 590.540 ;
        RECT 1545.670 590.340 1698.250 590.480 ;
        RECT 1545.670 590.280 1545.990 590.340 ;
        RECT 1697.930 590.280 1698.250 590.340 ;
        RECT 1697.930 2.960 1698.250 3.020 ;
        RECT 1703.450 2.960 1703.770 3.020 ;
        RECT 1697.930 2.820 1703.770 2.960 ;
        RECT 1697.930 2.760 1698.250 2.820 ;
        RECT 1703.450 2.760 1703.770 2.820 ;
      LAYER via ;
        RECT 1545.700 590.280 1545.960 590.540 ;
        RECT 1697.960 590.280 1698.220 590.540 ;
        RECT 1697.960 2.760 1698.220 3.020 ;
        RECT 1703.480 2.760 1703.740 3.020 ;
      LAYER met2 ;
        RECT 1545.010 600.000 1545.290 604.000 ;
        RECT 1545.070 598.810 1545.210 600.000 ;
        RECT 1545.070 598.670 1545.440 598.810 ;
        RECT 1545.300 591.330 1545.440 598.670 ;
        RECT 1545.300 591.190 1545.900 591.330 ;
        RECT 1545.760 590.570 1545.900 591.190 ;
        RECT 1545.700 590.250 1545.960 590.570 ;
        RECT 1697.960 590.250 1698.220 590.570 ;
        RECT 1698.020 3.050 1698.160 590.250 ;
        RECT 1697.960 2.730 1698.220 3.050 ;
        RECT 1703.480 2.730 1703.740 3.050 ;
        RECT 1703.540 2.400 1703.680 2.730 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1555.790 591.840 1556.110 591.900 ;
        RECT 1606.850 591.840 1607.170 591.900 ;
        RECT 1555.790 591.700 1607.170 591.840 ;
        RECT 1555.790 591.640 1556.110 591.700 ;
        RECT 1606.850 591.640 1607.170 591.700 ;
        RECT 1698.390 590.480 1698.710 590.540 ;
        RECT 1718.630 590.480 1718.950 590.540 ;
        RECT 1698.390 590.340 1718.950 590.480 ;
        RECT 1698.390 590.280 1698.710 590.340 ;
        RECT 1718.630 590.280 1718.950 590.340 ;
        RECT 1606.850 590.140 1607.170 590.200 ;
        RECT 1655.150 590.140 1655.470 590.200 ;
        RECT 1606.850 590.000 1655.470 590.140 ;
        RECT 1606.850 589.940 1607.170 590.000 ;
        RECT 1655.150 589.940 1655.470 590.000 ;
        RECT 1698.390 589.460 1698.710 589.520 ;
        RECT 1657.540 589.320 1698.710 589.460 ;
        RECT 1655.150 588.780 1655.470 588.840 ;
        RECT 1657.540 588.780 1657.680 589.320 ;
        RECT 1698.390 589.260 1698.710 589.320 ;
        RECT 1655.150 588.640 1657.680 588.780 ;
        RECT 1655.150 588.580 1655.470 588.640 ;
        RECT 1719.090 2.960 1719.410 3.020 ;
        RECT 1721.390 2.960 1721.710 3.020 ;
        RECT 1719.090 2.820 1721.710 2.960 ;
        RECT 1719.090 2.760 1719.410 2.820 ;
        RECT 1721.390 2.760 1721.710 2.820 ;
      LAYER via ;
        RECT 1555.820 591.640 1556.080 591.900 ;
        RECT 1606.880 591.640 1607.140 591.900 ;
        RECT 1698.420 590.280 1698.680 590.540 ;
        RECT 1718.660 590.280 1718.920 590.540 ;
        RECT 1606.880 589.940 1607.140 590.200 ;
        RECT 1655.180 589.940 1655.440 590.200 ;
        RECT 1655.180 588.580 1655.440 588.840 ;
        RECT 1698.420 589.260 1698.680 589.520 ;
        RECT 1719.120 2.760 1719.380 3.020 ;
        RECT 1721.420 2.760 1721.680 3.020 ;
      LAYER met2 ;
        RECT 1554.210 600.170 1554.490 604.000 ;
        RECT 1554.210 600.030 1556.020 600.170 ;
        RECT 1554.210 600.000 1554.490 600.030 ;
        RECT 1555.880 591.930 1556.020 600.030 ;
        RECT 1555.820 591.610 1556.080 591.930 ;
        RECT 1606.880 591.610 1607.140 591.930 ;
        RECT 1606.940 590.230 1607.080 591.610 ;
        RECT 1718.720 590.570 1719.320 590.650 ;
        RECT 1698.420 590.250 1698.680 590.570 ;
        RECT 1718.660 590.510 1719.320 590.570 ;
        RECT 1718.660 590.250 1718.920 590.510 ;
        RECT 1606.880 589.910 1607.140 590.230 ;
        RECT 1655.180 589.910 1655.440 590.230 ;
        RECT 1655.240 588.870 1655.380 589.910 ;
        RECT 1698.480 589.550 1698.620 590.250 ;
        RECT 1698.420 589.230 1698.680 589.550 ;
        RECT 1655.180 588.550 1655.440 588.870 ;
        RECT 1719.180 3.050 1719.320 590.510 ;
        RECT 1719.120 2.730 1719.380 3.050 ;
        RECT 1721.420 2.730 1721.680 3.050 ;
        RECT 1721.480 2.400 1721.620 2.730 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1739.790 590.480 1740.110 590.540 ;
        RECT 1719.180 590.340 1740.110 590.480 ;
        RECT 1719.180 589.800 1719.320 590.340 ;
        RECT 1739.790 590.280 1740.110 590.340 ;
        RECT 1581.180 589.660 1655.380 589.800 ;
        RECT 1564.990 589.120 1565.310 589.180 ;
        RECT 1581.180 589.120 1581.320 589.660 ;
        RECT 1564.990 588.980 1581.320 589.120 ;
        RECT 1655.240 589.120 1655.380 589.660 ;
        RECT 1657.080 589.660 1719.320 589.800 ;
        RECT 1657.080 589.120 1657.220 589.660 ;
        RECT 1655.240 588.980 1657.220 589.120 ;
        RECT 1564.990 588.920 1565.310 588.980 ;
      LAYER via ;
        RECT 1739.820 590.280 1740.080 590.540 ;
        RECT 1565.020 588.920 1565.280 589.180 ;
      LAYER met2 ;
        RECT 1563.410 600.170 1563.690 604.000 ;
        RECT 1563.410 600.030 1565.220 600.170 ;
        RECT 1563.410 600.000 1563.690 600.030 ;
        RECT 1565.080 589.210 1565.220 600.030 ;
        RECT 1739.820 590.250 1740.080 590.570 ;
        RECT 1565.020 588.890 1565.280 589.210 ;
        RECT 1739.880 3.130 1740.020 590.250 ;
        RECT 1739.420 2.990 1740.020 3.130 ;
        RECT 1739.420 2.400 1739.560 2.990 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.350 32.880 1572.670 32.940 ;
        RECT 1755.430 32.880 1755.750 32.940 ;
        RECT 1572.350 32.740 1755.750 32.880 ;
        RECT 1572.350 32.680 1572.670 32.740 ;
        RECT 1755.430 32.680 1755.750 32.740 ;
      LAYER via ;
        RECT 1572.380 32.680 1572.640 32.940 ;
        RECT 1755.460 32.680 1755.720 32.940 ;
      LAYER met2 ;
        RECT 1572.610 600.000 1572.890 604.000 ;
        RECT 1572.670 598.810 1572.810 600.000 ;
        RECT 1572.440 598.670 1572.810 598.810 ;
        RECT 1572.440 32.970 1572.580 598.670 ;
        RECT 1572.380 32.650 1572.640 32.970 ;
        RECT 1755.460 32.650 1755.720 32.970 ;
        RECT 1755.520 32.370 1755.660 32.650 ;
        RECT 1755.520 32.230 1757.040 32.370 ;
        RECT 1756.900 2.400 1757.040 32.230 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1583.390 586.740 1583.710 586.800 ;
        RECT 1586.610 586.740 1586.930 586.800 ;
        RECT 1583.390 586.600 1586.930 586.740 ;
        RECT 1583.390 586.540 1583.710 586.600 ;
        RECT 1586.610 586.540 1586.930 586.600 ;
        RECT 1586.610 29.480 1586.930 29.540 ;
        RECT 1774.750 29.480 1775.070 29.540 ;
        RECT 1586.610 29.340 1775.070 29.480 ;
        RECT 1586.610 29.280 1586.930 29.340 ;
        RECT 1774.750 29.280 1775.070 29.340 ;
      LAYER via ;
        RECT 1583.420 586.540 1583.680 586.800 ;
        RECT 1586.640 586.540 1586.900 586.800 ;
        RECT 1586.640 29.280 1586.900 29.540 ;
        RECT 1774.780 29.280 1775.040 29.540 ;
      LAYER met2 ;
        RECT 1581.810 600.170 1582.090 604.000 ;
        RECT 1581.810 600.030 1583.620 600.170 ;
        RECT 1581.810 600.000 1582.090 600.030 ;
        RECT 1583.480 586.830 1583.620 600.030 ;
        RECT 1583.420 586.510 1583.680 586.830 ;
        RECT 1586.640 586.510 1586.900 586.830 ;
        RECT 1586.700 29.570 1586.840 586.510 ;
        RECT 1586.640 29.250 1586.900 29.570 ;
        RECT 1774.780 29.250 1775.040 29.570 ;
        RECT 1774.840 2.400 1774.980 29.250 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1592.130 524.180 1592.450 524.240 ;
        RECT 1592.590 524.180 1592.910 524.240 ;
        RECT 1592.130 524.040 1592.910 524.180 ;
        RECT 1592.130 523.980 1592.450 524.040 ;
        RECT 1592.590 523.980 1592.910 524.040 ;
        RECT 1592.130 476.240 1592.450 476.300 ;
        RECT 1593.510 476.240 1593.830 476.300 ;
        RECT 1592.130 476.100 1593.830 476.240 ;
        RECT 1592.130 476.040 1592.450 476.100 ;
        RECT 1593.510 476.040 1593.830 476.100 ;
        RECT 1592.130 366.080 1592.450 366.140 ;
        RECT 1592.590 366.080 1592.910 366.140 ;
        RECT 1592.130 365.940 1592.910 366.080 ;
        RECT 1592.130 365.880 1592.450 365.940 ;
        RECT 1592.590 365.880 1592.910 365.940 ;
        RECT 1592.130 290.260 1592.450 290.320 ;
        RECT 1592.590 290.260 1592.910 290.320 ;
        RECT 1592.130 290.120 1592.910 290.260 ;
        RECT 1592.130 290.060 1592.450 290.120 ;
        RECT 1592.590 290.060 1592.910 290.120 ;
        RECT 1592.130 289.580 1592.450 289.640 ;
        RECT 1592.590 289.580 1592.910 289.640 ;
        RECT 1592.130 289.440 1592.910 289.580 ;
        RECT 1592.130 289.380 1592.450 289.440 ;
        RECT 1592.590 289.380 1592.910 289.440 ;
        RECT 1592.130 241.640 1592.450 241.700 ;
        RECT 1593.050 241.640 1593.370 241.700 ;
        RECT 1592.130 241.500 1593.370 241.640 ;
        RECT 1592.130 241.440 1592.450 241.500 ;
        RECT 1593.050 241.440 1593.370 241.500 ;
        RECT 1591.670 234.500 1591.990 234.560 ;
        RECT 1593.050 234.500 1593.370 234.560 ;
        RECT 1591.670 234.360 1593.370 234.500 ;
        RECT 1591.670 234.300 1591.990 234.360 ;
        RECT 1593.050 234.300 1593.370 234.360 ;
        RECT 1591.670 186.560 1591.990 186.620 ;
        RECT 1592.590 186.560 1592.910 186.620 ;
        RECT 1591.670 186.420 1592.910 186.560 ;
        RECT 1591.670 186.360 1591.990 186.420 ;
        RECT 1592.590 186.360 1592.910 186.420 ;
        RECT 1593.510 111.420 1593.830 111.480 ;
        RECT 1593.140 111.280 1593.830 111.420 ;
        RECT 1593.140 111.140 1593.280 111.280 ;
        RECT 1593.510 111.220 1593.830 111.280 ;
        RECT 1593.050 110.880 1593.370 111.140 ;
        RECT 1591.670 96.460 1591.990 96.520 ;
        RECT 1592.590 96.460 1592.910 96.520 ;
        RECT 1591.670 96.320 1592.910 96.460 ;
        RECT 1591.670 96.260 1591.990 96.320 ;
        RECT 1592.590 96.260 1592.910 96.320 ;
        RECT 1591.670 48.520 1591.990 48.580 ;
        RECT 1593.050 48.520 1593.370 48.580 ;
        RECT 1591.670 48.380 1593.370 48.520 ;
        RECT 1591.670 48.320 1591.990 48.380 ;
        RECT 1593.050 48.320 1593.370 48.380 ;
        RECT 1593.050 29.820 1593.370 29.880 ;
        RECT 1792.690 29.820 1793.010 29.880 ;
        RECT 1593.050 29.680 1793.010 29.820 ;
        RECT 1593.050 29.620 1593.370 29.680 ;
        RECT 1792.690 29.620 1793.010 29.680 ;
      LAYER via ;
        RECT 1592.160 523.980 1592.420 524.240 ;
        RECT 1592.620 523.980 1592.880 524.240 ;
        RECT 1592.160 476.040 1592.420 476.300 ;
        RECT 1593.540 476.040 1593.800 476.300 ;
        RECT 1592.160 365.880 1592.420 366.140 ;
        RECT 1592.620 365.880 1592.880 366.140 ;
        RECT 1592.160 290.060 1592.420 290.320 ;
        RECT 1592.620 290.060 1592.880 290.320 ;
        RECT 1592.160 289.380 1592.420 289.640 ;
        RECT 1592.620 289.380 1592.880 289.640 ;
        RECT 1592.160 241.440 1592.420 241.700 ;
        RECT 1593.080 241.440 1593.340 241.700 ;
        RECT 1591.700 234.300 1591.960 234.560 ;
        RECT 1593.080 234.300 1593.340 234.560 ;
        RECT 1591.700 186.360 1591.960 186.620 ;
        RECT 1592.620 186.360 1592.880 186.620 ;
        RECT 1593.540 111.220 1593.800 111.480 ;
        RECT 1593.080 110.880 1593.340 111.140 ;
        RECT 1591.700 96.260 1591.960 96.520 ;
        RECT 1592.620 96.260 1592.880 96.520 ;
        RECT 1591.700 48.320 1591.960 48.580 ;
        RECT 1593.080 48.320 1593.340 48.580 ;
        RECT 1593.080 29.620 1593.340 29.880 ;
        RECT 1792.720 29.620 1792.980 29.880 ;
      LAYER met2 ;
        RECT 1591.010 600.000 1591.290 604.000 ;
        RECT 1591.070 598.810 1591.210 600.000 ;
        RECT 1591.070 598.670 1591.440 598.810 ;
        RECT 1591.300 580.565 1591.440 598.670 ;
        RECT 1591.230 580.195 1591.510 580.565 ;
        RECT 1593.070 579.515 1593.350 579.885 ;
        RECT 1593.140 532.285 1593.280 579.515 ;
        RECT 1593.070 531.915 1593.350 532.285 ;
        RECT 1592.610 531.235 1592.890 531.605 ;
        RECT 1592.680 524.270 1592.820 531.235 ;
        RECT 1592.160 523.950 1592.420 524.270 ;
        RECT 1592.620 523.950 1592.880 524.270 ;
        RECT 1592.220 476.330 1592.360 523.950 ;
        RECT 1592.160 476.010 1592.420 476.330 ;
        RECT 1593.540 476.010 1593.800 476.330 ;
        RECT 1593.600 445.130 1593.740 476.010 ;
        RECT 1592.680 444.990 1593.740 445.130 ;
        RECT 1592.680 366.170 1592.820 444.990 ;
        RECT 1592.160 365.850 1592.420 366.170 ;
        RECT 1592.620 365.850 1592.880 366.170 ;
        RECT 1592.220 290.350 1592.360 365.850 ;
        RECT 1592.160 290.030 1592.420 290.350 ;
        RECT 1592.620 290.030 1592.880 290.350 ;
        RECT 1592.680 289.670 1592.820 290.030 ;
        RECT 1592.160 289.350 1592.420 289.670 ;
        RECT 1592.620 289.350 1592.880 289.670 ;
        RECT 1592.220 241.730 1592.360 289.350 ;
        RECT 1592.160 241.410 1592.420 241.730 ;
        RECT 1593.080 241.410 1593.340 241.730 ;
        RECT 1593.140 234.590 1593.280 241.410 ;
        RECT 1591.700 234.270 1591.960 234.590 ;
        RECT 1593.080 234.270 1593.340 234.590 ;
        RECT 1591.760 186.650 1591.900 234.270 ;
        RECT 1591.700 186.330 1591.960 186.650 ;
        RECT 1592.620 186.330 1592.880 186.650 ;
        RECT 1592.680 169.730 1592.820 186.330 ;
        RECT 1592.680 169.590 1593.280 169.730 ;
        RECT 1593.140 144.570 1593.280 169.590 ;
        RECT 1593.140 144.430 1593.740 144.570 ;
        RECT 1593.600 111.510 1593.740 144.430 ;
        RECT 1593.540 111.190 1593.800 111.510 ;
        RECT 1593.080 110.850 1593.340 111.170 ;
        RECT 1593.140 96.970 1593.280 110.850 ;
        RECT 1592.680 96.830 1593.280 96.970 ;
        RECT 1592.680 96.550 1592.820 96.830 ;
        RECT 1591.700 96.230 1591.960 96.550 ;
        RECT 1592.620 96.230 1592.880 96.550 ;
        RECT 1591.760 48.610 1591.900 96.230 ;
        RECT 1591.700 48.290 1591.960 48.610 ;
        RECT 1593.080 48.290 1593.340 48.610 ;
        RECT 1593.140 29.910 1593.280 48.290 ;
        RECT 1593.080 29.590 1593.340 29.910 ;
        RECT 1792.720 29.590 1792.980 29.910 ;
        RECT 1792.780 2.400 1792.920 29.590 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
      LAYER via2 ;
        RECT 1591.230 580.240 1591.510 580.520 ;
        RECT 1593.070 579.560 1593.350 579.840 ;
        RECT 1593.070 531.960 1593.350 532.240 ;
        RECT 1592.610 531.280 1592.890 531.560 ;
      LAYER met3 ;
        RECT 1591.205 580.530 1591.535 580.545 ;
        RECT 1591.205 580.230 1593.130 580.530 ;
        RECT 1591.205 580.215 1591.535 580.230 ;
        RECT 1592.830 579.865 1593.130 580.230 ;
        RECT 1592.830 579.550 1593.375 579.865 ;
        RECT 1593.045 579.535 1593.375 579.550 ;
        RECT 1593.045 532.250 1593.375 532.265 ;
        RECT 1591.910 531.950 1593.375 532.250 ;
        RECT 1591.910 531.570 1592.210 531.950 ;
        RECT 1593.045 531.935 1593.375 531.950 ;
        RECT 1592.585 531.570 1592.915 531.585 ;
        RECT 1591.910 531.270 1592.915 531.570 ;
        RECT 1592.585 531.255 1592.915 531.270 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1599.950 34.240 1600.270 34.300 ;
        RECT 1810.630 34.240 1810.950 34.300 ;
        RECT 1599.950 34.100 1810.950 34.240 ;
        RECT 1599.950 34.040 1600.270 34.100 ;
        RECT 1810.630 34.040 1810.950 34.100 ;
      LAYER via ;
        RECT 1599.980 34.040 1600.240 34.300 ;
        RECT 1810.660 34.040 1810.920 34.300 ;
      LAYER met2 ;
        RECT 1600.210 600.000 1600.490 604.000 ;
        RECT 1600.270 598.810 1600.410 600.000 ;
        RECT 1600.040 598.670 1600.410 598.810 ;
        RECT 1600.040 34.330 1600.180 598.670 ;
        RECT 1599.980 34.010 1600.240 34.330 ;
        RECT 1810.660 34.010 1810.920 34.330 ;
        RECT 1810.720 2.400 1810.860 34.010 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1610.530 586.740 1610.850 586.800 ;
        RECT 1614.210 586.740 1614.530 586.800 ;
        RECT 1610.530 586.600 1614.530 586.740 ;
        RECT 1610.530 586.540 1610.850 586.600 ;
        RECT 1614.210 586.540 1614.530 586.600 ;
        RECT 1613.290 41.720 1613.610 41.780 ;
        RECT 1614.210 41.720 1614.530 41.780 ;
        RECT 1613.290 41.580 1614.530 41.720 ;
        RECT 1613.290 41.520 1613.610 41.580 ;
        RECT 1614.210 41.520 1614.530 41.580 ;
        RECT 1613.290 21.320 1613.610 21.380 ;
        RECT 1828.570 21.320 1828.890 21.380 ;
        RECT 1613.290 21.180 1828.890 21.320 ;
        RECT 1613.290 21.120 1613.610 21.180 ;
        RECT 1828.570 21.120 1828.890 21.180 ;
      LAYER via ;
        RECT 1610.560 586.540 1610.820 586.800 ;
        RECT 1614.240 586.540 1614.500 586.800 ;
        RECT 1613.320 41.520 1613.580 41.780 ;
        RECT 1614.240 41.520 1614.500 41.780 ;
        RECT 1613.320 21.120 1613.580 21.380 ;
        RECT 1828.600 21.120 1828.860 21.380 ;
      LAYER met2 ;
        RECT 1608.950 600.170 1609.230 604.000 ;
        RECT 1608.950 600.030 1610.760 600.170 ;
        RECT 1608.950 600.000 1609.230 600.030 ;
        RECT 1610.620 586.830 1610.760 600.030 ;
        RECT 1610.560 586.510 1610.820 586.830 ;
        RECT 1614.240 586.510 1614.500 586.830 ;
        RECT 1614.300 41.810 1614.440 586.510 ;
        RECT 1613.320 41.490 1613.580 41.810 ;
        RECT 1614.240 41.490 1614.500 41.810 ;
        RECT 1613.380 21.410 1613.520 41.490 ;
        RECT 1613.320 21.090 1613.580 21.410 ;
        RECT 1828.600 21.090 1828.860 21.410 ;
        RECT 1828.660 2.400 1828.800 21.090 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1619.270 579.600 1619.590 579.660 ;
        RECT 1620.650 579.600 1620.970 579.660 ;
        RECT 1619.270 579.460 1620.970 579.600 ;
        RECT 1619.270 579.400 1619.590 579.460 ;
        RECT 1620.650 579.400 1620.970 579.460 ;
        RECT 1620.650 531.320 1620.970 531.380 ;
        RECT 1621.110 531.320 1621.430 531.380 ;
        RECT 1620.650 531.180 1621.430 531.320 ;
        RECT 1620.650 531.120 1620.970 531.180 ;
        RECT 1621.110 531.120 1621.430 531.180 ;
        RECT 1621.110 496.980 1621.430 497.040 ;
        RECT 1620.740 496.840 1621.430 496.980 ;
        RECT 1620.740 496.700 1620.880 496.840 ;
        RECT 1621.110 496.780 1621.430 496.840 ;
        RECT 1620.650 496.440 1620.970 496.700 ;
        RECT 1619.730 462.300 1620.050 462.360 ;
        RECT 1621.110 462.300 1621.430 462.360 ;
        RECT 1619.730 462.160 1621.430 462.300 ;
        RECT 1619.730 462.100 1620.050 462.160 ;
        RECT 1621.110 462.100 1621.430 462.160 ;
        RECT 1619.270 414.360 1619.590 414.420 ;
        RECT 1619.730 414.360 1620.050 414.420 ;
        RECT 1619.270 414.220 1620.050 414.360 ;
        RECT 1619.270 414.160 1619.590 414.220 ;
        RECT 1619.730 414.160 1620.050 414.220 ;
        RECT 1621.570 283.120 1621.890 283.180 ;
        RECT 1622.490 283.120 1622.810 283.180 ;
        RECT 1621.570 282.980 1622.810 283.120 ;
        RECT 1621.570 282.920 1621.890 282.980 ;
        RECT 1622.490 282.920 1622.810 282.980 ;
        RECT 1620.650 234.500 1620.970 234.560 ;
        RECT 1621.570 234.500 1621.890 234.560 ;
        RECT 1620.650 234.360 1621.890 234.500 ;
        RECT 1620.650 234.300 1620.970 234.360 ;
        RECT 1621.570 234.300 1621.890 234.360 ;
        RECT 1620.650 186.560 1620.970 186.620 ;
        RECT 1621.570 186.560 1621.890 186.620 ;
        RECT 1620.650 186.420 1621.890 186.560 ;
        RECT 1620.650 186.360 1620.970 186.420 ;
        RECT 1621.570 186.360 1621.890 186.420 ;
        RECT 1620.190 90.000 1620.510 90.060 ;
        RECT 1620.650 90.000 1620.970 90.060 ;
        RECT 1620.190 89.860 1620.970 90.000 ;
        RECT 1620.190 89.800 1620.510 89.860 ;
        RECT 1620.650 89.800 1620.970 89.860 ;
        RECT 1620.190 62.120 1620.510 62.180 ;
        RECT 1621.110 62.120 1621.430 62.180 ;
        RECT 1620.190 61.980 1621.430 62.120 ;
        RECT 1620.190 61.920 1620.510 61.980 ;
        RECT 1621.110 61.920 1621.430 61.980 ;
        RECT 1621.110 21.660 1621.430 21.720 ;
        RECT 1846.050 21.660 1846.370 21.720 ;
        RECT 1621.110 21.520 1846.370 21.660 ;
        RECT 1621.110 21.460 1621.430 21.520 ;
        RECT 1846.050 21.460 1846.370 21.520 ;
      LAYER via ;
        RECT 1619.300 579.400 1619.560 579.660 ;
        RECT 1620.680 579.400 1620.940 579.660 ;
        RECT 1620.680 531.120 1620.940 531.380 ;
        RECT 1621.140 531.120 1621.400 531.380 ;
        RECT 1621.140 496.780 1621.400 497.040 ;
        RECT 1620.680 496.440 1620.940 496.700 ;
        RECT 1619.760 462.100 1620.020 462.360 ;
        RECT 1621.140 462.100 1621.400 462.360 ;
        RECT 1619.300 414.160 1619.560 414.420 ;
        RECT 1619.760 414.160 1620.020 414.420 ;
        RECT 1621.600 282.920 1621.860 283.180 ;
        RECT 1622.520 282.920 1622.780 283.180 ;
        RECT 1620.680 234.300 1620.940 234.560 ;
        RECT 1621.600 234.300 1621.860 234.560 ;
        RECT 1620.680 186.360 1620.940 186.620 ;
        RECT 1621.600 186.360 1621.860 186.620 ;
        RECT 1620.220 89.800 1620.480 90.060 ;
        RECT 1620.680 89.800 1620.940 90.060 ;
        RECT 1620.220 61.920 1620.480 62.180 ;
        RECT 1621.140 61.920 1621.400 62.180 ;
        RECT 1621.140 21.460 1621.400 21.720 ;
        RECT 1846.080 21.460 1846.340 21.720 ;
      LAYER met2 ;
        RECT 1618.150 600.850 1618.430 604.000 ;
        RECT 1618.150 600.710 1619.500 600.850 ;
        RECT 1618.150 600.000 1618.430 600.710 ;
        RECT 1619.360 579.690 1619.500 600.710 ;
        RECT 1619.300 579.370 1619.560 579.690 ;
        RECT 1620.680 579.370 1620.940 579.690 ;
        RECT 1620.740 531.410 1620.880 579.370 ;
        RECT 1620.680 531.090 1620.940 531.410 ;
        RECT 1621.140 531.090 1621.400 531.410 ;
        RECT 1621.200 497.070 1621.340 531.090 ;
        RECT 1621.140 496.750 1621.400 497.070 ;
        RECT 1620.680 496.410 1620.940 496.730 ;
        RECT 1620.740 483.210 1620.880 496.410 ;
        RECT 1620.740 483.070 1621.340 483.210 ;
        RECT 1621.200 462.390 1621.340 483.070 ;
        RECT 1619.760 462.070 1620.020 462.390 ;
        RECT 1621.140 462.070 1621.400 462.390 ;
        RECT 1619.820 414.450 1619.960 462.070 ;
        RECT 1619.300 414.130 1619.560 414.450 ;
        RECT 1619.760 414.130 1620.020 414.450 ;
        RECT 1619.360 413.965 1619.500 414.130 ;
        RECT 1619.290 413.595 1619.570 413.965 ;
        RECT 1619.290 412.915 1619.570 413.285 ;
        RECT 1619.360 371.805 1619.500 412.915 ;
        RECT 1619.290 371.435 1619.570 371.805 ;
        RECT 1622.510 371.435 1622.790 371.805 ;
        RECT 1622.580 283.210 1622.720 371.435 ;
        RECT 1621.600 282.890 1621.860 283.210 ;
        RECT 1622.520 282.890 1622.780 283.210 ;
        RECT 1621.660 241.640 1621.800 282.890 ;
        RECT 1620.740 241.500 1621.800 241.640 ;
        RECT 1620.740 234.590 1620.880 241.500 ;
        RECT 1620.680 234.270 1620.940 234.590 ;
        RECT 1621.600 234.270 1621.860 234.590 ;
        RECT 1621.660 186.650 1621.800 234.270 ;
        RECT 1620.680 186.330 1620.940 186.650 ;
        RECT 1621.600 186.330 1621.860 186.650 ;
        RECT 1620.740 90.090 1620.880 186.330 ;
        RECT 1620.220 89.770 1620.480 90.090 ;
        RECT 1620.680 89.770 1620.940 90.090 ;
        RECT 1620.280 62.210 1620.420 89.770 ;
        RECT 1620.220 61.890 1620.480 62.210 ;
        RECT 1621.140 61.890 1621.400 62.210 ;
        RECT 1621.200 21.750 1621.340 61.890 ;
        RECT 1621.140 21.430 1621.400 21.750 ;
        RECT 1846.080 21.430 1846.340 21.750 ;
        RECT 1846.140 2.400 1846.280 21.430 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
      LAYER via2 ;
        RECT 1619.290 413.640 1619.570 413.920 ;
        RECT 1619.290 412.960 1619.570 413.240 ;
        RECT 1619.290 371.480 1619.570 371.760 ;
        RECT 1622.510 371.480 1622.790 371.760 ;
      LAYER met3 ;
        RECT 1619.265 413.615 1619.595 413.945 ;
        RECT 1619.280 413.265 1619.580 413.615 ;
        RECT 1619.265 412.935 1619.595 413.265 ;
        RECT 1619.265 371.770 1619.595 371.785 ;
        RECT 1622.485 371.770 1622.815 371.785 ;
        RECT 1619.265 371.470 1622.815 371.770 ;
        RECT 1619.265 371.455 1619.595 371.470 ;
        RECT 1622.485 371.455 1622.815 371.470 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1627.550 22.340 1627.870 22.400 ;
        RECT 1863.990 22.340 1864.310 22.400 ;
        RECT 1627.550 22.200 1864.310 22.340 ;
        RECT 1627.550 22.140 1627.870 22.200 ;
        RECT 1863.990 22.140 1864.310 22.200 ;
      LAYER via ;
        RECT 1627.580 22.140 1627.840 22.400 ;
        RECT 1864.020 22.140 1864.280 22.400 ;
      LAYER met2 ;
        RECT 1627.350 600.000 1627.630 604.000 ;
        RECT 1627.410 598.810 1627.550 600.000 ;
        RECT 1627.410 598.670 1627.780 598.810 ;
        RECT 1627.640 22.430 1627.780 598.670 ;
        RECT 1627.580 22.110 1627.840 22.430 ;
        RECT 1864.020 22.110 1864.280 22.430 ;
        RECT 1864.080 2.400 1864.220 22.110 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 955.490 588.780 955.810 588.840 ;
        RECT 1049.330 588.780 1049.650 588.840 ;
        RECT 955.490 588.640 1049.650 588.780 ;
        RECT 955.490 588.580 955.810 588.640 ;
        RECT 1049.330 588.580 1049.650 588.640 ;
        RECT 876.370 20.640 876.690 20.700 ;
        RECT 889.250 20.640 889.570 20.700 ;
        RECT 876.370 20.500 889.570 20.640 ;
        RECT 876.370 20.440 876.690 20.500 ;
        RECT 889.250 20.440 889.570 20.500 ;
        RECT 811.050 20.300 811.370 20.360 ;
        RECT 799.180 20.160 811.370 20.300 ;
        RECT 740.210 19.620 740.530 19.680 ;
        RECT 799.180 19.620 799.320 20.160 ;
        RECT 811.050 20.100 811.370 20.160 ;
        RECT 740.210 19.480 799.320 19.620 ;
        RECT 740.210 19.420 740.530 19.480 ;
        RECT 811.050 18.940 811.370 19.000 ;
        RECT 876.370 18.940 876.690 19.000 ;
        RECT 811.050 18.800 876.690 18.940 ;
        RECT 811.050 18.740 811.370 18.800 ;
        RECT 876.370 18.740 876.690 18.800 ;
        RECT 889.250 16.900 889.570 16.960 ;
        RECT 889.250 16.760 943.760 16.900 ;
        RECT 889.250 16.700 889.570 16.760 ;
        RECT 943.620 16.560 943.760 16.760 ;
        RECT 955.490 16.560 955.810 16.620 ;
        RECT 943.620 16.420 955.810 16.560 ;
        RECT 955.490 16.360 955.810 16.420 ;
      LAYER via ;
        RECT 955.520 588.580 955.780 588.840 ;
        RECT 1049.360 588.580 1049.620 588.840 ;
        RECT 876.400 20.440 876.660 20.700 ;
        RECT 889.280 20.440 889.540 20.700 ;
        RECT 740.240 19.420 740.500 19.680 ;
        RECT 811.080 20.100 811.340 20.360 ;
        RECT 811.080 18.740 811.340 19.000 ;
        RECT 876.400 18.740 876.660 19.000 ;
        RECT 889.280 16.700 889.540 16.960 ;
        RECT 955.520 16.360 955.780 16.620 ;
      LAYER met2 ;
        RECT 1050.050 600.170 1050.330 604.000 ;
        RECT 1049.420 600.030 1050.330 600.170 ;
        RECT 1049.420 588.870 1049.560 600.030 ;
        RECT 1050.050 600.000 1050.330 600.030 ;
        RECT 955.520 588.550 955.780 588.870 ;
        RECT 1049.360 588.550 1049.620 588.870 ;
        RECT 876.400 20.410 876.660 20.730 ;
        RECT 889.280 20.410 889.540 20.730 ;
        RECT 811.080 20.070 811.340 20.390 ;
        RECT 740.240 19.390 740.500 19.710 ;
        RECT 740.300 2.400 740.440 19.390 ;
        RECT 811.140 19.030 811.280 20.070 ;
        RECT 876.460 19.030 876.600 20.410 ;
        RECT 811.080 18.710 811.340 19.030 ;
        RECT 876.400 18.710 876.660 19.030 ;
        RECT 889.340 16.990 889.480 20.410 ;
        RECT 889.280 16.670 889.540 16.990 ;
        RECT 955.580 16.650 955.720 588.550 ;
        RECT 955.520 16.330 955.780 16.650 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1638.130 586.740 1638.450 586.800 ;
        RECT 1641.810 586.740 1642.130 586.800 ;
        RECT 1638.130 586.600 1642.130 586.740 ;
        RECT 1638.130 586.540 1638.450 586.600 ;
        RECT 1641.810 586.540 1642.130 586.600 ;
        RECT 1641.810 22.000 1642.130 22.060 ;
        RECT 1881.930 22.000 1882.250 22.060 ;
        RECT 1641.810 21.860 1882.250 22.000 ;
        RECT 1641.810 21.800 1642.130 21.860 ;
        RECT 1881.930 21.800 1882.250 21.860 ;
      LAYER via ;
        RECT 1638.160 586.540 1638.420 586.800 ;
        RECT 1641.840 586.540 1642.100 586.800 ;
        RECT 1641.840 21.800 1642.100 22.060 ;
        RECT 1881.960 21.800 1882.220 22.060 ;
      LAYER met2 ;
        RECT 1636.550 600.170 1636.830 604.000 ;
        RECT 1636.550 600.030 1638.360 600.170 ;
        RECT 1636.550 600.000 1636.830 600.030 ;
        RECT 1638.220 586.830 1638.360 600.030 ;
        RECT 1638.160 586.510 1638.420 586.830 ;
        RECT 1641.840 586.510 1642.100 586.830 ;
        RECT 1641.900 22.090 1642.040 586.510 ;
        RECT 1641.840 21.770 1642.100 22.090 ;
        RECT 1881.960 21.770 1882.220 22.090 ;
        RECT 1882.020 2.400 1882.160 21.770 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1648.250 22.680 1648.570 22.740 ;
        RECT 1899.870 22.680 1900.190 22.740 ;
        RECT 1648.250 22.540 1900.190 22.680 ;
        RECT 1648.250 22.480 1648.570 22.540 ;
        RECT 1899.870 22.480 1900.190 22.540 ;
      LAYER via ;
        RECT 1648.280 22.480 1648.540 22.740 ;
        RECT 1899.900 22.480 1900.160 22.740 ;
      LAYER met2 ;
        RECT 1645.750 600.170 1646.030 604.000 ;
        RECT 1645.750 600.030 1648.480 600.170 ;
        RECT 1645.750 600.000 1646.030 600.030 ;
        RECT 1648.340 22.770 1648.480 600.030 ;
        RECT 1648.280 22.450 1648.540 22.770 ;
        RECT 1899.900 22.450 1900.160 22.770 ;
        RECT 1899.960 2.400 1900.100 22.450 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1655.610 23.020 1655.930 23.080 ;
        RECT 1917.810 23.020 1918.130 23.080 ;
        RECT 1655.610 22.880 1918.130 23.020 ;
        RECT 1655.610 22.820 1655.930 22.880 ;
        RECT 1917.810 22.820 1918.130 22.880 ;
      LAYER via ;
        RECT 1655.640 22.820 1655.900 23.080 ;
        RECT 1917.840 22.820 1918.100 23.080 ;
      LAYER met2 ;
        RECT 1654.950 600.170 1655.230 604.000 ;
        RECT 1654.950 600.030 1655.840 600.170 ;
        RECT 1654.950 600.000 1655.230 600.030 ;
        RECT 1655.700 23.110 1655.840 600.030 ;
        RECT 1655.640 22.790 1655.900 23.110 ;
        RECT 1917.840 22.790 1918.100 23.110 ;
        RECT 1917.900 2.400 1918.040 22.790 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1665.730 586.740 1666.050 586.800 ;
        RECT 1669.410 586.740 1669.730 586.800 ;
        RECT 1665.730 586.600 1669.730 586.740 ;
        RECT 1665.730 586.540 1666.050 586.600 ;
        RECT 1669.410 586.540 1669.730 586.600 ;
        RECT 1669.410 23.360 1669.730 23.420 ;
        RECT 1935.290 23.360 1935.610 23.420 ;
        RECT 1669.410 23.220 1935.610 23.360 ;
        RECT 1669.410 23.160 1669.730 23.220 ;
        RECT 1935.290 23.160 1935.610 23.220 ;
      LAYER via ;
        RECT 1665.760 586.540 1666.020 586.800 ;
        RECT 1669.440 586.540 1669.700 586.800 ;
        RECT 1669.440 23.160 1669.700 23.420 ;
        RECT 1935.320 23.160 1935.580 23.420 ;
      LAYER met2 ;
        RECT 1664.150 600.170 1664.430 604.000 ;
        RECT 1664.150 600.030 1665.960 600.170 ;
        RECT 1664.150 600.000 1664.430 600.030 ;
        RECT 1665.820 586.830 1665.960 600.030 ;
        RECT 1665.760 586.510 1666.020 586.830 ;
        RECT 1669.440 586.510 1669.700 586.830 ;
        RECT 1669.500 23.450 1669.640 586.510 ;
        RECT 1669.440 23.130 1669.700 23.450 ;
        RECT 1935.320 23.130 1935.580 23.450 ;
        RECT 1935.380 2.400 1935.520 23.130 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1675.850 531.320 1676.170 531.380 ;
        RECT 1676.310 531.320 1676.630 531.380 ;
        RECT 1675.850 531.180 1676.630 531.320 ;
        RECT 1675.850 531.120 1676.170 531.180 ;
        RECT 1676.310 531.120 1676.630 531.180 ;
        RECT 1676.310 496.980 1676.630 497.040 ;
        RECT 1675.940 496.840 1676.630 496.980 ;
        RECT 1675.940 496.700 1676.080 496.840 ;
        RECT 1676.310 496.780 1676.630 496.840 ;
        RECT 1675.850 496.440 1676.170 496.700 ;
        RECT 1675.390 444.960 1675.710 445.020 ;
        RECT 1676.310 444.960 1676.630 445.020 ;
        RECT 1675.390 444.820 1676.630 444.960 ;
        RECT 1675.390 444.760 1675.710 444.820 ;
        RECT 1676.310 444.760 1676.630 444.820 ;
        RECT 1675.390 386.480 1675.710 386.540 ;
        RECT 1675.850 386.480 1676.170 386.540 ;
        RECT 1675.390 386.340 1676.170 386.480 ;
        RECT 1675.390 386.280 1675.710 386.340 ;
        RECT 1675.850 386.280 1676.170 386.340 ;
        RECT 1675.390 379.680 1675.710 379.740 ;
        RECT 1675.850 379.680 1676.170 379.740 ;
        RECT 1675.390 379.540 1676.170 379.680 ;
        RECT 1675.390 379.480 1675.710 379.540 ;
        RECT 1675.850 379.480 1676.170 379.540 ;
        RECT 1675.850 331.060 1676.170 331.120 ;
        RECT 1676.770 331.060 1677.090 331.120 ;
        RECT 1675.850 330.920 1677.090 331.060 ;
        RECT 1675.850 330.860 1676.170 330.920 ;
        RECT 1676.770 330.860 1677.090 330.920 ;
        RECT 1675.850 283.120 1676.170 283.180 ;
        RECT 1676.770 283.120 1677.090 283.180 ;
        RECT 1675.850 282.980 1677.090 283.120 ;
        RECT 1675.850 282.920 1676.170 282.980 ;
        RECT 1676.770 282.920 1677.090 282.980 ;
        RECT 1675.390 158.680 1675.710 158.740 ;
        RECT 1676.310 158.680 1676.630 158.740 ;
        RECT 1675.390 158.540 1676.630 158.680 ;
        RECT 1675.390 158.480 1675.710 158.540 ;
        RECT 1676.310 158.480 1676.630 158.540 ;
        RECT 1676.310 137.940 1676.630 138.000 ;
        RECT 1677.230 137.940 1677.550 138.000 ;
        RECT 1676.310 137.800 1677.550 137.940 ;
        RECT 1676.310 137.740 1676.630 137.800 ;
        RECT 1677.230 137.740 1677.550 137.800 ;
        RECT 1675.390 90.000 1675.710 90.060 ;
        RECT 1677.230 90.000 1677.550 90.060 ;
        RECT 1675.390 89.860 1677.550 90.000 ;
        RECT 1675.390 89.800 1675.710 89.860 ;
        RECT 1677.230 89.800 1677.550 89.860 ;
        RECT 1675.390 62.600 1675.710 62.860 ;
        RECT 1675.480 61.840 1675.620 62.600 ;
        RECT 1675.390 61.580 1675.710 61.840 ;
        RECT 1675.390 23.700 1675.710 23.760 ;
        RECT 1953.230 23.700 1953.550 23.760 ;
        RECT 1675.390 23.560 1953.550 23.700 ;
        RECT 1675.390 23.500 1675.710 23.560 ;
        RECT 1953.230 23.500 1953.550 23.560 ;
      LAYER via ;
        RECT 1675.880 531.120 1676.140 531.380 ;
        RECT 1676.340 531.120 1676.600 531.380 ;
        RECT 1676.340 496.780 1676.600 497.040 ;
        RECT 1675.880 496.440 1676.140 496.700 ;
        RECT 1675.420 444.760 1675.680 445.020 ;
        RECT 1676.340 444.760 1676.600 445.020 ;
        RECT 1675.420 386.280 1675.680 386.540 ;
        RECT 1675.880 386.280 1676.140 386.540 ;
        RECT 1675.420 379.480 1675.680 379.740 ;
        RECT 1675.880 379.480 1676.140 379.740 ;
        RECT 1675.880 330.860 1676.140 331.120 ;
        RECT 1676.800 330.860 1677.060 331.120 ;
        RECT 1675.880 282.920 1676.140 283.180 ;
        RECT 1676.800 282.920 1677.060 283.180 ;
        RECT 1675.420 158.480 1675.680 158.740 ;
        RECT 1676.340 158.480 1676.600 158.740 ;
        RECT 1676.340 137.740 1676.600 138.000 ;
        RECT 1677.260 137.740 1677.520 138.000 ;
        RECT 1675.420 89.800 1675.680 90.060 ;
        RECT 1677.260 89.800 1677.520 90.060 ;
        RECT 1675.420 62.600 1675.680 62.860 ;
        RECT 1675.420 61.580 1675.680 61.840 ;
        RECT 1675.420 23.500 1675.680 23.760 ;
        RECT 1953.260 23.500 1953.520 23.760 ;
      LAYER met2 ;
        RECT 1673.350 600.170 1673.630 604.000 ;
        RECT 1673.350 600.030 1674.700 600.170 ;
        RECT 1673.350 600.000 1673.630 600.030 ;
        RECT 1674.560 579.885 1674.700 600.030 ;
        RECT 1674.490 579.515 1674.770 579.885 ;
        RECT 1675.410 579.515 1675.690 579.885 ;
        RECT 1675.480 545.090 1675.620 579.515 ;
        RECT 1675.480 544.950 1676.080 545.090 ;
        RECT 1675.940 531.410 1676.080 544.950 ;
        RECT 1675.880 531.090 1676.140 531.410 ;
        RECT 1676.340 531.090 1676.600 531.410 ;
        RECT 1676.400 497.070 1676.540 531.090 ;
        RECT 1676.340 496.750 1676.600 497.070 ;
        RECT 1675.880 496.410 1676.140 496.730 ;
        RECT 1675.940 483.210 1676.080 496.410 ;
        RECT 1675.940 483.070 1676.540 483.210 ;
        RECT 1676.400 445.050 1676.540 483.070 ;
        RECT 1675.420 444.730 1675.680 445.050 ;
        RECT 1676.340 444.730 1676.600 445.050 ;
        RECT 1675.480 386.570 1675.620 444.730 ;
        RECT 1675.420 386.250 1675.680 386.570 ;
        RECT 1675.880 386.250 1676.140 386.570 ;
        RECT 1675.940 379.770 1676.080 386.250 ;
        RECT 1675.420 379.450 1675.680 379.770 ;
        RECT 1675.880 379.450 1676.140 379.770 ;
        RECT 1675.480 338.370 1675.620 379.450 ;
        RECT 1675.480 338.230 1676.080 338.370 ;
        RECT 1675.940 331.150 1676.080 338.230 ;
        RECT 1675.880 330.830 1676.140 331.150 ;
        RECT 1676.800 330.830 1677.060 331.150 ;
        RECT 1676.860 283.210 1677.000 330.830 ;
        RECT 1675.880 282.890 1676.140 283.210 ;
        RECT 1676.800 282.890 1677.060 283.210 ;
        RECT 1675.940 255.410 1676.080 282.890 ;
        RECT 1675.480 255.270 1676.080 255.410 ;
        RECT 1675.480 158.770 1675.620 255.270 ;
        RECT 1675.420 158.450 1675.680 158.770 ;
        RECT 1676.340 158.450 1676.600 158.770 ;
        RECT 1676.400 138.030 1676.540 158.450 ;
        RECT 1676.340 137.710 1676.600 138.030 ;
        RECT 1677.260 137.710 1677.520 138.030 ;
        RECT 1677.320 90.090 1677.460 137.710 ;
        RECT 1675.420 89.770 1675.680 90.090 ;
        RECT 1677.260 89.770 1677.520 90.090 ;
        RECT 1675.480 62.890 1675.620 89.770 ;
        RECT 1675.420 62.570 1675.680 62.890 ;
        RECT 1675.420 61.550 1675.680 61.870 ;
        RECT 1675.480 23.790 1675.620 61.550 ;
        RECT 1675.420 23.470 1675.680 23.790 ;
        RECT 1953.260 23.470 1953.520 23.790 ;
        RECT 1953.320 2.400 1953.460 23.470 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
      LAYER via2 ;
        RECT 1674.490 579.560 1674.770 579.840 ;
        RECT 1675.410 579.560 1675.690 579.840 ;
      LAYER met3 ;
        RECT 1674.465 579.850 1674.795 579.865 ;
        RECT 1675.385 579.850 1675.715 579.865 ;
        RECT 1674.465 579.550 1675.715 579.850 ;
        RECT 1674.465 579.535 1674.795 579.550 ;
        RECT 1675.385 579.535 1675.715 579.550 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.210 27.440 1683.530 27.500 ;
        RECT 1971.170 27.440 1971.490 27.500 ;
        RECT 1683.210 27.300 1971.490 27.440 ;
        RECT 1683.210 27.240 1683.530 27.300 ;
        RECT 1971.170 27.240 1971.490 27.300 ;
      LAYER via ;
        RECT 1683.240 27.240 1683.500 27.500 ;
        RECT 1971.200 27.240 1971.460 27.500 ;
      LAYER met2 ;
        RECT 1682.550 600.170 1682.830 604.000 ;
        RECT 1682.550 600.030 1683.440 600.170 ;
        RECT 1682.550 600.000 1682.830 600.030 ;
        RECT 1683.300 27.530 1683.440 600.030 ;
        RECT 1683.240 27.210 1683.500 27.530 ;
        RECT 1971.200 27.210 1971.460 27.530 ;
        RECT 1971.260 2.400 1971.400 27.210 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1693.330 586.740 1693.650 586.800 ;
        RECT 1697.010 586.740 1697.330 586.800 ;
        RECT 1693.330 586.600 1697.330 586.740 ;
        RECT 1693.330 586.540 1693.650 586.600 ;
        RECT 1697.010 586.540 1697.330 586.600 ;
        RECT 1697.010 27.100 1697.330 27.160 ;
        RECT 1989.110 27.100 1989.430 27.160 ;
        RECT 1697.010 26.960 1989.430 27.100 ;
        RECT 1697.010 26.900 1697.330 26.960 ;
        RECT 1989.110 26.900 1989.430 26.960 ;
      LAYER via ;
        RECT 1693.360 586.540 1693.620 586.800 ;
        RECT 1697.040 586.540 1697.300 586.800 ;
        RECT 1697.040 26.900 1697.300 27.160 ;
        RECT 1989.140 26.900 1989.400 27.160 ;
      LAYER met2 ;
        RECT 1691.750 600.170 1692.030 604.000 ;
        RECT 1691.750 600.030 1693.560 600.170 ;
        RECT 1691.750 600.000 1692.030 600.030 ;
        RECT 1693.420 586.830 1693.560 600.030 ;
        RECT 1693.360 586.510 1693.620 586.830 ;
        RECT 1697.040 586.510 1697.300 586.830 ;
        RECT 1697.100 27.190 1697.240 586.510 ;
        RECT 1697.040 26.870 1697.300 27.190 ;
        RECT 1989.140 26.870 1989.400 27.190 ;
        RECT 1989.200 2.400 1989.340 26.870 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1702.530 586.740 1702.850 586.800 ;
        RECT 1703.910 586.740 1704.230 586.800 ;
        RECT 1702.530 586.600 1704.230 586.740 ;
        RECT 1702.530 586.540 1702.850 586.600 ;
        RECT 1703.910 586.540 1704.230 586.600 ;
        RECT 1703.910 26.760 1704.230 26.820 ;
        RECT 2006.590 26.760 2006.910 26.820 ;
        RECT 1703.910 26.620 2006.910 26.760 ;
        RECT 1703.910 26.560 1704.230 26.620 ;
        RECT 2006.590 26.560 2006.910 26.620 ;
      LAYER via ;
        RECT 1702.560 586.540 1702.820 586.800 ;
        RECT 1703.940 586.540 1704.200 586.800 ;
        RECT 1703.940 26.560 1704.200 26.820 ;
        RECT 2006.620 26.560 2006.880 26.820 ;
      LAYER met2 ;
        RECT 1700.950 600.170 1701.230 604.000 ;
        RECT 1700.950 600.030 1702.760 600.170 ;
        RECT 1700.950 600.000 1701.230 600.030 ;
        RECT 1702.620 586.830 1702.760 600.030 ;
        RECT 1702.560 586.510 1702.820 586.830 ;
        RECT 1703.940 586.510 1704.200 586.830 ;
        RECT 1704.000 26.850 1704.140 586.510 ;
        RECT 1703.940 26.530 1704.200 26.850 ;
        RECT 2006.620 26.530 2006.880 26.850 ;
        RECT 2006.680 2.400 2006.820 26.530 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 26.420 1711.130 26.480 ;
        RECT 2024.530 26.420 2024.850 26.480 ;
        RECT 1710.810 26.280 2024.850 26.420 ;
        RECT 1710.810 26.220 1711.130 26.280 ;
        RECT 2024.530 26.220 2024.850 26.280 ;
      LAYER via ;
        RECT 1710.840 26.220 1711.100 26.480 ;
        RECT 2024.560 26.220 2024.820 26.480 ;
      LAYER met2 ;
        RECT 1710.150 600.170 1710.430 604.000 ;
        RECT 1710.150 600.030 1711.040 600.170 ;
        RECT 1710.150 600.000 1710.430 600.030 ;
        RECT 1710.900 26.510 1711.040 600.030 ;
        RECT 1710.840 26.190 1711.100 26.510 ;
        RECT 2024.560 26.190 2024.820 26.510 ;
        RECT 2024.620 2.400 2024.760 26.190 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1720.930 589.800 1721.250 589.860 ;
        RECT 1724.610 589.800 1724.930 589.860 ;
        RECT 1720.930 589.660 1724.930 589.800 ;
        RECT 1720.930 589.600 1721.250 589.660 ;
        RECT 1724.610 589.600 1724.930 589.660 ;
        RECT 1724.610 26.080 1724.930 26.140 ;
        RECT 2042.470 26.080 2042.790 26.140 ;
        RECT 1724.610 25.940 2042.790 26.080 ;
        RECT 1724.610 25.880 1724.930 25.940 ;
        RECT 2042.470 25.880 2042.790 25.940 ;
      LAYER via ;
        RECT 1720.960 589.600 1721.220 589.860 ;
        RECT 1724.640 589.600 1724.900 589.860 ;
        RECT 1724.640 25.880 1724.900 26.140 ;
        RECT 2042.500 25.880 2042.760 26.140 ;
      LAYER met2 ;
        RECT 1719.350 600.170 1719.630 604.000 ;
        RECT 1719.350 600.030 1721.160 600.170 ;
        RECT 1719.350 600.000 1719.630 600.030 ;
        RECT 1721.020 589.890 1721.160 600.030 ;
        RECT 1720.960 589.570 1721.220 589.890 ;
        RECT 1724.640 589.570 1724.900 589.890 ;
        RECT 1724.700 26.170 1724.840 589.570 ;
        RECT 1724.640 25.850 1724.900 26.170 ;
        RECT 2042.500 25.850 2042.760 26.170 ;
        RECT 2042.560 2.400 2042.700 25.850 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 976.190 589.120 976.510 589.180 ;
        RECT 979.870 589.120 980.190 589.180 ;
        RECT 976.190 588.980 980.190 589.120 ;
        RECT 976.190 588.920 976.510 588.980 ;
        RECT 979.870 588.920 980.190 588.980 ;
        RECT 979.870 588.440 980.190 588.500 ;
        RECT 1057.610 588.440 1057.930 588.500 ;
        RECT 979.870 588.300 1057.930 588.440 ;
        RECT 979.870 588.240 980.190 588.300 ;
        RECT 1057.610 588.240 1057.930 588.300 ;
        RECT 757.690 18.600 758.010 18.660 ;
        RECT 976.190 18.600 976.510 18.660 ;
        RECT 757.690 18.460 976.510 18.600 ;
        RECT 757.690 18.400 758.010 18.460 ;
        RECT 976.190 18.400 976.510 18.460 ;
      LAYER via ;
        RECT 976.220 588.920 976.480 589.180 ;
        RECT 979.900 588.920 980.160 589.180 ;
        RECT 979.900 588.240 980.160 588.500 ;
        RECT 1057.640 588.240 1057.900 588.500 ;
        RECT 757.720 18.400 757.980 18.660 ;
        RECT 976.220 18.400 976.480 18.660 ;
      LAYER met2 ;
        RECT 1059.250 600.170 1059.530 604.000 ;
        RECT 1057.700 600.030 1059.530 600.170 ;
        RECT 976.220 588.890 976.480 589.210 ;
        RECT 979.900 588.890 980.160 589.210 ;
        RECT 976.280 18.690 976.420 588.890 ;
        RECT 979.960 588.530 980.100 588.890 ;
        RECT 1057.700 588.530 1057.840 600.030 ;
        RECT 1059.250 600.000 1059.530 600.030 ;
        RECT 979.900 588.210 980.160 588.530 ;
        RECT 1057.640 588.210 1057.900 588.530 ;
        RECT 757.720 18.370 757.980 18.690 ;
        RECT 976.220 18.370 976.480 18.690 ;
        RECT 757.780 2.400 757.920 18.370 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1729.670 586.740 1729.990 586.800 ;
        RECT 1731.510 586.740 1731.830 586.800 ;
        RECT 1729.670 586.600 1731.830 586.740 ;
        RECT 1729.670 586.540 1729.990 586.600 ;
        RECT 1731.510 586.540 1731.830 586.600 ;
        RECT 1731.510 25.740 1731.830 25.800 ;
        RECT 2060.410 25.740 2060.730 25.800 ;
        RECT 1731.510 25.600 2060.730 25.740 ;
        RECT 1731.510 25.540 1731.830 25.600 ;
        RECT 2060.410 25.540 2060.730 25.600 ;
      LAYER via ;
        RECT 1729.700 586.540 1729.960 586.800 ;
        RECT 1731.540 586.540 1731.800 586.800 ;
        RECT 1731.540 25.540 1731.800 25.800 ;
        RECT 2060.440 25.540 2060.700 25.800 ;
      LAYER met2 ;
        RECT 1728.090 600.170 1728.370 604.000 ;
        RECT 1728.090 600.030 1729.900 600.170 ;
        RECT 1728.090 600.000 1728.370 600.030 ;
        RECT 1729.760 586.830 1729.900 600.030 ;
        RECT 1729.700 586.510 1729.960 586.830 ;
        RECT 1731.540 586.510 1731.800 586.830 ;
        RECT 1731.600 25.830 1731.740 586.510 ;
        RECT 1731.540 25.510 1731.800 25.830 ;
        RECT 2060.440 25.510 2060.700 25.830 ;
        RECT 2060.500 2.400 2060.640 25.510 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1738.410 25.400 1738.730 25.460 ;
        RECT 2078.350 25.400 2078.670 25.460 ;
        RECT 1738.410 25.260 2078.670 25.400 ;
        RECT 1738.410 25.200 1738.730 25.260 ;
        RECT 2078.350 25.200 2078.670 25.260 ;
      LAYER via ;
        RECT 1738.440 25.200 1738.700 25.460 ;
        RECT 2078.380 25.200 2078.640 25.460 ;
      LAYER met2 ;
        RECT 1737.290 600.170 1737.570 604.000 ;
        RECT 1737.290 600.030 1738.640 600.170 ;
        RECT 1737.290 600.000 1737.570 600.030 ;
        RECT 1738.500 25.490 1738.640 600.030 ;
        RECT 1738.440 25.170 1738.700 25.490 ;
        RECT 2078.380 25.170 2078.640 25.490 ;
        RECT 2078.440 2.400 2078.580 25.170 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1748.070 592.180 1748.390 592.240 ;
        RECT 1752.210 592.180 1752.530 592.240 ;
        RECT 1748.070 592.040 1752.530 592.180 ;
        RECT 1748.070 591.980 1748.390 592.040 ;
        RECT 1752.210 591.980 1752.530 592.040 ;
        RECT 1752.210 25.060 1752.530 25.120 ;
        RECT 2095.830 25.060 2096.150 25.120 ;
        RECT 1752.210 24.920 2096.150 25.060 ;
        RECT 1752.210 24.860 1752.530 24.920 ;
        RECT 2095.830 24.860 2096.150 24.920 ;
      LAYER via ;
        RECT 1748.100 591.980 1748.360 592.240 ;
        RECT 1752.240 591.980 1752.500 592.240 ;
        RECT 1752.240 24.860 1752.500 25.120 ;
        RECT 2095.860 24.860 2096.120 25.120 ;
      LAYER met2 ;
        RECT 1746.490 600.170 1746.770 604.000 ;
        RECT 1746.490 600.030 1748.300 600.170 ;
        RECT 1746.490 600.000 1746.770 600.030 ;
        RECT 1748.160 592.270 1748.300 600.030 ;
        RECT 1748.100 591.950 1748.360 592.270 ;
        RECT 1752.240 591.950 1752.500 592.270 ;
        RECT 1752.300 25.150 1752.440 591.950 ;
        RECT 1752.240 24.830 1752.500 25.150 ;
        RECT 2095.860 24.830 2096.120 25.150 ;
        RECT 2095.920 2.400 2096.060 24.830 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1757.270 586.740 1757.590 586.800 ;
        RECT 1759.110 586.740 1759.430 586.800 ;
        RECT 1757.270 586.600 1759.430 586.740 ;
        RECT 1757.270 586.540 1757.590 586.600 ;
        RECT 1759.110 586.540 1759.430 586.600 ;
        RECT 1759.110 24.720 1759.430 24.780 ;
        RECT 2113.770 24.720 2114.090 24.780 ;
        RECT 1759.110 24.580 2114.090 24.720 ;
        RECT 1759.110 24.520 1759.430 24.580 ;
        RECT 2113.770 24.520 2114.090 24.580 ;
      LAYER via ;
        RECT 1757.300 586.540 1757.560 586.800 ;
        RECT 1759.140 586.540 1759.400 586.800 ;
        RECT 1759.140 24.520 1759.400 24.780 ;
        RECT 2113.800 24.520 2114.060 24.780 ;
      LAYER met2 ;
        RECT 1755.690 600.170 1755.970 604.000 ;
        RECT 1755.690 600.030 1757.500 600.170 ;
        RECT 1755.690 600.000 1755.970 600.030 ;
        RECT 1757.360 586.830 1757.500 600.030 ;
        RECT 1757.300 586.510 1757.560 586.830 ;
        RECT 1759.140 586.510 1759.400 586.830 ;
        RECT 1759.200 24.810 1759.340 586.510 ;
        RECT 1759.140 24.490 1759.400 24.810 ;
        RECT 2113.800 24.490 2114.060 24.810 ;
        RECT 2113.860 2.400 2114.000 24.490 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.010 24.380 1766.330 24.440 ;
        RECT 2131.710 24.380 2132.030 24.440 ;
        RECT 1766.010 24.240 2132.030 24.380 ;
        RECT 1766.010 24.180 1766.330 24.240 ;
        RECT 2131.710 24.180 2132.030 24.240 ;
      LAYER via ;
        RECT 1766.040 24.180 1766.300 24.440 ;
        RECT 2131.740 24.180 2132.000 24.440 ;
      LAYER met2 ;
        RECT 1764.890 600.170 1765.170 604.000 ;
        RECT 1764.890 600.030 1766.240 600.170 ;
        RECT 1764.890 600.000 1765.170 600.030 ;
        RECT 1766.100 24.470 1766.240 600.030 ;
        RECT 1766.040 24.150 1766.300 24.470 ;
        RECT 2131.740 24.150 2132.000 24.470 ;
        RECT 2131.800 2.400 2131.940 24.150 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1775.670 590.140 1775.990 590.200 ;
        RECT 1779.810 590.140 1780.130 590.200 ;
        RECT 1775.670 590.000 1780.130 590.140 ;
        RECT 1775.670 589.940 1775.990 590.000 ;
        RECT 1779.810 589.940 1780.130 590.000 ;
        RECT 1779.810 24.040 1780.130 24.100 ;
        RECT 2149.650 24.040 2149.970 24.100 ;
        RECT 1779.810 23.900 2149.970 24.040 ;
        RECT 1779.810 23.840 1780.130 23.900 ;
        RECT 2149.650 23.840 2149.970 23.900 ;
      LAYER via ;
        RECT 1775.700 589.940 1775.960 590.200 ;
        RECT 1779.840 589.940 1780.100 590.200 ;
        RECT 1779.840 23.840 1780.100 24.100 ;
        RECT 2149.680 23.840 2149.940 24.100 ;
      LAYER met2 ;
        RECT 1774.090 600.170 1774.370 604.000 ;
        RECT 1774.090 600.030 1775.900 600.170 ;
        RECT 1774.090 600.000 1774.370 600.030 ;
        RECT 1775.760 590.230 1775.900 600.030 ;
        RECT 1775.700 589.910 1775.960 590.230 ;
        RECT 1779.840 589.910 1780.100 590.230 ;
        RECT 1779.900 24.130 1780.040 589.910 ;
        RECT 1779.840 23.810 1780.100 24.130 ;
        RECT 2149.680 23.810 2149.940 24.130 ;
        RECT 2149.740 2.400 2149.880 23.810 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1784.870 586.740 1785.190 586.800 ;
        RECT 1786.710 586.740 1787.030 586.800 ;
        RECT 1784.870 586.600 1787.030 586.740 ;
        RECT 1784.870 586.540 1785.190 586.600 ;
        RECT 1786.710 586.540 1787.030 586.600 ;
        RECT 1786.710 36.280 1787.030 36.340 ;
        RECT 2167.590 36.280 2167.910 36.340 ;
        RECT 1786.710 36.140 2167.910 36.280 ;
        RECT 1786.710 36.080 1787.030 36.140 ;
        RECT 2167.590 36.080 2167.910 36.140 ;
      LAYER via ;
        RECT 1784.900 586.540 1785.160 586.800 ;
        RECT 1786.740 586.540 1787.000 586.800 ;
        RECT 1786.740 36.080 1787.000 36.340 ;
        RECT 2167.620 36.080 2167.880 36.340 ;
      LAYER met2 ;
        RECT 1783.290 600.170 1783.570 604.000 ;
        RECT 1783.290 600.030 1785.100 600.170 ;
        RECT 1783.290 600.000 1783.570 600.030 ;
        RECT 1784.960 586.830 1785.100 600.030 ;
        RECT 1784.900 586.510 1785.160 586.830 ;
        RECT 1786.740 586.510 1787.000 586.830 ;
        RECT 1786.800 36.370 1786.940 586.510 ;
        RECT 1786.740 36.050 1787.000 36.370 ;
        RECT 2167.620 36.050 2167.880 36.370 ;
        RECT 2167.680 2.400 2167.820 36.050 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 43.080 1793.930 43.140 ;
        RECT 2185.070 43.080 2185.390 43.140 ;
        RECT 1793.610 42.940 2185.390 43.080 ;
        RECT 1793.610 42.880 1793.930 42.940 ;
        RECT 2185.070 42.880 2185.390 42.940 ;
      LAYER via ;
        RECT 1793.640 42.880 1793.900 43.140 ;
        RECT 2185.100 42.880 2185.360 43.140 ;
      LAYER met2 ;
        RECT 1792.490 600.170 1792.770 604.000 ;
        RECT 1792.490 600.030 1793.840 600.170 ;
        RECT 1792.490 600.000 1792.770 600.030 ;
        RECT 1793.700 43.170 1793.840 600.030 ;
        RECT 1793.640 42.850 1793.900 43.170 ;
        RECT 2185.100 42.850 2185.360 43.170 ;
        RECT 2185.160 2.400 2185.300 42.850 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1803.270 590.140 1803.590 590.200 ;
        RECT 1807.410 590.140 1807.730 590.200 ;
        RECT 1803.270 590.000 1807.730 590.140 ;
        RECT 1803.270 589.940 1803.590 590.000 ;
        RECT 1807.410 589.940 1807.730 590.000 ;
        RECT 1807.410 43.420 1807.730 43.480 ;
        RECT 2203.010 43.420 2203.330 43.480 ;
        RECT 1807.410 43.280 2203.330 43.420 ;
        RECT 1807.410 43.220 1807.730 43.280 ;
        RECT 2203.010 43.220 2203.330 43.280 ;
      LAYER via ;
        RECT 1803.300 589.940 1803.560 590.200 ;
        RECT 1807.440 589.940 1807.700 590.200 ;
        RECT 1807.440 43.220 1807.700 43.480 ;
        RECT 2203.040 43.220 2203.300 43.480 ;
      LAYER met2 ;
        RECT 1801.690 600.170 1801.970 604.000 ;
        RECT 1801.690 600.030 1803.500 600.170 ;
        RECT 1801.690 600.000 1801.970 600.030 ;
        RECT 1803.360 590.230 1803.500 600.030 ;
        RECT 1803.300 589.910 1803.560 590.230 ;
        RECT 1807.440 589.910 1807.700 590.230 ;
        RECT 1807.500 43.510 1807.640 589.910 ;
        RECT 1807.440 43.190 1807.700 43.510 ;
        RECT 2203.040 43.190 2203.300 43.510 ;
        RECT 2203.100 2.400 2203.240 43.190 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1812.470 586.740 1812.790 586.800 ;
        RECT 1814.310 586.740 1814.630 586.800 ;
        RECT 1812.470 586.600 1814.630 586.740 ;
        RECT 1812.470 586.540 1812.790 586.600 ;
        RECT 1814.310 586.540 1814.630 586.600 ;
        RECT 1814.310 43.760 1814.630 43.820 ;
        RECT 2220.950 43.760 2221.270 43.820 ;
        RECT 1814.310 43.620 2221.270 43.760 ;
        RECT 1814.310 43.560 1814.630 43.620 ;
        RECT 2220.950 43.560 2221.270 43.620 ;
      LAYER via ;
        RECT 1812.500 586.540 1812.760 586.800 ;
        RECT 1814.340 586.540 1814.600 586.800 ;
        RECT 1814.340 43.560 1814.600 43.820 ;
        RECT 2220.980 43.560 2221.240 43.820 ;
      LAYER met2 ;
        RECT 1810.890 600.170 1811.170 604.000 ;
        RECT 1810.890 600.030 1812.700 600.170 ;
        RECT 1810.890 600.000 1811.170 600.030 ;
        RECT 1812.560 586.830 1812.700 600.030 ;
        RECT 1812.500 586.510 1812.760 586.830 ;
        RECT 1814.340 586.510 1814.600 586.830 ;
        RECT 1814.400 43.850 1814.540 586.510 ;
        RECT 1814.340 43.530 1814.600 43.850 ;
        RECT 2220.980 43.530 2221.240 43.850 ;
        RECT 2221.040 2.400 2221.180 43.530 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1063.130 569.400 1063.450 569.460 ;
        RECT 1066.810 569.400 1067.130 569.460 ;
        RECT 1063.130 569.260 1067.130 569.400 ;
        RECT 1063.130 569.200 1063.450 569.260 ;
        RECT 1066.810 569.200 1067.130 569.260 ;
        RECT 858.890 27.100 859.210 27.160 ;
        RECT 1063.130 27.100 1063.450 27.160 ;
        RECT 858.890 26.960 1063.450 27.100 ;
        RECT 858.890 26.900 859.210 26.960 ;
        RECT 1063.130 26.900 1063.450 26.960 ;
        RECT 775.630 18.260 775.950 18.320 ;
        RECT 858.890 18.260 859.210 18.320 ;
        RECT 775.630 18.120 859.210 18.260 ;
        RECT 775.630 18.060 775.950 18.120 ;
        RECT 858.890 18.060 859.210 18.120 ;
      LAYER via ;
        RECT 1063.160 569.200 1063.420 569.460 ;
        RECT 1066.840 569.200 1067.100 569.460 ;
        RECT 858.920 26.900 859.180 27.160 ;
        RECT 1063.160 26.900 1063.420 27.160 ;
        RECT 775.660 18.060 775.920 18.320 ;
        RECT 858.920 18.060 859.180 18.320 ;
      LAYER met2 ;
        RECT 1068.450 600.170 1068.730 604.000 ;
        RECT 1066.900 600.030 1068.730 600.170 ;
        RECT 1066.900 569.490 1067.040 600.030 ;
        RECT 1068.450 600.000 1068.730 600.030 ;
        RECT 1063.160 569.170 1063.420 569.490 ;
        RECT 1066.840 569.170 1067.100 569.490 ;
        RECT 1063.220 27.190 1063.360 569.170 ;
        RECT 858.920 26.870 859.180 27.190 ;
        RECT 1063.160 26.870 1063.420 27.190 ;
        RECT 858.980 18.350 859.120 26.870 ;
        RECT 775.660 18.030 775.920 18.350 ;
        RECT 858.920 18.030 859.180 18.350 ;
        RECT 775.720 2.400 775.860 18.030 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.210 44.100 1821.530 44.160 ;
        RECT 2238.890 44.100 2239.210 44.160 ;
        RECT 1821.210 43.960 2239.210 44.100 ;
        RECT 1821.210 43.900 1821.530 43.960 ;
        RECT 2238.890 43.900 2239.210 43.960 ;
      LAYER via ;
        RECT 1821.240 43.900 1821.500 44.160 ;
        RECT 2238.920 43.900 2239.180 44.160 ;
      LAYER met2 ;
        RECT 1820.090 600.170 1820.370 604.000 ;
        RECT 1820.090 600.030 1821.440 600.170 ;
        RECT 1820.090 600.000 1820.370 600.030 ;
        RECT 1821.300 44.190 1821.440 600.030 ;
        RECT 1821.240 43.870 1821.500 44.190 ;
        RECT 2238.920 43.870 2239.180 44.190 ;
        RECT 2238.980 2.400 2239.120 43.870 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1830.870 590.140 1831.190 590.200 ;
        RECT 1835.010 590.140 1835.330 590.200 ;
        RECT 1830.870 590.000 1835.330 590.140 ;
        RECT 1830.870 589.940 1831.190 590.000 ;
        RECT 1835.010 589.940 1835.330 590.000 ;
        RECT 1835.010 44.440 1835.330 44.500 ;
        RECT 2256.830 44.440 2257.150 44.500 ;
        RECT 1835.010 44.300 2257.150 44.440 ;
        RECT 1835.010 44.240 1835.330 44.300 ;
        RECT 2256.830 44.240 2257.150 44.300 ;
      LAYER via ;
        RECT 1830.900 589.940 1831.160 590.200 ;
        RECT 1835.040 589.940 1835.300 590.200 ;
        RECT 1835.040 44.240 1835.300 44.500 ;
        RECT 2256.860 44.240 2257.120 44.500 ;
      LAYER met2 ;
        RECT 1829.290 600.170 1829.570 604.000 ;
        RECT 1829.290 600.030 1831.100 600.170 ;
        RECT 1829.290 600.000 1829.570 600.030 ;
        RECT 1830.960 590.230 1831.100 600.030 ;
        RECT 1830.900 589.910 1831.160 590.230 ;
        RECT 1835.040 589.910 1835.300 590.230 ;
        RECT 1835.100 44.530 1835.240 589.910 ;
        RECT 1835.040 44.210 1835.300 44.530 ;
        RECT 2256.860 44.210 2257.120 44.530 ;
        RECT 2256.920 7.210 2257.060 44.210 ;
        RECT 2256.460 7.070 2257.060 7.210 ;
        RECT 2256.460 2.400 2256.600 7.070 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1840.070 586.740 1840.390 586.800 ;
        RECT 1841.910 586.740 1842.230 586.800 ;
        RECT 1840.070 586.600 1842.230 586.740 ;
        RECT 1840.070 586.540 1840.390 586.600 ;
        RECT 1841.910 586.540 1842.230 586.600 ;
        RECT 1841.910 48.180 1842.230 48.240 ;
        RECT 2274.310 48.180 2274.630 48.240 ;
        RECT 1841.910 48.040 2274.630 48.180 ;
        RECT 1841.910 47.980 1842.230 48.040 ;
        RECT 2274.310 47.980 2274.630 48.040 ;
      LAYER via ;
        RECT 1840.100 586.540 1840.360 586.800 ;
        RECT 1841.940 586.540 1842.200 586.800 ;
        RECT 1841.940 47.980 1842.200 48.240 ;
        RECT 2274.340 47.980 2274.600 48.240 ;
      LAYER met2 ;
        RECT 1838.490 600.170 1838.770 604.000 ;
        RECT 1838.490 600.030 1840.300 600.170 ;
        RECT 1838.490 600.000 1838.770 600.030 ;
        RECT 1840.160 586.830 1840.300 600.030 ;
        RECT 1840.100 586.510 1840.360 586.830 ;
        RECT 1841.940 586.510 1842.200 586.830 ;
        RECT 1842.000 48.270 1842.140 586.510 ;
        RECT 1841.940 47.950 1842.200 48.270 ;
        RECT 2274.340 47.950 2274.600 48.270 ;
        RECT 2274.400 2.400 2274.540 47.950 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.350 47.500 1848.670 47.560 ;
        RECT 2292.250 47.500 2292.570 47.560 ;
        RECT 1848.350 47.360 2292.570 47.500 ;
        RECT 1848.350 47.300 1848.670 47.360 ;
        RECT 2292.250 47.300 2292.570 47.360 ;
      LAYER via ;
        RECT 1848.380 47.300 1848.640 47.560 ;
        RECT 2292.280 47.300 2292.540 47.560 ;
      LAYER met2 ;
        RECT 1847.230 600.170 1847.510 604.000 ;
        RECT 1847.230 600.030 1848.580 600.170 ;
        RECT 1847.230 600.000 1847.510 600.030 ;
        RECT 1848.440 47.590 1848.580 600.030 ;
        RECT 1848.380 47.270 1848.640 47.590 ;
        RECT 2292.280 47.270 2292.540 47.590 ;
        RECT 2292.340 2.400 2292.480 47.270 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1858.010 586.740 1858.330 586.800 ;
        RECT 1862.610 586.740 1862.930 586.800 ;
        RECT 1858.010 586.600 1862.930 586.740 ;
        RECT 1858.010 586.540 1858.330 586.600 ;
        RECT 1862.610 586.540 1862.930 586.600 ;
        RECT 1862.610 47.840 1862.930 47.900 ;
        RECT 2310.190 47.840 2310.510 47.900 ;
        RECT 1862.610 47.700 2310.510 47.840 ;
        RECT 1862.610 47.640 1862.930 47.700 ;
        RECT 2310.190 47.640 2310.510 47.700 ;
      LAYER via ;
        RECT 1858.040 586.540 1858.300 586.800 ;
        RECT 1862.640 586.540 1862.900 586.800 ;
        RECT 1862.640 47.640 1862.900 47.900 ;
        RECT 2310.220 47.640 2310.480 47.900 ;
      LAYER met2 ;
        RECT 1856.430 600.170 1856.710 604.000 ;
        RECT 1856.430 600.030 1858.240 600.170 ;
        RECT 1856.430 600.000 1856.710 600.030 ;
        RECT 1858.100 586.830 1858.240 600.030 ;
        RECT 1858.040 586.510 1858.300 586.830 ;
        RECT 1862.640 586.510 1862.900 586.830 ;
        RECT 1862.700 47.930 1862.840 586.510 ;
        RECT 1862.640 47.610 1862.900 47.930 ;
        RECT 2310.220 47.610 2310.480 47.930 ;
        RECT 2310.280 2.400 2310.420 47.610 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1867.210 586.740 1867.530 586.800 ;
        RECT 1869.050 586.740 1869.370 586.800 ;
        RECT 1867.210 586.600 1869.370 586.740 ;
        RECT 1867.210 586.540 1867.530 586.600 ;
        RECT 1869.050 586.540 1869.370 586.600 ;
        RECT 1869.050 28.120 1869.370 28.180 ;
        RECT 2328.130 28.120 2328.450 28.180 ;
        RECT 1869.050 27.980 2328.450 28.120 ;
        RECT 1869.050 27.920 1869.370 27.980 ;
        RECT 2328.130 27.920 2328.450 27.980 ;
      LAYER via ;
        RECT 1867.240 586.540 1867.500 586.800 ;
        RECT 1869.080 586.540 1869.340 586.800 ;
        RECT 1869.080 27.920 1869.340 28.180 ;
        RECT 2328.160 27.920 2328.420 28.180 ;
      LAYER met2 ;
        RECT 1865.630 600.170 1865.910 604.000 ;
        RECT 1865.630 600.030 1867.440 600.170 ;
        RECT 1865.630 600.000 1865.910 600.030 ;
        RECT 1867.300 586.830 1867.440 600.030 ;
        RECT 1867.240 586.510 1867.500 586.830 ;
        RECT 1869.080 586.510 1869.340 586.830 ;
        RECT 1869.140 28.210 1869.280 586.510 ;
        RECT 1869.080 27.890 1869.340 28.210 ;
        RECT 2328.160 27.890 2328.420 28.210 ;
        RECT 2328.220 2.400 2328.360 27.890 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.410 28.460 1876.730 28.520 ;
        RECT 2345.610 28.460 2345.930 28.520 ;
        RECT 1876.410 28.320 2345.930 28.460 ;
        RECT 1876.410 28.260 1876.730 28.320 ;
        RECT 2345.610 28.260 2345.930 28.320 ;
      LAYER via ;
        RECT 1876.440 28.260 1876.700 28.520 ;
        RECT 2345.640 28.260 2345.900 28.520 ;
      LAYER met2 ;
        RECT 1874.830 600.170 1875.110 604.000 ;
        RECT 1874.830 600.030 1876.640 600.170 ;
        RECT 1874.830 600.000 1875.110 600.030 ;
        RECT 1876.500 28.550 1876.640 600.030 ;
        RECT 1876.440 28.230 1876.700 28.550 ;
        RECT 2345.640 28.230 2345.900 28.550 ;
        RECT 2345.700 2.400 2345.840 28.230 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1885.610 586.740 1885.930 586.800 ;
        RECT 1890.210 586.740 1890.530 586.800 ;
        RECT 1885.610 586.600 1890.530 586.740 ;
        RECT 1885.610 586.540 1885.930 586.600 ;
        RECT 1890.210 586.540 1890.530 586.600 ;
        RECT 1890.210 28.800 1890.530 28.860 ;
        RECT 2363.550 28.800 2363.870 28.860 ;
        RECT 1890.210 28.660 2363.870 28.800 ;
        RECT 1890.210 28.600 1890.530 28.660 ;
        RECT 2363.550 28.600 2363.870 28.660 ;
      LAYER via ;
        RECT 1885.640 586.540 1885.900 586.800 ;
        RECT 1890.240 586.540 1890.500 586.800 ;
        RECT 1890.240 28.600 1890.500 28.860 ;
        RECT 2363.580 28.600 2363.840 28.860 ;
      LAYER met2 ;
        RECT 1884.030 600.170 1884.310 604.000 ;
        RECT 1884.030 600.030 1885.840 600.170 ;
        RECT 1884.030 600.000 1884.310 600.030 ;
        RECT 1885.700 586.830 1885.840 600.030 ;
        RECT 1885.640 586.510 1885.900 586.830 ;
        RECT 1890.240 586.510 1890.500 586.830 ;
        RECT 1890.300 28.890 1890.440 586.510 ;
        RECT 1890.240 28.570 1890.500 28.890 ;
        RECT 2363.580 28.570 2363.840 28.890 ;
        RECT 2363.640 2.400 2363.780 28.570 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1894.810 586.740 1895.130 586.800 ;
        RECT 1897.110 586.740 1897.430 586.800 ;
        RECT 1894.810 586.600 1897.430 586.740 ;
        RECT 1894.810 586.540 1895.130 586.600 ;
        RECT 1897.110 586.540 1897.430 586.600 ;
        RECT 1897.110 29.140 1897.430 29.200 ;
        RECT 2381.490 29.140 2381.810 29.200 ;
        RECT 1897.110 29.000 2381.810 29.140 ;
        RECT 1897.110 28.940 1897.430 29.000 ;
        RECT 2381.490 28.940 2381.810 29.000 ;
      LAYER via ;
        RECT 1894.840 586.540 1895.100 586.800 ;
        RECT 1897.140 586.540 1897.400 586.800 ;
        RECT 1897.140 28.940 1897.400 29.200 ;
        RECT 2381.520 28.940 2381.780 29.200 ;
      LAYER met2 ;
        RECT 1893.230 600.170 1893.510 604.000 ;
        RECT 1893.230 600.030 1895.040 600.170 ;
        RECT 1893.230 600.000 1893.510 600.030 ;
        RECT 1894.900 586.830 1895.040 600.030 ;
        RECT 1894.840 586.510 1895.100 586.830 ;
        RECT 1897.140 586.510 1897.400 586.830 ;
        RECT 1897.200 29.230 1897.340 586.510 ;
        RECT 1897.140 28.910 1897.400 29.230 ;
        RECT 2381.520 28.910 2381.780 29.230 ;
        RECT 2381.580 2.400 2381.720 28.910 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1903.550 29.480 1903.870 29.540 ;
        RECT 2399.430 29.480 2399.750 29.540 ;
        RECT 1903.550 29.340 2399.750 29.480 ;
        RECT 1903.550 29.280 1903.870 29.340 ;
        RECT 2399.430 29.280 2399.750 29.340 ;
      LAYER via ;
        RECT 1903.580 29.280 1903.840 29.540 ;
        RECT 2399.460 29.280 2399.720 29.540 ;
      LAYER met2 ;
        RECT 1902.430 600.170 1902.710 604.000 ;
        RECT 1902.430 600.030 1903.780 600.170 ;
        RECT 1902.430 600.000 1902.710 600.030 ;
        RECT 1903.640 29.570 1903.780 600.030 ;
        RECT 1903.580 29.250 1903.840 29.570 ;
        RECT 2399.460 29.250 2399.720 29.570 ;
        RECT 2399.520 2.400 2399.660 29.250 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.570 25.740 793.890 25.800 ;
        RECT 1076.470 25.740 1076.790 25.800 ;
        RECT 793.570 25.600 1076.790 25.740 ;
        RECT 793.570 25.540 793.890 25.600 ;
        RECT 1076.470 25.540 1076.790 25.600 ;
      LAYER via ;
        RECT 793.600 25.540 793.860 25.800 ;
        RECT 1076.500 25.540 1076.760 25.800 ;
      LAYER met2 ;
        RECT 1077.650 600.170 1077.930 604.000 ;
        RECT 1076.560 600.030 1077.930 600.170 ;
        RECT 1076.560 25.830 1076.700 600.030 ;
        RECT 1077.650 600.000 1077.930 600.030 ;
        RECT 793.600 25.510 793.860 25.830 ;
        RECT 1076.500 25.510 1076.760 25.830 ;
        RECT 793.660 2.400 793.800 25.510 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 994.590 476.240 994.910 476.300 ;
        RECT 995.970 476.240 996.290 476.300 ;
        RECT 994.590 476.100 996.290 476.240 ;
        RECT 994.590 476.040 994.910 476.100 ;
        RECT 995.970 476.040 996.290 476.100 ;
        RECT 994.590 434.420 994.910 434.480 ;
        RECT 995.970 434.420 996.290 434.480 ;
        RECT 994.590 434.280 996.290 434.420 ;
        RECT 994.590 434.220 994.910 434.280 ;
        RECT 995.970 434.220 996.290 434.280 ;
        RECT 995.050 420.820 995.370 420.880 ;
        RECT 995.970 420.820 996.290 420.880 ;
        RECT 995.050 420.680 996.290 420.820 ;
        RECT 995.050 420.620 995.370 420.680 ;
        RECT 995.970 420.620 996.290 420.680 ;
        RECT 995.050 414.020 995.370 414.080 ;
        RECT 995.970 414.020 996.290 414.080 ;
        RECT 995.050 413.880 996.290 414.020 ;
        RECT 995.050 413.820 995.370 413.880 ;
        RECT 995.970 413.820 996.290 413.880 ;
        RECT 994.130 366.080 994.450 366.140 ;
        RECT 995.970 366.080 996.290 366.140 ;
        RECT 994.130 365.940 996.290 366.080 ;
        RECT 994.130 365.880 994.450 365.940 ;
        RECT 995.970 365.880 996.290 365.940 ;
        RECT 994.130 338.540 994.450 338.600 ;
        RECT 994.130 338.400 994.820 338.540 ;
        RECT 994.130 338.340 994.450 338.400 ;
        RECT 994.680 337.580 994.820 338.400 ;
        RECT 994.590 337.320 994.910 337.580 ;
        RECT 994.590 234.500 994.910 234.560 ;
        RECT 995.970 234.500 996.290 234.560 ;
        RECT 994.590 234.360 996.290 234.500 ;
        RECT 994.590 234.300 994.910 234.360 ;
        RECT 995.970 234.300 996.290 234.360 ;
        RECT 994.590 144.740 994.910 144.800 ;
        RECT 995.050 144.740 995.370 144.800 ;
        RECT 994.590 144.600 995.370 144.740 ;
        RECT 994.590 144.540 994.910 144.600 ;
        RECT 995.050 144.540 995.370 144.600 ;
        RECT 994.590 96.800 994.910 96.860 ;
        RECT 995.050 96.800 995.370 96.860 ;
        RECT 994.590 96.660 995.370 96.800 ;
        RECT 994.590 96.600 994.910 96.660 ;
        RECT 995.050 96.600 995.370 96.660 ;
        RECT 639.010 36.620 639.330 36.680 ;
        RECT 995.050 36.620 995.370 36.680 ;
        RECT 639.010 36.480 995.370 36.620 ;
        RECT 639.010 36.420 639.330 36.480 ;
        RECT 995.050 36.420 995.370 36.480 ;
      LAYER via ;
        RECT 994.620 476.040 994.880 476.300 ;
        RECT 996.000 476.040 996.260 476.300 ;
        RECT 994.620 434.220 994.880 434.480 ;
        RECT 996.000 434.220 996.260 434.480 ;
        RECT 995.080 420.620 995.340 420.880 ;
        RECT 996.000 420.620 996.260 420.880 ;
        RECT 995.080 413.820 995.340 414.080 ;
        RECT 996.000 413.820 996.260 414.080 ;
        RECT 994.160 365.880 994.420 366.140 ;
        RECT 996.000 365.880 996.260 366.140 ;
        RECT 994.160 338.340 994.420 338.600 ;
        RECT 994.620 337.320 994.880 337.580 ;
        RECT 994.620 234.300 994.880 234.560 ;
        RECT 996.000 234.300 996.260 234.560 ;
        RECT 994.620 144.540 994.880 144.800 ;
        RECT 995.080 144.540 995.340 144.800 ;
        RECT 994.620 96.600 994.880 96.860 ;
        RECT 995.080 96.600 995.340 96.860 ;
        RECT 639.040 36.420 639.300 36.680 ;
        RECT 995.080 36.420 995.340 36.680 ;
      LAYER met2 ;
        RECT 998.070 600.000 998.350 604.000 ;
        RECT 998.130 598.810 998.270 600.000 ;
        RECT 997.900 598.670 998.270 598.810 ;
        RECT 997.900 579.885 998.040 598.670 ;
        RECT 995.990 579.515 996.270 579.885 ;
        RECT 997.830 579.515 998.110 579.885 ;
        RECT 996.060 476.330 996.200 579.515 ;
        RECT 994.620 476.010 994.880 476.330 ;
        RECT 996.000 476.010 996.260 476.330 ;
        RECT 994.680 434.510 994.820 476.010 ;
        RECT 994.620 434.190 994.880 434.510 ;
        RECT 996.000 434.190 996.260 434.510 ;
        RECT 996.060 420.910 996.200 434.190 ;
        RECT 995.080 420.590 995.340 420.910 ;
        RECT 996.000 420.590 996.260 420.910 ;
        RECT 995.140 414.110 995.280 420.590 ;
        RECT 995.080 413.790 995.340 414.110 ;
        RECT 996.000 413.790 996.260 414.110 ;
        RECT 996.060 366.170 996.200 413.790 ;
        RECT 994.160 365.850 994.420 366.170 ;
        RECT 996.000 365.850 996.260 366.170 ;
        RECT 994.220 338.630 994.360 365.850 ;
        RECT 994.160 338.310 994.420 338.630 ;
        RECT 994.620 337.290 994.880 337.610 ;
        RECT 994.680 317.290 994.820 337.290 ;
        RECT 994.680 317.150 995.280 317.290 ;
        RECT 995.140 241.810 995.280 317.150 ;
        RECT 994.680 241.670 995.280 241.810 ;
        RECT 994.680 234.590 994.820 241.670 ;
        RECT 994.620 234.270 994.880 234.590 ;
        RECT 996.000 234.270 996.260 234.590 ;
        RECT 996.060 145.365 996.200 234.270 ;
        RECT 995.070 144.995 995.350 145.365 ;
        RECT 995.990 144.995 996.270 145.365 ;
        RECT 995.140 144.830 995.280 144.995 ;
        RECT 994.620 144.510 994.880 144.830 ;
        RECT 995.080 144.510 995.340 144.830 ;
        RECT 994.680 96.890 994.820 144.510 ;
        RECT 994.620 96.570 994.880 96.890 ;
        RECT 995.080 96.570 995.340 96.890 ;
        RECT 995.140 36.710 995.280 96.570 ;
        RECT 639.040 36.390 639.300 36.710 ;
        RECT 995.080 36.390 995.340 36.710 ;
        RECT 639.100 2.400 639.240 36.390 ;
        RECT 638.890 -4.800 639.450 2.400 ;
      LAYER via2 ;
        RECT 995.990 579.560 996.270 579.840 ;
        RECT 997.830 579.560 998.110 579.840 ;
        RECT 995.070 145.040 995.350 145.320 ;
        RECT 995.990 145.040 996.270 145.320 ;
      LAYER met3 ;
        RECT 995.965 579.850 996.295 579.865 ;
        RECT 997.805 579.850 998.135 579.865 ;
        RECT 995.965 579.550 998.135 579.850 ;
        RECT 995.965 579.535 996.295 579.550 ;
        RECT 997.805 579.535 998.135 579.550 ;
        RECT 995.045 145.330 995.375 145.345 ;
        RECT 995.965 145.330 996.295 145.345 ;
        RECT 995.045 145.030 996.295 145.330 ;
        RECT 995.045 145.015 995.375 145.030 ;
        RECT 995.965 145.015 996.295 145.030 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1916.430 586.740 1916.750 586.800 ;
        RECT 1917.810 586.740 1918.130 586.800 ;
        RECT 1916.430 586.600 1918.130 586.740 ;
        RECT 1916.430 586.540 1916.750 586.600 ;
        RECT 1917.810 586.540 1918.130 586.600 ;
        RECT 1917.810 29.820 1918.130 29.880 ;
        RECT 2422.890 29.820 2423.210 29.880 ;
        RECT 1917.810 29.680 2423.210 29.820 ;
        RECT 1917.810 29.620 1918.130 29.680 ;
        RECT 2422.890 29.620 2423.210 29.680 ;
      LAYER via ;
        RECT 1916.460 586.540 1916.720 586.800 ;
        RECT 1917.840 586.540 1918.100 586.800 ;
        RECT 1917.840 29.620 1918.100 29.880 ;
        RECT 2422.920 29.620 2423.180 29.880 ;
      LAYER met2 ;
        RECT 1914.850 600.170 1915.130 604.000 ;
        RECT 1914.850 600.030 1916.660 600.170 ;
        RECT 1914.850 600.000 1915.130 600.030 ;
        RECT 1916.520 586.830 1916.660 600.030 ;
        RECT 1916.460 586.510 1916.720 586.830 ;
        RECT 1917.840 586.510 1918.100 586.830 ;
        RECT 1917.900 29.910 1918.040 586.510 ;
        RECT 1917.840 29.590 1918.100 29.910 ;
        RECT 2422.920 29.590 2423.180 29.910 ;
        RECT 2422.980 2.400 2423.120 29.590 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1924.710 30.160 1925.030 30.220 ;
        RECT 2440.830 30.160 2441.150 30.220 ;
        RECT 1924.710 30.020 2441.150 30.160 ;
        RECT 1924.710 29.960 1925.030 30.020 ;
        RECT 2440.830 29.960 2441.150 30.020 ;
      LAYER via ;
        RECT 1924.740 29.960 1925.000 30.220 ;
        RECT 2440.860 29.960 2441.120 30.220 ;
      LAYER met2 ;
        RECT 1924.050 600.170 1924.330 604.000 ;
        RECT 1924.050 600.030 1924.940 600.170 ;
        RECT 1924.050 600.000 1924.330 600.030 ;
        RECT 1924.800 30.250 1924.940 600.030 ;
        RECT 1924.740 29.930 1925.000 30.250 ;
        RECT 2440.860 29.930 2441.120 30.250 ;
        RECT 2440.920 2.400 2441.060 29.930 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1934.370 586.740 1934.690 586.800 ;
        RECT 1938.510 586.740 1938.830 586.800 ;
        RECT 1934.370 586.600 1938.830 586.740 ;
        RECT 1934.370 586.540 1934.690 586.600 ;
        RECT 1938.510 586.540 1938.830 586.600 ;
        RECT 1938.510 30.500 1938.830 30.560 ;
        RECT 2458.770 30.500 2459.090 30.560 ;
        RECT 1938.510 30.360 2459.090 30.500 ;
        RECT 1938.510 30.300 1938.830 30.360 ;
        RECT 2458.770 30.300 2459.090 30.360 ;
      LAYER via ;
        RECT 1934.400 586.540 1934.660 586.800 ;
        RECT 1938.540 586.540 1938.800 586.800 ;
        RECT 1938.540 30.300 1938.800 30.560 ;
        RECT 2458.800 30.300 2459.060 30.560 ;
      LAYER met2 ;
        RECT 1932.790 600.170 1933.070 604.000 ;
        RECT 1932.790 600.030 1934.600 600.170 ;
        RECT 1932.790 600.000 1933.070 600.030 ;
        RECT 1934.460 586.830 1934.600 600.030 ;
        RECT 1934.400 586.510 1934.660 586.830 ;
        RECT 1938.540 586.510 1938.800 586.830 ;
        RECT 1938.600 30.590 1938.740 586.510 ;
        RECT 1938.540 30.270 1938.800 30.590 ;
        RECT 2458.800 30.270 2459.060 30.590 ;
        RECT 2458.860 2.400 2459.000 30.270 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1943.570 586.740 1943.890 586.800 ;
        RECT 1945.410 586.740 1945.730 586.800 ;
        RECT 1943.570 586.600 1945.730 586.740 ;
        RECT 1943.570 586.540 1943.890 586.600 ;
        RECT 1945.410 586.540 1945.730 586.600 ;
        RECT 1945.410 34.240 1945.730 34.300 ;
        RECT 2476.710 34.240 2477.030 34.300 ;
        RECT 1945.410 34.100 2477.030 34.240 ;
        RECT 1945.410 34.040 1945.730 34.100 ;
        RECT 2476.710 34.040 2477.030 34.100 ;
      LAYER via ;
        RECT 1943.600 586.540 1943.860 586.800 ;
        RECT 1945.440 586.540 1945.700 586.800 ;
        RECT 1945.440 34.040 1945.700 34.300 ;
        RECT 2476.740 34.040 2477.000 34.300 ;
      LAYER met2 ;
        RECT 1941.990 600.170 1942.270 604.000 ;
        RECT 1941.990 600.030 1943.800 600.170 ;
        RECT 1941.990 600.000 1942.270 600.030 ;
        RECT 1943.660 586.830 1943.800 600.030 ;
        RECT 1943.600 586.510 1943.860 586.830 ;
        RECT 1945.440 586.510 1945.700 586.830 ;
        RECT 1945.500 34.330 1945.640 586.510 ;
        RECT 1945.440 34.010 1945.700 34.330 ;
        RECT 2476.740 34.010 2477.000 34.330 ;
        RECT 2476.800 2.400 2476.940 34.010 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1952.310 33.900 1952.630 33.960 ;
        RECT 2494.650 33.900 2494.970 33.960 ;
        RECT 1952.310 33.760 2494.970 33.900 ;
        RECT 1952.310 33.700 1952.630 33.760 ;
        RECT 2494.650 33.700 2494.970 33.760 ;
      LAYER via ;
        RECT 1952.340 33.700 1952.600 33.960 ;
        RECT 2494.680 33.700 2494.940 33.960 ;
      LAYER met2 ;
        RECT 1951.190 600.170 1951.470 604.000 ;
        RECT 1951.190 600.030 1952.540 600.170 ;
        RECT 1951.190 600.000 1951.470 600.030 ;
        RECT 1952.400 33.990 1952.540 600.030 ;
        RECT 1952.340 33.670 1952.600 33.990 ;
        RECT 2494.680 33.670 2494.940 33.990 ;
        RECT 2494.740 2.400 2494.880 33.670 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1961.970 586.740 1962.290 586.800 ;
        RECT 1966.110 586.740 1966.430 586.800 ;
        RECT 1961.970 586.600 1966.430 586.740 ;
        RECT 1961.970 586.540 1962.290 586.600 ;
        RECT 1966.110 586.540 1966.430 586.600 ;
        RECT 1966.110 33.560 1966.430 33.620 ;
        RECT 2512.130 33.560 2512.450 33.620 ;
        RECT 1966.110 33.420 2512.450 33.560 ;
        RECT 1966.110 33.360 1966.430 33.420 ;
        RECT 2512.130 33.360 2512.450 33.420 ;
      LAYER via ;
        RECT 1962.000 586.540 1962.260 586.800 ;
        RECT 1966.140 586.540 1966.400 586.800 ;
        RECT 1966.140 33.360 1966.400 33.620 ;
        RECT 2512.160 33.360 2512.420 33.620 ;
      LAYER met2 ;
        RECT 1960.390 600.170 1960.670 604.000 ;
        RECT 1960.390 600.030 1962.200 600.170 ;
        RECT 1960.390 600.000 1960.670 600.030 ;
        RECT 1962.060 586.830 1962.200 600.030 ;
        RECT 1962.000 586.510 1962.260 586.830 ;
        RECT 1966.140 586.510 1966.400 586.830 ;
        RECT 1966.200 33.650 1966.340 586.510 ;
        RECT 1966.140 33.330 1966.400 33.650 ;
        RECT 2512.160 33.330 2512.420 33.650 ;
        RECT 2512.220 2.400 2512.360 33.330 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1971.170 586.740 1971.490 586.800 ;
        RECT 1973.010 586.740 1973.330 586.800 ;
        RECT 1971.170 586.600 1973.330 586.740 ;
        RECT 1971.170 586.540 1971.490 586.600 ;
        RECT 1973.010 586.540 1973.330 586.600 ;
        RECT 1973.010 33.220 1973.330 33.280 ;
        RECT 2530.070 33.220 2530.390 33.280 ;
        RECT 1973.010 33.080 2530.390 33.220 ;
        RECT 1973.010 33.020 1973.330 33.080 ;
        RECT 2530.070 33.020 2530.390 33.080 ;
      LAYER via ;
        RECT 1971.200 586.540 1971.460 586.800 ;
        RECT 1973.040 586.540 1973.300 586.800 ;
        RECT 1973.040 33.020 1973.300 33.280 ;
        RECT 2530.100 33.020 2530.360 33.280 ;
      LAYER met2 ;
        RECT 1969.590 600.170 1969.870 604.000 ;
        RECT 1969.590 600.030 1971.400 600.170 ;
        RECT 1969.590 600.000 1969.870 600.030 ;
        RECT 1971.260 586.830 1971.400 600.030 ;
        RECT 1971.200 586.510 1971.460 586.830 ;
        RECT 1973.040 586.510 1973.300 586.830 ;
        RECT 1973.100 33.310 1973.240 586.510 ;
        RECT 1973.040 32.990 1973.300 33.310 ;
        RECT 2530.100 32.990 2530.360 33.310 ;
        RECT 2530.160 2.400 2530.300 32.990 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1979.910 32.880 1980.230 32.940 ;
        RECT 2548.010 32.880 2548.330 32.940 ;
        RECT 1979.910 32.740 2548.330 32.880 ;
        RECT 1979.910 32.680 1980.230 32.740 ;
        RECT 2548.010 32.680 2548.330 32.740 ;
      LAYER via ;
        RECT 1979.940 32.680 1980.200 32.940 ;
        RECT 2548.040 32.680 2548.300 32.940 ;
      LAYER met2 ;
        RECT 1978.790 600.170 1979.070 604.000 ;
        RECT 1978.790 600.030 1980.140 600.170 ;
        RECT 1978.790 600.000 1979.070 600.030 ;
        RECT 1980.000 32.970 1980.140 600.030 ;
        RECT 1979.940 32.650 1980.200 32.970 ;
        RECT 2548.040 32.650 2548.300 32.970 ;
        RECT 2548.100 2.400 2548.240 32.650 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1989.570 586.740 1989.890 586.800 ;
        RECT 1993.710 586.740 1994.030 586.800 ;
        RECT 1989.570 586.600 1994.030 586.740 ;
        RECT 1989.570 586.540 1989.890 586.600 ;
        RECT 1993.710 586.540 1994.030 586.600 ;
        RECT 1993.710 32.540 1994.030 32.600 ;
        RECT 2565.950 32.540 2566.270 32.600 ;
        RECT 1993.710 32.400 2566.270 32.540 ;
        RECT 1993.710 32.340 1994.030 32.400 ;
        RECT 2565.950 32.340 2566.270 32.400 ;
      LAYER via ;
        RECT 1989.600 586.540 1989.860 586.800 ;
        RECT 1993.740 586.540 1994.000 586.800 ;
        RECT 1993.740 32.340 1994.000 32.600 ;
        RECT 2565.980 32.340 2566.240 32.600 ;
      LAYER met2 ;
        RECT 1987.990 600.170 1988.270 604.000 ;
        RECT 1987.990 600.030 1989.800 600.170 ;
        RECT 1987.990 600.000 1988.270 600.030 ;
        RECT 1989.660 586.830 1989.800 600.030 ;
        RECT 1989.600 586.510 1989.860 586.830 ;
        RECT 1993.740 586.510 1994.000 586.830 ;
        RECT 1993.800 32.630 1993.940 586.510 ;
        RECT 1993.740 32.310 1994.000 32.630 ;
        RECT 2565.980 32.310 2566.240 32.630 ;
        RECT 2566.040 2.400 2566.180 32.310 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1998.770 579.940 1999.090 580.000 ;
        RECT 1999.230 579.940 1999.550 580.000 ;
        RECT 1998.770 579.800 1999.550 579.940 ;
        RECT 1998.770 579.740 1999.090 579.800 ;
        RECT 1999.230 579.740 1999.550 579.800 ;
        RECT 1999.690 531.320 2000.010 531.380 ;
        RECT 2000.150 531.320 2000.470 531.380 ;
        RECT 1999.690 531.180 2000.470 531.320 ;
        RECT 1999.690 531.120 2000.010 531.180 ;
        RECT 2000.150 531.120 2000.470 531.180 ;
        RECT 2000.150 496.980 2000.470 497.040 ;
        RECT 1999.780 496.840 2000.470 496.980 ;
        RECT 1999.780 496.700 1999.920 496.840 ;
        RECT 2000.150 496.780 2000.470 496.840 ;
        RECT 1999.690 496.440 2000.010 496.700 ;
        RECT 1999.230 448.700 1999.550 448.760 ;
        RECT 2000.150 448.700 2000.470 448.760 ;
        RECT 1999.230 448.560 2000.470 448.700 ;
        RECT 1999.230 448.500 1999.550 448.560 ;
        RECT 2000.150 448.500 2000.470 448.560 ;
        RECT 1998.770 434.760 1999.090 434.820 ;
        RECT 1999.690 434.760 2000.010 434.820 ;
        RECT 1998.770 434.620 2000.010 434.760 ;
        RECT 1998.770 434.560 1999.090 434.620 ;
        RECT 1999.690 434.560 2000.010 434.620 ;
        RECT 1998.770 386.480 1999.090 386.540 ;
        RECT 2000.150 386.480 2000.470 386.540 ;
        RECT 1998.770 386.340 2000.470 386.480 ;
        RECT 1998.770 386.280 1999.090 386.340 ;
        RECT 2000.150 386.280 2000.470 386.340 ;
        RECT 1998.770 379.340 1999.090 379.400 ;
        RECT 2000.150 379.340 2000.470 379.400 ;
        RECT 1998.770 379.200 2000.470 379.340 ;
        RECT 1998.770 379.140 1999.090 379.200 ;
        RECT 2000.150 379.140 2000.470 379.200 ;
        RECT 1999.690 234.840 2000.010 234.900 ;
        RECT 2000.150 234.840 2000.470 234.900 ;
        RECT 1999.690 234.700 2000.470 234.840 ;
        RECT 1999.690 234.640 2000.010 234.700 ;
        RECT 2000.150 234.640 2000.470 234.700 ;
        RECT 1999.230 186.560 1999.550 186.620 ;
        RECT 2000.150 186.560 2000.470 186.620 ;
        RECT 1999.230 186.420 2000.470 186.560 ;
        RECT 1999.230 186.360 1999.550 186.420 ;
        RECT 2000.150 186.360 2000.470 186.420 ;
        RECT 1999.230 32.200 1999.550 32.260 ;
        RECT 2583.890 32.200 2584.210 32.260 ;
        RECT 1999.230 32.060 2584.210 32.200 ;
        RECT 1999.230 32.000 1999.550 32.060 ;
        RECT 2583.890 32.000 2584.210 32.060 ;
      LAYER via ;
        RECT 1998.800 579.740 1999.060 580.000 ;
        RECT 1999.260 579.740 1999.520 580.000 ;
        RECT 1999.720 531.120 1999.980 531.380 ;
        RECT 2000.180 531.120 2000.440 531.380 ;
        RECT 2000.180 496.780 2000.440 497.040 ;
        RECT 1999.720 496.440 1999.980 496.700 ;
        RECT 1999.260 448.500 1999.520 448.760 ;
        RECT 2000.180 448.500 2000.440 448.760 ;
        RECT 1998.800 434.560 1999.060 434.820 ;
        RECT 1999.720 434.560 1999.980 434.820 ;
        RECT 1998.800 386.280 1999.060 386.540 ;
        RECT 2000.180 386.280 2000.440 386.540 ;
        RECT 1998.800 379.140 1999.060 379.400 ;
        RECT 2000.180 379.140 2000.440 379.400 ;
        RECT 1999.720 234.640 1999.980 234.900 ;
        RECT 2000.180 234.640 2000.440 234.900 ;
        RECT 1999.260 186.360 1999.520 186.620 ;
        RECT 2000.180 186.360 2000.440 186.620 ;
        RECT 1999.260 32.000 1999.520 32.260 ;
        RECT 2583.920 32.000 2584.180 32.260 ;
      LAYER met2 ;
        RECT 1997.190 600.170 1997.470 604.000 ;
        RECT 1997.190 600.030 1999.000 600.170 ;
        RECT 1997.190 600.000 1997.470 600.030 ;
        RECT 1998.860 580.030 1999.000 600.030 ;
        RECT 1998.800 579.710 1999.060 580.030 ;
        RECT 1999.260 579.710 1999.520 580.030 ;
        RECT 1999.320 545.090 1999.460 579.710 ;
        RECT 1999.320 544.950 1999.920 545.090 ;
        RECT 1999.780 531.410 1999.920 544.950 ;
        RECT 1999.720 531.090 1999.980 531.410 ;
        RECT 2000.180 531.090 2000.440 531.410 ;
        RECT 2000.240 497.070 2000.380 531.090 ;
        RECT 2000.180 496.750 2000.440 497.070 ;
        RECT 1999.720 496.410 1999.980 496.730 ;
        RECT 1999.780 483.210 1999.920 496.410 ;
        RECT 1999.780 483.070 2000.380 483.210 ;
        RECT 2000.240 448.790 2000.380 483.070 ;
        RECT 1999.260 448.530 1999.520 448.790 ;
        RECT 1999.260 448.470 1999.920 448.530 ;
        RECT 2000.180 448.470 2000.440 448.790 ;
        RECT 1999.320 448.390 1999.920 448.470 ;
        RECT 1999.780 434.850 1999.920 448.390 ;
        RECT 1998.800 434.530 1999.060 434.850 ;
        RECT 1999.720 434.530 1999.980 434.850 ;
        RECT 1998.860 386.570 1999.000 434.530 ;
        RECT 1998.800 386.250 1999.060 386.570 ;
        RECT 2000.180 386.250 2000.440 386.570 ;
        RECT 2000.240 379.430 2000.380 386.250 ;
        RECT 1998.800 379.110 1999.060 379.430 ;
        RECT 2000.180 379.110 2000.440 379.430 ;
        RECT 1998.860 351.290 1999.000 379.110 ;
        RECT 1998.860 351.150 1999.920 351.290 ;
        RECT 1999.780 303.690 1999.920 351.150 ;
        RECT 1999.780 303.550 2000.380 303.690 ;
        RECT 2000.240 234.930 2000.380 303.550 ;
        RECT 1999.720 234.610 1999.980 234.930 ;
        RECT 2000.180 234.610 2000.440 234.930 ;
        RECT 1999.780 234.330 1999.920 234.610 ;
        RECT 1999.320 234.190 1999.920 234.330 ;
        RECT 1999.320 186.650 1999.460 234.190 ;
        RECT 1999.260 186.330 1999.520 186.650 ;
        RECT 2000.180 186.330 2000.440 186.650 ;
        RECT 2000.240 158.850 2000.380 186.330 ;
        RECT 1999.320 158.710 2000.380 158.850 ;
        RECT 1999.320 158.170 1999.460 158.710 ;
        RECT 1999.320 158.030 1999.920 158.170 ;
        RECT 1999.780 62.290 1999.920 158.030 ;
        RECT 1999.320 62.150 1999.920 62.290 ;
        RECT 1999.320 32.290 1999.460 62.150 ;
        RECT 1999.260 31.970 1999.520 32.290 ;
        RECT 2583.920 31.970 2584.180 32.290 ;
        RECT 2583.980 2.400 2584.120 31.970 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1083.830 552.400 1084.150 552.460 ;
        RECT 1087.970 552.400 1088.290 552.460 ;
        RECT 1083.830 552.260 1088.290 552.400 ;
        RECT 1083.830 552.200 1084.150 552.260 ;
        RECT 1087.970 552.200 1088.290 552.260 ;
        RECT 817.490 26.080 817.810 26.140 ;
        RECT 1083.830 26.080 1084.150 26.140 ;
        RECT 817.490 25.940 1084.150 26.080 ;
        RECT 817.490 25.880 817.810 25.940 ;
        RECT 1083.830 25.880 1084.150 25.940 ;
      LAYER via ;
        RECT 1083.860 552.200 1084.120 552.460 ;
        RECT 1088.000 552.200 1088.260 552.460 ;
        RECT 817.520 25.880 817.780 26.140 ;
        RECT 1083.860 25.880 1084.120 26.140 ;
      LAYER met2 ;
        RECT 1089.610 600.170 1089.890 604.000 ;
        RECT 1088.060 600.030 1089.890 600.170 ;
        RECT 1088.060 552.490 1088.200 600.030 ;
        RECT 1089.610 600.000 1089.890 600.030 ;
        RECT 1083.860 552.170 1084.120 552.490 ;
        RECT 1088.000 552.170 1088.260 552.490 ;
        RECT 1083.920 26.170 1084.060 552.170 ;
        RECT 817.520 25.850 817.780 26.170 ;
        RECT 1083.860 25.850 1084.120 26.170 ;
        RECT 817.580 2.400 817.720 25.850 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2007.050 31.520 2007.370 31.580 ;
        RECT 2601.370 31.520 2601.690 31.580 ;
        RECT 2007.050 31.380 2601.690 31.520 ;
        RECT 2007.050 31.320 2007.370 31.380 ;
        RECT 2601.370 31.320 2601.690 31.380 ;
      LAYER via ;
        RECT 2007.080 31.320 2007.340 31.580 ;
        RECT 2601.400 31.320 2601.660 31.580 ;
      LAYER met2 ;
        RECT 2006.390 600.170 2006.670 604.000 ;
        RECT 2006.390 600.030 2007.280 600.170 ;
        RECT 2006.390 600.000 2006.670 600.030 ;
        RECT 2007.140 31.610 2007.280 600.030 ;
        RECT 2007.080 31.290 2007.340 31.610 ;
        RECT 2601.400 31.290 2601.660 31.610 ;
        RECT 2601.460 2.400 2601.600 31.290 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2017.170 586.740 2017.490 586.800 ;
        RECT 2021.310 586.740 2021.630 586.800 ;
        RECT 2017.170 586.600 2021.630 586.740 ;
        RECT 2017.170 586.540 2017.490 586.600 ;
        RECT 2021.310 586.540 2021.630 586.600 ;
        RECT 2021.310 31.860 2021.630 31.920 ;
        RECT 2619.310 31.860 2619.630 31.920 ;
        RECT 2021.310 31.720 2619.630 31.860 ;
        RECT 2021.310 31.660 2021.630 31.720 ;
        RECT 2619.310 31.660 2619.630 31.720 ;
      LAYER via ;
        RECT 2017.200 586.540 2017.460 586.800 ;
        RECT 2021.340 586.540 2021.600 586.800 ;
        RECT 2021.340 31.660 2021.600 31.920 ;
        RECT 2619.340 31.660 2619.600 31.920 ;
      LAYER met2 ;
        RECT 2015.590 600.170 2015.870 604.000 ;
        RECT 2015.590 600.030 2017.400 600.170 ;
        RECT 2015.590 600.000 2015.870 600.030 ;
        RECT 2017.260 586.830 2017.400 600.030 ;
        RECT 2017.200 586.510 2017.460 586.830 ;
        RECT 2021.340 586.510 2021.600 586.830 ;
        RECT 2021.400 31.950 2021.540 586.510 ;
        RECT 2021.340 31.630 2021.600 31.950 ;
        RECT 2619.340 31.630 2619.600 31.950 ;
        RECT 2619.400 2.400 2619.540 31.630 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2025.450 579.940 2025.770 580.000 ;
        RECT 2025.910 579.940 2026.230 580.000 ;
        RECT 2025.450 579.800 2026.230 579.940 ;
        RECT 2025.450 579.740 2025.770 579.800 ;
        RECT 2025.910 579.740 2026.230 579.800 ;
        RECT 2027.290 531.320 2027.610 531.380 ;
        RECT 2027.750 531.320 2028.070 531.380 ;
        RECT 2027.290 531.180 2028.070 531.320 ;
        RECT 2027.290 531.120 2027.610 531.180 ;
        RECT 2027.750 531.120 2028.070 531.180 ;
        RECT 2027.750 496.980 2028.070 497.040 ;
        RECT 2027.380 496.840 2028.070 496.980 ;
        RECT 2027.380 496.700 2027.520 496.840 ;
        RECT 2027.750 496.780 2028.070 496.840 ;
        RECT 2027.290 496.440 2027.610 496.700 ;
        RECT 2026.830 448.360 2027.150 448.420 ;
        RECT 2027.750 448.360 2028.070 448.420 ;
        RECT 2026.830 448.220 2028.070 448.360 ;
        RECT 2026.830 448.160 2027.150 448.220 ;
        RECT 2027.750 448.160 2028.070 448.220 ;
        RECT 2026.830 403.820 2027.150 403.880 ;
        RECT 2028.670 403.820 2028.990 403.880 ;
        RECT 2026.830 403.680 2028.990 403.820 ;
        RECT 2026.830 403.620 2027.150 403.680 ;
        RECT 2028.670 403.620 2028.990 403.680 ;
        RECT 2025.910 379.340 2026.230 379.400 ;
        RECT 2026.830 379.340 2027.150 379.400 ;
        RECT 2025.910 379.200 2027.150 379.340 ;
        RECT 2025.910 379.140 2026.230 379.200 ;
        RECT 2026.830 379.140 2027.150 379.200 ;
        RECT 2025.910 331.400 2026.230 331.460 ;
        RECT 2027.290 331.400 2027.610 331.460 ;
        RECT 2025.910 331.260 2027.610 331.400 ;
        RECT 2025.910 331.200 2026.230 331.260 ;
        RECT 2027.290 331.200 2027.610 331.260 ;
        RECT 2027.290 303.860 2027.610 303.920 ;
        RECT 2026.920 303.720 2027.610 303.860 ;
        RECT 2026.920 303.580 2027.060 303.720 ;
        RECT 2027.290 303.660 2027.610 303.720 ;
        RECT 2026.830 303.320 2027.150 303.580 ;
        RECT 2025.910 282.780 2026.230 282.840 ;
        RECT 2026.830 282.780 2027.150 282.840 ;
        RECT 2025.910 282.640 2027.150 282.780 ;
        RECT 2025.910 282.580 2026.230 282.640 ;
        RECT 2026.830 282.580 2027.150 282.640 ;
        RECT 2026.830 186.020 2027.150 186.280 ;
        RECT 2026.920 185.600 2027.060 186.020 ;
        RECT 2026.830 185.340 2027.150 185.600 ;
        RECT 2026.830 138.280 2027.150 138.340 ;
        RECT 2027.750 138.280 2028.070 138.340 ;
        RECT 2026.830 138.140 2028.070 138.280 ;
        RECT 2026.830 138.080 2027.150 138.140 ;
        RECT 2027.750 138.080 2028.070 138.140 ;
        RECT 2027.750 110.740 2028.070 110.800 ;
        RECT 2027.380 110.600 2028.070 110.740 ;
        RECT 2027.380 110.460 2027.520 110.600 ;
        RECT 2027.750 110.540 2028.070 110.600 ;
        RECT 2027.290 110.200 2027.610 110.460 ;
        RECT 2025.910 96.460 2026.230 96.520 ;
        RECT 2027.290 96.460 2027.610 96.520 ;
        RECT 2025.910 96.320 2027.610 96.460 ;
        RECT 2025.910 96.260 2026.230 96.320 ;
        RECT 2027.290 96.260 2027.610 96.320 ;
        RECT 2025.910 48.520 2026.230 48.580 ;
        RECT 2026.830 48.520 2027.150 48.580 ;
        RECT 2025.910 48.380 2027.150 48.520 ;
        RECT 2025.910 48.320 2026.230 48.380 ;
        RECT 2026.830 48.320 2027.150 48.380 ;
        RECT 2026.830 31.180 2027.150 31.240 ;
        RECT 2637.250 31.180 2637.570 31.240 ;
        RECT 2026.830 31.040 2637.570 31.180 ;
        RECT 2026.830 30.980 2027.150 31.040 ;
        RECT 2637.250 30.980 2637.570 31.040 ;
      LAYER via ;
        RECT 2025.480 579.740 2025.740 580.000 ;
        RECT 2025.940 579.740 2026.200 580.000 ;
        RECT 2027.320 531.120 2027.580 531.380 ;
        RECT 2027.780 531.120 2028.040 531.380 ;
        RECT 2027.780 496.780 2028.040 497.040 ;
        RECT 2027.320 496.440 2027.580 496.700 ;
        RECT 2026.860 448.160 2027.120 448.420 ;
        RECT 2027.780 448.160 2028.040 448.420 ;
        RECT 2026.860 403.620 2027.120 403.880 ;
        RECT 2028.700 403.620 2028.960 403.880 ;
        RECT 2025.940 379.140 2026.200 379.400 ;
        RECT 2026.860 379.140 2027.120 379.400 ;
        RECT 2025.940 331.200 2026.200 331.460 ;
        RECT 2027.320 331.200 2027.580 331.460 ;
        RECT 2027.320 303.660 2027.580 303.920 ;
        RECT 2026.860 303.320 2027.120 303.580 ;
        RECT 2025.940 282.580 2026.200 282.840 ;
        RECT 2026.860 282.580 2027.120 282.840 ;
        RECT 2026.860 186.020 2027.120 186.280 ;
        RECT 2026.860 185.340 2027.120 185.600 ;
        RECT 2026.860 138.080 2027.120 138.340 ;
        RECT 2027.780 138.080 2028.040 138.340 ;
        RECT 2027.780 110.540 2028.040 110.800 ;
        RECT 2027.320 110.200 2027.580 110.460 ;
        RECT 2025.940 96.260 2026.200 96.520 ;
        RECT 2027.320 96.260 2027.580 96.520 ;
        RECT 2025.940 48.320 2026.200 48.580 ;
        RECT 2026.860 48.320 2027.120 48.580 ;
        RECT 2026.860 30.980 2027.120 31.240 ;
        RECT 2637.280 30.980 2637.540 31.240 ;
      LAYER met2 ;
        RECT 2024.790 600.170 2025.070 604.000 ;
        RECT 2024.790 600.030 2025.680 600.170 ;
        RECT 2024.790 600.000 2025.070 600.030 ;
        RECT 2025.540 580.030 2025.680 600.030 ;
        RECT 2025.480 579.710 2025.740 580.030 ;
        RECT 2025.940 579.710 2026.200 580.030 ;
        RECT 2026.000 545.090 2026.140 579.710 ;
        RECT 2026.000 544.950 2027.060 545.090 ;
        RECT 2026.920 544.410 2027.060 544.950 ;
        RECT 2026.920 544.270 2027.520 544.410 ;
        RECT 2027.380 531.410 2027.520 544.270 ;
        RECT 2027.320 531.090 2027.580 531.410 ;
        RECT 2027.780 531.090 2028.040 531.410 ;
        RECT 2027.840 497.070 2027.980 531.090 ;
        RECT 2027.780 496.750 2028.040 497.070 ;
        RECT 2027.320 496.410 2027.580 496.730 ;
        RECT 2027.380 483.210 2027.520 496.410 ;
        RECT 2027.380 483.070 2027.980 483.210 ;
        RECT 2027.840 448.450 2027.980 483.070 ;
        RECT 2026.860 448.130 2027.120 448.450 ;
        RECT 2027.780 448.130 2028.040 448.450 ;
        RECT 2026.920 403.910 2027.060 448.130 ;
        RECT 2026.860 403.590 2027.120 403.910 ;
        RECT 2028.700 403.590 2028.960 403.910 ;
        RECT 2028.760 379.965 2028.900 403.590 ;
        RECT 2027.310 379.850 2027.590 379.965 ;
        RECT 2026.920 379.710 2027.590 379.850 ;
        RECT 2026.920 379.430 2027.060 379.710 ;
        RECT 2027.310 379.595 2027.590 379.710 ;
        RECT 2028.690 379.595 2028.970 379.965 ;
        RECT 2025.940 379.110 2026.200 379.430 ;
        RECT 2026.860 379.110 2027.120 379.430 ;
        RECT 2026.000 331.490 2026.140 379.110 ;
        RECT 2025.940 331.170 2026.200 331.490 ;
        RECT 2027.320 331.170 2027.580 331.490 ;
        RECT 2027.380 303.950 2027.520 331.170 ;
        RECT 2027.320 303.630 2027.580 303.950 ;
        RECT 2026.860 303.290 2027.120 303.610 ;
        RECT 2026.920 282.870 2027.060 303.290 ;
        RECT 2025.940 282.550 2026.200 282.870 ;
        RECT 2026.860 282.550 2027.120 282.870 ;
        RECT 2026.000 254.050 2026.140 282.550 ;
        RECT 2026.000 253.910 2027.060 254.050 ;
        RECT 2026.920 186.310 2027.060 253.910 ;
        RECT 2026.860 185.990 2027.120 186.310 ;
        RECT 2026.860 185.310 2027.120 185.630 ;
        RECT 2026.920 138.370 2027.060 185.310 ;
        RECT 2026.860 138.050 2027.120 138.370 ;
        RECT 2027.780 138.050 2028.040 138.370 ;
        RECT 2027.840 110.830 2027.980 138.050 ;
        RECT 2027.780 110.510 2028.040 110.830 ;
        RECT 2027.320 110.170 2027.580 110.490 ;
        RECT 2027.380 96.550 2027.520 110.170 ;
        RECT 2025.940 96.230 2026.200 96.550 ;
        RECT 2027.320 96.230 2027.580 96.550 ;
        RECT 2026.000 48.610 2026.140 96.230 ;
        RECT 2025.940 48.290 2026.200 48.610 ;
        RECT 2026.860 48.290 2027.120 48.610 ;
        RECT 2026.920 31.270 2027.060 48.290 ;
        RECT 2026.860 30.950 2027.120 31.270 ;
        RECT 2637.280 30.950 2637.540 31.270 ;
        RECT 2637.340 2.400 2637.480 30.950 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
      LAYER via2 ;
        RECT 2027.310 379.640 2027.590 379.920 ;
        RECT 2028.690 379.640 2028.970 379.920 ;
      LAYER met3 ;
        RECT 2027.285 379.930 2027.615 379.945 ;
        RECT 2028.665 379.930 2028.995 379.945 ;
        RECT 2027.285 379.630 2028.995 379.930 ;
        RECT 2027.285 379.615 2027.615 379.630 ;
        RECT 2028.665 379.615 2028.995 379.630 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2034.650 30.840 2034.970 30.900 ;
        RECT 2655.190 30.840 2655.510 30.900 ;
        RECT 2034.650 30.700 2655.510 30.840 ;
        RECT 2034.650 30.640 2034.970 30.700 ;
        RECT 2655.190 30.640 2655.510 30.700 ;
      LAYER via ;
        RECT 2034.680 30.640 2034.940 30.900 ;
        RECT 2655.220 30.640 2655.480 30.900 ;
      LAYER met2 ;
        RECT 2033.990 600.170 2034.270 604.000 ;
        RECT 2033.990 600.030 2034.880 600.170 ;
        RECT 2033.990 600.000 2034.270 600.030 ;
        RECT 2034.740 30.930 2034.880 600.030 ;
        RECT 2034.680 30.610 2034.940 30.930 ;
        RECT 2655.220 30.610 2655.480 30.930 ;
        RECT 2655.280 2.400 2655.420 30.610 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2044.770 586.740 2045.090 586.800 ;
        RECT 2048.910 586.740 2049.230 586.800 ;
        RECT 2044.770 586.600 2049.230 586.740 ;
        RECT 2044.770 586.540 2045.090 586.600 ;
        RECT 2048.910 586.540 2049.230 586.600 ;
        RECT 2048.910 41.380 2049.230 41.440 ;
        RECT 2672.670 41.380 2672.990 41.440 ;
        RECT 2048.910 41.240 2672.990 41.380 ;
        RECT 2048.910 41.180 2049.230 41.240 ;
        RECT 2672.670 41.180 2672.990 41.240 ;
      LAYER via ;
        RECT 2044.800 586.540 2045.060 586.800 ;
        RECT 2048.940 586.540 2049.200 586.800 ;
        RECT 2048.940 41.180 2049.200 41.440 ;
        RECT 2672.700 41.180 2672.960 41.440 ;
      LAYER met2 ;
        RECT 2043.190 600.170 2043.470 604.000 ;
        RECT 2043.190 600.030 2045.000 600.170 ;
        RECT 2043.190 600.000 2043.470 600.030 ;
        RECT 2044.860 586.830 2045.000 600.030 ;
        RECT 2044.800 586.510 2045.060 586.830 ;
        RECT 2048.940 586.510 2049.200 586.830 ;
        RECT 2049.000 41.470 2049.140 586.510 ;
        RECT 2048.940 41.150 2049.200 41.470 ;
        RECT 2672.700 41.150 2672.960 41.470 ;
        RECT 2672.760 2.400 2672.900 41.150 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2052.590 579.940 2052.910 580.000 ;
        RECT 2053.510 579.940 2053.830 580.000 ;
        RECT 2052.590 579.800 2053.830 579.940 ;
        RECT 2052.590 579.740 2052.910 579.800 ;
        RECT 2053.510 579.740 2053.830 579.800 ;
        RECT 2054.430 497.120 2054.750 497.380 ;
        RECT 2054.520 496.700 2054.660 497.120 ;
        RECT 2054.430 496.440 2054.750 496.700 ;
        RECT 2054.890 483.040 2055.210 483.100 ;
        RECT 2056.270 483.040 2056.590 483.100 ;
        RECT 2054.890 482.900 2056.590 483.040 ;
        RECT 2054.890 482.840 2055.210 482.900 ;
        RECT 2056.270 482.840 2056.590 482.900 ;
        RECT 2053.510 434.760 2053.830 434.820 ;
        RECT 2054.430 434.760 2054.750 434.820 ;
        RECT 2053.510 434.620 2054.750 434.760 ;
        RECT 2053.510 434.560 2053.830 434.620 ;
        RECT 2054.430 434.560 2054.750 434.620 ;
        RECT 2053.510 386.480 2053.830 386.540 ;
        RECT 2053.970 386.480 2054.290 386.540 ;
        RECT 2053.510 386.340 2054.290 386.480 ;
        RECT 2053.510 386.280 2053.830 386.340 ;
        RECT 2053.970 386.280 2054.290 386.340 ;
        RECT 2052.590 324.260 2052.910 324.320 ;
        RECT 2053.510 324.260 2053.830 324.320 ;
        RECT 2052.590 324.120 2053.830 324.260 ;
        RECT 2052.590 324.060 2052.910 324.120 ;
        RECT 2053.510 324.060 2053.830 324.120 ;
        RECT 2052.590 276.320 2052.910 276.380 ;
        RECT 2054.430 276.320 2054.750 276.380 ;
        RECT 2052.590 276.180 2054.750 276.320 ;
        RECT 2052.590 276.120 2052.910 276.180 ;
        RECT 2054.430 276.120 2054.750 276.180 ;
        RECT 2053.970 158.820 2054.290 159.080 ;
        RECT 2054.060 158.340 2054.200 158.820 ;
        RECT 2054.430 158.340 2054.750 158.400 ;
        RECT 2054.060 158.200 2054.750 158.340 ;
        RECT 2054.430 158.140 2054.750 158.200 ;
        RECT 2054.430 41.040 2054.750 41.100 ;
        RECT 2690.610 41.040 2690.930 41.100 ;
        RECT 2054.430 40.900 2690.930 41.040 ;
        RECT 2054.430 40.840 2054.750 40.900 ;
        RECT 2690.610 40.840 2690.930 40.900 ;
      LAYER via ;
        RECT 2052.620 579.740 2052.880 580.000 ;
        RECT 2053.540 579.740 2053.800 580.000 ;
        RECT 2054.460 497.120 2054.720 497.380 ;
        RECT 2054.460 496.440 2054.720 496.700 ;
        RECT 2054.920 482.840 2055.180 483.100 ;
        RECT 2056.300 482.840 2056.560 483.100 ;
        RECT 2053.540 434.560 2053.800 434.820 ;
        RECT 2054.460 434.560 2054.720 434.820 ;
        RECT 2053.540 386.280 2053.800 386.540 ;
        RECT 2054.000 386.280 2054.260 386.540 ;
        RECT 2052.620 324.060 2052.880 324.320 ;
        RECT 2053.540 324.060 2053.800 324.320 ;
        RECT 2052.620 276.120 2052.880 276.380 ;
        RECT 2054.460 276.120 2054.720 276.380 ;
        RECT 2054.000 158.820 2054.260 159.080 ;
        RECT 2054.460 158.140 2054.720 158.400 ;
        RECT 2054.460 40.840 2054.720 41.100 ;
        RECT 2690.640 40.840 2690.900 41.100 ;
      LAYER met2 ;
        RECT 2051.930 600.170 2052.210 604.000 ;
        RECT 2051.930 600.030 2052.820 600.170 ;
        RECT 2051.930 600.000 2052.210 600.030 ;
        RECT 2052.680 580.030 2052.820 600.030 ;
        RECT 2052.620 579.710 2052.880 580.030 ;
        RECT 2053.540 579.710 2053.800 580.030 ;
        RECT 2053.600 545.090 2053.740 579.710 ;
        RECT 2053.600 544.950 2054.660 545.090 ;
        RECT 2054.520 497.410 2054.660 544.950 ;
        RECT 2054.460 497.090 2054.720 497.410 ;
        RECT 2054.460 496.410 2054.720 496.730 ;
        RECT 2054.520 483.210 2054.660 496.410 ;
        RECT 2054.520 483.130 2055.120 483.210 ;
        RECT 2054.520 483.070 2055.180 483.130 ;
        RECT 2054.920 482.810 2055.180 483.070 ;
        RECT 2056.300 482.810 2056.560 483.130 ;
        RECT 2054.980 482.655 2055.120 482.810 ;
        RECT 2056.360 435.045 2056.500 482.810 ;
        RECT 2054.910 434.930 2055.190 435.045 ;
        RECT 2054.520 434.850 2055.190 434.930 ;
        RECT 2053.540 434.530 2053.800 434.850 ;
        RECT 2054.460 434.790 2055.190 434.850 ;
        RECT 2054.460 434.530 2054.720 434.790 ;
        RECT 2054.910 434.675 2055.190 434.790 ;
        RECT 2056.290 434.675 2056.570 435.045 ;
        RECT 2053.600 386.570 2053.740 434.530 ;
        RECT 2053.540 386.250 2053.800 386.570 ;
        RECT 2054.000 386.250 2054.260 386.570 ;
        RECT 2054.060 331.570 2054.200 386.250 ;
        RECT 2053.600 331.430 2054.200 331.570 ;
        RECT 2053.600 324.350 2053.740 331.430 ;
        RECT 2052.620 324.030 2052.880 324.350 ;
        RECT 2053.540 324.030 2053.800 324.350 ;
        RECT 2052.680 276.410 2052.820 324.030 ;
        RECT 2052.620 276.090 2052.880 276.410 ;
        RECT 2054.460 276.090 2054.720 276.410 ;
        RECT 2054.520 241.130 2054.660 276.090 ;
        RECT 2053.600 240.990 2054.660 241.130 ;
        RECT 2053.600 234.445 2053.740 240.990 ;
        RECT 2053.530 234.075 2053.810 234.445 ;
        RECT 2053.990 233.395 2054.270 233.765 ;
        RECT 2054.060 159.110 2054.200 233.395 ;
        RECT 2054.000 158.790 2054.260 159.110 ;
        RECT 2054.460 158.110 2054.720 158.430 ;
        RECT 2054.520 110.570 2054.660 158.110 ;
        RECT 2054.520 110.430 2055.120 110.570 ;
        RECT 2054.980 62.290 2055.120 110.430 ;
        RECT 2054.520 62.150 2055.120 62.290 ;
        RECT 2054.520 41.130 2054.660 62.150 ;
        RECT 2054.460 40.810 2054.720 41.130 ;
        RECT 2690.640 40.810 2690.900 41.130 ;
        RECT 2690.700 2.400 2690.840 40.810 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
      LAYER via2 ;
        RECT 2054.910 434.720 2055.190 435.000 ;
        RECT 2056.290 434.720 2056.570 435.000 ;
        RECT 2053.530 234.120 2053.810 234.400 ;
        RECT 2053.990 233.440 2054.270 233.720 ;
      LAYER met3 ;
        RECT 2054.885 435.010 2055.215 435.025 ;
        RECT 2056.265 435.010 2056.595 435.025 ;
        RECT 2054.885 434.710 2056.595 435.010 ;
        RECT 2054.885 434.695 2055.215 434.710 ;
        RECT 2056.265 434.695 2056.595 434.710 ;
        RECT 2053.505 234.410 2053.835 234.425 ;
        RECT 2052.830 234.110 2053.835 234.410 ;
        RECT 2052.830 233.730 2053.130 234.110 ;
        RECT 2053.505 234.095 2053.835 234.110 ;
        RECT 2053.965 233.730 2054.295 233.745 ;
        RECT 2052.830 233.430 2054.295 233.730 ;
        RECT 2053.965 233.415 2054.295 233.430 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2062.250 40.700 2062.570 40.760 ;
        RECT 2708.550 40.700 2708.870 40.760 ;
        RECT 2062.250 40.560 2708.870 40.700 ;
        RECT 2062.250 40.500 2062.570 40.560 ;
        RECT 2708.550 40.500 2708.870 40.560 ;
      LAYER via ;
        RECT 2062.280 40.500 2062.540 40.760 ;
        RECT 2708.580 40.500 2708.840 40.760 ;
      LAYER met2 ;
        RECT 2061.130 600.170 2061.410 604.000 ;
        RECT 2061.130 600.030 2062.480 600.170 ;
        RECT 2061.130 600.000 2061.410 600.030 ;
        RECT 2062.340 40.790 2062.480 600.030 ;
        RECT 2062.280 40.470 2062.540 40.790 ;
        RECT 2708.580 40.470 2708.840 40.790 ;
        RECT 2708.640 2.400 2708.780 40.470 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2071.910 586.740 2072.230 586.800 ;
        RECT 2076.050 586.740 2076.370 586.800 ;
        RECT 2071.910 586.600 2076.370 586.740 ;
        RECT 2071.910 586.540 2072.230 586.600 ;
        RECT 2076.050 586.540 2076.370 586.600 ;
        RECT 2076.050 40.360 2076.370 40.420 ;
        RECT 2726.490 40.360 2726.810 40.420 ;
        RECT 2076.050 40.220 2726.810 40.360 ;
        RECT 2076.050 40.160 2076.370 40.220 ;
        RECT 2726.490 40.160 2726.810 40.220 ;
      LAYER via ;
        RECT 2071.940 586.540 2072.200 586.800 ;
        RECT 2076.080 586.540 2076.340 586.800 ;
        RECT 2076.080 40.160 2076.340 40.420 ;
        RECT 2726.520 40.160 2726.780 40.420 ;
      LAYER met2 ;
        RECT 2070.330 600.170 2070.610 604.000 ;
        RECT 2070.330 600.030 2072.140 600.170 ;
        RECT 2070.330 600.000 2070.610 600.030 ;
        RECT 2072.000 586.830 2072.140 600.030 ;
        RECT 2071.940 586.510 2072.200 586.830 ;
        RECT 2076.080 586.510 2076.340 586.830 ;
        RECT 2076.140 40.450 2076.280 586.510 ;
        RECT 2076.080 40.130 2076.340 40.450 ;
        RECT 2726.520 40.130 2726.780 40.450 ;
        RECT 2726.580 2.400 2726.720 40.130 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2082.490 496.780 2082.810 497.040 ;
        RECT 2082.580 496.640 2082.720 496.780 ;
        RECT 2082.950 496.640 2083.270 496.700 ;
        RECT 2082.580 496.500 2083.270 496.640 ;
        RECT 2082.950 496.440 2083.270 496.500 ;
        RECT 2082.490 421.160 2082.810 421.220 ;
        RECT 2082.950 421.160 2083.270 421.220 ;
        RECT 2082.490 421.020 2083.270 421.160 ;
        RECT 2082.490 420.960 2082.810 421.020 ;
        RECT 2082.950 420.960 2083.270 421.020 ;
        RECT 2081.570 372.880 2081.890 372.940 ;
        RECT 2082.030 372.880 2082.350 372.940 ;
        RECT 2081.570 372.740 2082.350 372.880 ;
        RECT 2081.570 372.680 2081.890 372.740 ;
        RECT 2082.030 372.680 2082.350 372.740 ;
        RECT 2080.650 324.600 2080.970 324.660 ;
        RECT 2082.490 324.600 2082.810 324.660 ;
        RECT 2080.650 324.460 2082.810 324.600 ;
        RECT 2080.650 324.400 2080.970 324.460 ;
        RECT 2082.490 324.400 2082.810 324.460 ;
        RECT 2082.490 303.860 2082.810 303.920 ;
        RECT 2082.120 303.720 2082.810 303.860 ;
        RECT 2082.120 303.580 2082.260 303.720 ;
        RECT 2082.490 303.660 2082.810 303.720 ;
        RECT 2082.030 303.320 2082.350 303.580 ;
        RECT 2081.110 275.980 2081.430 276.040 ;
        RECT 2082.030 275.980 2082.350 276.040 ;
        RECT 2081.110 275.840 2082.350 275.980 ;
        RECT 2081.110 275.780 2081.430 275.840 ;
        RECT 2082.030 275.780 2082.350 275.840 ;
        RECT 2081.110 228.040 2081.430 228.100 ;
        RECT 2082.490 228.040 2082.810 228.100 ;
        RECT 2081.110 227.900 2082.810 228.040 ;
        RECT 2081.110 227.840 2081.430 227.900 ;
        RECT 2082.490 227.840 2082.810 227.900 ;
        RECT 2082.490 144.400 2082.810 144.460 ;
        RECT 2083.870 144.400 2084.190 144.460 ;
        RECT 2082.490 144.260 2084.190 144.400 ;
        RECT 2082.490 144.200 2082.810 144.260 ;
        RECT 2083.870 144.200 2084.190 144.260 ;
        RECT 2082.490 110.740 2082.810 110.800 ;
        RECT 2082.950 110.740 2083.270 110.800 ;
        RECT 2082.490 110.600 2083.270 110.740 ;
        RECT 2082.490 110.540 2082.810 110.600 ;
        RECT 2082.950 110.540 2083.270 110.600 ;
        RECT 2082.950 62.460 2083.270 62.520 ;
        RECT 2082.580 62.320 2083.270 62.460 ;
        RECT 2082.580 62.180 2082.720 62.320 ;
        RECT 2082.950 62.260 2083.270 62.320 ;
        RECT 2082.490 61.920 2082.810 62.180 ;
        RECT 2082.490 40.020 2082.810 40.080 ;
        RECT 2744.430 40.020 2744.750 40.080 ;
        RECT 2082.490 39.880 2744.750 40.020 ;
        RECT 2082.490 39.820 2082.810 39.880 ;
        RECT 2744.430 39.820 2744.750 39.880 ;
      LAYER via ;
        RECT 2082.520 496.780 2082.780 497.040 ;
        RECT 2082.980 496.440 2083.240 496.700 ;
        RECT 2082.520 420.960 2082.780 421.220 ;
        RECT 2082.980 420.960 2083.240 421.220 ;
        RECT 2081.600 372.680 2081.860 372.940 ;
        RECT 2082.060 372.680 2082.320 372.940 ;
        RECT 2080.680 324.400 2080.940 324.660 ;
        RECT 2082.520 324.400 2082.780 324.660 ;
        RECT 2082.520 303.660 2082.780 303.920 ;
        RECT 2082.060 303.320 2082.320 303.580 ;
        RECT 2081.140 275.780 2081.400 276.040 ;
        RECT 2082.060 275.780 2082.320 276.040 ;
        RECT 2081.140 227.840 2081.400 228.100 ;
        RECT 2082.520 227.840 2082.780 228.100 ;
        RECT 2082.520 144.200 2082.780 144.460 ;
        RECT 2083.900 144.200 2084.160 144.460 ;
        RECT 2082.520 110.540 2082.780 110.800 ;
        RECT 2082.980 110.540 2083.240 110.800 ;
        RECT 2082.980 62.260 2083.240 62.520 ;
        RECT 2082.520 61.920 2082.780 62.180 ;
        RECT 2082.520 39.820 2082.780 40.080 ;
        RECT 2744.460 39.820 2744.720 40.080 ;
      LAYER met2 ;
        RECT 2079.530 601.530 2079.810 604.000 ;
        RECT 2079.530 601.390 2081.340 601.530 ;
        RECT 2079.530 600.000 2079.810 601.390 ;
        RECT 2081.200 545.090 2081.340 601.390 ;
        RECT 2081.200 544.950 2082.260 545.090 ;
        RECT 2082.120 544.410 2082.260 544.950 ;
        RECT 2082.120 544.270 2082.720 544.410 ;
        RECT 2082.580 497.070 2082.720 544.270 ;
        RECT 2082.520 496.750 2082.780 497.070 ;
        RECT 2082.980 496.410 2083.240 496.730 ;
        RECT 2083.040 421.250 2083.180 496.410 ;
        RECT 2082.520 420.930 2082.780 421.250 ;
        RECT 2082.980 420.930 2083.240 421.250 ;
        RECT 2082.580 401.610 2082.720 420.930 ;
        RECT 2082.120 401.470 2082.720 401.610 ;
        RECT 2082.120 372.970 2082.260 401.470 ;
        RECT 2081.600 372.650 2081.860 372.970 ;
        RECT 2082.060 372.650 2082.320 372.970 ;
        RECT 2081.660 353.330 2081.800 372.650 ;
        RECT 2080.740 353.190 2081.800 353.330 ;
        RECT 2080.740 324.690 2080.880 353.190 ;
        RECT 2080.680 324.370 2080.940 324.690 ;
        RECT 2082.520 324.370 2082.780 324.690 ;
        RECT 2082.580 303.950 2082.720 324.370 ;
        RECT 2082.520 303.630 2082.780 303.950 ;
        RECT 2082.060 303.290 2082.320 303.610 ;
        RECT 2082.120 276.070 2082.260 303.290 ;
        RECT 2081.140 275.750 2081.400 276.070 ;
        RECT 2082.060 275.750 2082.320 276.070 ;
        RECT 2081.200 228.130 2081.340 275.750 ;
        RECT 2081.140 227.810 2081.400 228.130 ;
        RECT 2082.520 227.810 2082.780 228.130 ;
        RECT 2082.580 227.645 2082.720 227.810 ;
        RECT 2082.510 227.275 2082.790 227.645 ;
        RECT 2083.890 226.595 2084.170 226.965 ;
        RECT 2083.960 144.490 2084.100 226.595 ;
        RECT 2082.520 144.170 2082.780 144.490 ;
        RECT 2083.900 144.170 2084.160 144.490 ;
        RECT 2082.580 110.830 2082.720 144.170 ;
        RECT 2082.520 110.510 2082.780 110.830 ;
        RECT 2082.980 110.510 2083.240 110.830 ;
        RECT 2083.040 62.550 2083.180 110.510 ;
        RECT 2082.980 62.230 2083.240 62.550 ;
        RECT 2082.520 61.890 2082.780 62.210 ;
        RECT 2082.580 40.110 2082.720 61.890 ;
        RECT 2082.520 39.790 2082.780 40.110 ;
        RECT 2744.460 39.790 2744.720 40.110 ;
        RECT 2744.520 2.400 2744.660 39.790 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
      LAYER via2 ;
        RECT 2082.510 227.320 2082.790 227.600 ;
        RECT 2083.890 226.640 2084.170 226.920 ;
      LAYER met3 ;
        RECT 2082.485 227.295 2082.815 227.625 ;
        RECT 2082.500 226.930 2082.800 227.295 ;
        RECT 2083.865 226.930 2084.195 226.945 ;
        RECT 2082.500 226.630 2084.195 226.930 ;
        RECT 2083.865 226.615 2084.195 226.630 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2089.850 39.680 2090.170 39.740 ;
        RECT 2761.910 39.680 2762.230 39.740 ;
        RECT 2089.850 39.540 2762.230 39.680 ;
        RECT 2089.850 39.480 2090.170 39.540 ;
        RECT 2761.910 39.480 2762.230 39.540 ;
      LAYER via ;
        RECT 2089.880 39.480 2090.140 39.740 ;
        RECT 2761.940 39.480 2762.200 39.740 ;
      LAYER met2 ;
        RECT 2088.730 600.170 2089.010 604.000 ;
        RECT 2088.730 600.030 2090.080 600.170 ;
        RECT 2088.730 600.000 2089.010 600.030 ;
        RECT 2089.940 39.770 2090.080 600.030 ;
        RECT 2089.880 39.450 2090.140 39.770 ;
        RECT 2761.940 39.450 2762.200 39.770 ;
        RECT 2762.000 2.400 2762.140 39.450 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 835.430 26.420 835.750 26.480 ;
        RECT 1097.170 26.420 1097.490 26.480 ;
        RECT 835.430 26.280 1097.490 26.420 ;
        RECT 835.430 26.220 835.750 26.280 ;
        RECT 1097.170 26.220 1097.490 26.280 ;
      LAYER via ;
        RECT 835.460 26.220 835.720 26.480 ;
        RECT 1097.200 26.220 1097.460 26.480 ;
      LAYER met2 ;
        RECT 1098.810 600.170 1099.090 604.000 ;
        RECT 1097.260 600.030 1099.090 600.170 ;
        RECT 1097.260 26.510 1097.400 600.030 ;
        RECT 1098.810 600.000 1099.090 600.030 ;
        RECT 835.460 26.190 835.720 26.510 ;
        RECT 1097.200 26.190 1097.460 26.510 ;
        RECT 835.520 2.400 835.660 26.190 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2099.510 586.740 2099.830 586.800 ;
        RECT 2103.650 586.740 2103.970 586.800 ;
        RECT 2099.510 586.600 2103.970 586.740 ;
        RECT 2099.510 586.540 2099.830 586.600 ;
        RECT 2103.650 586.540 2103.970 586.600 ;
        RECT 2103.650 39.340 2103.970 39.400 ;
        RECT 2779.850 39.340 2780.170 39.400 ;
        RECT 2103.650 39.200 2780.170 39.340 ;
        RECT 2103.650 39.140 2103.970 39.200 ;
        RECT 2779.850 39.140 2780.170 39.200 ;
      LAYER via ;
        RECT 2099.540 586.540 2099.800 586.800 ;
        RECT 2103.680 586.540 2103.940 586.800 ;
        RECT 2103.680 39.140 2103.940 39.400 ;
        RECT 2779.880 39.140 2780.140 39.400 ;
      LAYER met2 ;
        RECT 2097.930 600.170 2098.210 604.000 ;
        RECT 2097.930 600.030 2099.740 600.170 ;
        RECT 2097.930 600.000 2098.210 600.030 ;
        RECT 2099.600 586.830 2099.740 600.030 ;
        RECT 2099.540 586.510 2099.800 586.830 ;
        RECT 2103.680 586.510 2103.940 586.830 ;
        RECT 2103.740 39.430 2103.880 586.510 ;
        RECT 2103.680 39.110 2103.940 39.430 ;
        RECT 2779.880 39.110 2780.140 39.430 ;
        RECT 2779.940 2.400 2780.080 39.110 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2107.790 579.940 2108.110 580.000 ;
        RECT 2108.710 579.940 2109.030 580.000 ;
        RECT 2107.790 579.800 2109.030 579.940 ;
        RECT 2107.790 579.740 2108.110 579.800 ;
        RECT 2108.710 579.740 2109.030 579.800 ;
        RECT 2110.090 531.320 2110.410 531.380 ;
        RECT 2110.550 531.320 2110.870 531.380 ;
        RECT 2110.090 531.180 2110.870 531.320 ;
        RECT 2110.090 531.120 2110.410 531.180 ;
        RECT 2110.550 531.120 2110.870 531.180 ;
        RECT 2110.550 496.980 2110.870 497.040 ;
        RECT 2110.180 496.840 2110.870 496.980 ;
        RECT 2110.180 496.700 2110.320 496.840 ;
        RECT 2110.550 496.780 2110.870 496.840 ;
        RECT 2110.090 496.440 2110.410 496.700 ;
        RECT 2109.630 421.160 2109.950 421.220 ;
        RECT 2110.550 421.160 2110.870 421.220 ;
        RECT 2109.630 421.020 2110.870 421.160 ;
        RECT 2109.630 420.960 2109.950 421.020 ;
        RECT 2110.550 420.960 2110.870 421.020 ;
        RECT 2109.630 414.020 2109.950 414.080 ;
        RECT 2110.550 414.020 2110.870 414.080 ;
        RECT 2109.630 413.880 2110.870 414.020 ;
        RECT 2109.630 413.820 2109.950 413.880 ;
        RECT 2110.550 413.820 2110.870 413.880 ;
        RECT 2110.550 304.540 2110.870 304.600 ;
        RECT 2110.180 304.400 2110.870 304.540 ;
        RECT 2110.180 304.260 2110.320 304.400 ;
        RECT 2110.550 304.340 2110.870 304.400 ;
        RECT 2110.090 304.000 2110.410 304.260 ;
        RECT 2109.630 228.040 2109.950 228.100 ;
        RECT 2110.550 228.040 2110.870 228.100 ;
        RECT 2109.630 227.900 2110.870 228.040 ;
        RECT 2109.630 227.840 2109.950 227.900 ;
        RECT 2110.550 227.840 2110.870 227.900 ;
        RECT 2108.710 220.560 2109.030 220.620 ;
        RECT 2109.630 220.560 2109.950 220.620 ;
        RECT 2108.710 220.420 2109.950 220.560 ;
        RECT 2108.710 220.360 2109.030 220.420 ;
        RECT 2109.630 220.360 2109.950 220.420 ;
        RECT 2108.710 172.620 2109.030 172.680 ;
        RECT 2110.090 172.620 2110.410 172.680 ;
        RECT 2108.710 172.480 2110.410 172.620 ;
        RECT 2108.710 172.420 2109.030 172.480 ;
        RECT 2110.090 172.420 2110.410 172.480 ;
        RECT 2109.170 76.060 2109.490 76.120 ;
        RECT 2109.630 76.060 2109.950 76.120 ;
        RECT 2109.170 75.920 2109.950 76.060 ;
        RECT 2109.170 75.860 2109.490 75.920 ;
        RECT 2109.630 75.860 2109.950 75.920 ;
        RECT 2109.170 48.520 2109.490 48.580 ;
        RECT 2110.090 48.520 2110.410 48.580 ;
        RECT 2109.170 48.380 2110.410 48.520 ;
        RECT 2109.170 48.320 2109.490 48.380 ;
        RECT 2110.090 48.320 2110.410 48.380 ;
        RECT 2110.090 39.000 2110.410 39.060 ;
        RECT 2797.790 39.000 2798.110 39.060 ;
        RECT 2110.090 38.860 2798.110 39.000 ;
        RECT 2110.090 38.800 2110.410 38.860 ;
        RECT 2797.790 38.800 2798.110 38.860 ;
      LAYER via ;
        RECT 2107.820 579.740 2108.080 580.000 ;
        RECT 2108.740 579.740 2109.000 580.000 ;
        RECT 2110.120 531.120 2110.380 531.380 ;
        RECT 2110.580 531.120 2110.840 531.380 ;
        RECT 2110.580 496.780 2110.840 497.040 ;
        RECT 2110.120 496.440 2110.380 496.700 ;
        RECT 2109.660 420.960 2109.920 421.220 ;
        RECT 2110.580 420.960 2110.840 421.220 ;
        RECT 2109.660 413.820 2109.920 414.080 ;
        RECT 2110.580 413.820 2110.840 414.080 ;
        RECT 2110.580 304.340 2110.840 304.600 ;
        RECT 2110.120 304.000 2110.380 304.260 ;
        RECT 2109.660 227.840 2109.920 228.100 ;
        RECT 2110.580 227.840 2110.840 228.100 ;
        RECT 2108.740 220.360 2109.000 220.620 ;
        RECT 2109.660 220.360 2109.920 220.620 ;
        RECT 2108.740 172.420 2109.000 172.680 ;
        RECT 2110.120 172.420 2110.380 172.680 ;
        RECT 2109.200 75.860 2109.460 76.120 ;
        RECT 2109.660 75.860 2109.920 76.120 ;
        RECT 2109.200 48.320 2109.460 48.580 ;
        RECT 2110.120 48.320 2110.380 48.580 ;
        RECT 2110.120 38.800 2110.380 39.060 ;
        RECT 2797.820 38.800 2798.080 39.060 ;
      LAYER met2 ;
        RECT 2107.130 600.170 2107.410 604.000 ;
        RECT 2107.130 600.030 2108.020 600.170 ;
        RECT 2107.130 600.000 2107.410 600.030 ;
        RECT 2107.880 580.030 2108.020 600.030 ;
        RECT 2107.820 579.710 2108.080 580.030 ;
        RECT 2108.740 579.710 2109.000 580.030 ;
        RECT 2108.800 545.090 2108.940 579.710 ;
        RECT 2108.800 544.950 2109.860 545.090 ;
        RECT 2109.720 544.410 2109.860 544.950 ;
        RECT 2109.720 544.270 2110.320 544.410 ;
        RECT 2110.180 531.410 2110.320 544.270 ;
        RECT 2110.120 531.090 2110.380 531.410 ;
        RECT 2110.580 531.090 2110.840 531.410 ;
        RECT 2110.640 497.070 2110.780 531.090 ;
        RECT 2110.580 496.750 2110.840 497.070 ;
        RECT 2110.120 496.410 2110.380 496.730 ;
        RECT 2110.180 483.210 2110.320 496.410 ;
        RECT 2110.180 483.070 2110.780 483.210 ;
        RECT 2110.640 421.250 2110.780 483.070 ;
        RECT 2109.660 420.930 2109.920 421.250 ;
        RECT 2110.580 420.930 2110.840 421.250 ;
        RECT 2109.720 414.110 2109.860 420.930 ;
        RECT 2109.660 413.790 2109.920 414.110 ;
        RECT 2110.580 413.790 2110.840 414.110 ;
        RECT 2110.640 304.630 2110.780 413.790 ;
        RECT 2110.580 304.310 2110.840 304.630 ;
        RECT 2110.120 303.970 2110.380 304.290 ;
        RECT 2110.180 283.290 2110.320 303.970 ;
        RECT 2109.720 283.150 2110.320 283.290 ;
        RECT 2109.720 240.450 2109.860 283.150 ;
        RECT 2109.720 240.310 2110.780 240.450 ;
        RECT 2110.640 228.130 2110.780 240.310 ;
        RECT 2109.660 227.810 2109.920 228.130 ;
        RECT 2110.580 227.810 2110.840 228.130 ;
        RECT 2109.720 220.650 2109.860 227.810 ;
        RECT 2108.740 220.330 2109.000 220.650 ;
        RECT 2109.660 220.330 2109.920 220.650 ;
        RECT 2108.800 172.710 2108.940 220.330 ;
        RECT 2108.740 172.390 2109.000 172.710 ;
        RECT 2110.120 172.390 2110.380 172.710 ;
        RECT 2110.180 111.250 2110.320 172.390 ;
        RECT 2109.720 111.110 2110.320 111.250 ;
        RECT 2109.720 76.150 2109.860 111.110 ;
        RECT 2109.200 75.830 2109.460 76.150 ;
        RECT 2109.660 75.830 2109.920 76.150 ;
        RECT 2109.260 48.610 2109.400 75.830 ;
        RECT 2109.200 48.290 2109.460 48.610 ;
        RECT 2110.120 48.290 2110.380 48.610 ;
        RECT 2110.180 39.090 2110.320 48.290 ;
        RECT 2110.120 38.770 2110.380 39.090 ;
        RECT 2797.820 38.770 2798.080 39.090 ;
        RECT 2797.880 2.400 2798.020 38.770 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2117.450 38.660 2117.770 38.720 ;
        RECT 2815.730 38.660 2816.050 38.720 ;
        RECT 2117.450 38.520 2816.050 38.660 ;
        RECT 2117.450 38.460 2117.770 38.520 ;
        RECT 2815.730 38.460 2816.050 38.520 ;
      LAYER via ;
        RECT 2117.480 38.460 2117.740 38.720 ;
        RECT 2815.760 38.460 2816.020 38.720 ;
      LAYER met2 ;
        RECT 2116.330 600.170 2116.610 604.000 ;
        RECT 2116.330 600.030 2117.680 600.170 ;
        RECT 2116.330 600.000 2116.610 600.030 ;
        RECT 2117.540 38.750 2117.680 600.030 ;
        RECT 2117.480 38.430 2117.740 38.750 ;
        RECT 2815.760 38.430 2816.020 38.750 ;
        RECT 2815.820 2.400 2815.960 38.430 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2127.110 588.100 2127.430 588.160 ;
        RECT 2130.790 588.100 2131.110 588.160 ;
        RECT 2127.110 587.960 2131.110 588.100 ;
        RECT 2127.110 587.900 2127.430 587.960 ;
        RECT 2130.790 587.900 2131.110 587.960 ;
        RECT 2130.790 38.320 2131.110 38.380 ;
        RECT 2833.670 38.320 2833.990 38.380 ;
        RECT 2130.790 38.180 2833.990 38.320 ;
        RECT 2130.790 38.120 2131.110 38.180 ;
        RECT 2833.670 38.120 2833.990 38.180 ;
      LAYER via ;
        RECT 2127.140 587.900 2127.400 588.160 ;
        RECT 2130.820 587.900 2131.080 588.160 ;
        RECT 2130.820 38.120 2131.080 38.380 ;
        RECT 2833.700 38.120 2833.960 38.380 ;
      LAYER met2 ;
        RECT 2125.530 600.170 2125.810 604.000 ;
        RECT 2125.530 600.030 2127.340 600.170 ;
        RECT 2125.530 600.000 2125.810 600.030 ;
        RECT 2127.200 588.190 2127.340 600.030 ;
        RECT 2127.140 587.870 2127.400 588.190 ;
        RECT 2130.820 587.870 2131.080 588.190 ;
        RECT 2130.880 38.410 2131.020 587.870 ;
        RECT 2130.820 38.090 2131.080 38.410 ;
        RECT 2833.700 38.090 2833.960 38.410 ;
        RECT 2833.760 2.400 2833.900 38.090 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2136.310 586.740 2136.630 586.800 ;
        RECT 2138.610 586.740 2138.930 586.800 ;
        RECT 2136.310 586.600 2138.930 586.740 ;
        RECT 2136.310 586.540 2136.630 586.600 ;
        RECT 2138.610 586.540 2138.930 586.600 ;
        RECT 2138.610 37.980 2138.930 38.040 ;
        RECT 2851.150 37.980 2851.470 38.040 ;
        RECT 2138.610 37.840 2851.470 37.980 ;
        RECT 2138.610 37.780 2138.930 37.840 ;
        RECT 2851.150 37.780 2851.470 37.840 ;
      LAYER via ;
        RECT 2136.340 586.540 2136.600 586.800 ;
        RECT 2138.640 586.540 2138.900 586.800 ;
        RECT 2138.640 37.780 2138.900 38.040 ;
        RECT 2851.180 37.780 2851.440 38.040 ;
      LAYER met2 ;
        RECT 2134.730 600.170 2135.010 604.000 ;
        RECT 2134.730 600.030 2136.540 600.170 ;
        RECT 2134.730 600.000 2135.010 600.030 ;
        RECT 2136.400 586.830 2136.540 600.030 ;
        RECT 2136.340 586.510 2136.600 586.830 ;
        RECT 2138.640 586.510 2138.900 586.830 ;
        RECT 2138.700 38.070 2138.840 586.510 ;
        RECT 2138.640 37.750 2138.900 38.070 ;
        RECT 2851.180 37.750 2851.440 38.070 ;
        RECT 2851.240 2.400 2851.380 37.750 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2145.050 45.460 2145.370 45.520 ;
        RECT 2869.090 45.460 2869.410 45.520 ;
        RECT 2145.050 45.320 2869.410 45.460 ;
        RECT 2145.050 45.260 2145.370 45.320 ;
        RECT 2869.090 45.260 2869.410 45.320 ;
      LAYER via ;
        RECT 2145.080 45.260 2145.340 45.520 ;
        RECT 2869.120 45.260 2869.380 45.520 ;
      LAYER met2 ;
        RECT 2143.930 600.170 2144.210 604.000 ;
        RECT 2143.930 600.030 2145.280 600.170 ;
        RECT 2143.930 600.000 2144.210 600.030 ;
        RECT 2145.140 45.550 2145.280 600.030 ;
        RECT 2145.080 45.230 2145.340 45.550 ;
        RECT 2869.120 45.230 2869.380 45.550 ;
        RECT 2869.180 2.400 2869.320 45.230 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2154.710 586.740 2155.030 586.800 ;
        RECT 2158.850 586.740 2159.170 586.800 ;
        RECT 2154.710 586.600 2159.170 586.740 ;
        RECT 2154.710 586.540 2155.030 586.600 ;
        RECT 2158.850 586.540 2159.170 586.600 ;
        RECT 2158.850 45.120 2159.170 45.180 ;
        RECT 2887.030 45.120 2887.350 45.180 ;
        RECT 2158.850 44.980 2887.350 45.120 ;
        RECT 2158.850 44.920 2159.170 44.980 ;
        RECT 2887.030 44.920 2887.350 44.980 ;
      LAYER via ;
        RECT 2154.740 586.540 2155.000 586.800 ;
        RECT 2158.880 586.540 2159.140 586.800 ;
        RECT 2158.880 44.920 2159.140 45.180 ;
        RECT 2887.060 44.920 2887.320 45.180 ;
      LAYER met2 ;
        RECT 2153.130 600.170 2153.410 604.000 ;
        RECT 2153.130 600.030 2154.940 600.170 ;
        RECT 2153.130 600.000 2153.410 600.030 ;
        RECT 2154.800 586.830 2154.940 600.030 ;
        RECT 2154.740 586.510 2155.000 586.830 ;
        RECT 2158.880 586.510 2159.140 586.830 ;
        RECT 2158.940 45.210 2159.080 586.510 ;
        RECT 2158.880 44.890 2159.140 45.210 ;
        RECT 2887.060 44.890 2887.320 45.210 ;
        RECT 2887.120 2.400 2887.260 44.890 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2165.290 545.400 2165.610 545.660 ;
        RECT 2165.380 544.980 2165.520 545.400 ;
        RECT 2165.290 544.720 2165.610 544.980 ;
        RECT 2163.450 379.340 2163.770 379.400 ;
        RECT 2165.290 379.340 2165.610 379.400 ;
        RECT 2163.450 379.200 2165.610 379.340 ;
        RECT 2163.450 379.140 2163.770 379.200 ;
        RECT 2165.290 379.140 2165.610 379.200 ;
        RECT 2163.450 331.740 2163.770 331.800 ;
        RECT 2163.910 331.740 2164.230 331.800 ;
        RECT 2163.450 331.600 2164.230 331.740 ;
        RECT 2163.450 331.540 2163.770 331.600 ;
        RECT 2163.910 331.540 2164.230 331.600 ;
        RECT 2163.450 324.260 2163.770 324.320 ;
        RECT 2164.370 324.260 2164.690 324.320 ;
        RECT 2163.450 324.120 2164.690 324.260 ;
        RECT 2163.450 324.060 2163.770 324.120 ;
        RECT 2164.370 324.060 2164.690 324.120 ;
        RECT 2163.450 276.320 2163.770 276.380 ;
        RECT 2164.830 276.320 2165.150 276.380 ;
        RECT 2163.450 276.180 2165.150 276.320 ;
        RECT 2163.450 276.120 2163.770 276.180 ;
        RECT 2164.830 276.120 2165.150 276.180 ;
        RECT 2164.370 234.840 2164.690 234.900 ;
        RECT 2164.830 234.840 2165.150 234.900 ;
        RECT 2164.370 234.700 2165.150 234.840 ;
        RECT 2164.370 234.640 2164.690 234.700 ;
        RECT 2164.830 234.640 2165.150 234.700 ;
        RECT 2164.830 145.080 2165.150 145.140 ;
        RECT 2165.750 145.080 2166.070 145.140 ;
        RECT 2164.830 144.940 2166.070 145.080 ;
        RECT 2164.830 144.880 2165.150 144.940 ;
        RECT 2165.750 144.880 2166.070 144.940 ;
        RECT 2163.910 96.460 2164.230 96.520 ;
        RECT 2164.830 96.460 2165.150 96.520 ;
        RECT 2163.910 96.320 2165.150 96.460 ;
        RECT 2163.910 96.260 2164.230 96.320 ;
        RECT 2164.830 96.260 2165.150 96.320 ;
        RECT 2163.910 48.520 2164.230 48.580 ;
        RECT 2165.290 48.520 2165.610 48.580 ;
        RECT 2163.910 48.380 2165.610 48.520 ;
        RECT 2163.910 48.320 2164.230 48.380 ;
        RECT 2165.290 48.320 2165.610 48.380 ;
        RECT 2164.830 44.780 2165.150 44.840 ;
        RECT 2904.970 44.780 2905.290 44.840 ;
        RECT 2164.830 44.640 2905.290 44.780 ;
        RECT 2164.830 44.580 2165.150 44.640 ;
        RECT 2904.970 44.580 2905.290 44.640 ;
      LAYER via ;
        RECT 2165.320 545.400 2165.580 545.660 ;
        RECT 2165.320 544.720 2165.580 544.980 ;
        RECT 2163.480 379.140 2163.740 379.400 ;
        RECT 2165.320 379.140 2165.580 379.400 ;
        RECT 2163.480 331.540 2163.740 331.800 ;
        RECT 2163.940 331.540 2164.200 331.800 ;
        RECT 2163.480 324.060 2163.740 324.320 ;
        RECT 2164.400 324.060 2164.660 324.320 ;
        RECT 2163.480 276.120 2163.740 276.380 ;
        RECT 2164.860 276.120 2165.120 276.380 ;
        RECT 2164.400 234.640 2164.660 234.900 ;
        RECT 2164.860 234.640 2165.120 234.900 ;
        RECT 2164.860 144.880 2165.120 145.140 ;
        RECT 2165.780 144.880 2166.040 145.140 ;
        RECT 2163.940 96.260 2164.200 96.520 ;
        RECT 2164.860 96.260 2165.120 96.520 ;
        RECT 2163.940 48.320 2164.200 48.580 ;
        RECT 2165.320 48.320 2165.580 48.580 ;
        RECT 2164.860 44.580 2165.120 44.840 ;
        RECT 2905.000 44.580 2905.260 44.840 ;
      LAYER met2 ;
        RECT 2162.330 600.170 2162.610 604.000 ;
        RECT 2162.330 600.030 2164.140 600.170 ;
        RECT 2162.330 600.000 2162.610 600.030 ;
        RECT 2164.000 596.770 2164.140 600.030 ;
        RECT 2164.000 596.630 2165.060 596.770 ;
        RECT 2164.920 593.370 2165.060 596.630 ;
        RECT 2164.920 593.230 2165.520 593.370 ;
        RECT 2165.380 545.690 2165.520 593.230 ;
        RECT 2165.320 545.370 2165.580 545.690 ;
        RECT 2165.320 544.690 2165.580 545.010 ;
        RECT 2165.380 507.010 2165.520 544.690 ;
        RECT 2164.920 506.870 2165.520 507.010 ;
        RECT 2164.920 448.530 2165.060 506.870 ;
        RECT 2164.920 448.390 2165.520 448.530 ;
        RECT 2165.380 401.045 2165.520 448.390 ;
        RECT 2165.310 400.675 2165.590 401.045 ;
        RECT 2165.310 399.315 2165.590 399.685 ;
        RECT 2165.380 379.430 2165.520 399.315 ;
        RECT 2163.480 379.110 2163.740 379.430 ;
        RECT 2165.320 379.110 2165.580 379.430 ;
        RECT 2163.540 331.830 2163.680 379.110 ;
        RECT 2163.480 331.510 2163.740 331.830 ;
        RECT 2163.940 331.570 2164.200 331.830 ;
        RECT 2163.940 331.510 2164.600 331.570 ;
        RECT 2164.000 331.430 2164.600 331.510 ;
        RECT 2164.460 324.350 2164.600 331.430 ;
        RECT 2163.480 324.030 2163.740 324.350 ;
        RECT 2164.400 324.030 2164.660 324.350 ;
        RECT 2163.540 276.410 2163.680 324.030 ;
        RECT 2163.480 276.090 2163.740 276.410 ;
        RECT 2164.860 276.090 2165.120 276.410 ;
        RECT 2164.920 234.930 2165.060 276.090 ;
        RECT 2164.400 234.610 2164.660 234.930 ;
        RECT 2164.860 234.610 2165.120 234.930 ;
        RECT 2164.460 207.245 2164.600 234.610 ;
        RECT 2164.390 206.875 2164.670 207.245 ;
        RECT 2164.390 206.195 2164.670 206.565 ;
        RECT 2164.460 169.050 2164.600 206.195 ;
        RECT 2164.460 168.910 2165.060 169.050 ;
        RECT 2164.920 145.170 2165.060 168.910 ;
        RECT 2164.860 144.850 2165.120 145.170 ;
        RECT 2165.780 144.850 2166.040 145.170 ;
        RECT 2165.840 110.570 2165.980 144.850 ;
        RECT 2164.920 110.430 2165.980 110.570 ;
        RECT 2164.920 96.550 2165.060 110.430 ;
        RECT 2163.940 96.230 2164.200 96.550 ;
        RECT 2164.860 96.230 2165.120 96.550 ;
        RECT 2164.000 48.610 2164.140 96.230 ;
        RECT 2163.940 48.290 2164.200 48.610 ;
        RECT 2165.320 48.290 2165.580 48.610 ;
        RECT 2165.380 48.010 2165.520 48.290 ;
        RECT 2164.920 47.870 2165.520 48.010 ;
        RECT 2164.920 44.870 2165.060 47.870 ;
        RECT 2164.860 44.550 2165.120 44.870 ;
        RECT 2905.000 44.550 2905.260 44.870 ;
        RECT 2905.060 2.400 2905.200 44.550 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 2165.310 400.720 2165.590 401.000 ;
        RECT 2165.310 399.360 2165.590 399.640 ;
        RECT 2164.390 206.920 2164.670 207.200 ;
        RECT 2164.390 206.240 2164.670 206.520 ;
      LAYER met3 ;
        RECT 2165.285 401.010 2165.615 401.025 ;
        RECT 2165.070 400.695 2165.615 401.010 ;
        RECT 2165.070 399.665 2165.370 400.695 ;
        RECT 2165.070 399.350 2165.615 399.665 ;
        RECT 2165.285 399.335 2165.615 399.350 ;
        RECT 2164.365 207.210 2164.695 207.225 ;
        RECT 2164.150 206.895 2164.695 207.210 ;
        RECT 2164.150 206.545 2164.450 206.895 ;
        RECT 2164.150 206.230 2164.695 206.545 ;
        RECT 2164.365 206.215 2164.695 206.230 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1105.910 572.460 1106.230 572.520 ;
        RECT 1106.830 572.460 1107.150 572.520 ;
        RECT 1105.910 572.320 1107.150 572.460 ;
        RECT 1105.910 572.260 1106.230 572.320 ;
        RECT 1106.830 572.260 1107.150 572.320 ;
        RECT 1105.910 524.520 1106.230 524.580 ;
        RECT 1106.830 524.520 1107.150 524.580 ;
        RECT 1105.910 524.380 1107.150 524.520 ;
        RECT 1105.910 524.320 1106.230 524.380 ;
        RECT 1106.830 524.320 1107.150 524.380 ;
        RECT 1104.990 476.240 1105.310 476.300 ;
        RECT 1105.910 476.240 1106.230 476.300 ;
        RECT 1104.990 476.100 1106.230 476.240 ;
        RECT 1104.990 476.040 1105.310 476.100 ;
        RECT 1105.910 476.040 1106.230 476.100 ;
        RECT 1104.990 427.620 1105.310 427.680 ;
        RECT 1106.370 427.620 1106.690 427.680 ;
        RECT 1104.990 427.480 1106.690 427.620 ;
        RECT 1104.990 427.420 1105.310 427.480 ;
        RECT 1106.370 427.420 1106.690 427.480 ;
        RECT 1105.450 379.680 1105.770 379.740 ;
        RECT 1106.370 379.680 1106.690 379.740 ;
        RECT 1105.450 379.540 1106.690 379.680 ;
        RECT 1105.450 379.480 1105.770 379.540 ;
        RECT 1106.370 379.480 1106.690 379.540 ;
        RECT 1104.990 338.200 1105.310 338.260 ;
        RECT 1105.450 338.200 1105.770 338.260 ;
        RECT 1104.990 338.060 1105.770 338.200 ;
        RECT 1104.990 338.000 1105.310 338.060 ;
        RECT 1105.450 338.000 1105.770 338.060 ;
        RECT 1104.530 331.060 1104.850 331.120 ;
        RECT 1104.990 331.060 1105.310 331.120 ;
        RECT 1104.530 330.920 1105.310 331.060 ;
        RECT 1104.530 330.860 1104.850 330.920 ;
        RECT 1104.990 330.860 1105.310 330.920 ;
        RECT 1104.530 283.120 1104.850 283.180 ;
        RECT 1105.450 283.120 1105.770 283.180 ;
        RECT 1104.530 282.980 1105.770 283.120 ;
        RECT 1104.530 282.920 1104.850 282.980 ;
        RECT 1105.450 282.920 1105.770 282.980 ;
        RECT 1104.530 282.440 1104.850 282.500 ;
        RECT 1105.450 282.440 1105.770 282.500 ;
        RECT 1104.530 282.300 1105.770 282.440 ;
        RECT 1104.530 282.240 1104.850 282.300 ;
        RECT 1105.450 282.240 1105.770 282.300 ;
        RECT 1104.530 234.840 1104.850 234.900 ;
        RECT 1105.910 234.840 1106.230 234.900 ;
        RECT 1104.530 234.700 1106.230 234.840 ;
        RECT 1104.530 234.640 1104.850 234.700 ;
        RECT 1105.910 234.640 1106.230 234.700 ;
        RECT 1104.990 206.620 1105.310 206.680 ;
        RECT 1105.910 206.620 1106.230 206.680 ;
        RECT 1104.990 206.480 1106.230 206.620 ;
        RECT 1104.990 206.420 1105.310 206.480 ;
        RECT 1105.910 206.420 1106.230 206.480 ;
        RECT 1104.530 138.280 1104.850 138.340 ;
        RECT 1105.450 138.280 1105.770 138.340 ;
        RECT 1104.530 138.140 1105.770 138.280 ;
        RECT 1104.530 138.080 1104.850 138.140 ;
        RECT 1105.450 138.080 1105.770 138.140 ;
        RECT 1105.450 110.740 1105.770 110.800 ;
        RECT 1105.080 110.600 1105.770 110.740 ;
        RECT 1105.080 110.460 1105.220 110.600 ;
        RECT 1105.450 110.540 1105.770 110.600 ;
        RECT 1104.990 110.200 1105.310 110.460 ;
        RECT 852.910 26.760 853.230 26.820 ;
        RECT 1104.530 26.760 1104.850 26.820 ;
        RECT 852.910 26.620 1104.850 26.760 ;
        RECT 852.910 26.560 853.230 26.620 ;
        RECT 1104.530 26.560 1104.850 26.620 ;
      LAYER via ;
        RECT 1105.940 572.260 1106.200 572.520 ;
        RECT 1106.860 572.260 1107.120 572.520 ;
        RECT 1105.940 524.320 1106.200 524.580 ;
        RECT 1106.860 524.320 1107.120 524.580 ;
        RECT 1105.020 476.040 1105.280 476.300 ;
        RECT 1105.940 476.040 1106.200 476.300 ;
        RECT 1105.020 427.420 1105.280 427.680 ;
        RECT 1106.400 427.420 1106.660 427.680 ;
        RECT 1105.480 379.480 1105.740 379.740 ;
        RECT 1106.400 379.480 1106.660 379.740 ;
        RECT 1105.020 338.000 1105.280 338.260 ;
        RECT 1105.480 338.000 1105.740 338.260 ;
        RECT 1104.560 330.860 1104.820 331.120 ;
        RECT 1105.020 330.860 1105.280 331.120 ;
        RECT 1104.560 282.920 1104.820 283.180 ;
        RECT 1105.480 282.920 1105.740 283.180 ;
        RECT 1104.560 282.240 1104.820 282.500 ;
        RECT 1105.480 282.240 1105.740 282.500 ;
        RECT 1104.560 234.640 1104.820 234.900 ;
        RECT 1105.940 234.640 1106.200 234.900 ;
        RECT 1105.020 206.420 1105.280 206.680 ;
        RECT 1105.940 206.420 1106.200 206.680 ;
        RECT 1104.560 138.080 1104.820 138.340 ;
        RECT 1105.480 138.080 1105.740 138.340 ;
        RECT 1105.480 110.540 1105.740 110.800 ;
        RECT 1105.020 110.200 1105.280 110.460 ;
        RECT 852.940 26.560 853.200 26.820 ;
        RECT 1104.560 26.560 1104.820 26.820 ;
      LAYER met2 ;
        RECT 1108.010 600.170 1108.290 604.000 ;
        RECT 1107.380 600.030 1108.290 600.170 ;
        RECT 1107.380 573.765 1107.520 600.030 ;
        RECT 1108.010 600.000 1108.290 600.030 ;
        RECT 1107.310 573.395 1107.590 573.765 ;
        RECT 1105.930 572.715 1106.210 573.085 ;
        RECT 1106.000 572.550 1106.140 572.715 ;
        RECT 1105.940 572.230 1106.200 572.550 ;
        RECT 1106.860 572.230 1107.120 572.550 ;
        RECT 1106.920 524.610 1107.060 572.230 ;
        RECT 1105.940 524.290 1106.200 524.610 ;
        RECT 1106.860 524.290 1107.120 524.610 ;
        RECT 1106.000 476.330 1106.140 524.290 ;
        RECT 1105.020 476.010 1105.280 476.330 ;
        RECT 1105.940 476.010 1106.200 476.330 ;
        RECT 1105.080 441.730 1105.220 476.010 ;
        RECT 1104.620 441.590 1105.220 441.730 ;
        RECT 1104.620 434.250 1104.760 441.590 ;
        RECT 1104.620 434.110 1105.220 434.250 ;
        RECT 1105.080 427.710 1105.220 434.110 ;
        RECT 1105.020 427.390 1105.280 427.710 ;
        RECT 1106.400 427.390 1106.660 427.710 ;
        RECT 1106.460 379.770 1106.600 427.390 ;
        RECT 1105.480 379.450 1105.740 379.770 ;
        RECT 1106.400 379.450 1106.660 379.770 ;
        RECT 1105.540 338.290 1105.680 379.450 ;
        RECT 1105.020 337.970 1105.280 338.290 ;
        RECT 1105.480 337.970 1105.740 338.290 ;
        RECT 1105.080 331.150 1105.220 337.970 ;
        RECT 1104.560 330.830 1104.820 331.150 ;
        RECT 1105.020 330.830 1105.280 331.150 ;
        RECT 1104.620 283.210 1104.760 330.830 ;
        RECT 1104.560 282.890 1104.820 283.210 ;
        RECT 1105.480 282.890 1105.740 283.210 ;
        RECT 1105.540 282.530 1105.680 282.890 ;
        RECT 1104.560 282.210 1104.820 282.530 ;
        RECT 1105.480 282.210 1105.740 282.530 ;
        RECT 1104.620 234.930 1104.760 282.210 ;
        RECT 1104.560 234.610 1104.820 234.930 ;
        RECT 1105.940 234.610 1106.200 234.930 ;
        RECT 1106.000 206.710 1106.140 234.610 ;
        RECT 1105.020 206.390 1105.280 206.710 ;
        RECT 1105.940 206.390 1106.200 206.710 ;
        RECT 1105.080 162.250 1105.220 206.390 ;
        RECT 1104.620 162.110 1105.220 162.250 ;
        RECT 1104.620 138.370 1104.760 162.110 ;
        RECT 1104.560 138.050 1104.820 138.370 ;
        RECT 1105.480 138.050 1105.740 138.370 ;
        RECT 1105.540 110.830 1105.680 138.050 ;
        RECT 1105.480 110.510 1105.740 110.830 ;
        RECT 1105.020 110.170 1105.280 110.490 ;
        RECT 1105.080 73.170 1105.220 110.170 ;
        RECT 1105.080 73.030 1105.680 73.170 ;
        RECT 1105.540 71.810 1105.680 73.030 ;
        RECT 1104.620 71.670 1105.680 71.810 ;
        RECT 1104.620 26.850 1104.760 71.670 ;
        RECT 852.940 26.530 853.200 26.850 ;
        RECT 1104.560 26.530 1104.820 26.850 ;
        RECT 853.000 2.400 853.140 26.530 ;
        RECT 852.790 -4.800 853.350 2.400 ;
      LAYER via2 ;
        RECT 1107.310 573.440 1107.590 573.720 ;
        RECT 1105.930 572.760 1106.210 573.040 ;
      LAYER met3 ;
        RECT 1107.285 573.730 1107.615 573.745 ;
        RECT 1105.230 573.430 1107.615 573.730 ;
        RECT 1105.230 573.050 1105.530 573.430 ;
        RECT 1107.285 573.415 1107.615 573.430 ;
        RECT 1105.905 573.050 1106.235 573.065 ;
        RECT 1105.230 572.750 1106.235 573.050 ;
        RECT 1105.905 572.735 1106.235 572.750 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 875.910 590.480 876.230 590.540 ;
        RECT 1115.570 590.480 1115.890 590.540 ;
        RECT 875.910 590.340 1115.890 590.480 ;
        RECT 875.910 590.280 876.230 590.340 ;
        RECT 1115.570 590.280 1115.890 590.340 ;
        RECT 870.850 20.640 871.170 20.700 ;
        RECT 875.910 20.640 876.230 20.700 ;
        RECT 870.850 20.500 876.230 20.640 ;
        RECT 870.850 20.440 871.170 20.500 ;
        RECT 875.910 20.440 876.230 20.500 ;
      LAYER via ;
        RECT 875.940 590.280 876.200 590.540 ;
        RECT 1115.600 590.280 1115.860 590.540 ;
        RECT 870.880 20.440 871.140 20.700 ;
        RECT 875.940 20.440 876.200 20.700 ;
      LAYER met2 ;
        RECT 1117.210 600.170 1117.490 604.000 ;
        RECT 1115.660 600.030 1117.490 600.170 ;
        RECT 1115.660 590.570 1115.800 600.030 ;
        RECT 1117.210 600.000 1117.490 600.030 ;
        RECT 875.940 590.250 876.200 590.570 ;
        RECT 1115.600 590.250 1115.860 590.570 ;
        RECT 876.000 20.730 876.140 590.250 ;
        RECT 870.880 20.410 871.140 20.730 ;
        RECT 875.940 20.410 876.200 20.730 ;
        RECT 870.940 2.400 871.080 20.410 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 889.710 589.800 890.030 589.860 ;
        RECT 1124.770 589.800 1125.090 589.860 ;
        RECT 889.710 589.660 1125.090 589.800 ;
        RECT 889.710 589.600 890.030 589.660 ;
        RECT 1124.770 589.600 1125.090 589.660 ;
      LAYER via ;
        RECT 889.740 589.600 890.000 589.860 ;
        RECT 1124.800 589.600 1125.060 589.860 ;
      LAYER met2 ;
        RECT 1126.410 600.170 1126.690 604.000 ;
        RECT 1124.860 600.030 1126.690 600.170 ;
        RECT 1124.860 589.890 1125.000 600.030 ;
        RECT 1126.410 600.000 1126.690 600.030 ;
        RECT 889.740 589.570 890.000 589.890 ;
        RECT 1124.800 589.570 1125.060 589.890 ;
        RECT 889.800 3.130 889.940 589.570 ;
        RECT 888.880 2.990 889.940 3.130 ;
        RECT 888.880 2.400 889.020 2.990 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 910.410 590.140 910.730 590.200 ;
        RECT 1133.970 590.140 1134.290 590.200 ;
        RECT 910.410 590.000 1134.290 590.140 ;
        RECT 910.410 589.940 910.730 590.000 ;
        RECT 1133.970 589.940 1134.290 590.000 ;
        RECT 906.730 20.640 907.050 20.700 ;
        RECT 910.410 20.640 910.730 20.700 ;
        RECT 906.730 20.500 910.730 20.640 ;
        RECT 906.730 20.440 907.050 20.500 ;
        RECT 910.410 20.440 910.730 20.500 ;
      LAYER via ;
        RECT 910.440 589.940 910.700 590.200 ;
        RECT 1134.000 589.940 1134.260 590.200 ;
        RECT 906.760 20.440 907.020 20.700 ;
        RECT 910.440 20.440 910.700 20.700 ;
      LAYER met2 ;
        RECT 1135.610 600.170 1135.890 604.000 ;
        RECT 1134.060 600.030 1135.890 600.170 ;
        RECT 1134.060 590.230 1134.200 600.030 ;
        RECT 1135.610 600.000 1135.890 600.030 ;
        RECT 910.440 589.910 910.700 590.230 ;
        RECT 1134.000 589.910 1134.260 590.230 ;
        RECT 910.500 20.730 910.640 589.910 ;
        RECT 906.760 20.410 907.020 20.730 ;
        RECT 910.440 20.410 910.700 20.730 ;
        RECT 906.820 2.400 906.960 20.410 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 592.180 924.530 592.240 ;
        RECT 1143.170 592.180 1143.490 592.240 ;
        RECT 924.210 592.040 1143.490 592.180 ;
        RECT 924.210 591.980 924.530 592.040 ;
        RECT 1143.170 591.980 1143.490 592.040 ;
      LAYER via ;
        RECT 924.240 591.980 924.500 592.240 ;
        RECT 1143.200 591.980 1143.460 592.240 ;
      LAYER met2 ;
        RECT 1144.810 600.170 1145.090 604.000 ;
        RECT 1143.260 600.030 1145.090 600.170 ;
        RECT 1143.260 592.270 1143.400 600.030 ;
        RECT 1144.810 600.000 1145.090 600.030 ;
        RECT 924.240 591.950 924.500 592.270 ;
        RECT 1143.200 591.950 1143.460 592.270 ;
        RECT 924.300 2.400 924.440 591.950 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 944.910 592.520 945.230 592.580 ;
        RECT 1152.370 592.520 1152.690 592.580 ;
        RECT 944.910 592.380 1152.690 592.520 ;
        RECT 944.910 592.320 945.230 592.380 ;
        RECT 1152.370 592.320 1152.690 592.380 ;
        RECT 942.150 19.960 942.470 20.020 ;
        RECT 944.910 19.960 945.230 20.020 ;
        RECT 942.150 19.820 945.230 19.960 ;
        RECT 942.150 19.760 942.470 19.820 ;
        RECT 944.910 19.760 945.230 19.820 ;
      LAYER via ;
        RECT 944.940 592.320 945.200 592.580 ;
        RECT 1152.400 592.320 1152.660 592.580 ;
        RECT 942.180 19.760 942.440 20.020 ;
        RECT 944.940 19.760 945.200 20.020 ;
      LAYER met2 ;
        RECT 1154.010 600.170 1154.290 604.000 ;
        RECT 1152.460 600.030 1154.290 600.170 ;
        RECT 1152.460 592.610 1152.600 600.030 ;
        RECT 1154.010 600.000 1154.290 600.030 ;
        RECT 944.940 592.290 945.200 592.610 ;
        RECT 1152.400 592.290 1152.660 592.610 ;
        RECT 945.000 20.050 945.140 592.290 ;
        RECT 942.180 19.730 942.440 20.050 ;
        RECT 944.940 19.730 945.200 20.050 ;
        RECT 942.240 2.400 942.380 19.730 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1155.590 586.740 1155.910 586.800 ;
        RECT 1161.570 586.740 1161.890 586.800 ;
        RECT 1155.590 586.600 1161.890 586.740 ;
        RECT 1155.590 586.540 1155.910 586.600 ;
        RECT 1161.570 586.540 1161.890 586.600 ;
        RECT 960.090 18.940 960.410 19.000 ;
        RECT 1081.070 18.940 1081.390 19.000 ;
        RECT 960.090 18.800 1081.390 18.940 ;
        RECT 960.090 18.740 960.410 18.800 ;
        RECT 1081.070 18.740 1081.390 18.800 ;
        RECT 1081.070 16.560 1081.390 16.620 ;
        RECT 1155.590 16.560 1155.910 16.620 ;
        RECT 1081.070 16.420 1155.910 16.560 ;
        RECT 1081.070 16.360 1081.390 16.420 ;
        RECT 1155.590 16.360 1155.910 16.420 ;
      LAYER via ;
        RECT 1155.620 586.540 1155.880 586.800 ;
        RECT 1161.600 586.540 1161.860 586.800 ;
        RECT 960.120 18.740 960.380 19.000 ;
        RECT 1081.100 18.740 1081.360 19.000 ;
        RECT 1081.100 16.360 1081.360 16.620 ;
        RECT 1155.620 16.360 1155.880 16.620 ;
      LAYER met2 ;
        RECT 1163.210 600.170 1163.490 604.000 ;
        RECT 1161.660 600.030 1163.490 600.170 ;
        RECT 1161.660 586.830 1161.800 600.030 ;
        RECT 1163.210 600.000 1163.490 600.030 ;
        RECT 1155.620 586.510 1155.880 586.830 ;
        RECT 1161.600 586.510 1161.860 586.830 ;
        RECT 960.120 18.710 960.380 19.030 ;
        RECT 1081.100 18.710 1081.360 19.030 ;
        RECT 960.180 2.400 960.320 18.710 ;
        RECT 1081.160 16.650 1081.300 18.710 ;
        RECT 1155.680 16.650 1155.820 586.510 ;
        RECT 1081.100 16.330 1081.360 16.650 ;
        RECT 1155.620 16.330 1155.880 16.650 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1162.490 572.800 1162.810 572.860 ;
        RECT 1170.770 572.800 1171.090 572.860 ;
        RECT 1162.490 572.660 1171.090 572.800 ;
        RECT 1162.490 572.600 1162.810 572.660 ;
        RECT 1170.770 572.600 1171.090 572.660 ;
        RECT 1160.650 30.500 1160.970 30.560 ;
        RECT 1162.490 30.500 1162.810 30.560 ;
        RECT 1160.650 30.360 1162.810 30.500 ;
        RECT 1160.650 30.300 1160.970 30.360 ;
        RECT 1162.490 30.300 1162.810 30.360 ;
        RECT 1014.830 19.960 1015.150 20.020 ;
        RECT 1014.830 19.820 1147.540 19.960 ;
        RECT 1014.830 19.760 1015.150 19.820 ;
        RECT 1147.400 19.280 1147.540 19.820 ;
        RECT 1160.650 19.280 1160.970 19.340 ;
        RECT 1147.400 19.140 1160.970 19.280 ;
        RECT 1160.650 19.080 1160.970 19.140 ;
        RECT 978.030 18.600 978.350 18.660 ;
        RECT 1014.830 18.600 1015.150 18.660 ;
        RECT 978.030 18.460 1015.150 18.600 ;
        RECT 978.030 18.400 978.350 18.460 ;
        RECT 1014.830 18.400 1015.150 18.460 ;
      LAYER via ;
        RECT 1162.520 572.600 1162.780 572.860 ;
        RECT 1170.800 572.600 1171.060 572.860 ;
        RECT 1160.680 30.300 1160.940 30.560 ;
        RECT 1162.520 30.300 1162.780 30.560 ;
        RECT 1014.860 19.760 1015.120 20.020 ;
        RECT 1160.680 19.080 1160.940 19.340 ;
        RECT 978.060 18.400 978.320 18.660 ;
        RECT 1014.860 18.400 1015.120 18.660 ;
      LAYER met2 ;
        RECT 1172.410 600.170 1172.690 604.000 ;
        RECT 1170.860 600.030 1172.690 600.170 ;
        RECT 1170.860 572.890 1171.000 600.030 ;
        RECT 1172.410 600.000 1172.690 600.030 ;
        RECT 1162.520 572.570 1162.780 572.890 ;
        RECT 1170.800 572.570 1171.060 572.890 ;
        RECT 1162.580 30.590 1162.720 572.570 ;
        RECT 1160.680 30.270 1160.940 30.590 ;
        RECT 1162.520 30.270 1162.780 30.590 ;
        RECT 1014.860 19.730 1015.120 20.050 ;
        RECT 1014.920 18.690 1015.060 19.730 ;
        RECT 1160.740 19.370 1160.880 30.270 ;
        RECT 1160.680 19.050 1160.940 19.370 ;
        RECT 978.060 18.370 978.320 18.690 ;
        RECT 1014.860 18.370 1015.120 18.690 ;
        RECT 978.120 2.400 978.260 18.370 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 43.420 657.270 43.480 ;
        RECT 1007.930 43.420 1008.250 43.480 ;
        RECT 656.950 43.280 1008.250 43.420 ;
        RECT 656.950 43.220 657.270 43.280 ;
        RECT 1007.930 43.220 1008.250 43.280 ;
      LAYER via ;
        RECT 656.980 43.220 657.240 43.480 ;
        RECT 1007.960 43.220 1008.220 43.480 ;
      LAYER met2 ;
        RECT 1007.270 600.170 1007.550 604.000 ;
        RECT 1007.270 600.030 1008.160 600.170 ;
        RECT 1007.270 600.000 1007.550 600.030 ;
        RECT 1008.020 43.510 1008.160 600.030 ;
        RECT 656.980 43.190 657.240 43.510 ;
        RECT 1007.960 43.190 1008.220 43.510 ;
        RECT 657.040 2.400 657.180 43.190 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1000.110 592.860 1000.430 592.920 ;
        RECT 1179.970 592.860 1180.290 592.920 ;
        RECT 1000.110 592.720 1180.290 592.860 ;
        RECT 1000.110 592.660 1000.430 592.720 ;
        RECT 1179.970 592.660 1180.290 592.720 ;
        RECT 995.970 20.640 996.290 20.700 ;
        RECT 1000.110 20.640 1000.430 20.700 ;
        RECT 995.970 20.500 1000.430 20.640 ;
        RECT 995.970 20.440 996.290 20.500 ;
        RECT 1000.110 20.440 1000.430 20.500 ;
      LAYER via ;
        RECT 1000.140 592.660 1000.400 592.920 ;
        RECT 1180.000 592.660 1180.260 592.920 ;
        RECT 996.000 20.440 996.260 20.700 ;
        RECT 1000.140 20.440 1000.400 20.700 ;
      LAYER met2 ;
        RECT 1181.610 600.170 1181.890 604.000 ;
        RECT 1180.060 600.030 1181.890 600.170 ;
        RECT 1180.060 592.950 1180.200 600.030 ;
        RECT 1181.610 600.000 1181.890 600.030 ;
        RECT 1000.140 592.630 1000.400 592.950 ;
        RECT 1180.000 592.630 1180.260 592.950 ;
        RECT 1000.200 20.730 1000.340 592.630 ;
        RECT 996.000 20.410 996.260 20.730 ;
        RECT 1000.140 20.410 1000.400 20.730 ;
        RECT 996.060 2.400 996.200 20.410 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1186.870 569.400 1187.190 569.460 ;
        RECT 1189.170 569.400 1189.490 569.460 ;
        RECT 1186.870 569.260 1189.490 569.400 ;
        RECT 1186.870 569.200 1187.190 569.260 ;
        RECT 1189.170 569.200 1189.490 569.260 ;
        RECT 1124.770 19.620 1125.090 19.680 ;
        RECT 1124.770 19.480 1147.080 19.620 ;
        RECT 1124.770 19.420 1125.090 19.480 ;
        RECT 1146.940 18.940 1147.080 19.480 ;
        RECT 1186.870 18.940 1187.190 19.000 ;
        RECT 1146.940 18.800 1187.190 18.940 ;
        RECT 1186.870 18.740 1187.190 18.800 ;
        RECT 1015.290 18.600 1015.610 18.660 ;
        RECT 1124.770 18.600 1125.090 18.660 ;
        RECT 1015.290 18.460 1125.090 18.600 ;
        RECT 1015.290 18.400 1015.610 18.460 ;
        RECT 1124.770 18.400 1125.090 18.460 ;
      LAYER via ;
        RECT 1186.900 569.200 1187.160 569.460 ;
        RECT 1189.200 569.200 1189.460 569.460 ;
        RECT 1124.800 19.420 1125.060 19.680 ;
        RECT 1186.900 18.740 1187.160 19.000 ;
        RECT 1015.320 18.400 1015.580 18.660 ;
        RECT 1124.800 18.400 1125.060 18.660 ;
      LAYER met2 ;
        RECT 1190.810 600.170 1191.090 604.000 ;
        RECT 1189.260 600.030 1191.090 600.170 ;
        RECT 1189.260 569.490 1189.400 600.030 ;
        RECT 1190.810 600.000 1191.090 600.030 ;
        RECT 1186.900 569.170 1187.160 569.490 ;
        RECT 1189.200 569.170 1189.460 569.490 ;
        RECT 1124.800 19.390 1125.060 19.710 ;
        RECT 1124.860 18.690 1125.000 19.390 ;
        RECT 1186.960 19.030 1187.100 569.170 ;
        RECT 1186.900 18.710 1187.160 19.030 ;
        RECT 1015.320 18.370 1015.580 18.690 ;
        RECT 1124.800 18.370 1125.060 18.690 ;
        RECT 1015.380 18.090 1015.520 18.370 ;
        RECT 1013.540 17.950 1015.520 18.090 ;
        RECT 1013.540 2.400 1013.680 17.950 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1194.690 592.860 1195.010 592.920 ;
        RECT 1197.910 592.860 1198.230 592.920 ;
        RECT 1194.690 592.720 1198.230 592.860 ;
        RECT 1194.690 592.660 1195.010 592.720 ;
        RECT 1197.910 592.660 1198.230 592.720 ;
        RECT 1148.690 591.160 1149.010 591.220 ;
        RECT 1194.690 591.160 1195.010 591.220 ;
        RECT 1148.690 591.020 1195.010 591.160 ;
        RECT 1148.690 590.960 1149.010 591.020 ;
        RECT 1194.690 590.960 1195.010 591.020 ;
        RECT 1034.610 589.460 1034.930 589.520 ;
        RECT 1148.690 589.460 1149.010 589.520 ;
        RECT 1034.610 589.320 1149.010 589.460 ;
        RECT 1034.610 589.260 1034.930 589.320 ;
        RECT 1148.690 589.260 1149.010 589.320 ;
        RECT 1031.390 20.640 1031.710 20.700 ;
        RECT 1034.610 20.640 1034.930 20.700 ;
        RECT 1031.390 20.500 1034.930 20.640 ;
        RECT 1031.390 20.440 1031.710 20.500 ;
        RECT 1034.610 20.440 1034.930 20.500 ;
      LAYER via ;
        RECT 1194.720 592.660 1194.980 592.920 ;
        RECT 1197.940 592.660 1198.200 592.920 ;
        RECT 1148.720 590.960 1148.980 591.220 ;
        RECT 1194.720 590.960 1194.980 591.220 ;
        RECT 1034.640 589.260 1034.900 589.520 ;
        RECT 1148.720 589.260 1148.980 589.520 ;
        RECT 1031.420 20.440 1031.680 20.700 ;
        RECT 1034.640 20.440 1034.900 20.700 ;
      LAYER met2 ;
        RECT 1199.550 600.170 1199.830 604.000 ;
        RECT 1198.000 600.030 1199.830 600.170 ;
        RECT 1198.000 592.950 1198.140 600.030 ;
        RECT 1199.550 600.000 1199.830 600.030 ;
        RECT 1194.720 592.630 1194.980 592.950 ;
        RECT 1197.940 592.630 1198.200 592.950 ;
        RECT 1194.780 591.250 1194.920 592.630 ;
        RECT 1148.720 590.930 1148.980 591.250 ;
        RECT 1194.720 590.930 1194.980 591.250 ;
        RECT 1148.780 589.550 1148.920 590.930 ;
        RECT 1034.640 589.230 1034.900 589.550 ;
        RECT 1148.720 589.230 1148.980 589.550 ;
        RECT 1034.700 20.730 1034.840 589.230 ;
        RECT 1031.420 20.410 1031.680 20.730 ;
        RECT 1034.640 20.410 1034.900 20.730 ;
        RECT 1031.480 2.400 1031.620 20.410 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1049.330 20.300 1049.650 20.360 ;
        RECT 1208.030 20.300 1208.350 20.360 ;
        RECT 1049.330 20.160 1208.350 20.300 ;
        RECT 1049.330 20.100 1049.650 20.160 ;
        RECT 1208.030 20.100 1208.350 20.160 ;
      LAYER via ;
        RECT 1049.360 20.100 1049.620 20.360 ;
        RECT 1208.060 20.100 1208.320 20.360 ;
      LAYER met2 ;
        RECT 1208.750 600.170 1209.030 604.000 ;
        RECT 1208.120 600.030 1209.030 600.170 ;
        RECT 1208.120 20.390 1208.260 600.030 ;
        RECT 1208.750 600.000 1209.030 600.030 ;
        RECT 1049.360 20.070 1049.620 20.390 ;
        RECT 1208.060 20.070 1208.320 20.390 ;
        RECT 1049.420 2.400 1049.560 20.070 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1214.470 563.960 1214.790 564.020 ;
        RECT 1216.310 563.960 1216.630 564.020 ;
        RECT 1214.470 563.820 1216.630 563.960 ;
        RECT 1214.470 563.760 1214.790 563.820 ;
        RECT 1216.310 563.760 1216.630 563.820 ;
        RECT 1067.270 20.640 1067.590 20.700 ;
        RECT 1173.530 20.640 1173.850 20.700 ;
        RECT 1067.270 20.500 1173.850 20.640 ;
        RECT 1067.270 20.440 1067.590 20.500 ;
        RECT 1173.530 20.440 1173.850 20.500 ;
        RECT 1173.530 19.960 1173.850 20.020 ;
        RECT 1214.470 19.960 1214.790 20.020 ;
        RECT 1173.530 19.820 1214.790 19.960 ;
        RECT 1173.530 19.760 1173.850 19.820 ;
        RECT 1214.470 19.760 1214.790 19.820 ;
      LAYER via ;
        RECT 1214.500 563.760 1214.760 564.020 ;
        RECT 1216.340 563.760 1216.600 564.020 ;
        RECT 1067.300 20.440 1067.560 20.700 ;
        RECT 1173.560 20.440 1173.820 20.700 ;
        RECT 1173.560 19.760 1173.820 20.020 ;
        RECT 1214.500 19.760 1214.760 20.020 ;
      LAYER met2 ;
        RECT 1217.950 600.170 1218.230 604.000 ;
        RECT 1216.400 600.030 1218.230 600.170 ;
        RECT 1216.400 564.050 1216.540 600.030 ;
        RECT 1217.950 600.000 1218.230 600.030 ;
        RECT 1214.500 563.730 1214.760 564.050 ;
        RECT 1216.340 563.730 1216.600 564.050 ;
        RECT 1067.300 20.410 1067.560 20.730 ;
        RECT 1173.560 20.410 1173.820 20.730 ;
        RECT 1067.360 2.400 1067.500 20.410 ;
        RECT 1173.620 20.050 1173.760 20.410 ;
        RECT 1214.560 20.050 1214.700 563.730 ;
        RECT 1173.560 19.730 1173.820 20.050 ;
        RECT 1214.500 19.730 1214.760 20.050 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 588.440 1090.130 588.500 ;
        RECT 1225.510 588.440 1225.830 588.500 ;
        RECT 1089.810 588.300 1225.830 588.440 ;
        RECT 1089.810 588.240 1090.130 588.300 ;
        RECT 1225.510 588.240 1225.830 588.300 ;
        RECT 1085.210 19.620 1085.530 19.680 ;
        RECT 1089.810 19.620 1090.130 19.680 ;
        RECT 1085.210 19.480 1090.130 19.620 ;
        RECT 1085.210 19.420 1085.530 19.480 ;
        RECT 1089.810 19.420 1090.130 19.480 ;
      LAYER via ;
        RECT 1089.840 588.240 1090.100 588.500 ;
        RECT 1225.540 588.240 1225.800 588.500 ;
        RECT 1085.240 19.420 1085.500 19.680 ;
        RECT 1089.840 19.420 1090.100 19.680 ;
      LAYER met2 ;
        RECT 1227.150 600.170 1227.430 604.000 ;
        RECT 1225.600 600.030 1227.430 600.170 ;
        RECT 1225.600 588.530 1225.740 600.030 ;
        RECT 1227.150 600.000 1227.430 600.030 ;
        RECT 1089.840 588.210 1090.100 588.530 ;
        RECT 1225.540 588.210 1225.800 588.530 ;
        RECT 1089.900 19.710 1090.040 588.210 ;
        RECT 1085.240 19.390 1085.500 19.710 ;
        RECT 1089.840 19.390 1090.100 19.710 ;
        RECT 1085.300 2.400 1085.440 19.390 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1109.130 588.780 1109.450 588.840 ;
        RECT 1235.170 588.780 1235.490 588.840 ;
        RECT 1109.130 588.640 1235.490 588.780 ;
        RECT 1109.130 588.580 1109.450 588.640 ;
        RECT 1235.170 588.580 1235.490 588.640 ;
        RECT 1103.610 566.000 1103.930 566.060 ;
        RECT 1109.130 566.000 1109.450 566.060 ;
        RECT 1103.610 565.860 1109.450 566.000 ;
        RECT 1103.610 565.800 1103.930 565.860 ;
        RECT 1109.130 565.800 1109.450 565.860 ;
        RECT 1103.610 517.720 1103.930 517.780 ;
        RECT 1104.990 517.720 1105.310 517.780 ;
        RECT 1103.610 517.580 1105.310 517.720 ;
        RECT 1103.610 517.520 1103.930 517.580 ;
        RECT 1104.990 517.520 1105.310 517.580 ;
        RECT 1103.610 469.100 1103.930 469.160 ;
        RECT 1105.450 469.100 1105.770 469.160 ;
        RECT 1103.610 468.960 1105.770 469.100 ;
        RECT 1103.610 468.900 1103.930 468.960 ;
        RECT 1105.450 468.900 1105.770 468.960 ;
        RECT 1103.150 420.820 1103.470 420.880 ;
        RECT 1103.610 420.820 1103.930 420.880 ;
        RECT 1103.150 420.680 1103.930 420.820 ;
        RECT 1103.150 420.620 1103.470 420.680 ;
        RECT 1103.610 420.620 1103.930 420.680 ;
        RECT 1103.150 386.480 1103.470 386.540 ;
        RECT 1103.610 386.480 1103.930 386.540 ;
        RECT 1103.150 386.340 1103.930 386.480 ;
        RECT 1103.150 386.280 1103.470 386.340 ;
        RECT 1103.610 386.280 1103.930 386.340 ;
        RECT 1102.690 234.500 1103.010 234.560 ;
        RECT 1103.610 234.500 1103.930 234.560 ;
        RECT 1102.690 234.360 1103.930 234.500 ;
        RECT 1102.690 234.300 1103.010 234.360 ;
        RECT 1103.610 234.300 1103.930 234.360 ;
        RECT 1102.690 186.560 1103.010 186.620 ;
        RECT 1103.610 186.560 1103.930 186.620 ;
        RECT 1102.690 186.420 1103.930 186.560 ;
        RECT 1102.690 186.360 1103.010 186.420 ;
        RECT 1103.610 186.360 1103.930 186.420 ;
        RECT 1101.770 96.460 1102.090 96.520 ;
        RECT 1103.610 96.460 1103.930 96.520 ;
        RECT 1101.770 96.320 1103.930 96.460 ;
        RECT 1101.770 96.260 1102.090 96.320 ;
        RECT 1103.610 96.260 1103.930 96.320 ;
        RECT 1101.770 48.520 1102.090 48.580 ;
        RECT 1102.690 48.520 1103.010 48.580 ;
        RECT 1101.770 48.380 1103.010 48.520 ;
        RECT 1101.770 48.320 1102.090 48.380 ;
        RECT 1102.690 48.320 1103.010 48.380 ;
      LAYER via ;
        RECT 1109.160 588.580 1109.420 588.840 ;
        RECT 1235.200 588.580 1235.460 588.840 ;
        RECT 1103.640 565.800 1103.900 566.060 ;
        RECT 1109.160 565.800 1109.420 566.060 ;
        RECT 1103.640 517.520 1103.900 517.780 ;
        RECT 1105.020 517.520 1105.280 517.780 ;
        RECT 1103.640 468.900 1103.900 469.160 ;
        RECT 1105.480 468.900 1105.740 469.160 ;
        RECT 1103.180 420.620 1103.440 420.880 ;
        RECT 1103.640 420.620 1103.900 420.880 ;
        RECT 1103.180 386.280 1103.440 386.540 ;
        RECT 1103.640 386.280 1103.900 386.540 ;
        RECT 1102.720 234.300 1102.980 234.560 ;
        RECT 1103.640 234.300 1103.900 234.560 ;
        RECT 1102.720 186.360 1102.980 186.620 ;
        RECT 1103.640 186.360 1103.900 186.620 ;
        RECT 1101.800 96.260 1102.060 96.520 ;
        RECT 1103.640 96.260 1103.900 96.520 ;
        RECT 1101.800 48.320 1102.060 48.580 ;
        RECT 1102.720 48.320 1102.980 48.580 ;
      LAYER met2 ;
        RECT 1236.350 600.170 1236.630 604.000 ;
        RECT 1235.260 600.030 1236.630 600.170 ;
        RECT 1235.260 588.870 1235.400 600.030 ;
        RECT 1236.350 600.000 1236.630 600.030 ;
        RECT 1109.160 588.550 1109.420 588.870 ;
        RECT 1235.200 588.550 1235.460 588.870 ;
        RECT 1109.220 566.090 1109.360 588.550 ;
        RECT 1103.640 565.770 1103.900 566.090 ;
        RECT 1109.160 565.770 1109.420 566.090 ;
        RECT 1103.700 565.605 1103.840 565.770 ;
        RECT 1103.630 565.235 1103.910 565.605 ;
        RECT 1105.010 565.235 1105.290 565.605 ;
        RECT 1105.080 517.810 1105.220 565.235 ;
        RECT 1103.640 517.490 1103.900 517.810 ;
        RECT 1105.020 517.490 1105.280 517.810 ;
        RECT 1103.700 469.190 1103.840 517.490 ;
        RECT 1103.640 468.870 1103.900 469.190 ;
        RECT 1105.480 468.870 1105.740 469.190 ;
        RECT 1105.540 421.445 1105.680 468.870 ;
        RECT 1103.630 421.075 1103.910 421.445 ;
        RECT 1105.470 421.075 1105.750 421.445 ;
        RECT 1103.700 420.910 1103.840 421.075 ;
        RECT 1103.180 420.590 1103.440 420.910 ;
        RECT 1103.640 420.590 1103.900 420.910 ;
        RECT 1103.240 386.570 1103.380 420.590 ;
        RECT 1103.180 386.250 1103.440 386.570 ;
        RECT 1103.640 386.250 1103.900 386.570 ;
        RECT 1103.700 234.590 1103.840 386.250 ;
        RECT 1102.720 234.270 1102.980 234.590 ;
        RECT 1103.640 234.270 1103.900 234.590 ;
        RECT 1102.780 186.650 1102.920 234.270 ;
        RECT 1102.720 186.330 1102.980 186.650 ;
        RECT 1103.640 186.330 1103.900 186.650 ;
        RECT 1103.700 96.550 1103.840 186.330 ;
        RECT 1101.800 96.230 1102.060 96.550 ;
        RECT 1103.640 96.230 1103.900 96.550 ;
        RECT 1101.860 48.610 1102.000 96.230 ;
        RECT 1101.800 48.290 1102.060 48.610 ;
        RECT 1102.720 48.290 1102.980 48.610 ;
        RECT 1102.780 2.400 1102.920 48.290 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
      LAYER via2 ;
        RECT 1103.630 565.280 1103.910 565.560 ;
        RECT 1105.010 565.280 1105.290 565.560 ;
        RECT 1103.630 421.120 1103.910 421.400 ;
        RECT 1105.470 421.120 1105.750 421.400 ;
      LAYER met3 ;
        RECT 1103.605 565.570 1103.935 565.585 ;
        RECT 1104.985 565.570 1105.315 565.585 ;
        RECT 1103.605 565.270 1105.315 565.570 ;
        RECT 1103.605 565.255 1103.935 565.270 ;
        RECT 1104.985 565.255 1105.315 565.270 ;
        RECT 1103.605 421.410 1103.935 421.425 ;
        RECT 1105.445 421.410 1105.775 421.425 ;
        RECT 1103.605 421.110 1105.775 421.410 ;
        RECT 1103.605 421.095 1103.935 421.110 ;
        RECT 1105.445 421.095 1105.775 421.110 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1196.990 590.480 1197.310 590.540 ;
        RECT 1243.910 590.480 1244.230 590.540 ;
        RECT 1196.990 590.340 1244.230 590.480 ;
        RECT 1196.990 590.280 1197.310 590.340 ;
        RECT 1243.910 590.280 1244.230 590.340 ;
        RECT 1149.150 589.460 1149.470 589.520 ;
        RECT 1196.990 589.460 1197.310 589.520 ;
        RECT 1149.150 589.320 1197.310 589.460 ;
        RECT 1149.150 589.260 1149.470 589.320 ;
        RECT 1196.990 589.260 1197.310 589.320 ;
        RECT 1124.310 582.320 1124.630 582.380 ;
        RECT 1149.150 582.320 1149.470 582.380 ;
        RECT 1124.310 582.180 1149.470 582.320 ;
        RECT 1124.310 582.120 1124.630 582.180 ;
        RECT 1149.150 582.120 1149.470 582.180 ;
        RECT 1120.630 19.620 1120.950 19.680 ;
        RECT 1124.310 19.620 1124.630 19.680 ;
        RECT 1120.630 19.480 1124.630 19.620 ;
        RECT 1120.630 19.420 1120.950 19.480 ;
        RECT 1124.310 19.420 1124.630 19.480 ;
      LAYER via ;
        RECT 1197.020 590.280 1197.280 590.540 ;
        RECT 1243.940 590.280 1244.200 590.540 ;
        RECT 1149.180 589.260 1149.440 589.520 ;
        RECT 1197.020 589.260 1197.280 589.520 ;
        RECT 1124.340 582.120 1124.600 582.380 ;
        RECT 1149.180 582.120 1149.440 582.380 ;
        RECT 1120.660 19.420 1120.920 19.680 ;
        RECT 1124.340 19.420 1124.600 19.680 ;
      LAYER met2 ;
        RECT 1245.550 600.170 1245.830 604.000 ;
        RECT 1244.000 600.030 1245.830 600.170 ;
        RECT 1244.000 590.570 1244.140 600.030 ;
        RECT 1245.550 600.000 1245.830 600.030 ;
        RECT 1197.020 590.250 1197.280 590.570 ;
        RECT 1243.940 590.250 1244.200 590.570 ;
        RECT 1197.080 589.550 1197.220 590.250 ;
        RECT 1149.180 589.230 1149.440 589.550 ;
        RECT 1197.020 589.230 1197.280 589.550 ;
        RECT 1149.240 582.410 1149.380 589.230 ;
        RECT 1124.340 582.090 1124.600 582.410 ;
        RECT 1149.180 582.090 1149.440 582.410 ;
        RECT 1124.400 19.710 1124.540 582.090 ;
        RECT 1120.660 19.390 1120.920 19.710 ;
        RECT 1124.340 19.390 1124.600 19.710 ;
        RECT 1120.720 2.400 1120.860 19.390 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1144.550 590.140 1144.870 590.200 ;
        RECT 1253.110 590.140 1253.430 590.200 ;
        RECT 1144.550 590.000 1253.430 590.140 ;
        RECT 1144.550 589.940 1144.870 590.000 ;
        RECT 1253.110 589.940 1253.430 590.000 ;
        RECT 1144.550 62.260 1144.870 62.520 ;
        RECT 1144.640 61.840 1144.780 62.260 ;
        RECT 1144.550 61.580 1144.870 61.840 ;
        RECT 1138.570 14.520 1138.890 14.580 ;
        RECT 1144.550 14.520 1144.870 14.580 ;
        RECT 1138.570 14.380 1144.870 14.520 ;
        RECT 1138.570 14.320 1138.890 14.380 ;
        RECT 1144.550 14.320 1144.870 14.380 ;
      LAYER via ;
        RECT 1144.580 589.940 1144.840 590.200 ;
        RECT 1253.140 589.940 1253.400 590.200 ;
        RECT 1144.580 62.260 1144.840 62.520 ;
        RECT 1144.580 61.580 1144.840 61.840 ;
        RECT 1138.600 14.320 1138.860 14.580 ;
        RECT 1144.580 14.320 1144.840 14.580 ;
      LAYER met2 ;
        RECT 1254.750 600.170 1255.030 604.000 ;
        RECT 1253.200 600.030 1255.030 600.170 ;
        RECT 1253.200 590.230 1253.340 600.030 ;
        RECT 1254.750 600.000 1255.030 600.030 ;
        RECT 1144.580 589.910 1144.840 590.230 ;
        RECT 1253.140 589.910 1253.400 590.230 ;
        RECT 1144.640 62.550 1144.780 589.910 ;
        RECT 1144.580 62.230 1144.840 62.550 ;
        RECT 1144.580 61.550 1144.840 61.870 ;
        RECT 1144.640 14.610 1144.780 61.550 ;
        RECT 1138.600 14.290 1138.860 14.610 ;
        RECT 1144.580 14.290 1144.840 14.610 ;
        RECT 1138.660 2.400 1138.800 14.290 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.810 590.820 1159.130 590.880 ;
        RECT 1262.770 590.820 1263.090 590.880 ;
        RECT 1158.810 590.680 1263.090 590.820 ;
        RECT 1158.810 590.620 1159.130 590.680 ;
        RECT 1262.770 590.620 1263.090 590.680 ;
        RECT 1156.510 19.960 1156.830 20.020 ;
        RECT 1158.810 19.960 1159.130 20.020 ;
        RECT 1156.510 19.820 1159.130 19.960 ;
        RECT 1156.510 19.760 1156.830 19.820 ;
        RECT 1158.810 19.760 1159.130 19.820 ;
      LAYER via ;
        RECT 1158.840 590.620 1159.100 590.880 ;
        RECT 1262.800 590.620 1263.060 590.880 ;
        RECT 1156.540 19.760 1156.800 20.020 ;
        RECT 1158.840 19.760 1159.100 20.020 ;
      LAYER met2 ;
        RECT 1263.950 600.170 1264.230 604.000 ;
        RECT 1262.860 600.030 1264.230 600.170 ;
        RECT 1262.860 590.910 1263.000 600.030 ;
        RECT 1263.950 600.000 1264.230 600.030 ;
        RECT 1158.840 590.590 1159.100 590.910 ;
        RECT 1262.800 590.590 1263.060 590.910 ;
        RECT 1158.900 20.050 1159.040 590.590 ;
        RECT 1156.540 19.730 1156.800 20.050 ;
        RECT 1158.840 19.730 1159.100 20.050 ;
        RECT 1156.600 2.400 1156.740 19.730 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 674.430 43.080 674.750 43.140 ;
        RECT 1014.370 43.080 1014.690 43.140 ;
        RECT 674.430 42.940 1014.690 43.080 ;
        RECT 674.430 42.880 674.750 42.940 ;
        RECT 1014.370 42.880 1014.690 42.940 ;
      LAYER via ;
        RECT 674.460 42.880 674.720 43.140 ;
        RECT 1014.400 42.880 1014.660 43.140 ;
      LAYER met2 ;
        RECT 1016.470 600.170 1016.750 604.000 ;
        RECT 1014.460 600.030 1016.750 600.170 ;
        RECT 1014.460 43.170 1014.600 600.030 ;
        RECT 1016.470 600.000 1016.750 600.030 ;
        RECT 674.460 42.850 674.720 43.170 ;
        RECT 1014.400 42.850 1014.660 43.170 ;
        RECT 674.520 2.400 674.660 42.850 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1202.050 592.180 1202.370 592.240 ;
        RECT 1271.510 592.180 1271.830 592.240 ;
        RECT 1202.050 592.040 1271.830 592.180 ;
        RECT 1202.050 591.980 1202.370 592.040 ;
        RECT 1271.510 591.980 1271.830 592.040 ;
        RECT 1179.510 588.100 1179.830 588.160 ;
        RECT 1202.050 588.100 1202.370 588.160 ;
        RECT 1179.510 587.960 1202.370 588.100 ;
        RECT 1179.510 587.900 1179.830 587.960 ;
        RECT 1202.050 587.900 1202.370 587.960 ;
        RECT 1173.990 20.640 1174.310 20.700 ;
        RECT 1179.510 20.640 1179.830 20.700 ;
        RECT 1173.990 20.500 1179.830 20.640 ;
        RECT 1173.990 20.440 1174.310 20.500 ;
        RECT 1179.510 20.440 1179.830 20.500 ;
      LAYER via ;
        RECT 1202.080 591.980 1202.340 592.240 ;
        RECT 1271.540 591.980 1271.800 592.240 ;
        RECT 1179.540 587.900 1179.800 588.160 ;
        RECT 1202.080 587.900 1202.340 588.160 ;
        RECT 1174.020 20.440 1174.280 20.700 ;
        RECT 1179.540 20.440 1179.800 20.700 ;
      LAYER met2 ;
        RECT 1273.150 600.170 1273.430 604.000 ;
        RECT 1271.600 600.030 1273.430 600.170 ;
        RECT 1271.600 592.270 1271.740 600.030 ;
        RECT 1273.150 600.000 1273.430 600.030 ;
        RECT 1202.080 591.950 1202.340 592.270 ;
        RECT 1271.540 591.950 1271.800 592.270 ;
        RECT 1202.140 588.190 1202.280 591.950 ;
        RECT 1179.540 587.870 1179.800 588.190 ;
        RECT 1202.080 587.870 1202.340 588.190 ;
        RECT 1179.600 20.730 1179.740 587.870 ;
        RECT 1174.020 20.410 1174.280 20.730 ;
        RECT 1179.540 20.410 1179.800 20.730 ;
        RECT 1174.080 2.400 1174.220 20.410 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1193.310 593.200 1193.630 593.260 ;
        RECT 1280.710 593.200 1281.030 593.260 ;
        RECT 1193.310 593.060 1281.030 593.200 ;
        RECT 1193.310 593.000 1193.630 593.060 ;
        RECT 1280.710 593.000 1281.030 593.060 ;
        RECT 1191.930 2.960 1192.250 3.020 ;
        RECT 1193.310 2.960 1193.630 3.020 ;
        RECT 1191.930 2.820 1193.630 2.960 ;
        RECT 1191.930 2.760 1192.250 2.820 ;
        RECT 1193.310 2.760 1193.630 2.820 ;
      LAYER via ;
        RECT 1193.340 593.000 1193.600 593.260 ;
        RECT 1280.740 593.000 1281.000 593.260 ;
        RECT 1191.960 2.760 1192.220 3.020 ;
        RECT 1193.340 2.760 1193.600 3.020 ;
      LAYER met2 ;
        RECT 1282.350 600.170 1282.630 604.000 ;
        RECT 1280.800 600.030 1282.630 600.170 ;
        RECT 1280.800 593.290 1280.940 600.030 ;
        RECT 1282.350 600.000 1282.630 600.030 ;
        RECT 1193.340 592.970 1193.600 593.290 ;
        RECT 1280.740 592.970 1281.000 593.290 ;
        RECT 1193.400 3.050 1193.540 592.970 ;
        RECT 1191.960 2.730 1192.220 3.050 ;
        RECT 1193.340 2.730 1193.600 3.050 ;
        RECT 1192.020 2.400 1192.160 2.730 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1214.010 588.100 1214.330 588.160 ;
        RECT 1290.830 588.100 1291.150 588.160 ;
        RECT 1214.010 587.960 1291.150 588.100 ;
        RECT 1214.010 587.900 1214.330 587.960 ;
        RECT 1290.830 587.900 1291.150 587.960 ;
        RECT 1209.870 16.220 1210.190 16.280 ;
        RECT 1214.010 16.220 1214.330 16.280 ;
        RECT 1209.870 16.080 1214.330 16.220 ;
        RECT 1209.870 16.020 1210.190 16.080 ;
        RECT 1214.010 16.020 1214.330 16.080 ;
      LAYER via ;
        RECT 1214.040 587.900 1214.300 588.160 ;
        RECT 1290.860 587.900 1291.120 588.160 ;
        RECT 1209.900 16.020 1210.160 16.280 ;
        RECT 1214.040 16.020 1214.300 16.280 ;
      LAYER met2 ;
        RECT 1291.550 600.170 1291.830 604.000 ;
        RECT 1290.920 600.030 1291.830 600.170 ;
        RECT 1290.920 588.190 1291.060 600.030 ;
        RECT 1291.550 600.000 1291.830 600.030 ;
        RECT 1214.040 587.870 1214.300 588.190 ;
        RECT 1290.860 587.870 1291.120 588.190 ;
        RECT 1214.100 16.310 1214.240 587.870 ;
        RECT 1209.900 15.990 1210.160 16.310 ;
        RECT 1214.040 15.990 1214.300 16.310 ;
        RECT 1209.960 2.400 1210.100 15.990 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 588.440 1228.130 588.500 ;
        RECT 1299.110 588.440 1299.430 588.500 ;
        RECT 1227.810 588.300 1299.430 588.440 ;
        RECT 1227.810 588.240 1228.130 588.300 ;
        RECT 1299.110 588.240 1299.430 588.300 ;
      LAYER via ;
        RECT 1227.840 588.240 1228.100 588.500 ;
        RECT 1299.140 588.240 1299.400 588.500 ;
      LAYER met2 ;
        RECT 1300.750 600.170 1301.030 604.000 ;
        RECT 1299.200 600.030 1301.030 600.170 ;
        RECT 1299.200 588.530 1299.340 600.030 ;
        RECT 1300.750 600.000 1301.030 600.030 ;
        RECT 1227.840 588.210 1228.100 588.530 ;
        RECT 1299.140 588.210 1299.400 588.530 ;
        RECT 1227.900 2.400 1228.040 588.210 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 590.480 1248.830 590.540 ;
        RECT 1308.310 590.480 1308.630 590.540 ;
        RECT 1248.510 590.340 1308.630 590.480 ;
        RECT 1248.510 590.280 1248.830 590.340 ;
        RECT 1308.310 590.280 1308.630 590.340 ;
        RECT 1245.750 16.560 1246.070 16.620 ;
        RECT 1248.510 16.560 1248.830 16.620 ;
        RECT 1245.750 16.420 1248.830 16.560 ;
        RECT 1245.750 16.360 1246.070 16.420 ;
        RECT 1248.510 16.360 1248.830 16.420 ;
      LAYER via ;
        RECT 1248.540 590.280 1248.800 590.540 ;
        RECT 1308.340 590.280 1308.600 590.540 ;
        RECT 1245.780 16.360 1246.040 16.620 ;
        RECT 1248.540 16.360 1248.800 16.620 ;
      LAYER met2 ;
        RECT 1309.950 600.170 1310.230 604.000 ;
        RECT 1308.400 600.030 1310.230 600.170 ;
        RECT 1308.400 590.570 1308.540 600.030 ;
        RECT 1309.950 600.000 1310.230 600.030 ;
        RECT 1248.540 590.250 1248.800 590.570 ;
        RECT 1308.340 590.250 1308.600 590.570 ;
        RECT 1248.600 16.650 1248.740 590.250 ;
        RECT 1245.780 16.330 1246.040 16.650 ;
        RECT 1248.540 16.330 1248.800 16.650 ;
        RECT 1245.840 2.400 1245.980 16.330 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1269.210 591.500 1269.530 591.560 ;
        RECT 1317.970 591.500 1318.290 591.560 ;
        RECT 1269.210 591.360 1318.290 591.500 ;
        RECT 1269.210 591.300 1269.530 591.360 ;
        RECT 1317.970 591.300 1318.290 591.360 ;
        RECT 1263.230 16.560 1263.550 16.620 ;
        RECT 1269.210 16.560 1269.530 16.620 ;
        RECT 1263.230 16.420 1269.530 16.560 ;
        RECT 1263.230 16.360 1263.550 16.420 ;
        RECT 1269.210 16.360 1269.530 16.420 ;
      LAYER via ;
        RECT 1269.240 591.300 1269.500 591.560 ;
        RECT 1318.000 591.300 1318.260 591.560 ;
        RECT 1263.260 16.360 1263.520 16.620 ;
        RECT 1269.240 16.360 1269.500 16.620 ;
      LAYER met2 ;
        RECT 1319.150 600.170 1319.430 604.000 ;
        RECT 1318.060 600.030 1319.430 600.170 ;
        RECT 1318.060 591.590 1318.200 600.030 ;
        RECT 1319.150 600.000 1319.430 600.030 ;
        RECT 1269.240 591.270 1269.500 591.590 ;
        RECT 1318.000 591.270 1318.260 591.590 ;
        RECT 1269.300 16.650 1269.440 591.270 ;
        RECT 1263.260 16.330 1263.520 16.650 ;
        RECT 1269.240 16.330 1269.500 16.650 ;
        RECT 1263.320 2.400 1263.460 16.330 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 591.840 1283.330 591.900 ;
        RECT 1326.250 591.840 1326.570 591.900 ;
        RECT 1283.010 591.700 1326.570 591.840 ;
        RECT 1283.010 591.640 1283.330 591.700 ;
        RECT 1326.250 591.640 1326.570 591.700 ;
      LAYER via ;
        RECT 1283.040 591.640 1283.300 591.900 ;
        RECT 1326.280 591.640 1326.540 591.900 ;
      LAYER met2 ;
        RECT 1327.890 600.170 1328.170 604.000 ;
        RECT 1326.340 600.030 1328.170 600.170 ;
        RECT 1326.340 591.930 1326.480 600.030 ;
        RECT 1327.890 600.000 1328.170 600.030 ;
        RECT 1283.040 591.610 1283.300 591.930 ;
        RECT 1326.280 591.610 1326.540 591.930 ;
        RECT 1283.100 16.730 1283.240 591.610 ;
        RECT 1281.260 16.590 1283.240 16.730 ;
        RECT 1281.260 2.400 1281.400 16.590 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.710 586.740 1304.030 586.800 ;
        RECT 1335.450 586.740 1335.770 586.800 ;
        RECT 1303.710 586.600 1335.770 586.740 ;
        RECT 1303.710 586.540 1304.030 586.600 ;
        RECT 1335.450 586.540 1335.770 586.600 ;
        RECT 1299.110 17.580 1299.430 17.640 ;
        RECT 1303.710 17.580 1304.030 17.640 ;
        RECT 1299.110 17.440 1304.030 17.580 ;
        RECT 1299.110 17.380 1299.430 17.440 ;
        RECT 1303.710 17.380 1304.030 17.440 ;
      LAYER via ;
        RECT 1303.740 586.540 1304.000 586.800 ;
        RECT 1335.480 586.540 1335.740 586.800 ;
        RECT 1299.140 17.380 1299.400 17.640 ;
        RECT 1303.740 17.380 1304.000 17.640 ;
      LAYER met2 ;
        RECT 1337.090 600.170 1337.370 604.000 ;
        RECT 1335.540 600.030 1337.370 600.170 ;
        RECT 1335.540 586.830 1335.680 600.030 ;
        RECT 1337.090 600.000 1337.370 600.030 ;
        RECT 1303.740 586.510 1304.000 586.830 ;
        RECT 1335.480 586.510 1335.740 586.830 ;
        RECT 1303.800 17.670 1303.940 586.510 ;
        RECT 1299.140 17.350 1299.400 17.670 ;
        RECT 1303.740 17.350 1304.000 17.670 ;
        RECT 1299.200 2.400 1299.340 17.350 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.990 590.140 1335.310 590.200 ;
        RECT 1345.570 590.140 1345.890 590.200 ;
        RECT 1334.990 590.000 1345.890 590.140 ;
        RECT 1334.990 589.940 1335.310 590.000 ;
        RECT 1345.570 589.940 1345.890 590.000 ;
        RECT 1317.050 17.920 1317.370 17.980 ;
        RECT 1334.990 17.920 1335.310 17.980 ;
        RECT 1317.050 17.780 1335.310 17.920 ;
        RECT 1317.050 17.720 1317.370 17.780 ;
        RECT 1334.990 17.720 1335.310 17.780 ;
      LAYER via ;
        RECT 1335.020 589.940 1335.280 590.200 ;
        RECT 1345.600 589.940 1345.860 590.200 ;
        RECT 1317.080 17.720 1317.340 17.980 ;
        RECT 1335.020 17.720 1335.280 17.980 ;
      LAYER met2 ;
        RECT 1346.290 600.170 1346.570 604.000 ;
        RECT 1345.660 600.030 1346.570 600.170 ;
        RECT 1345.660 590.230 1345.800 600.030 ;
        RECT 1346.290 600.000 1346.570 600.030 ;
        RECT 1335.020 589.910 1335.280 590.230 ;
        RECT 1345.600 589.910 1345.860 590.230 ;
        RECT 1335.080 18.010 1335.220 589.910 ;
        RECT 1317.080 17.690 1317.340 18.010 ;
        RECT 1335.020 17.690 1335.280 18.010 ;
        RECT 1317.140 2.400 1317.280 17.690 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 590.820 1338.530 590.880 ;
        RECT 1353.850 590.820 1354.170 590.880 ;
        RECT 1338.210 590.680 1354.170 590.820 ;
        RECT 1338.210 590.620 1338.530 590.680 ;
        RECT 1353.850 590.620 1354.170 590.680 ;
        RECT 1334.990 17.240 1335.310 17.300 ;
        RECT 1338.210 17.240 1338.530 17.300 ;
        RECT 1334.990 17.100 1338.530 17.240 ;
        RECT 1334.990 17.040 1335.310 17.100 ;
        RECT 1338.210 17.040 1338.530 17.100 ;
      LAYER via ;
        RECT 1338.240 590.620 1338.500 590.880 ;
        RECT 1353.880 590.620 1354.140 590.880 ;
        RECT 1335.020 17.040 1335.280 17.300 ;
        RECT 1338.240 17.040 1338.500 17.300 ;
      LAYER met2 ;
        RECT 1355.490 600.170 1355.770 604.000 ;
        RECT 1353.940 600.030 1355.770 600.170 ;
        RECT 1353.940 590.910 1354.080 600.030 ;
        RECT 1355.490 600.000 1355.770 600.030 ;
        RECT 1338.240 590.590 1338.500 590.910 ;
        RECT 1353.880 590.590 1354.140 590.910 ;
        RECT 1338.300 17.330 1338.440 590.590 ;
        RECT 1335.020 17.010 1335.280 17.330 ;
        RECT 1338.240 17.010 1338.500 17.330 ;
        RECT 1335.080 2.400 1335.220 17.010 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1021.270 569.400 1021.590 569.460 ;
        RECT 1024.030 569.400 1024.350 569.460 ;
        RECT 1021.270 569.260 1024.350 569.400 ;
        RECT 1021.270 569.200 1021.590 569.260 ;
        RECT 1024.030 569.200 1024.350 569.260 ;
        RECT 692.370 24.040 692.690 24.100 ;
        RECT 1021.270 24.040 1021.590 24.100 ;
        RECT 692.370 23.900 1021.590 24.040 ;
        RECT 692.370 23.840 692.690 23.900 ;
        RECT 1021.270 23.840 1021.590 23.900 ;
      LAYER via ;
        RECT 1021.300 569.200 1021.560 569.460 ;
        RECT 1024.060 569.200 1024.320 569.460 ;
        RECT 692.400 23.840 692.660 24.100 ;
        RECT 1021.300 23.840 1021.560 24.100 ;
      LAYER met2 ;
        RECT 1025.670 600.170 1025.950 604.000 ;
        RECT 1024.120 600.030 1025.950 600.170 ;
        RECT 1024.120 569.490 1024.260 600.030 ;
        RECT 1025.670 600.000 1025.950 600.030 ;
        RECT 1021.300 569.170 1021.560 569.490 ;
        RECT 1024.060 569.170 1024.320 569.490 ;
        RECT 1021.360 24.130 1021.500 569.170 ;
        RECT 692.400 23.810 692.660 24.130 ;
        RECT 1021.300 23.810 1021.560 24.130 ;
        RECT 692.460 2.400 692.600 23.810 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1358.450 586.740 1358.770 586.800 ;
        RECT 1363.050 586.740 1363.370 586.800 ;
        RECT 1358.450 586.600 1363.370 586.740 ;
        RECT 1358.450 586.540 1358.770 586.600 ;
        RECT 1363.050 586.540 1363.370 586.600 ;
        RECT 1352.470 20.640 1352.790 20.700 ;
        RECT 1357.990 20.640 1358.310 20.700 ;
        RECT 1352.470 20.500 1358.310 20.640 ;
        RECT 1352.470 20.440 1352.790 20.500 ;
        RECT 1357.990 20.440 1358.310 20.500 ;
      LAYER via ;
        RECT 1358.480 586.540 1358.740 586.800 ;
        RECT 1363.080 586.540 1363.340 586.800 ;
        RECT 1352.500 20.440 1352.760 20.700 ;
        RECT 1358.020 20.440 1358.280 20.700 ;
      LAYER met2 ;
        RECT 1364.690 600.170 1364.970 604.000 ;
        RECT 1363.140 600.030 1364.970 600.170 ;
        RECT 1363.140 586.830 1363.280 600.030 ;
        RECT 1364.690 600.000 1364.970 600.030 ;
        RECT 1358.480 586.510 1358.740 586.830 ;
        RECT 1363.080 586.510 1363.340 586.830 ;
        RECT 1358.540 24.890 1358.680 586.510 ;
        RECT 1358.080 24.750 1358.680 24.890 ;
        RECT 1358.080 20.730 1358.220 24.750 ;
        RECT 1352.500 20.410 1352.760 20.730 ;
        RECT 1358.020 20.410 1358.280 20.730 ;
        RECT 1352.560 2.400 1352.700 20.410 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.410 20.640 1370.730 20.700 ;
        RECT 1373.630 20.640 1373.950 20.700 ;
        RECT 1370.410 20.500 1373.950 20.640 ;
        RECT 1370.410 20.440 1370.730 20.500 ;
        RECT 1373.630 20.440 1373.950 20.500 ;
      LAYER via ;
        RECT 1370.440 20.440 1370.700 20.700 ;
        RECT 1373.660 20.440 1373.920 20.700 ;
      LAYER met2 ;
        RECT 1373.890 600.000 1374.170 604.000 ;
        RECT 1373.950 598.810 1374.090 600.000 ;
        RECT 1373.720 598.670 1374.090 598.810 ;
        RECT 1373.720 20.730 1373.860 598.670 ;
        RECT 1370.440 20.410 1370.700 20.730 ;
        RECT 1373.660 20.410 1373.920 20.730 ;
        RECT 1370.500 2.400 1370.640 20.410 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1384.670 586.740 1384.990 586.800 ;
        RECT 1386.510 586.740 1386.830 586.800 ;
        RECT 1384.670 586.600 1386.830 586.740 ;
        RECT 1384.670 586.540 1384.990 586.600 ;
        RECT 1386.510 586.540 1386.830 586.600 ;
        RECT 1386.510 20.640 1386.830 20.700 ;
        RECT 1388.350 20.640 1388.670 20.700 ;
        RECT 1386.510 20.500 1388.670 20.640 ;
        RECT 1386.510 20.440 1386.830 20.500 ;
        RECT 1388.350 20.440 1388.670 20.500 ;
      LAYER via ;
        RECT 1384.700 586.540 1384.960 586.800 ;
        RECT 1386.540 586.540 1386.800 586.800 ;
        RECT 1386.540 20.440 1386.800 20.700 ;
        RECT 1388.380 20.440 1388.640 20.700 ;
      LAYER met2 ;
        RECT 1383.090 600.170 1383.370 604.000 ;
        RECT 1383.090 600.030 1384.900 600.170 ;
        RECT 1383.090 600.000 1383.370 600.030 ;
        RECT 1384.760 586.830 1384.900 600.030 ;
        RECT 1384.700 586.510 1384.960 586.830 ;
        RECT 1386.540 586.510 1386.800 586.830 ;
        RECT 1386.600 20.730 1386.740 586.510 ;
        RECT 1386.540 20.410 1386.800 20.730 ;
        RECT 1388.380 20.410 1388.640 20.730 ;
        RECT 1388.440 2.400 1388.580 20.410 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1392.950 589.120 1393.270 589.180 ;
        RECT 1401.690 589.120 1402.010 589.180 ;
        RECT 1392.950 588.980 1402.010 589.120 ;
        RECT 1392.950 588.920 1393.270 588.980 ;
        RECT 1401.690 588.920 1402.010 588.980 ;
        RECT 1401.690 2.960 1402.010 3.020 ;
        RECT 1406.290 2.960 1406.610 3.020 ;
        RECT 1401.690 2.820 1406.610 2.960 ;
        RECT 1401.690 2.760 1402.010 2.820 ;
        RECT 1406.290 2.760 1406.610 2.820 ;
      LAYER via ;
        RECT 1392.980 588.920 1393.240 589.180 ;
        RECT 1401.720 588.920 1401.980 589.180 ;
        RECT 1401.720 2.760 1401.980 3.020 ;
        RECT 1406.320 2.760 1406.580 3.020 ;
      LAYER met2 ;
        RECT 1392.290 600.170 1392.570 604.000 ;
        RECT 1392.290 600.030 1393.180 600.170 ;
        RECT 1392.290 600.000 1392.570 600.030 ;
        RECT 1393.040 589.210 1393.180 600.030 ;
        RECT 1392.980 588.890 1393.240 589.210 ;
        RECT 1401.720 588.890 1401.980 589.210 ;
        RECT 1401.780 3.050 1401.920 588.890 ;
        RECT 1401.720 2.730 1401.980 3.050 ;
        RECT 1406.320 2.730 1406.580 3.050 ;
        RECT 1406.380 2.400 1406.520 2.730 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1403.070 587.420 1403.390 587.480 ;
        RECT 1406.750 587.420 1407.070 587.480 ;
        RECT 1403.070 587.280 1407.070 587.420 ;
        RECT 1403.070 587.220 1403.390 587.280 ;
        RECT 1406.750 587.220 1407.070 587.280 ;
        RECT 1406.750 15.880 1407.070 15.940 ;
        RECT 1423.770 15.880 1424.090 15.940 ;
        RECT 1406.750 15.740 1424.090 15.880 ;
        RECT 1406.750 15.680 1407.070 15.740 ;
        RECT 1423.770 15.680 1424.090 15.740 ;
      LAYER via ;
        RECT 1403.100 587.220 1403.360 587.480 ;
        RECT 1406.780 587.220 1407.040 587.480 ;
        RECT 1406.780 15.680 1407.040 15.940 ;
        RECT 1423.800 15.680 1424.060 15.940 ;
      LAYER met2 ;
        RECT 1401.490 600.170 1401.770 604.000 ;
        RECT 1401.490 600.030 1403.300 600.170 ;
        RECT 1401.490 600.000 1401.770 600.030 ;
        RECT 1403.160 587.510 1403.300 600.030 ;
        RECT 1403.100 587.190 1403.360 587.510 ;
        RECT 1406.780 587.190 1407.040 587.510 ;
        RECT 1406.840 15.970 1406.980 587.190 ;
        RECT 1406.780 15.650 1407.040 15.970 ;
        RECT 1423.800 15.650 1424.060 15.970 ;
        RECT 1423.860 2.400 1424.000 15.650 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1413.650 18.940 1413.970 19.000 ;
        RECT 1441.710 18.940 1442.030 19.000 ;
        RECT 1413.650 18.800 1442.030 18.940 ;
        RECT 1413.650 18.740 1413.970 18.800 ;
        RECT 1441.710 18.740 1442.030 18.800 ;
      LAYER via ;
        RECT 1413.680 18.740 1413.940 19.000 ;
        RECT 1441.740 18.740 1442.000 19.000 ;
      LAYER met2 ;
        RECT 1410.690 600.170 1410.970 604.000 ;
        RECT 1410.690 600.030 1412.960 600.170 ;
        RECT 1410.690 600.000 1410.970 600.030 ;
        RECT 1412.820 587.250 1412.960 600.030 ;
        RECT 1412.820 587.110 1413.880 587.250 ;
        RECT 1413.740 19.030 1413.880 587.110 ;
        RECT 1413.680 18.710 1413.940 19.030 ;
        RECT 1441.740 18.710 1442.000 19.030 ;
        RECT 1441.800 2.400 1441.940 18.710 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1420.550 19.280 1420.870 19.340 ;
        RECT 1430.670 19.280 1430.990 19.340 ;
        RECT 1420.550 19.140 1430.990 19.280 ;
        RECT 1420.550 19.080 1420.870 19.140 ;
        RECT 1430.670 19.080 1430.990 19.140 ;
        RECT 1430.670 17.580 1430.990 17.640 ;
        RECT 1459.650 17.580 1459.970 17.640 ;
        RECT 1430.670 17.440 1459.970 17.580 ;
        RECT 1430.670 17.380 1430.990 17.440 ;
        RECT 1459.650 17.380 1459.970 17.440 ;
      LAYER via ;
        RECT 1420.580 19.080 1420.840 19.340 ;
        RECT 1430.700 19.080 1430.960 19.340 ;
        RECT 1430.700 17.380 1430.960 17.640 ;
        RECT 1459.680 17.380 1459.940 17.640 ;
      LAYER met2 ;
        RECT 1419.890 600.170 1420.170 604.000 ;
        RECT 1419.890 600.030 1420.780 600.170 ;
        RECT 1419.890 600.000 1420.170 600.030 ;
        RECT 1420.640 19.370 1420.780 600.030 ;
        RECT 1420.580 19.050 1420.840 19.370 ;
        RECT 1430.700 19.050 1430.960 19.370 ;
        RECT 1430.760 17.670 1430.900 19.050 ;
        RECT 1430.700 17.350 1430.960 17.670 ;
        RECT 1459.680 17.350 1459.940 17.670 ;
        RECT 1459.740 2.400 1459.880 17.350 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1430.670 586.740 1430.990 586.800 ;
        RECT 1434.810 586.740 1435.130 586.800 ;
        RECT 1430.670 586.600 1435.130 586.740 ;
        RECT 1430.670 586.540 1430.990 586.600 ;
        RECT 1434.810 586.540 1435.130 586.600 ;
        RECT 1434.810 20.300 1435.130 20.360 ;
        RECT 1477.590 20.300 1477.910 20.360 ;
        RECT 1434.810 20.160 1477.910 20.300 ;
        RECT 1434.810 20.100 1435.130 20.160 ;
        RECT 1477.590 20.100 1477.910 20.160 ;
      LAYER via ;
        RECT 1430.700 586.540 1430.960 586.800 ;
        RECT 1434.840 586.540 1435.100 586.800 ;
        RECT 1434.840 20.100 1435.100 20.360 ;
        RECT 1477.620 20.100 1477.880 20.360 ;
      LAYER met2 ;
        RECT 1429.090 600.170 1429.370 604.000 ;
        RECT 1429.090 600.030 1430.900 600.170 ;
        RECT 1429.090 600.000 1429.370 600.030 ;
        RECT 1430.760 586.830 1430.900 600.030 ;
        RECT 1430.700 586.510 1430.960 586.830 ;
        RECT 1434.840 586.510 1435.100 586.830 ;
        RECT 1434.900 20.390 1435.040 586.510 ;
        RECT 1434.840 20.070 1435.100 20.390 ;
        RECT 1477.620 20.070 1477.880 20.390 ;
        RECT 1477.680 2.400 1477.820 20.070 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.250 19.280 1441.570 19.340 ;
        RECT 1495.530 19.280 1495.850 19.340 ;
        RECT 1441.250 19.140 1495.850 19.280 ;
        RECT 1441.250 19.080 1441.570 19.140 ;
        RECT 1495.530 19.080 1495.850 19.140 ;
      LAYER via ;
        RECT 1441.280 19.080 1441.540 19.340 ;
        RECT 1495.560 19.080 1495.820 19.340 ;
      LAYER met2 ;
        RECT 1438.290 600.170 1438.570 604.000 ;
        RECT 1438.290 600.030 1440.560 600.170 ;
        RECT 1438.290 600.000 1438.570 600.030 ;
        RECT 1440.420 587.250 1440.560 600.030 ;
        RECT 1440.420 587.110 1441.480 587.250 ;
        RECT 1441.340 19.370 1441.480 587.110 ;
        RECT 1441.280 19.050 1441.540 19.370 ;
        RECT 1495.560 19.050 1495.820 19.370 ;
        RECT 1495.620 2.400 1495.760 19.050 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1448.610 18.940 1448.930 19.000 ;
        RECT 1513.010 18.940 1513.330 19.000 ;
        RECT 1448.610 18.800 1513.330 18.940 ;
        RECT 1448.610 18.740 1448.930 18.800 ;
        RECT 1513.010 18.740 1513.330 18.800 ;
      LAYER via ;
        RECT 1448.640 18.740 1448.900 19.000 ;
        RECT 1513.040 18.740 1513.300 19.000 ;
      LAYER met2 ;
        RECT 1447.030 600.170 1447.310 604.000 ;
        RECT 1447.030 600.030 1448.840 600.170 ;
        RECT 1447.030 600.000 1447.310 600.030 ;
        RECT 1448.700 19.030 1448.840 600.030 ;
        RECT 1448.640 18.710 1448.900 19.030 ;
        RECT 1513.040 18.710 1513.300 19.030 ;
        RECT 1513.100 2.400 1513.240 18.710 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 710.310 24.380 710.630 24.440 ;
        RECT 1035.070 24.380 1035.390 24.440 ;
        RECT 710.310 24.240 1035.390 24.380 ;
        RECT 710.310 24.180 710.630 24.240 ;
        RECT 1035.070 24.180 1035.390 24.240 ;
      LAYER via ;
        RECT 710.340 24.180 710.600 24.440 ;
        RECT 1035.100 24.180 1035.360 24.440 ;
      LAYER met2 ;
        RECT 1034.870 600.000 1035.150 604.000 ;
        RECT 1034.930 598.810 1035.070 600.000 ;
        RECT 1034.930 598.670 1035.300 598.810 ;
        RECT 1035.160 24.470 1035.300 598.670 ;
        RECT 710.340 24.150 710.600 24.470 ;
        RECT 1035.100 24.150 1035.360 24.470 ;
        RECT 710.400 2.400 710.540 24.150 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1457.810 586.740 1458.130 586.800 ;
        RECT 1462.410 586.740 1462.730 586.800 ;
        RECT 1457.810 586.600 1462.730 586.740 ;
        RECT 1457.810 586.540 1458.130 586.600 ;
        RECT 1462.410 586.540 1462.730 586.600 ;
        RECT 1462.410 20.640 1462.730 20.700 ;
        RECT 1530.950 20.640 1531.270 20.700 ;
        RECT 1462.410 20.500 1531.270 20.640 ;
        RECT 1462.410 20.440 1462.730 20.500 ;
        RECT 1530.950 20.440 1531.270 20.500 ;
      LAYER via ;
        RECT 1457.840 586.540 1458.100 586.800 ;
        RECT 1462.440 586.540 1462.700 586.800 ;
        RECT 1462.440 20.440 1462.700 20.700 ;
        RECT 1530.980 20.440 1531.240 20.700 ;
      LAYER met2 ;
        RECT 1456.230 600.170 1456.510 604.000 ;
        RECT 1456.230 600.030 1458.040 600.170 ;
        RECT 1456.230 600.000 1456.510 600.030 ;
        RECT 1457.900 586.830 1458.040 600.030 ;
        RECT 1457.840 586.510 1458.100 586.830 ;
        RECT 1462.440 586.510 1462.700 586.830 ;
        RECT 1462.500 20.730 1462.640 586.510 ;
        RECT 1462.440 20.410 1462.700 20.730 ;
        RECT 1530.980 20.410 1531.240 20.730 ;
        RECT 1531.040 2.400 1531.180 20.410 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1466.090 565.660 1466.410 565.720 ;
        RECT 1467.010 565.660 1467.330 565.720 ;
        RECT 1466.090 565.520 1467.330 565.660 ;
        RECT 1466.090 565.460 1466.410 565.520 ;
        RECT 1467.010 565.460 1467.330 565.520 ;
        RECT 1466.090 517.720 1466.410 517.780 ;
        RECT 1467.470 517.720 1467.790 517.780 ;
        RECT 1466.090 517.580 1467.790 517.720 ;
        RECT 1466.090 517.520 1466.410 517.580 ;
        RECT 1467.470 517.520 1467.790 517.580 ;
        RECT 1467.470 475.900 1467.790 475.960 ;
        RECT 1467.930 475.900 1468.250 475.960 ;
        RECT 1467.470 475.760 1468.250 475.900 ;
        RECT 1467.470 475.700 1467.790 475.760 ;
        RECT 1467.930 475.700 1468.250 475.760 ;
        RECT 1467.470 427.960 1467.790 428.020 ;
        RECT 1467.930 427.960 1468.250 428.020 ;
        RECT 1467.470 427.820 1468.250 427.960 ;
        RECT 1467.470 427.760 1467.790 427.820 ;
        RECT 1467.930 427.760 1468.250 427.820 ;
        RECT 1467.470 372.540 1467.790 372.600 ;
        RECT 1467.930 372.540 1468.250 372.600 ;
        RECT 1467.470 372.400 1468.250 372.540 ;
        RECT 1467.470 372.340 1467.790 372.400 ;
        RECT 1467.930 372.340 1468.250 372.400 ;
        RECT 1467.470 324.600 1467.790 324.660 ;
        RECT 1468.390 324.600 1468.710 324.660 ;
        RECT 1467.470 324.460 1468.710 324.600 ;
        RECT 1467.470 324.400 1467.790 324.460 ;
        RECT 1468.390 324.400 1468.710 324.460 ;
        RECT 1468.390 304.200 1468.710 304.260 ;
        RECT 1468.020 304.060 1468.710 304.200 ;
        RECT 1468.020 303.580 1468.160 304.060 ;
        RECT 1468.390 304.000 1468.710 304.060 ;
        RECT 1467.930 303.320 1468.250 303.580 ;
        RECT 1467.010 275.980 1467.330 276.040 ;
        RECT 1467.930 275.980 1468.250 276.040 ;
        RECT 1467.010 275.840 1468.250 275.980 ;
        RECT 1467.010 275.780 1467.330 275.840 ;
        RECT 1467.930 275.780 1468.250 275.840 ;
        RECT 1467.010 228.040 1467.330 228.100 ;
        RECT 1467.470 228.040 1467.790 228.100 ;
        RECT 1467.010 227.900 1467.790 228.040 ;
        RECT 1467.010 227.840 1467.330 227.900 ;
        RECT 1467.470 227.840 1467.790 227.900 ;
        RECT 1467.470 138.280 1467.790 138.340 ;
        RECT 1468.390 138.280 1468.710 138.340 ;
        RECT 1467.470 138.140 1468.710 138.280 ;
        RECT 1467.470 138.080 1467.790 138.140 ;
        RECT 1468.390 138.080 1468.710 138.140 ;
        RECT 1467.010 131.140 1467.330 131.200 ;
        RECT 1468.390 131.140 1468.710 131.200 ;
        RECT 1467.010 131.000 1468.710 131.140 ;
        RECT 1467.010 130.940 1467.330 131.000 ;
        RECT 1468.390 130.940 1468.710 131.000 ;
        RECT 1467.010 83.200 1467.330 83.260 ;
        RECT 1467.930 83.200 1468.250 83.260 ;
        RECT 1467.010 83.060 1468.250 83.200 ;
        RECT 1467.010 83.000 1467.330 83.060 ;
        RECT 1467.930 83.000 1468.250 83.060 ;
        RECT 1468.850 17.920 1469.170 17.980 ;
        RECT 1548.890 17.920 1549.210 17.980 ;
        RECT 1468.850 17.780 1549.210 17.920 ;
        RECT 1468.850 17.720 1469.170 17.780 ;
        RECT 1548.890 17.720 1549.210 17.780 ;
      LAYER via ;
        RECT 1466.120 565.460 1466.380 565.720 ;
        RECT 1467.040 565.460 1467.300 565.720 ;
        RECT 1466.120 517.520 1466.380 517.780 ;
        RECT 1467.500 517.520 1467.760 517.780 ;
        RECT 1467.500 475.700 1467.760 475.960 ;
        RECT 1467.960 475.700 1468.220 475.960 ;
        RECT 1467.500 427.760 1467.760 428.020 ;
        RECT 1467.960 427.760 1468.220 428.020 ;
        RECT 1467.500 372.340 1467.760 372.600 ;
        RECT 1467.960 372.340 1468.220 372.600 ;
        RECT 1467.500 324.400 1467.760 324.660 ;
        RECT 1468.420 324.400 1468.680 324.660 ;
        RECT 1468.420 304.000 1468.680 304.260 ;
        RECT 1467.960 303.320 1468.220 303.580 ;
        RECT 1467.040 275.780 1467.300 276.040 ;
        RECT 1467.960 275.780 1468.220 276.040 ;
        RECT 1467.040 227.840 1467.300 228.100 ;
        RECT 1467.500 227.840 1467.760 228.100 ;
        RECT 1467.500 138.080 1467.760 138.340 ;
        RECT 1468.420 138.080 1468.680 138.340 ;
        RECT 1467.040 130.940 1467.300 131.200 ;
        RECT 1468.420 130.940 1468.680 131.200 ;
        RECT 1467.040 83.000 1467.300 83.260 ;
        RECT 1467.960 83.000 1468.220 83.260 ;
        RECT 1468.880 17.720 1469.140 17.980 ;
        RECT 1548.920 17.720 1549.180 17.980 ;
      LAYER met2 ;
        RECT 1465.430 600.850 1465.710 604.000 ;
        RECT 1465.430 600.710 1466.320 600.850 ;
        RECT 1465.430 600.000 1465.710 600.710 ;
        RECT 1466.180 589.970 1466.320 600.710 ;
        RECT 1466.180 589.830 1467.240 589.970 ;
        RECT 1467.100 565.750 1467.240 589.830 ;
        RECT 1466.120 565.430 1466.380 565.750 ;
        RECT 1467.040 565.430 1467.300 565.750 ;
        RECT 1466.180 517.810 1466.320 565.430 ;
        RECT 1466.120 517.490 1466.380 517.810 ;
        RECT 1467.500 517.490 1467.760 517.810 ;
        RECT 1467.560 475.990 1467.700 517.490 ;
        RECT 1467.500 475.670 1467.760 475.990 ;
        RECT 1467.960 475.670 1468.220 475.990 ;
        RECT 1468.020 428.050 1468.160 475.670 ;
        RECT 1467.500 427.730 1467.760 428.050 ;
        RECT 1467.960 427.730 1468.220 428.050 ;
        RECT 1467.560 399.570 1467.700 427.730 ;
        RECT 1467.560 399.430 1468.160 399.570 ;
        RECT 1468.020 372.630 1468.160 399.430 ;
        RECT 1467.500 372.310 1467.760 372.630 ;
        RECT 1467.960 372.310 1468.220 372.630 ;
        RECT 1467.560 324.690 1467.700 372.310 ;
        RECT 1467.500 324.370 1467.760 324.690 ;
        RECT 1468.420 324.370 1468.680 324.690 ;
        RECT 1468.480 304.290 1468.620 324.370 ;
        RECT 1468.420 303.970 1468.680 304.290 ;
        RECT 1467.960 303.290 1468.220 303.610 ;
        RECT 1468.020 276.070 1468.160 303.290 ;
        RECT 1467.040 275.750 1467.300 276.070 ;
        RECT 1467.960 275.750 1468.220 276.070 ;
        RECT 1467.100 228.130 1467.240 275.750 ;
        RECT 1467.040 227.810 1467.300 228.130 ;
        RECT 1467.500 227.810 1467.760 228.130 ;
        RECT 1467.560 138.370 1467.700 227.810 ;
        RECT 1467.500 138.050 1467.760 138.370 ;
        RECT 1468.420 138.050 1468.680 138.370 ;
        RECT 1468.480 131.230 1468.620 138.050 ;
        RECT 1467.040 130.910 1467.300 131.230 ;
        RECT 1468.420 130.910 1468.680 131.230 ;
        RECT 1467.100 83.290 1467.240 130.910 ;
        RECT 1467.040 82.970 1467.300 83.290 ;
        RECT 1467.960 82.970 1468.220 83.290 ;
        RECT 1468.020 62.290 1468.160 82.970 ;
        RECT 1468.020 62.150 1469.080 62.290 ;
        RECT 1468.940 18.010 1469.080 62.150 ;
        RECT 1468.880 17.690 1469.140 18.010 ;
        RECT 1548.920 17.690 1549.180 18.010 ;
        RECT 1548.980 2.400 1549.120 17.690 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1476.210 17.240 1476.530 17.300 ;
        RECT 1566.830 17.240 1567.150 17.300 ;
        RECT 1476.210 17.100 1567.150 17.240 ;
        RECT 1476.210 17.040 1476.530 17.100 ;
        RECT 1566.830 17.040 1567.150 17.100 ;
      LAYER via ;
        RECT 1476.240 17.040 1476.500 17.300 ;
        RECT 1566.860 17.040 1567.120 17.300 ;
      LAYER met2 ;
        RECT 1474.630 600.170 1474.910 604.000 ;
        RECT 1474.630 600.030 1476.440 600.170 ;
        RECT 1474.630 600.000 1474.910 600.030 ;
        RECT 1476.300 17.330 1476.440 600.030 ;
        RECT 1476.240 17.010 1476.500 17.330 ;
        RECT 1566.860 17.010 1567.120 17.330 ;
        RECT 1566.920 2.400 1567.060 17.010 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1485.410 589.800 1485.730 589.860 ;
        RECT 1580.170 589.800 1580.490 589.860 ;
        RECT 1485.410 589.660 1580.490 589.800 ;
        RECT 1485.410 589.600 1485.730 589.660 ;
        RECT 1580.170 589.600 1580.490 589.660 ;
        RECT 1580.170 579.600 1580.490 579.660 ;
        RECT 1581.090 579.600 1581.410 579.660 ;
        RECT 1580.170 579.460 1581.410 579.600 ;
        RECT 1580.170 579.400 1580.490 579.460 ;
        RECT 1581.090 579.400 1581.410 579.460 ;
        RECT 1580.170 531.660 1580.490 531.720 ;
        RECT 1581.090 531.660 1581.410 531.720 ;
        RECT 1580.170 531.520 1581.410 531.660 ;
        RECT 1580.170 531.460 1580.490 531.520 ;
        RECT 1581.090 531.460 1581.410 531.520 ;
        RECT 1580.170 193.020 1580.490 193.080 ;
        RECT 1581.090 193.020 1581.410 193.080 ;
        RECT 1580.170 192.880 1581.410 193.020 ;
        RECT 1580.170 192.820 1580.490 192.880 ;
        RECT 1581.090 192.820 1581.410 192.880 ;
        RECT 1580.170 145.080 1580.490 145.140 ;
        RECT 1581.090 145.080 1581.410 145.140 ;
        RECT 1580.170 144.940 1581.410 145.080 ;
        RECT 1580.170 144.880 1580.490 144.940 ;
        RECT 1581.090 144.880 1581.410 144.940 ;
        RECT 1580.170 96.460 1580.490 96.520 ;
        RECT 1581.090 96.460 1581.410 96.520 ;
        RECT 1580.170 96.320 1581.410 96.460 ;
        RECT 1580.170 96.260 1580.490 96.320 ;
        RECT 1581.090 96.260 1581.410 96.320 ;
        RECT 1580.170 48.520 1580.490 48.580 ;
        RECT 1581.090 48.520 1581.410 48.580 ;
        RECT 1580.170 48.380 1581.410 48.520 ;
        RECT 1580.170 48.320 1580.490 48.380 ;
        RECT 1581.090 48.320 1581.410 48.380 ;
        RECT 1579.710 2.960 1580.030 3.020 ;
        RECT 1584.770 2.960 1585.090 3.020 ;
        RECT 1579.710 2.820 1585.090 2.960 ;
        RECT 1579.710 2.760 1580.030 2.820 ;
        RECT 1584.770 2.760 1585.090 2.820 ;
      LAYER via ;
        RECT 1485.440 589.600 1485.700 589.860 ;
        RECT 1580.200 589.600 1580.460 589.860 ;
        RECT 1580.200 579.400 1580.460 579.660 ;
        RECT 1581.120 579.400 1581.380 579.660 ;
        RECT 1580.200 531.460 1580.460 531.720 ;
        RECT 1581.120 531.460 1581.380 531.720 ;
        RECT 1580.200 192.820 1580.460 193.080 ;
        RECT 1581.120 192.820 1581.380 193.080 ;
        RECT 1580.200 144.880 1580.460 145.140 ;
        RECT 1581.120 144.880 1581.380 145.140 ;
        RECT 1580.200 96.260 1580.460 96.520 ;
        RECT 1581.120 96.260 1581.380 96.520 ;
        RECT 1580.200 48.320 1580.460 48.580 ;
        RECT 1581.120 48.320 1581.380 48.580 ;
        RECT 1579.740 2.760 1580.000 3.020 ;
        RECT 1584.800 2.760 1585.060 3.020 ;
      LAYER met2 ;
        RECT 1483.830 600.170 1484.110 604.000 ;
        RECT 1483.830 600.030 1485.640 600.170 ;
        RECT 1483.830 600.000 1484.110 600.030 ;
        RECT 1485.500 589.890 1485.640 600.030 ;
        RECT 1485.440 589.570 1485.700 589.890 ;
        RECT 1580.200 589.570 1580.460 589.890 ;
        RECT 1580.260 579.690 1580.400 589.570 ;
        RECT 1580.200 579.370 1580.460 579.690 ;
        RECT 1581.120 579.370 1581.380 579.690 ;
        RECT 1581.180 531.750 1581.320 579.370 ;
        RECT 1580.200 531.430 1580.460 531.750 ;
        RECT 1581.120 531.430 1581.380 531.750 ;
        RECT 1580.260 193.110 1580.400 531.430 ;
        RECT 1580.200 192.790 1580.460 193.110 ;
        RECT 1581.120 192.790 1581.380 193.110 ;
        RECT 1581.180 145.170 1581.320 192.790 ;
        RECT 1580.200 144.850 1580.460 145.170 ;
        RECT 1581.120 144.850 1581.380 145.170 ;
        RECT 1580.260 96.550 1580.400 144.850 ;
        RECT 1580.200 96.230 1580.460 96.550 ;
        RECT 1581.120 96.230 1581.380 96.550 ;
        RECT 1581.180 48.610 1581.320 96.230 ;
        RECT 1580.200 48.290 1580.460 48.610 ;
        RECT 1581.120 48.290 1581.380 48.610 ;
        RECT 1580.260 14.690 1580.400 48.290 ;
        RECT 1579.800 14.550 1580.400 14.690 ;
        RECT 1579.800 3.050 1579.940 14.550 ;
        RECT 1579.740 2.730 1580.000 3.050 ;
        RECT 1584.800 2.730 1585.060 3.050 ;
        RECT 1584.860 2.400 1585.000 2.730 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1494.610 593.200 1494.930 593.260 ;
        RECT 1601.790 593.200 1602.110 593.260 ;
        RECT 1494.610 593.060 1602.110 593.200 ;
        RECT 1494.610 593.000 1494.930 593.060 ;
        RECT 1601.790 593.000 1602.110 593.060 ;
        RECT 1601.790 96.460 1602.110 96.520 ;
        RECT 1602.710 96.460 1603.030 96.520 ;
        RECT 1601.790 96.320 1603.030 96.460 ;
        RECT 1601.790 96.260 1602.110 96.320 ;
        RECT 1602.710 96.260 1603.030 96.320 ;
        RECT 1601.790 48.520 1602.110 48.580 ;
        RECT 1602.710 48.520 1603.030 48.580 ;
        RECT 1601.790 48.380 1603.030 48.520 ;
        RECT 1601.790 48.320 1602.110 48.380 ;
        RECT 1602.710 48.320 1603.030 48.380 ;
        RECT 1601.790 13.980 1602.110 14.240 ;
        RECT 1601.880 13.560 1602.020 13.980 ;
        RECT 1601.790 13.300 1602.110 13.560 ;
        RECT 1601.790 2.960 1602.110 3.020 ;
        RECT 1602.250 2.960 1602.570 3.020 ;
        RECT 1601.790 2.820 1602.570 2.960 ;
        RECT 1601.790 2.760 1602.110 2.820 ;
        RECT 1602.250 2.760 1602.570 2.820 ;
      LAYER via ;
        RECT 1494.640 593.000 1494.900 593.260 ;
        RECT 1601.820 593.000 1602.080 593.260 ;
        RECT 1601.820 96.260 1602.080 96.520 ;
        RECT 1602.740 96.260 1603.000 96.520 ;
        RECT 1601.820 48.320 1602.080 48.580 ;
        RECT 1602.740 48.320 1603.000 48.580 ;
        RECT 1601.820 13.980 1602.080 14.240 ;
        RECT 1601.820 13.300 1602.080 13.560 ;
        RECT 1601.820 2.760 1602.080 3.020 ;
        RECT 1602.280 2.760 1602.540 3.020 ;
      LAYER met2 ;
        RECT 1493.030 600.170 1493.310 604.000 ;
        RECT 1493.030 600.030 1494.840 600.170 ;
        RECT 1493.030 600.000 1493.310 600.030 ;
        RECT 1494.700 593.290 1494.840 600.030 ;
        RECT 1494.640 592.970 1494.900 593.290 ;
        RECT 1601.820 592.970 1602.080 593.290 ;
        RECT 1601.880 96.550 1602.020 592.970 ;
        RECT 1601.820 96.230 1602.080 96.550 ;
        RECT 1602.740 96.230 1603.000 96.550 ;
        RECT 1602.800 48.610 1602.940 96.230 ;
        RECT 1601.820 48.290 1602.080 48.610 ;
        RECT 1602.740 48.290 1603.000 48.610 ;
        RECT 1601.880 14.270 1602.020 48.290 ;
        RECT 1601.820 13.950 1602.080 14.270 ;
        RECT 1601.820 13.270 1602.080 13.590 ;
        RECT 1601.880 3.050 1602.020 13.270 ;
        RECT 1601.820 2.730 1602.080 3.050 ;
        RECT 1602.280 2.730 1602.540 3.050 ;
        RECT 1602.340 2.400 1602.480 2.730 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1503.810 592.180 1504.130 592.240 ;
        RECT 1615.590 592.180 1615.910 592.240 ;
        RECT 1503.810 592.040 1615.910 592.180 ;
        RECT 1503.810 591.980 1504.130 592.040 ;
        RECT 1615.590 591.980 1615.910 592.040 ;
        RECT 1615.590 62.120 1615.910 62.180 ;
        RECT 1619.730 62.120 1620.050 62.180 ;
        RECT 1615.590 61.980 1620.050 62.120 ;
        RECT 1615.590 61.920 1615.910 61.980 ;
        RECT 1619.730 61.920 1620.050 61.980 ;
      LAYER via ;
        RECT 1503.840 591.980 1504.100 592.240 ;
        RECT 1615.620 591.980 1615.880 592.240 ;
        RECT 1615.620 61.920 1615.880 62.180 ;
        RECT 1619.760 61.920 1620.020 62.180 ;
      LAYER met2 ;
        RECT 1502.230 600.170 1502.510 604.000 ;
        RECT 1502.230 600.030 1504.040 600.170 ;
        RECT 1502.230 600.000 1502.510 600.030 ;
        RECT 1503.900 592.270 1504.040 600.030 ;
        RECT 1503.840 591.950 1504.100 592.270 ;
        RECT 1615.620 591.950 1615.880 592.270 ;
        RECT 1615.680 62.210 1615.820 591.950 ;
        RECT 1615.620 61.890 1615.880 62.210 ;
        RECT 1619.760 61.890 1620.020 62.210 ;
        RECT 1619.820 61.610 1619.960 61.890 ;
        RECT 1619.820 61.470 1620.420 61.610 ;
        RECT 1620.280 2.400 1620.420 61.470 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1513.010 590.820 1513.330 590.880 ;
        RECT 1517.610 590.820 1517.930 590.880 ;
        RECT 1513.010 590.680 1517.930 590.820 ;
        RECT 1513.010 590.620 1513.330 590.680 ;
        RECT 1517.610 590.620 1517.930 590.680 ;
        RECT 1517.610 26.080 1517.930 26.140 ;
        RECT 1638.130 26.080 1638.450 26.140 ;
        RECT 1517.610 25.940 1638.450 26.080 ;
        RECT 1517.610 25.880 1517.930 25.940 ;
        RECT 1638.130 25.880 1638.450 25.940 ;
      LAYER via ;
        RECT 1513.040 590.620 1513.300 590.880 ;
        RECT 1517.640 590.620 1517.900 590.880 ;
        RECT 1517.640 25.880 1517.900 26.140 ;
        RECT 1638.160 25.880 1638.420 26.140 ;
      LAYER met2 ;
        RECT 1511.430 600.170 1511.710 604.000 ;
        RECT 1511.430 600.030 1513.240 600.170 ;
        RECT 1511.430 600.000 1511.710 600.030 ;
        RECT 1513.100 590.910 1513.240 600.030 ;
        RECT 1513.040 590.590 1513.300 590.910 ;
        RECT 1517.640 590.590 1517.900 590.910 ;
        RECT 1517.700 26.170 1517.840 590.590 ;
        RECT 1517.640 25.850 1517.900 26.170 ;
        RECT 1638.160 25.850 1638.420 26.170 ;
        RECT 1638.220 2.400 1638.360 25.850 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1522.210 586.740 1522.530 586.800 ;
        RECT 1524.510 586.740 1524.830 586.800 ;
        RECT 1522.210 586.600 1524.830 586.740 ;
        RECT 1522.210 586.540 1522.530 586.600 ;
        RECT 1524.510 586.540 1524.830 586.600 ;
        RECT 1524.510 25.740 1524.830 25.800 ;
        RECT 1656.070 25.740 1656.390 25.800 ;
        RECT 1524.510 25.600 1656.390 25.740 ;
        RECT 1524.510 25.540 1524.830 25.600 ;
        RECT 1656.070 25.540 1656.390 25.600 ;
      LAYER via ;
        RECT 1522.240 586.540 1522.500 586.800 ;
        RECT 1524.540 586.540 1524.800 586.800 ;
        RECT 1524.540 25.540 1524.800 25.800 ;
        RECT 1656.100 25.540 1656.360 25.800 ;
      LAYER met2 ;
        RECT 1520.630 600.170 1520.910 604.000 ;
        RECT 1520.630 600.030 1522.440 600.170 ;
        RECT 1520.630 600.000 1520.910 600.030 ;
        RECT 1522.300 586.830 1522.440 600.030 ;
        RECT 1522.240 586.510 1522.500 586.830 ;
        RECT 1524.540 586.510 1524.800 586.830 ;
        RECT 1524.600 25.830 1524.740 586.510 ;
        RECT 1524.540 25.510 1524.800 25.830 ;
        RECT 1656.100 25.510 1656.360 25.830 ;
        RECT 1656.160 2.400 1656.300 25.510 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1531.410 25.400 1531.730 25.460 ;
        RECT 1673.550 25.400 1673.870 25.460 ;
        RECT 1531.410 25.260 1673.870 25.400 ;
        RECT 1531.410 25.200 1531.730 25.260 ;
        RECT 1673.550 25.200 1673.870 25.260 ;
      LAYER via ;
        RECT 1531.440 25.200 1531.700 25.460 ;
        RECT 1673.580 25.200 1673.840 25.460 ;
      LAYER met2 ;
        RECT 1529.830 600.170 1530.110 604.000 ;
        RECT 1529.830 600.030 1531.640 600.170 ;
        RECT 1529.830 600.000 1530.110 600.030 ;
        RECT 1531.500 25.490 1531.640 600.030 ;
        RECT 1531.440 25.170 1531.700 25.490 ;
        RECT 1673.580 25.170 1673.840 25.490 ;
        RECT 1673.640 2.400 1673.780 25.170 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1540.610 583.340 1540.930 583.400 ;
        RECT 1544.750 583.340 1545.070 583.400 ;
        RECT 1540.610 583.200 1545.070 583.340 ;
        RECT 1540.610 583.140 1540.930 583.200 ;
        RECT 1544.750 583.140 1545.070 583.200 ;
        RECT 1544.750 25.060 1545.070 25.120 ;
        RECT 1691.490 25.060 1691.810 25.120 ;
        RECT 1544.750 24.920 1691.810 25.060 ;
        RECT 1544.750 24.860 1545.070 24.920 ;
        RECT 1691.490 24.860 1691.810 24.920 ;
      LAYER via ;
        RECT 1540.640 583.140 1540.900 583.400 ;
        RECT 1544.780 583.140 1545.040 583.400 ;
        RECT 1544.780 24.860 1545.040 25.120 ;
        RECT 1691.520 24.860 1691.780 25.120 ;
      LAYER met2 ;
        RECT 1539.030 600.170 1539.310 604.000 ;
        RECT 1539.030 600.030 1540.840 600.170 ;
        RECT 1539.030 600.000 1539.310 600.030 ;
        RECT 1540.700 583.430 1540.840 600.030 ;
        RECT 1540.640 583.110 1540.900 583.430 ;
        RECT 1544.780 583.110 1545.040 583.430 ;
        RECT 1544.840 25.150 1544.980 583.110 ;
        RECT 1544.780 24.830 1545.040 25.150 ;
        RECT 1691.520 24.830 1691.780 25.150 ;
        RECT 1691.580 2.400 1691.720 24.830 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1041.970 469.920 1042.290 470.180 ;
        RECT 1042.060 468.480 1042.200 469.920 ;
        RECT 1041.970 468.220 1042.290 468.480 ;
        RECT 728.250 24.720 728.570 24.780 ;
        RECT 1041.970 24.720 1042.290 24.780 ;
        RECT 728.250 24.580 1042.290 24.720 ;
        RECT 728.250 24.520 728.570 24.580 ;
        RECT 1041.970 24.520 1042.290 24.580 ;
      LAYER via ;
        RECT 1042.000 469.920 1042.260 470.180 ;
        RECT 1042.000 468.220 1042.260 468.480 ;
        RECT 728.280 24.520 728.540 24.780 ;
        RECT 1042.000 24.520 1042.260 24.780 ;
      LAYER met2 ;
        RECT 1044.070 600.170 1044.350 604.000 ;
        RECT 1042.060 600.030 1044.350 600.170 ;
        RECT 1042.060 470.210 1042.200 600.030 ;
        RECT 1044.070 600.000 1044.350 600.030 ;
        RECT 1042.000 469.890 1042.260 470.210 ;
        RECT 1042.000 468.190 1042.260 468.510 ;
        RECT 1042.060 24.810 1042.200 468.190 ;
        RECT 728.280 24.490 728.540 24.810 ;
        RECT 1042.000 24.490 1042.260 24.810 ;
        RECT 728.340 2.400 728.480 24.490 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1548.890 572.800 1549.210 572.860 ;
        RECT 1550.730 572.800 1551.050 572.860 ;
        RECT 1548.890 572.660 1551.050 572.800 ;
        RECT 1548.890 572.600 1549.210 572.660 ;
        RECT 1550.730 572.600 1551.050 572.660 ;
        RECT 1550.270 496.780 1550.590 497.040 ;
        RECT 1550.360 496.640 1550.500 496.780 ;
        RECT 1550.730 496.640 1551.050 496.700 ;
        RECT 1550.360 496.500 1551.050 496.640 ;
        RECT 1550.730 496.440 1551.050 496.500 ;
        RECT 1550.730 475.900 1551.050 475.960 ;
        RECT 1551.650 475.900 1551.970 475.960 ;
        RECT 1550.730 475.760 1551.970 475.900 ;
        RECT 1550.730 475.700 1551.050 475.760 ;
        RECT 1551.650 475.700 1551.970 475.760 ;
        RECT 1549.810 379.340 1550.130 379.400 ;
        RECT 1550.730 379.340 1551.050 379.400 ;
        RECT 1549.810 379.200 1551.050 379.340 ;
        RECT 1549.810 379.140 1550.130 379.200 ;
        RECT 1550.730 379.140 1551.050 379.200 ;
        RECT 1549.810 337.860 1550.130 337.920 ;
        RECT 1551.190 337.860 1551.510 337.920 ;
        RECT 1549.810 337.720 1551.510 337.860 ;
        RECT 1549.810 337.660 1550.130 337.720 ;
        RECT 1551.190 337.660 1551.510 337.720 ;
        RECT 1550.730 289.920 1551.050 289.980 ;
        RECT 1551.190 289.920 1551.510 289.980 ;
        RECT 1550.730 289.780 1551.510 289.920 ;
        RECT 1550.730 289.720 1551.050 289.780 ;
        RECT 1551.190 289.720 1551.510 289.780 ;
        RECT 1549.810 282.780 1550.130 282.840 ;
        RECT 1550.730 282.780 1551.050 282.840 ;
        RECT 1549.810 282.640 1551.050 282.780 ;
        RECT 1549.810 282.580 1550.130 282.640 ;
        RECT 1550.730 282.580 1551.050 282.640 ;
        RECT 1549.810 234.840 1550.130 234.900 ;
        RECT 1551.190 234.840 1551.510 234.900 ;
        RECT 1549.810 234.700 1551.510 234.840 ;
        RECT 1549.810 234.640 1550.130 234.700 ;
        RECT 1551.190 234.640 1551.510 234.700 ;
        RECT 1550.270 193.160 1550.590 193.420 ;
        RECT 1550.360 192.740 1550.500 193.160 ;
        RECT 1550.270 192.480 1550.590 192.740 ;
        RECT 1550.270 145.080 1550.590 145.140 ;
        RECT 1551.650 145.080 1551.970 145.140 ;
        RECT 1550.270 144.940 1551.970 145.080 ;
        RECT 1550.270 144.880 1550.590 144.940 ;
        RECT 1551.650 144.880 1551.970 144.940 ;
        RECT 1550.730 144.060 1551.050 144.120 ;
        RECT 1551.650 144.060 1551.970 144.120 ;
        RECT 1550.730 143.920 1551.970 144.060 ;
        RECT 1550.730 143.860 1551.050 143.920 ;
        RECT 1551.650 143.860 1551.970 143.920 ;
        RECT 1551.650 24.720 1551.970 24.780 ;
        RECT 1709.430 24.720 1709.750 24.780 ;
        RECT 1551.650 24.580 1709.750 24.720 ;
        RECT 1551.650 24.520 1551.970 24.580 ;
        RECT 1709.430 24.520 1709.750 24.580 ;
      LAYER via ;
        RECT 1548.920 572.600 1549.180 572.860 ;
        RECT 1550.760 572.600 1551.020 572.860 ;
        RECT 1550.300 496.780 1550.560 497.040 ;
        RECT 1550.760 496.440 1551.020 496.700 ;
        RECT 1550.760 475.700 1551.020 475.960 ;
        RECT 1551.680 475.700 1551.940 475.960 ;
        RECT 1549.840 379.140 1550.100 379.400 ;
        RECT 1550.760 379.140 1551.020 379.400 ;
        RECT 1549.840 337.660 1550.100 337.920 ;
        RECT 1551.220 337.660 1551.480 337.920 ;
        RECT 1550.760 289.720 1551.020 289.980 ;
        RECT 1551.220 289.720 1551.480 289.980 ;
        RECT 1549.840 282.580 1550.100 282.840 ;
        RECT 1550.760 282.580 1551.020 282.840 ;
        RECT 1549.840 234.640 1550.100 234.900 ;
        RECT 1551.220 234.640 1551.480 234.900 ;
        RECT 1550.300 193.160 1550.560 193.420 ;
        RECT 1550.300 192.480 1550.560 192.740 ;
        RECT 1550.300 144.880 1550.560 145.140 ;
        RECT 1551.680 144.880 1551.940 145.140 ;
        RECT 1550.760 143.860 1551.020 144.120 ;
        RECT 1551.680 143.860 1551.940 144.120 ;
        RECT 1551.680 24.520 1551.940 24.780 ;
        RECT 1709.460 24.520 1709.720 24.780 ;
      LAYER met2 ;
        RECT 1548.230 600.170 1548.510 604.000 ;
        RECT 1548.230 600.030 1549.120 600.170 ;
        RECT 1548.230 600.000 1548.510 600.030 ;
        RECT 1548.980 572.890 1549.120 600.030 ;
        RECT 1548.920 572.570 1549.180 572.890 ;
        RECT 1550.760 572.570 1551.020 572.890 ;
        RECT 1550.820 531.490 1550.960 572.570 ;
        RECT 1550.360 531.350 1550.960 531.490 ;
        RECT 1550.360 497.070 1550.500 531.350 ;
        RECT 1550.300 496.750 1550.560 497.070 ;
        RECT 1550.760 496.410 1551.020 496.730 ;
        RECT 1550.820 475.990 1550.960 496.410 ;
        RECT 1550.760 475.670 1551.020 475.990 ;
        RECT 1551.680 475.670 1551.940 475.990 ;
        RECT 1551.740 447.850 1551.880 475.670 ;
        RECT 1550.820 447.710 1551.880 447.850 ;
        RECT 1550.820 400.365 1550.960 447.710 ;
        RECT 1550.750 399.995 1551.030 400.365 ;
        RECT 1550.750 399.315 1551.030 399.685 ;
        RECT 1550.820 379.430 1550.960 399.315 ;
        RECT 1549.840 379.110 1550.100 379.430 ;
        RECT 1550.760 379.110 1551.020 379.430 ;
        RECT 1549.900 337.950 1550.040 379.110 ;
        RECT 1549.840 337.630 1550.100 337.950 ;
        RECT 1551.220 337.630 1551.480 337.950 ;
        RECT 1551.280 290.010 1551.420 337.630 ;
        RECT 1550.760 289.690 1551.020 290.010 ;
        RECT 1551.220 289.690 1551.480 290.010 ;
        RECT 1550.820 282.870 1550.960 289.690 ;
        RECT 1549.840 282.550 1550.100 282.870 ;
        RECT 1550.760 282.550 1551.020 282.870 ;
        RECT 1549.900 234.930 1550.040 282.550 ;
        RECT 1549.840 234.610 1550.100 234.930 ;
        RECT 1551.220 234.610 1551.480 234.930 ;
        RECT 1551.280 209.170 1551.420 234.610 ;
        RECT 1550.360 209.030 1551.420 209.170 ;
        RECT 1550.360 193.450 1550.500 209.030 ;
        RECT 1550.300 193.130 1550.560 193.450 ;
        RECT 1550.300 192.450 1550.560 192.770 ;
        RECT 1550.360 145.170 1550.500 192.450 ;
        RECT 1550.300 144.850 1550.560 145.170 ;
        RECT 1551.680 144.850 1551.940 145.170 ;
        RECT 1551.740 144.150 1551.880 144.850 ;
        RECT 1550.760 143.830 1551.020 144.150 ;
        RECT 1551.680 143.830 1551.940 144.150 ;
        RECT 1550.820 62.290 1550.960 143.830 ;
        RECT 1550.820 62.150 1551.880 62.290 ;
        RECT 1551.740 24.810 1551.880 62.150 ;
        RECT 1551.680 24.490 1551.940 24.810 ;
        RECT 1709.460 24.490 1709.720 24.810 ;
        RECT 1709.520 2.400 1709.660 24.490 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
      LAYER via2 ;
        RECT 1550.750 400.040 1551.030 400.320 ;
        RECT 1550.750 399.360 1551.030 399.640 ;
      LAYER met3 ;
        RECT 1550.725 400.330 1551.055 400.345 ;
        RECT 1550.510 400.015 1551.055 400.330 ;
        RECT 1550.510 399.665 1550.810 400.015 ;
        RECT 1550.510 399.350 1551.055 399.665 ;
        RECT 1550.725 399.335 1551.055 399.350 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1559.010 24.380 1559.330 24.440 ;
        RECT 1727.370 24.380 1727.690 24.440 ;
        RECT 1559.010 24.240 1727.690 24.380 ;
        RECT 1559.010 24.180 1559.330 24.240 ;
        RECT 1727.370 24.180 1727.690 24.240 ;
      LAYER via ;
        RECT 1559.040 24.180 1559.300 24.440 ;
        RECT 1727.400 24.180 1727.660 24.440 ;
      LAYER met2 ;
        RECT 1557.430 600.170 1557.710 604.000 ;
        RECT 1557.430 600.030 1559.240 600.170 ;
        RECT 1557.430 600.000 1557.710 600.030 ;
        RECT 1559.100 24.470 1559.240 600.030 ;
        RECT 1559.040 24.150 1559.300 24.470 ;
        RECT 1727.400 24.150 1727.660 24.470 ;
        RECT 1727.460 2.400 1727.600 24.150 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1567.750 588.780 1568.070 588.840 ;
        RECT 1572.810 588.780 1573.130 588.840 ;
        RECT 1567.750 588.640 1573.130 588.780 ;
        RECT 1567.750 588.580 1568.070 588.640 ;
        RECT 1572.810 588.580 1573.130 588.640 ;
        RECT 1572.810 24.040 1573.130 24.100 ;
        RECT 1745.310 24.040 1745.630 24.100 ;
        RECT 1572.810 23.900 1745.630 24.040 ;
        RECT 1572.810 23.840 1573.130 23.900 ;
        RECT 1745.310 23.840 1745.630 23.900 ;
      LAYER via ;
        RECT 1567.780 588.580 1568.040 588.840 ;
        RECT 1572.840 588.580 1573.100 588.840 ;
        RECT 1572.840 23.840 1573.100 24.100 ;
        RECT 1745.340 23.840 1745.600 24.100 ;
      LAYER met2 ;
        RECT 1566.170 600.170 1566.450 604.000 ;
        RECT 1566.170 600.030 1567.980 600.170 ;
        RECT 1566.170 600.000 1566.450 600.030 ;
        RECT 1567.840 588.870 1567.980 600.030 ;
        RECT 1567.780 588.550 1568.040 588.870 ;
        RECT 1572.840 588.550 1573.100 588.870 ;
        RECT 1572.900 24.130 1573.040 588.550 ;
        RECT 1572.840 23.810 1573.100 24.130 ;
        RECT 1745.340 23.810 1745.600 24.130 ;
        RECT 1745.400 2.400 1745.540 23.810 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1576.950 586.740 1577.270 586.800 ;
        RECT 1579.250 586.740 1579.570 586.800 ;
        RECT 1576.950 586.600 1579.570 586.740 ;
        RECT 1576.950 586.540 1577.270 586.600 ;
        RECT 1579.250 586.540 1579.570 586.600 ;
        RECT 1579.250 29.140 1579.570 29.200 ;
        RECT 1762.790 29.140 1763.110 29.200 ;
        RECT 1579.250 29.000 1763.110 29.140 ;
        RECT 1579.250 28.940 1579.570 29.000 ;
        RECT 1762.790 28.940 1763.110 29.000 ;
      LAYER via ;
        RECT 1576.980 586.540 1577.240 586.800 ;
        RECT 1579.280 586.540 1579.540 586.800 ;
        RECT 1579.280 28.940 1579.540 29.200 ;
        RECT 1762.820 28.940 1763.080 29.200 ;
      LAYER met2 ;
        RECT 1575.370 600.170 1575.650 604.000 ;
        RECT 1575.370 600.030 1577.180 600.170 ;
        RECT 1575.370 600.000 1575.650 600.030 ;
        RECT 1577.040 586.830 1577.180 600.030 ;
        RECT 1576.980 586.510 1577.240 586.830 ;
        RECT 1579.280 586.510 1579.540 586.830 ;
        RECT 1579.340 29.230 1579.480 586.510 ;
        RECT 1579.280 28.910 1579.540 29.230 ;
        RECT 1762.820 28.910 1763.080 29.230 ;
        RECT 1762.880 2.400 1763.020 28.910 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1586.150 30.500 1586.470 30.560 ;
        RECT 1780.730 30.500 1781.050 30.560 ;
        RECT 1586.150 30.360 1781.050 30.500 ;
        RECT 1586.150 30.300 1586.470 30.360 ;
        RECT 1780.730 30.300 1781.050 30.360 ;
      LAYER via ;
        RECT 1586.180 30.300 1586.440 30.560 ;
        RECT 1780.760 30.300 1781.020 30.560 ;
      LAYER met2 ;
        RECT 1584.570 600.170 1584.850 604.000 ;
        RECT 1584.570 600.030 1586.380 600.170 ;
        RECT 1584.570 600.000 1584.850 600.030 ;
        RECT 1586.240 30.590 1586.380 600.030 ;
        RECT 1586.180 30.270 1586.440 30.590 ;
        RECT 1780.760 30.270 1781.020 30.590 ;
        RECT 1780.820 2.400 1780.960 30.270 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1595.350 588.780 1595.670 588.840 ;
        RECT 1600.410 588.780 1600.730 588.840 ;
        RECT 1595.350 588.640 1600.730 588.780 ;
        RECT 1595.350 588.580 1595.670 588.640 ;
        RECT 1600.410 588.580 1600.730 588.640 ;
        RECT 1600.410 30.160 1600.730 30.220 ;
        RECT 1798.670 30.160 1798.990 30.220 ;
        RECT 1600.410 30.020 1798.990 30.160 ;
        RECT 1600.410 29.960 1600.730 30.020 ;
        RECT 1798.670 29.960 1798.990 30.020 ;
      LAYER via ;
        RECT 1595.380 588.580 1595.640 588.840 ;
        RECT 1600.440 588.580 1600.700 588.840 ;
        RECT 1600.440 29.960 1600.700 30.220 ;
        RECT 1798.700 29.960 1798.960 30.220 ;
      LAYER met2 ;
        RECT 1593.770 600.170 1594.050 604.000 ;
        RECT 1593.770 600.030 1595.580 600.170 ;
        RECT 1593.770 600.000 1594.050 600.030 ;
        RECT 1595.440 588.870 1595.580 600.030 ;
        RECT 1595.380 588.550 1595.640 588.870 ;
        RECT 1600.440 588.550 1600.700 588.870 ;
        RECT 1600.500 30.250 1600.640 588.550 ;
        RECT 1600.440 29.930 1600.700 30.250 ;
        RECT 1798.700 29.930 1798.960 30.250 ;
        RECT 1798.760 2.400 1798.900 29.930 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1604.550 586.740 1604.870 586.800 ;
        RECT 1606.850 586.740 1607.170 586.800 ;
        RECT 1604.550 586.600 1607.170 586.740 ;
        RECT 1604.550 586.540 1604.870 586.600 ;
        RECT 1606.850 586.540 1607.170 586.600 ;
        RECT 1606.850 33.900 1607.170 33.960 ;
        RECT 1816.610 33.900 1816.930 33.960 ;
        RECT 1606.850 33.760 1816.930 33.900 ;
        RECT 1606.850 33.700 1607.170 33.760 ;
        RECT 1816.610 33.700 1816.930 33.760 ;
      LAYER via ;
        RECT 1604.580 586.540 1604.840 586.800 ;
        RECT 1606.880 586.540 1607.140 586.800 ;
        RECT 1606.880 33.700 1607.140 33.960 ;
        RECT 1816.640 33.700 1816.900 33.960 ;
      LAYER met2 ;
        RECT 1602.970 600.170 1603.250 604.000 ;
        RECT 1602.970 600.030 1604.780 600.170 ;
        RECT 1602.970 600.000 1603.250 600.030 ;
        RECT 1604.640 586.830 1604.780 600.030 ;
        RECT 1604.580 586.510 1604.840 586.830 ;
        RECT 1606.880 586.510 1607.140 586.830 ;
        RECT 1606.940 33.990 1607.080 586.510 ;
        RECT 1606.880 33.670 1607.140 33.990 ;
        RECT 1816.640 33.670 1816.900 33.990 ;
        RECT 1816.700 2.400 1816.840 33.670 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1613.750 33.220 1614.070 33.280 ;
        RECT 1834.550 33.220 1834.870 33.280 ;
        RECT 1613.750 33.080 1834.870 33.220 ;
        RECT 1613.750 33.020 1614.070 33.080 ;
        RECT 1834.550 33.020 1834.870 33.080 ;
      LAYER via ;
        RECT 1613.780 33.020 1614.040 33.280 ;
        RECT 1834.580 33.020 1834.840 33.280 ;
      LAYER met2 ;
        RECT 1612.170 600.170 1612.450 604.000 ;
        RECT 1612.170 600.030 1613.980 600.170 ;
        RECT 1612.170 600.000 1612.450 600.030 ;
        RECT 1613.840 33.310 1613.980 600.030 ;
        RECT 1613.780 32.990 1614.040 33.310 ;
        RECT 1834.580 32.990 1834.840 33.310 ;
        RECT 1834.640 2.400 1834.780 32.990 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1622.950 586.740 1623.270 586.800 ;
        RECT 1627.090 586.740 1627.410 586.800 ;
        RECT 1622.950 586.600 1627.410 586.740 ;
        RECT 1622.950 586.540 1623.270 586.600 ;
        RECT 1627.090 586.540 1627.410 586.600 ;
        RECT 1627.090 32.540 1627.410 32.600 ;
        RECT 1852.030 32.540 1852.350 32.600 ;
        RECT 1627.090 32.400 1852.350 32.540 ;
        RECT 1627.090 32.340 1627.410 32.400 ;
        RECT 1852.030 32.340 1852.350 32.400 ;
      LAYER via ;
        RECT 1622.980 586.540 1623.240 586.800 ;
        RECT 1627.120 586.540 1627.380 586.800 ;
        RECT 1627.120 32.340 1627.380 32.600 ;
        RECT 1852.060 32.340 1852.320 32.600 ;
      LAYER met2 ;
        RECT 1621.370 600.170 1621.650 604.000 ;
        RECT 1621.370 600.030 1623.180 600.170 ;
        RECT 1621.370 600.000 1621.650 600.030 ;
        RECT 1623.040 586.830 1623.180 600.030 ;
        RECT 1622.980 586.510 1623.240 586.830 ;
        RECT 1627.120 586.510 1627.380 586.830 ;
        RECT 1627.180 32.630 1627.320 586.510 ;
        RECT 1627.120 32.310 1627.380 32.630 ;
        RECT 1852.060 32.310 1852.320 32.630 ;
        RECT 1852.120 2.400 1852.260 32.310 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1632.150 586.740 1632.470 586.800 ;
        RECT 1634.910 586.740 1635.230 586.800 ;
        RECT 1632.150 586.600 1635.230 586.740 ;
        RECT 1632.150 586.540 1632.470 586.600 ;
        RECT 1634.910 586.540 1635.230 586.600 ;
        RECT 1634.910 32.200 1635.230 32.260 ;
        RECT 1869.970 32.200 1870.290 32.260 ;
        RECT 1634.910 32.060 1870.290 32.200 ;
        RECT 1634.910 32.000 1635.230 32.060 ;
        RECT 1869.970 32.000 1870.290 32.060 ;
      LAYER via ;
        RECT 1632.180 586.540 1632.440 586.800 ;
        RECT 1634.940 586.540 1635.200 586.800 ;
        RECT 1634.940 32.000 1635.200 32.260 ;
        RECT 1870.000 32.000 1870.260 32.260 ;
      LAYER met2 ;
        RECT 1630.570 600.170 1630.850 604.000 ;
        RECT 1630.570 600.030 1632.380 600.170 ;
        RECT 1630.570 600.000 1630.850 600.030 ;
        RECT 1632.240 586.830 1632.380 600.030 ;
        RECT 1632.180 586.510 1632.440 586.830 ;
        RECT 1634.940 586.510 1635.200 586.830 ;
        RECT 1635.000 32.290 1635.140 586.510 ;
        RECT 1634.940 31.970 1635.200 32.290 ;
        RECT 1870.000 31.970 1870.260 32.290 ;
        RECT 1870.060 2.400 1870.200 31.970 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1049.330 420.820 1049.650 420.880 ;
        RECT 1049.790 420.820 1050.110 420.880 ;
        RECT 1049.330 420.680 1050.110 420.820 ;
        RECT 1049.330 420.620 1049.650 420.680 ;
        RECT 1049.790 420.620 1050.110 420.680 ;
        RECT 1048.870 331.400 1049.190 331.460 ;
        RECT 1049.790 331.400 1050.110 331.460 ;
        RECT 1048.870 331.260 1050.110 331.400 ;
        RECT 1048.870 331.200 1049.190 331.260 ;
        RECT 1049.790 331.200 1050.110 331.260 ;
        RECT 1048.410 241.300 1048.730 241.360 ;
        RECT 1049.330 241.300 1049.650 241.360 ;
        RECT 1048.410 241.160 1049.650 241.300 ;
        RECT 1048.410 241.100 1048.730 241.160 ;
        RECT 1049.330 241.100 1049.650 241.160 ;
        RECT 1048.870 136.580 1049.190 136.640 ;
        RECT 1049.790 136.580 1050.110 136.640 ;
        RECT 1048.870 136.440 1050.110 136.580 ;
        RECT 1048.870 136.380 1049.190 136.440 ;
        RECT 1049.790 136.380 1050.110 136.440 ;
        RECT 1048.410 89.660 1048.730 89.720 ;
        RECT 1049.790 89.660 1050.110 89.720 ;
        RECT 1048.410 89.520 1050.110 89.660 ;
        RECT 1048.410 89.460 1048.730 89.520 ;
        RECT 1049.790 89.460 1050.110 89.520 ;
        RECT 1048.410 41.720 1048.730 41.780 ;
        RECT 1049.330 41.720 1049.650 41.780 ;
        RECT 1048.410 41.580 1049.650 41.720 ;
        RECT 1048.410 41.520 1048.730 41.580 ;
        RECT 1049.330 41.520 1049.650 41.580 ;
        RECT 746.190 25.400 746.510 25.460 ;
        RECT 1049.330 25.400 1049.650 25.460 ;
        RECT 746.190 25.260 1049.650 25.400 ;
        RECT 746.190 25.200 746.510 25.260 ;
        RECT 1049.330 25.200 1049.650 25.260 ;
      LAYER via ;
        RECT 1049.360 420.620 1049.620 420.880 ;
        RECT 1049.820 420.620 1050.080 420.880 ;
        RECT 1048.900 331.200 1049.160 331.460 ;
        RECT 1049.820 331.200 1050.080 331.460 ;
        RECT 1048.440 241.100 1048.700 241.360 ;
        RECT 1049.360 241.100 1049.620 241.360 ;
        RECT 1048.900 136.380 1049.160 136.640 ;
        RECT 1049.820 136.380 1050.080 136.640 ;
        RECT 1048.440 89.460 1048.700 89.720 ;
        RECT 1049.820 89.460 1050.080 89.720 ;
        RECT 1048.440 41.520 1048.700 41.780 ;
        RECT 1049.360 41.520 1049.620 41.780 ;
        RECT 746.220 25.200 746.480 25.460 ;
        RECT 1049.360 25.200 1049.620 25.460 ;
      LAYER met2 ;
        RECT 1053.270 600.170 1053.550 604.000 ;
        RECT 1051.260 600.030 1053.550 600.170 ;
        RECT 1051.260 569.570 1051.400 600.030 ;
        RECT 1053.270 600.000 1053.550 600.030 ;
        RECT 1049.420 569.430 1051.400 569.570 ;
        RECT 1049.420 498.170 1049.560 569.430 ;
        RECT 1048.960 498.030 1049.560 498.170 ;
        RECT 1048.960 493.410 1049.100 498.030 ;
        RECT 1048.960 493.270 1049.560 493.410 ;
        RECT 1049.420 420.910 1049.560 493.270 ;
        RECT 1049.360 420.590 1049.620 420.910 ;
        RECT 1049.820 420.590 1050.080 420.910 ;
        RECT 1049.880 331.490 1050.020 420.590 ;
        RECT 1048.900 331.170 1049.160 331.490 ;
        RECT 1049.820 331.170 1050.080 331.490 ;
        RECT 1048.960 306.410 1049.100 331.170 ;
        RECT 1048.960 306.270 1049.560 306.410 ;
        RECT 1049.420 241.390 1049.560 306.270 ;
        RECT 1048.440 241.070 1048.700 241.390 ;
        RECT 1049.360 241.070 1049.620 241.390 ;
        RECT 1048.500 193.530 1048.640 241.070 ;
        RECT 1048.500 193.390 1049.100 193.530 ;
        RECT 1048.960 159.530 1049.100 193.390 ;
        RECT 1048.500 159.390 1049.100 159.530 ;
        RECT 1048.500 144.740 1048.640 159.390 ;
        RECT 1048.500 144.600 1049.100 144.740 ;
        RECT 1048.960 136.670 1049.100 144.600 ;
        RECT 1048.900 136.350 1049.160 136.670 ;
        RECT 1049.820 136.350 1050.080 136.670 ;
        RECT 1049.880 89.750 1050.020 136.350 ;
        RECT 1048.440 89.430 1048.700 89.750 ;
        RECT 1049.820 89.430 1050.080 89.750 ;
        RECT 1048.500 41.810 1048.640 89.430 ;
        RECT 1048.440 41.490 1048.700 41.810 ;
        RECT 1049.360 41.490 1049.620 41.810 ;
        RECT 1049.420 25.490 1049.560 41.490 ;
        RECT 746.220 25.170 746.480 25.490 ;
        RECT 1049.360 25.170 1049.620 25.490 ;
        RECT 746.280 2.400 746.420 25.170 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1641.350 31.860 1641.670 31.920 ;
        RECT 1887.910 31.860 1888.230 31.920 ;
        RECT 1641.350 31.720 1888.230 31.860 ;
        RECT 1641.350 31.660 1641.670 31.720 ;
        RECT 1887.910 31.660 1888.230 31.720 ;
      LAYER via ;
        RECT 1641.380 31.660 1641.640 31.920 ;
        RECT 1887.940 31.660 1888.200 31.920 ;
      LAYER met2 ;
        RECT 1639.770 600.170 1640.050 604.000 ;
        RECT 1639.770 600.030 1641.580 600.170 ;
        RECT 1639.770 600.000 1640.050 600.030 ;
        RECT 1641.440 31.950 1641.580 600.030 ;
        RECT 1641.380 31.630 1641.640 31.950 ;
        RECT 1887.940 31.630 1888.200 31.950 ;
        RECT 1888.000 2.400 1888.140 31.630 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1650.550 586.740 1650.870 586.800 ;
        RECT 1655.150 586.740 1655.470 586.800 ;
        RECT 1650.550 586.600 1655.470 586.740 ;
        RECT 1650.550 586.540 1650.870 586.600 ;
        RECT 1655.150 586.540 1655.470 586.600 ;
        RECT 1655.150 31.520 1655.470 31.580 ;
        RECT 1905.850 31.520 1906.170 31.580 ;
        RECT 1655.150 31.380 1906.170 31.520 ;
        RECT 1655.150 31.320 1655.470 31.380 ;
        RECT 1905.850 31.320 1906.170 31.380 ;
      LAYER via ;
        RECT 1650.580 586.540 1650.840 586.800 ;
        RECT 1655.180 586.540 1655.440 586.800 ;
        RECT 1655.180 31.320 1655.440 31.580 ;
        RECT 1905.880 31.320 1906.140 31.580 ;
      LAYER met2 ;
        RECT 1648.970 600.170 1649.250 604.000 ;
        RECT 1648.970 600.030 1650.780 600.170 ;
        RECT 1648.970 600.000 1649.250 600.030 ;
        RECT 1650.640 586.830 1650.780 600.030 ;
        RECT 1650.580 586.510 1650.840 586.830 ;
        RECT 1655.180 586.510 1655.440 586.830 ;
        RECT 1655.240 31.610 1655.380 586.510 ;
        RECT 1655.180 31.290 1655.440 31.610 ;
        RECT 1905.880 31.290 1906.140 31.610 ;
        RECT 1905.940 2.400 1906.080 31.290 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1659.750 586.740 1660.070 586.800 ;
        RECT 1662.510 586.740 1662.830 586.800 ;
        RECT 1659.750 586.600 1662.830 586.740 ;
        RECT 1659.750 586.540 1660.070 586.600 ;
        RECT 1662.510 586.540 1662.830 586.600 ;
        RECT 1662.510 31.180 1662.830 31.240 ;
        RECT 1923.330 31.180 1923.650 31.240 ;
        RECT 1662.510 31.040 1923.650 31.180 ;
        RECT 1662.510 30.980 1662.830 31.040 ;
        RECT 1923.330 30.980 1923.650 31.040 ;
      LAYER via ;
        RECT 1659.780 586.540 1660.040 586.800 ;
        RECT 1662.540 586.540 1662.800 586.800 ;
        RECT 1662.540 30.980 1662.800 31.240 ;
        RECT 1923.360 30.980 1923.620 31.240 ;
      LAYER met2 ;
        RECT 1658.170 600.170 1658.450 604.000 ;
        RECT 1658.170 600.030 1659.980 600.170 ;
        RECT 1658.170 600.000 1658.450 600.030 ;
        RECT 1659.840 586.830 1659.980 600.030 ;
        RECT 1659.780 586.510 1660.040 586.830 ;
        RECT 1662.540 586.510 1662.800 586.830 ;
        RECT 1662.600 31.270 1662.740 586.510 ;
        RECT 1662.540 30.950 1662.800 31.270 ;
        RECT 1923.360 30.950 1923.620 31.270 ;
        RECT 1923.420 2.400 1923.560 30.950 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1668.950 30.840 1669.270 30.900 ;
        RECT 1941.270 30.840 1941.590 30.900 ;
        RECT 1668.950 30.700 1941.590 30.840 ;
        RECT 1668.950 30.640 1669.270 30.700 ;
        RECT 1941.270 30.640 1941.590 30.700 ;
      LAYER via ;
        RECT 1668.980 30.640 1669.240 30.900 ;
        RECT 1941.300 30.640 1941.560 30.900 ;
      LAYER met2 ;
        RECT 1667.370 600.170 1667.650 604.000 ;
        RECT 1667.370 600.030 1669.180 600.170 ;
        RECT 1667.370 600.000 1667.650 600.030 ;
        RECT 1669.040 30.930 1669.180 600.030 ;
        RECT 1668.980 30.610 1669.240 30.930 ;
        RECT 1941.300 30.610 1941.560 30.930 ;
        RECT 1941.360 2.400 1941.500 30.610 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1742.550 592.520 1742.870 592.580 ;
        RECT 1714.120 592.380 1742.870 592.520 ;
        RECT 1678.150 591.500 1678.470 591.560 ;
        RECT 1714.120 591.500 1714.260 592.380 ;
        RECT 1742.550 592.320 1742.870 592.380 ;
        RECT 1678.150 591.360 1714.260 591.500 ;
        RECT 1678.150 591.300 1678.470 591.360 ;
        RECT 1742.550 33.560 1742.870 33.620 ;
        RECT 1959.210 33.560 1959.530 33.620 ;
        RECT 1742.550 33.420 1959.530 33.560 ;
        RECT 1742.550 33.360 1742.870 33.420 ;
        RECT 1959.210 33.360 1959.530 33.420 ;
      LAYER via ;
        RECT 1678.180 591.300 1678.440 591.560 ;
        RECT 1742.580 592.320 1742.840 592.580 ;
        RECT 1742.580 33.360 1742.840 33.620 ;
        RECT 1959.240 33.360 1959.500 33.620 ;
      LAYER met2 ;
        RECT 1676.570 600.170 1676.850 604.000 ;
        RECT 1676.570 600.030 1678.380 600.170 ;
        RECT 1676.570 600.000 1676.850 600.030 ;
        RECT 1678.240 591.590 1678.380 600.030 ;
        RECT 1742.580 592.290 1742.840 592.610 ;
        RECT 1678.180 591.270 1678.440 591.590 ;
        RECT 1742.640 33.650 1742.780 592.290 ;
        RECT 1742.580 33.330 1742.840 33.650 ;
        RECT 1959.240 33.330 1959.500 33.650 ;
        RECT 1959.300 2.400 1959.440 33.330 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1686.890 591.160 1687.210 591.220 ;
        RECT 1755.890 591.160 1756.210 591.220 ;
        RECT 1686.890 591.020 1756.210 591.160 ;
        RECT 1686.890 590.960 1687.210 591.020 ;
        RECT 1755.890 590.960 1756.210 591.020 ;
        RECT 1755.890 32.880 1756.210 32.940 ;
        RECT 1977.150 32.880 1977.470 32.940 ;
        RECT 1755.890 32.740 1977.470 32.880 ;
        RECT 1755.890 32.680 1756.210 32.740 ;
        RECT 1977.150 32.680 1977.470 32.740 ;
      LAYER via ;
        RECT 1686.920 590.960 1687.180 591.220 ;
        RECT 1755.920 590.960 1756.180 591.220 ;
        RECT 1755.920 32.680 1756.180 32.940 ;
        RECT 1977.180 32.680 1977.440 32.940 ;
      LAYER met2 ;
        RECT 1685.310 600.170 1685.590 604.000 ;
        RECT 1685.310 600.030 1687.120 600.170 ;
        RECT 1685.310 600.000 1685.590 600.030 ;
        RECT 1686.980 591.250 1687.120 600.030 ;
        RECT 1686.920 590.930 1687.180 591.250 ;
        RECT 1755.920 590.930 1756.180 591.250 ;
        RECT 1755.980 32.970 1756.120 590.930 ;
        RECT 1755.920 32.650 1756.180 32.970 ;
        RECT 1977.180 32.650 1977.440 32.970 ;
        RECT 1977.240 2.400 1977.380 32.650 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1696.090 590.820 1696.410 590.880 ;
        RECT 1770.150 590.820 1770.470 590.880 ;
        RECT 1696.090 590.680 1770.470 590.820 ;
        RECT 1696.090 590.620 1696.410 590.680 ;
        RECT 1770.150 590.620 1770.470 590.680 ;
        RECT 1769.690 497.120 1770.010 497.380 ;
        RECT 1769.780 496.700 1769.920 497.120 ;
        RECT 1769.690 496.440 1770.010 496.700 ;
        RECT 1768.770 427.620 1769.090 427.680 ;
        RECT 1769.230 427.620 1769.550 427.680 ;
        RECT 1768.770 427.480 1769.550 427.620 ;
        RECT 1768.770 427.420 1769.090 427.480 ;
        RECT 1769.230 427.420 1769.550 427.480 ;
        RECT 1768.770 379.680 1769.090 379.740 ;
        RECT 1770.150 379.680 1770.470 379.740 ;
        RECT 1768.770 379.540 1770.470 379.680 ;
        RECT 1768.770 379.480 1769.090 379.540 ;
        RECT 1770.150 379.480 1770.470 379.540 ;
        RECT 1768.770 289.580 1769.090 289.640 ;
        RECT 1770.150 289.580 1770.470 289.640 ;
        RECT 1768.770 289.440 1770.470 289.580 ;
        RECT 1768.770 289.380 1769.090 289.440 ;
        RECT 1770.150 289.380 1770.470 289.440 ;
        RECT 1768.770 186.560 1769.090 186.620 ;
        RECT 1769.230 186.560 1769.550 186.620 ;
        RECT 1768.770 186.420 1769.550 186.560 ;
        RECT 1768.770 186.360 1769.090 186.420 ;
        RECT 1769.230 186.360 1769.550 186.420 ;
        RECT 1768.770 145.420 1769.090 145.480 ;
        RECT 1769.690 145.420 1770.010 145.480 ;
        RECT 1768.770 145.280 1770.010 145.420 ;
        RECT 1768.770 145.220 1769.090 145.280 ;
        RECT 1769.690 145.220 1770.010 145.280 ;
        RECT 1769.690 137.940 1770.010 138.000 ;
        RECT 1770.150 137.940 1770.470 138.000 ;
        RECT 1769.690 137.800 1770.470 137.940 ;
        RECT 1769.690 137.740 1770.010 137.800 ;
        RECT 1770.150 137.740 1770.470 137.800 ;
        RECT 1770.150 96.600 1770.470 96.860 ;
        RECT 1770.240 96.180 1770.380 96.600 ;
        RECT 1770.150 95.920 1770.470 96.180 ;
        RECT 1769.690 27.780 1770.010 27.840 ;
        RECT 1995.090 27.780 1995.410 27.840 ;
        RECT 1769.690 27.640 1995.410 27.780 ;
        RECT 1769.690 27.580 1770.010 27.640 ;
        RECT 1995.090 27.580 1995.410 27.640 ;
      LAYER via ;
        RECT 1696.120 590.620 1696.380 590.880 ;
        RECT 1770.180 590.620 1770.440 590.880 ;
        RECT 1769.720 497.120 1769.980 497.380 ;
        RECT 1769.720 496.440 1769.980 496.700 ;
        RECT 1768.800 427.420 1769.060 427.680 ;
        RECT 1769.260 427.420 1769.520 427.680 ;
        RECT 1768.800 379.480 1769.060 379.740 ;
        RECT 1770.180 379.480 1770.440 379.740 ;
        RECT 1768.800 289.380 1769.060 289.640 ;
        RECT 1770.180 289.380 1770.440 289.640 ;
        RECT 1768.800 186.360 1769.060 186.620 ;
        RECT 1769.260 186.360 1769.520 186.620 ;
        RECT 1768.800 145.220 1769.060 145.480 ;
        RECT 1769.720 145.220 1769.980 145.480 ;
        RECT 1769.720 137.740 1769.980 138.000 ;
        RECT 1770.180 137.740 1770.440 138.000 ;
        RECT 1770.180 96.600 1770.440 96.860 ;
        RECT 1770.180 95.920 1770.440 96.180 ;
        RECT 1769.720 27.580 1769.980 27.840 ;
        RECT 1995.120 27.580 1995.380 27.840 ;
      LAYER met2 ;
        RECT 1694.510 600.170 1694.790 604.000 ;
        RECT 1694.510 600.030 1696.320 600.170 ;
        RECT 1694.510 600.000 1694.790 600.030 ;
        RECT 1696.180 590.910 1696.320 600.030 ;
        RECT 1696.120 590.590 1696.380 590.910 ;
        RECT 1770.180 590.590 1770.440 590.910 ;
        RECT 1770.240 545.090 1770.380 590.590 ;
        RECT 1769.780 544.950 1770.380 545.090 ;
        RECT 1769.780 497.410 1769.920 544.950 ;
        RECT 1769.720 497.090 1769.980 497.410 ;
        RECT 1769.720 496.410 1769.980 496.730 ;
        RECT 1769.780 458.050 1769.920 496.410 ;
        RECT 1769.320 457.910 1769.920 458.050 ;
        RECT 1769.320 427.710 1769.460 457.910 ;
        RECT 1768.800 427.390 1769.060 427.710 ;
        RECT 1769.260 427.390 1769.520 427.710 ;
        RECT 1768.860 379.770 1769.000 427.390 ;
        RECT 1768.800 379.450 1769.060 379.770 ;
        RECT 1770.180 379.450 1770.440 379.770 ;
        RECT 1770.240 351.290 1770.380 379.450 ;
        RECT 1769.780 351.150 1770.380 351.290 ;
        RECT 1769.780 303.690 1769.920 351.150 ;
        RECT 1769.780 303.550 1770.380 303.690 ;
        RECT 1770.240 289.670 1770.380 303.550 ;
        RECT 1768.800 289.350 1769.060 289.670 ;
        RECT 1770.180 289.350 1770.440 289.670 ;
        RECT 1768.860 254.730 1769.000 289.350 ;
        RECT 1768.860 254.590 1769.920 254.730 ;
        RECT 1769.780 207.810 1769.920 254.590 ;
        RECT 1769.320 207.670 1769.920 207.810 ;
        RECT 1769.320 186.650 1769.460 207.670 ;
        RECT 1768.800 186.330 1769.060 186.650 ;
        RECT 1769.260 186.330 1769.520 186.650 ;
        RECT 1768.860 145.510 1769.000 186.330 ;
        RECT 1768.800 145.190 1769.060 145.510 ;
        RECT 1769.720 145.190 1769.980 145.510 ;
        RECT 1769.780 138.030 1769.920 145.190 ;
        RECT 1769.720 137.710 1769.980 138.030 ;
        RECT 1770.180 137.710 1770.440 138.030 ;
        RECT 1770.240 96.890 1770.380 137.710 ;
        RECT 1770.180 96.570 1770.440 96.890 ;
        RECT 1770.180 95.890 1770.440 96.210 ;
        RECT 1770.240 61.610 1770.380 95.890 ;
        RECT 1769.780 61.470 1770.380 61.610 ;
        RECT 1769.780 27.870 1769.920 61.470 ;
        RECT 1769.720 27.550 1769.980 27.870 ;
        RECT 1995.120 27.550 1995.380 27.870 ;
        RECT 1995.180 2.400 1995.320 27.550 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1703.450 40.020 1703.770 40.080 ;
        RECT 2012.570 40.020 2012.890 40.080 ;
        RECT 1703.450 39.880 2012.890 40.020 ;
        RECT 1703.450 39.820 1703.770 39.880 ;
        RECT 2012.570 39.820 2012.890 39.880 ;
      LAYER via ;
        RECT 1703.480 39.820 1703.740 40.080 ;
        RECT 2012.600 39.820 2012.860 40.080 ;
      LAYER met2 ;
        RECT 1703.710 600.000 1703.990 604.000 ;
        RECT 1703.770 598.810 1703.910 600.000 ;
        RECT 1703.540 598.670 1703.910 598.810 ;
        RECT 1703.540 40.110 1703.680 598.670 ;
        RECT 1703.480 39.790 1703.740 40.110 ;
        RECT 2012.600 39.790 2012.860 40.110 ;
        RECT 2012.660 2.400 2012.800 39.790 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1714.490 591.500 1714.810 591.560 ;
        RECT 1717.710 591.500 1718.030 591.560 ;
        RECT 1714.490 591.360 1718.030 591.500 ;
        RECT 1714.490 591.300 1714.810 591.360 ;
        RECT 1717.710 591.300 1718.030 591.360 ;
        RECT 1717.710 39.680 1718.030 39.740 ;
        RECT 2030.510 39.680 2030.830 39.740 ;
        RECT 1717.710 39.540 2030.830 39.680 ;
        RECT 1717.710 39.480 1718.030 39.540 ;
        RECT 2030.510 39.480 2030.830 39.540 ;
      LAYER via ;
        RECT 1714.520 591.300 1714.780 591.560 ;
        RECT 1717.740 591.300 1718.000 591.560 ;
        RECT 1717.740 39.480 1718.000 39.740 ;
        RECT 2030.540 39.480 2030.800 39.740 ;
      LAYER met2 ;
        RECT 1712.910 600.170 1713.190 604.000 ;
        RECT 1712.910 600.030 1714.720 600.170 ;
        RECT 1712.910 600.000 1713.190 600.030 ;
        RECT 1714.580 591.590 1714.720 600.030 ;
        RECT 1714.520 591.270 1714.780 591.590 ;
        RECT 1717.740 591.270 1718.000 591.590 ;
        RECT 1717.800 39.770 1717.940 591.270 ;
        RECT 1717.740 39.450 1718.000 39.770 ;
        RECT 2030.540 39.450 2030.800 39.770 ;
        RECT 2030.600 2.400 2030.740 39.450 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1724.150 39.340 1724.470 39.400 ;
        RECT 2048.450 39.340 2048.770 39.400 ;
        RECT 1724.150 39.200 2048.770 39.340 ;
        RECT 1724.150 39.140 1724.470 39.200 ;
        RECT 2048.450 39.140 2048.770 39.200 ;
      LAYER via ;
        RECT 1724.180 39.140 1724.440 39.400 ;
        RECT 2048.480 39.140 2048.740 39.400 ;
      LAYER met2 ;
        RECT 1722.110 600.170 1722.390 604.000 ;
        RECT 1722.110 600.030 1724.380 600.170 ;
        RECT 1722.110 600.000 1722.390 600.030 ;
        RECT 1724.240 39.430 1724.380 600.030 ;
        RECT 1724.180 39.110 1724.440 39.430 ;
        RECT 2048.480 39.110 2048.740 39.430 ;
        RECT 2048.540 2.400 2048.680 39.110 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 763.670 25.060 763.990 25.120 ;
        RECT 1062.670 25.060 1062.990 25.120 ;
        RECT 763.670 24.920 1062.990 25.060 ;
        RECT 763.670 24.860 763.990 24.920 ;
        RECT 1062.670 24.860 1062.990 24.920 ;
      LAYER via ;
        RECT 763.700 24.860 763.960 25.120 ;
        RECT 1062.700 24.860 1062.960 25.120 ;
      LAYER met2 ;
        RECT 1062.470 600.000 1062.750 604.000 ;
        RECT 1062.530 598.810 1062.670 600.000 ;
        RECT 1062.530 598.670 1062.900 598.810 ;
        RECT 1062.760 25.150 1062.900 598.670 ;
        RECT 763.700 24.830 763.960 25.150 ;
        RECT 1062.700 24.830 1062.960 25.150 ;
        RECT 763.760 2.400 763.900 24.830 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1731.050 39.000 1731.370 39.060 ;
        RECT 2066.390 39.000 2066.710 39.060 ;
        RECT 1731.050 38.860 2066.710 39.000 ;
        RECT 1731.050 38.800 1731.370 38.860 ;
        RECT 2066.390 38.800 2066.710 38.860 ;
      LAYER via ;
        RECT 1731.080 38.800 1731.340 39.060 ;
        RECT 2066.420 38.800 2066.680 39.060 ;
      LAYER met2 ;
        RECT 1731.310 600.000 1731.590 604.000 ;
        RECT 1731.370 598.810 1731.510 600.000 ;
        RECT 1731.140 598.670 1731.510 598.810 ;
        RECT 1731.140 39.090 1731.280 598.670 ;
        RECT 1731.080 38.770 1731.340 39.090 ;
        RECT 2066.420 38.770 2066.680 39.090 ;
        RECT 2066.480 2.400 2066.620 38.770 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1742.090 591.500 1742.410 591.560 ;
        RECT 1745.310 591.500 1745.630 591.560 ;
        RECT 1742.090 591.360 1745.630 591.500 ;
        RECT 1742.090 591.300 1742.410 591.360 ;
        RECT 1745.310 591.300 1745.630 591.360 ;
        RECT 1745.310 38.660 1745.630 38.720 ;
        RECT 2084.330 38.660 2084.650 38.720 ;
        RECT 1745.310 38.520 2084.650 38.660 ;
        RECT 1745.310 38.460 1745.630 38.520 ;
        RECT 2084.330 38.460 2084.650 38.520 ;
      LAYER via ;
        RECT 1742.120 591.300 1742.380 591.560 ;
        RECT 1745.340 591.300 1745.600 591.560 ;
        RECT 1745.340 38.460 1745.600 38.720 ;
        RECT 2084.360 38.460 2084.620 38.720 ;
      LAYER met2 ;
        RECT 1740.510 600.170 1740.790 604.000 ;
        RECT 1740.510 600.030 1742.320 600.170 ;
        RECT 1740.510 600.000 1740.790 600.030 ;
        RECT 1742.180 591.590 1742.320 600.030 ;
        RECT 1742.120 591.270 1742.380 591.590 ;
        RECT 1745.340 591.270 1745.600 591.590 ;
        RECT 1745.400 38.750 1745.540 591.270 ;
        RECT 1745.340 38.430 1745.600 38.750 ;
        RECT 2084.360 38.430 2084.620 38.750 ;
        RECT 2084.420 2.400 2084.560 38.430 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1751.750 38.320 1752.070 38.380 ;
        RECT 2101.810 38.320 2102.130 38.380 ;
        RECT 1751.750 38.180 2102.130 38.320 ;
        RECT 1751.750 38.120 1752.070 38.180 ;
        RECT 2101.810 38.120 2102.130 38.180 ;
      LAYER via ;
        RECT 1751.780 38.120 1752.040 38.380 ;
        RECT 2101.840 38.120 2102.100 38.380 ;
      LAYER met2 ;
        RECT 1749.710 600.170 1749.990 604.000 ;
        RECT 1749.710 600.030 1751.980 600.170 ;
        RECT 1749.710 600.000 1749.990 600.030 ;
        RECT 1751.840 38.410 1751.980 600.030 ;
        RECT 1751.780 38.090 1752.040 38.410 ;
        RECT 2101.840 38.090 2102.100 38.410 ;
        RECT 2101.900 2.400 2102.040 38.090 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1758.650 37.980 1758.970 38.040 ;
        RECT 2119.750 37.980 2120.070 38.040 ;
        RECT 1758.650 37.840 2120.070 37.980 ;
        RECT 1758.650 37.780 1758.970 37.840 ;
        RECT 2119.750 37.780 2120.070 37.840 ;
      LAYER via ;
        RECT 1758.680 37.780 1758.940 38.040 ;
        RECT 2119.780 37.780 2120.040 38.040 ;
      LAYER met2 ;
        RECT 1758.910 600.000 1759.190 604.000 ;
        RECT 1758.970 598.810 1759.110 600.000 ;
        RECT 1758.740 598.670 1759.110 598.810 ;
        RECT 1758.740 38.070 1758.880 598.670 ;
        RECT 1758.680 37.750 1758.940 38.070 ;
        RECT 2119.780 37.750 2120.040 38.070 ;
        RECT 2119.840 2.400 2119.980 37.750 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1769.690 591.500 1770.010 591.560 ;
        RECT 1772.910 591.500 1773.230 591.560 ;
        RECT 1769.690 591.360 1773.230 591.500 ;
        RECT 1769.690 591.300 1770.010 591.360 ;
        RECT 1772.910 591.300 1773.230 591.360 ;
        RECT 1772.910 35.940 1773.230 36.000 ;
        RECT 2137.690 35.940 2138.010 36.000 ;
        RECT 1772.910 35.800 2138.010 35.940 ;
        RECT 1772.910 35.740 1773.230 35.800 ;
        RECT 2137.690 35.740 2138.010 35.800 ;
      LAYER via ;
        RECT 1769.720 591.300 1769.980 591.560 ;
        RECT 1772.940 591.300 1773.200 591.560 ;
        RECT 1772.940 35.740 1773.200 36.000 ;
        RECT 2137.720 35.740 2137.980 36.000 ;
      LAYER met2 ;
        RECT 1768.110 600.170 1768.390 604.000 ;
        RECT 1768.110 600.030 1769.920 600.170 ;
        RECT 1768.110 600.000 1768.390 600.030 ;
        RECT 1769.780 591.590 1769.920 600.030 ;
        RECT 1769.720 591.270 1769.980 591.590 ;
        RECT 1772.940 591.270 1773.200 591.590 ;
        RECT 1773.000 36.030 1773.140 591.270 ;
        RECT 1772.940 35.710 1773.200 36.030 ;
        RECT 2137.720 35.710 2137.980 36.030 ;
        RECT 2137.780 2.400 2137.920 35.710 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.350 44.780 1779.670 44.840 ;
        RECT 2155.630 44.780 2155.950 44.840 ;
        RECT 1779.350 44.640 2155.950 44.780 ;
        RECT 1779.350 44.580 1779.670 44.640 ;
        RECT 2155.630 44.580 2155.950 44.640 ;
      LAYER via ;
        RECT 1779.380 44.580 1779.640 44.840 ;
        RECT 2155.660 44.580 2155.920 44.840 ;
      LAYER met2 ;
        RECT 1777.310 600.170 1777.590 604.000 ;
        RECT 1777.310 600.030 1779.580 600.170 ;
        RECT 1777.310 600.000 1777.590 600.030 ;
        RECT 1779.440 44.870 1779.580 600.030 ;
        RECT 1779.380 44.550 1779.640 44.870 ;
        RECT 2155.660 44.550 2155.920 44.870 ;
        RECT 2155.720 2.400 2155.860 44.550 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1786.250 42.740 1786.570 42.800 ;
        RECT 2173.110 42.740 2173.430 42.800 ;
        RECT 1786.250 42.600 2173.430 42.740 ;
        RECT 1786.250 42.540 1786.570 42.600 ;
        RECT 2173.110 42.540 2173.430 42.600 ;
      LAYER via ;
        RECT 1786.280 42.540 1786.540 42.800 ;
        RECT 2173.140 42.540 2173.400 42.800 ;
      LAYER met2 ;
        RECT 1786.510 600.000 1786.790 604.000 ;
        RECT 1786.570 598.810 1786.710 600.000 ;
        RECT 1786.340 598.670 1786.710 598.810 ;
        RECT 1786.340 42.830 1786.480 598.670 ;
        RECT 1786.280 42.510 1786.540 42.830 ;
        RECT 2173.140 42.510 2173.400 42.830 ;
        RECT 2173.200 2.400 2173.340 42.510 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1797.290 586.740 1797.610 586.800 ;
        RECT 1800.510 586.740 1800.830 586.800 ;
        RECT 1797.290 586.600 1800.830 586.740 ;
        RECT 1797.290 586.540 1797.610 586.600 ;
        RECT 1800.510 586.540 1800.830 586.600 ;
        RECT 1800.510 50.220 1800.830 50.280 ;
        RECT 2187.370 50.220 2187.690 50.280 ;
        RECT 1800.510 50.080 2187.690 50.220 ;
        RECT 1800.510 50.020 1800.830 50.080 ;
        RECT 2187.370 50.020 2187.690 50.080 ;
      LAYER via ;
        RECT 1797.320 586.540 1797.580 586.800 ;
        RECT 1800.540 586.540 1800.800 586.800 ;
        RECT 1800.540 50.020 1800.800 50.280 ;
        RECT 2187.400 50.020 2187.660 50.280 ;
      LAYER met2 ;
        RECT 1795.710 600.170 1795.990 604.000 ;
        RECT 1795.710 600.030 1797.520 600.170 ;
        RECT 1795.710 600.000 1795.990 600.030 ;
        RECT 1797.380 586.830 1797.520 600.030 ;
        RECT 1797.320 586.510 1797.580 586.830 ;
        RECT 1800.540 586.510 1800.800 586.830 ;
        RECT 1800.600 50.310 1800.740 586.510 ;
        RECT 1800.540 49.990 1800.800 50.310 ;
        RECT 2187.400 49.990 2187.660 50.310 ;
        RECT 2187.460 16.730 2187.600 49.990 ;
        RECT 2187.460 16.590 2191.280 16.730 ;
        RECT 2191.140 2.400 2191.280 16.590 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1806.950 50.560 1807.270 50.620 ;
        RECT 2208.070 50.560 2208.390 50.620 ;
        RECT 1806.950 50.420 2208.390 50.560 ;
        RECT 1806.950 50.360 1807.270 50.420 ;
        RECT 2208.070 50.360 2208.390 50.420 ;
      LAYER via ;
        RECT 1806.980 50.360 1807.240 50.620 ;
        RECT 2208.100 50.360 2208.360 50.620 ;
      LAYER met2 ;
        RECT 1804.910 600.170 1805.190 604.000 ;
        RECT 1804.910 600.030 1807.180 600.170 ;
        RECT 1804.910 600.000 1805.190 600.030 ;
        RECT 1807.040 50.650 1807.180 600.030 ;
        RECT 1806.980 50.330 1807.240 50.650 ;
        RECT 2208.100 50.330 2208.360 50.650 ;
        RECT 2208.160 17.410 2208.300 50.330 ;
        RECT 2208.160 17.270 2209.220 17.410 ;
        RECT 2209.080 2.400 2209.220 17.270 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1813.850 50.900 1814.170 50.960 ;
        RECT 2221.870 50.900 2222.190 50.960 ;
        RECT 1813.850 50.760 2222.190 50.900 ;
        RECT 1813.850 50.700 1814.170 50.760 ;
        RECT 2221.870 50.700 2222.190 50.760 ;
      LAYER via ;
        RECT 1813.880 50.700 1814.140 50.960 ;
        RECT 2221.900 50.700 2222.160 50.960 ;
      LAYER met2 ;
        RECT 1813.650 600.000 1813.930 604.000 ;
        RECT 1813.710 598.810 1813.850 600.000 ;
        RECT 1813.710 598.670 1814.080 598.810 ;
        RECT 1813.940 50.990 1814.080 598.670 ;
        RECT 1813.880 50.670 1814.140 50.990 ;
        RECT 2221.900 50.670 2222.160 50.990 ;
        RECT 2221.960 17.410 2222.100 50.670 ;
        RECT 2221.960 17.270 2227.160 17.410 ;
        RECT 2227.020 2.400 2227.160 17.270 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 814.270 22.680 814.590 22.740 ;
        RECT 1069.570 22.680 1069.890 22.740 ;
        RECT 814.270 22.540 1069.890 22.680 ;
        RECT 814.270 22.480 814.590 22.540 ;
        RECT 1069.570 22.480 1069.890 22.540 ;
        RECT 781.610 14.180 781.930 14.240 ;
        RECT 814.270 14.180 814.590 14.240 ;
        RECT 781.610 14.040 814.590 14.180 ;
        RECT 781.610 13.980 781.930 14.040 ;
        RECT 814.270 13.980 814.590 14.040 ;
      LAYER via ;
        RECT 814.300 22.480 814.560 22.740 ;
        RECT 1069.600 22.480 1069.860 22.740 ;
        RECT 781.640 13.980 781.900 14.240 ;
        RECT 814.300 13.980 814.560 14.240 ;
      LAYER met2 ;
        RECT 1071.670 600.170 1071.950 604.000 ;
        RECT 1069.660 600.030 1071.950 600.170 ;
        RECT 1069.660 22.770 1069.800 600.030 ;
        RECT 1071.670 600.000 1071.950 600.030 ;
        RECT 814.300 22.450 814.560 22.770 ;
        RECT 1069.600 22.450 1069.860 22.770 ;
        RECT 814.360 14.270 814.500 22.450 ;
        RECT 781.640 13.950 781.900 14.270 ;
        RECT 814.300 13.950 814.560 14.270 ;
        RECT 781.700 2.400 781.840 13.950 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1824.430 586.740 1824.750 586.800 ;
        RECT 1828.110 586.740 1828.430 586.800 ;
        RECT 1824.430 586.600 1828.430 586.740 ;
        RECT 1824.430 586.540 1824.750 586.600 ;
        RECT 1828.110 586.540 1828.430 586.600 ;
        RECT 1828.110 51.240 1828.430 51.300 ;
        RECT 2242.570 51.240 2242.890 51.300 ;
        RECT 1828.110 51.100 2242.890 51.240 ;
        RECT 1828.110 51.040 1828.430 51.100 ;
        RECT 2242.570 51.040 2242.890 51.100 ;
      LAYER via ;
        RECT 1824.460 586.540 1824.720 586.800 ;
        RECT 1828.140 586.540 1828.400 586.800 ;
        RECT 1828.140 51.040 1828.400 51.300 ;
        RECT 2242.600 51.040 2242.860 51.300 ;
      LAYER met2 ;
        RECT 1822.850 600.170 1823.130 604.000 ;
        RECT 1822.850 600.030 1824.660 600.170 ;
        RECT 1822.850 600.000 1823.130 600.030 ;
        RECT 1824.520 586.830 1824.660 600.030 ;
        RECT 1824.460 586.510 1824.720 586.830 ;
        RECT 1828.140 586.510 1828.400 586.830 ;
        RECT 1828.200 51.330 1828.340 586.510 ;
        RECT 1828.140 51.010 1828.400 51.330 ;
        RECT 2242.600 51.010 2242.860 51.330 ;
        RECT 2242.660 17.410 2242.800 51.010 ;
        RECT 2242.660 17.270 2245.100 17.410 ;
        RECT 2244.960 2.400 2245.100 17.270 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1834.550 54.980 1834.870 55.040 ;
        RECT 2256.370 54.980 2256.690 55.040 ;
        RECT 1834.550 54.840 2256.690 54.980 ;
        RECT 1834.550 54.780 1834.870 54.840 ;
        RECT 2256.370 54.780 2256.690 54.840 ;
        RECT 2256.370 15.880 2256.690 15.940 ;
        RECT 2262.350 15.880 2262.670 15.940 ;
        RECT 2256.370 15.740 2262.670 15.880 ;
        RECT 2256.370 15.680 2256.690 15.740 ;
        RECT 2262.350 15.680 2262.670 15.740 ;
      LAYER via ;
        RECT 1834.580 54.780 1834.840 55.040 ;
        RECT 2256.400 54.780 2256.660 55.040 ;
        RECT 2256.400 15.680 2256.660 15.940 ;
        RECT 2262.380 15.680 2262.640 15.940 ;
      LAYER met2 ;
        RECT 1832.050 600.170 1832.330 604.000 ;
        RECT 1832.050 600.030 1834.780 600.170 ;
        RECT 1832.050 600.000 1832.330 600.030 ;
        RECT 1834.640 55.070 1834.780 600.030 ;
        RECT 1834.580 54.750 1834.840 55.070 ;
        RECT 2256.400 54.750 2256.660 55.070 ;
        RECT 2256.460 15.970 2256.600 54.750 ;
        RECT 2256.400 15.650 2256.660 15.970 ;
        RECT 2262.380 15.650 2262.640 15.970 ;
        RECT 2262.440 2.400 2262.580 15.650 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1841.450 54.640 1841.770 54.700 ;
        RECT 2277.070 54.640 2277.390 54.700 ;
        RECT 1841.450 54.500 2277.390 54.640 ;
        RECT 1841.450 54.440 1841.770 54.500 ;
        RECT 2277.070 54.440 2277.390 54.500 ;
        RECT 2277.070 2.960 2277.390 3.020 ;
        RECT 2280.290 2.960 2280.610 3.020 ;
        RECT 2277.070 2.820 2280.610 2.960 ;
        RECT 2277.070 2.760 2277.390 2.820 ;
        RECT 2280.290 2.760 2280.610 2.820 ;
      LAYER via ;
        RECT 1841.480 54.440 1841.740 54.700 ;
        RECT 2277.100 54.440 2277.360 54.700 ;
        RECT 2277.100 2.760 2277.360 3.020 ;
        RECT 2280.320 2.760 2280.580 3.020 ;
      LAYER met2 ;
        RECT 1841.250 600.000 1841.530 604.000 ;
        RECT 1841.310 598.810 1841.450 600.000 ;
        RECT 1841.310 598.670 1841.680 598.810 ;
        RECT 1841.540 54.730 1841.680 598.670 ;
        RECT 1841.480 54.410 1841.740 54.730 ;
        RECT 2277.100 54.410 2277.360 54.730 ;
        RECT 2277.160 3.050 2277.300 54.410 ;
        RECT 2277.100 2.730 2277.360 3.050 ;
        RECT 2280.320 2.730 2280.580 3.050 ;
        RECT 2280.380 2.400 2280.520 2.730 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1852.030 586.740 1852.350 586.800 ;
        RECT 1855.710 586.740 1856.030 586.800 ;
        RECT 1852.030 586.600 1856.030 586.740 ;
        RECT 1852.030 586.540 1852.350 586.600 ;
        RECT 1855.710 586.540 1856.030 586.600 ;
        RECT 1855.710 54.300 1856.030 54.360 ;
        RECT 2298.230 54.300 2298.550 54.360 ;
        RECT 1855.710 54.160 2298.550 54.300 ;
        RECT 1855.710 54.100 1856.030 54.160 ;
        RECT 2298.230 54.100 2298.550 54.160 ;
      LAYER via ;
        RECT 1852.060 586.540 1852.320 586.800 ;
        RECT 1855.740 586.540 1856.000 586.800 ;
        RECT 1855.740 54.100 1856.000 54.360 ;
        RECT 2298.260 54.100 2298.520 54.360 ;
      LAYER met2 ;
        RECT 1850.450 600.170 1850.730 604.000 ;
        RECT 1850.450 600.030 1852.260 600.170 ;
        RECT 1850.450 600.000 1850.730 600.030 ;
        RECT 1852.120 586.830 1852.260 600.030 ;
        RECT 1852.060 586.510 1852.320 586.830 ;
        RECT 1855.740 586.510 1856.000 586.830 ;
        RECT 1855.800 54.390 1855.940 586.510 ;
        RECT 1855.740 54.070 1856.000 54.390 ;
        RECT 2298.260 54.070 2298.520 54.390 ;
        RECT 2298.320 2.400 2298.460 54.070 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1862.150 53.960 1862.470 54.020 ;
        RECT 2311.570 53.960 2311.890 54.020 ;
        RECT 1862.150 53.820 2311.890 53.960 ;
        RECT 1862.150 53.760 1862.470 53.820 ;
        RECT 2311.570 53.760 2311.890 53.820 ;
      LAYER via ;
        RECT 1862.180 53.760 1862.440 54.020 ;
        RECT 2311.600 53.760 2311.860 54.020 ;
      LAYER met2 ;
        RECT 1859.650 600.170 1859.930 604.000 ;
        RECT 1859.650 600.030 1862.380 600.170 ;
        RECT 1859.650 600.000 1859.930 600.030 ;
        RECT 1862.240 54.050 1862.380 600.030 ;
        RECT 1862.180 53.730 1862.440 54.050 ;
        RECT 2311.600 53.730 2311.860 54.050 ;
        RECT 2311.660 17.410 2311.800 53.730 ;
        RECT 2311.660 17.270 2316.400 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1868.590 53.280 1868.910 53.340 ;
        RECT 2332.270 53.280 2332.590 53.340 ;
        RECT 1868.590 53.140 2332.590 53.280 ;
        RECT 1868.590 53.080 1868.910 53.140 ;
        RECT 2332.270 53.080 2332.590 53.140 ;
      LAYER via ;
        RECT 1868.620 53.080 1868.880 53.340 ;
        RECT 2332.300 53.080 2332.560 53.340 ;
      LAYER met2 ;
        RECT 1868.850 600.000 1869.130 604.000 ;
        RECT 1868.910 598.810 1869.050 600.000 ;
        RECT 1868.680 598.670 1869.050 598.810 ;
        RECT 1868.680 53.370 1868.820 598.670 ;
        RECT 1868.620 53.050 1868.880 53.370 ;
        RECT 2332.300 53.050 2332.560 53.370 ;
        RECT 2332.360 17.410 2332.500 53.050 ;
        RECT 2332.360 17.270 2334.340 17.410 ;
        RECT 2334.200 2.400 2334.340 17.270 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1879.630 586.740 1879.950 586.800 ;
        RECT 1882.850 586.740 1883.170 586.800 ;
        RECT 1879.630 586.600 1883.170 586.740 ;
        RECT 1879.630 586.540 1879.950 586.600 ;
        RECT 1882.850 586.540 1883.170 586.600 ;
        RECT 1882.850 53.620 1883.170 53.680 ;
        RECT 2346.070 53.620 2346.390 53.680 ;
        RECT 1882.850 53.480 2346.390 53.620 ;
        RECT 1882.850 53.420 1883.170 53.480 ;
        RECT 2346.070 53.420 2346.390 53.480 ;
      LAYER via ;
        RECT 1879.660 586.540 1879.920 586.800 ;
        RECT 1882.880 586.540 1883.140 586.800 ;
        RECT 1882.880 53.420 1883.140 53.680 ;
        RECT 2346.100 53.420 2346.360 53.680 ;
      LAYER met2 ;
        RECT 1878.050 600.170 1878.330 604.000 ;
        RECT 1878.050 600.030 1879.860 600.170 ;
        RECT 1878.050 600.000 1878.330 600.030 ;
        RECT 1879.720 586.830 1879.860 600.030 ;
        RECT 1879.660 586.510 1879.920 586.830 ;
        RECT 1882.880 586.510 1883.140 586.830 ;
        RECT 1882.940 53.710 1883.080 586.510 ;
        RECT 1882.880 53.390 1883.140 53.710 ;
        RECT 2346.100 53.390 2346.360 53.710 ;
        RECT 2346.160 14.010 2346.300 53.390 ;
        RECT 2346.160 13.870 2351.820 14.010 ;
        RECT 2351.680 2.400 2351.820 13.870 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1888.830 579.600 1889.150 579.660 ;
        RECT 1889.290 579.600 1889.610 579.660 ;
        RECT 1888.830 579.460 1889.610 579.600 ;
        RECT 1888.830 579.400 1889.150 579.460 ;
        RECT 1889.290 579.400 1889.610 579.460 ;
        RECT 1888.830 545.060 1889.150 545.320 ;
        RECT 1888.920 544.920 1889.060 545.060 ;
        RECT 1889.290 544.920 1889.610 544.980 ;
        RECT 1888.920 544.780 1889.610 544.920 ;
        RECT 1889.290 544.720 1889.610 544.780 ;
        RECT 1888.830 531.120 1889.150 531.380 ;
        RECT 1888.920 530.640 1889.060 531.120 ;
        RECT 1889.750 530.640 1890.070 530.700 ;
        RECT 1888.920 530.500 1890.070 530.640 ;
        RECT 1889.750 530.440 1890.070 530.500 ;
        RECT 1888.830 448.700 1889.150 448.760 ;
        RECT 1889.750 448.700 1890.070 448.760 ;
        RECT 1888.830 448.560 1890.070 448.700 ;
        RECT 1888.830 448.500 1889.150 448.560 ;
        RECT 1889.750 448.500 1890.070 448.560 ;
        RECT 1888.370 434.760 1888.690 434.820 ;
        RECT 1889.290 434.760 1889.610 434.820 ;
        RECT 1888.370 434.620 1889.610 434.760 ;
        RECT 1888.370 434.560 1888.690 434.620 ;
        RECT 1889.290 434.560 1889.610 434.620 ;
        RECT 1888.370 386.480 1888.690 386.540 ;
        RECT 1889.750 386.480 1890.070 386.540 ;
        RECT 1888.370 386.340 1890.070 386.480 ;
        RECT 1888.370 386.280 1888.690 386.340 ;
        RECT 1889.750 386.280 1890.070 386.340 ;
        RECT 1888.370 282.780 1888.690 282.840 ;
        RECT 1889.750 282.780 1890.070 282.840 ;
        RECT 1888.370 282.640 1890.070 282.780 ;
        RECT 1888.370 282.580 1888.690 282.640 ;
        RECT 1889.750 282.580 1890.070 282.640 ;
        RECT 1889.290 96.460 1889.610 96.520 ;
        RECT 1889.750 96.460 1890.070 96.520 ;
        RECT 1889.290 96.320 1890.070 96.460 ;
        RECT 1889.290 96.260 1889.610 96.320 ;
        RECT 1889.750 96.260 1890.070 96.320 ;
        RECT 1889.750 52.940 1890.070 53.000 ;
        RECT 2366.770 52.940 2367.090 53.000 ;
        RECT 1889.750 52.800 2367.090 52.940 ;
        RECT 1889.750 52.740 1890.070 52.800 ;
        RECT 2366.770 52.740 2367.090 52.800 ;
        RECT 2366.770 2.960 2367.090 3.020 ;
        RECT 2369.530 2.960 2369.850 3.020 ;
        RECT 2366.770 2.820 2369.850 2.960 ;
        RECT 2366.770 2.760 2367.090 2.820 ;
        RECT 2369.530 2.760 2369.850 2.820 ;
      LAYER via ;
        RECT 1888.860 579.400 1889.120 579.660 ;
        RECT 1889.320 579.400 1889.580 579.660 ;
        RECT 1888.860 545.060 1889.120 545.320 ;
        RECT 1889.320 544.720 1889.580 544.980 ;
        RECT 1888.860 531.120 1889.120 531.380 ;
        RECT 1889.780 530.440 1890.040 530.700 ;
        RECT 1888.860 448.500 1889.120 448.760 ;
        RECT 1889.780 448.500 1890.040 448.760 ;
        RECT 1888.400 434.560 1888.660 434.820 ;
        RECT 1889.320 434.560 1889.580 434.820 ;
        RECT 1888.400 386.280 1888.660 386.540 ;
        RECT 1889.780 386.280 1890.040 386.540 ;
        RECT 1888.400 282.580 1888.660 282.840 ;
        RECT 1889.780 282.580 1890.040 282.840 ;
        RECT 1889.320 96.260 1889.580 96.520 ;
        RECT 1889.780 96.260 1890.040 96.520 ;
        RECT 1889.780 52.740 1890.040 53.000 ;
        RECT 2366.800 52.740 2367.060 53.000 ;
        RECT 2366.800 2.760 2367.060 3.020 ;
        RECT 2369.560 2.760 2369.820 3.020 ;
      LAYER met2 ;
        RECT 1887.250 601.530 1887.530 604.000 ;
        RECT 1887.250 601.390 1889.520 601.530 ;
        RECT 1887.250 600.000 1887.530 601.390 ;
        RECT 1889.380 579.690 1889.520 601.390 ;
        RECT 1888.860 579.370 1889.120 579.690 ;
        RECT 1889.320 579.370 1889.580 579.690 ;
        RECT 1888.920 545.350 1889.060 579.370 ;
        RECT 1888.860 545.030 1889.120 545.350 ;
        RECT 1889.320 544.690 1889.580 545.010 ;
        RECT 1889.380 531.490 1889.520 544.690 ;
        RECT 1888.920 531.410 1889.520 531.490 ;
        RECT 1888.860 531.350 1889.520 531.410 ;
        RECT 1888.860 531.090 1889.120 531.350 ;
        RECT 1889.780 530.410 1890.040 530.730 ;
        RECT 1889.840 448.790 1889.980 530.410 ;
        RECT 1888.860 448.530 1889.120 448.790 ;
        RECT 1888.860 448.470 1889.520 448.530 ;
        RECT 1889.780 448.470 1890.040 448.790 ;
        RECT 1888.920 448.390 1889.520 448.470 ;
        RECT 1889.380 434.850 1889.520 448.390 ;
        RECT 1888.400 434.530 1888.660 434.850 ;
        RECT 1889.320 434.530 1889.580 434.850 ;
        RECT 1888.460 386.570 1888.600 434.530 ;
        RECT 1888.400 386.250 1888.660 386.570 ;
        RECT 1889.780 386.250 1890.040 386.570 ;
        RECT 1889.840 351.970 1889.980 386.250 ;
        RECT 1889.380 351.830 1889.980 351.970 ;
        RECT 1889.380 303.690 1889.520 351.830 ;
        RECT 1889.380 303.550 1889.980 303.690 ;
        RECT 1889.840 282.870 1889.980 303.550 ;
        RECT 1888.400 282.550 1888.660 282.870 ;
        RECT 1889.780 282.550 1890.040 282.870 ;
        RECT 1888.460 254.730 1888.600 282.550 ;
        RECT 1888.460 254.590 1889.520 254.730 ;
        RECT 1889.380 207.130 1889.520 254.590 ;
        RECT 1889.380 206.990 1889.980 207.130 ;
        RECT 1889.840 158.850 1889.980 206.990 ;
        RECT 1888.920 158.710 1889.980 158.850 ;
        RECT 1888.920 158.170 1889.060 158.710 ;
        RECT 1888.920 158.030 1889.520 158.170 ;
        RECT 1889.380 96.550 1889.520 158.030 ;
        RECT 1889.320 96.230 1889.580 96.550 ;
        RECT 1889.780 96.230 1890.040 96.550 ;
        RECT 1889.840 53.030 1889.980 96.230 ;
        RECT 1889.780 52.710 1890.040 53.030 ;
        RECT 2366.800 52.710 2367.060 53.030 ;
        RECT 2366.860 3.050 2367.000 52.710 ;
        RECT 2366.800 2.730 2367.060 3.050 ;
        RECT 2369.560 2.730 2369.820 3.050 ;
        RECT 2369.620 2.400 2369.760 2.730 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1896.650 52.260 1896.970 52.320 ;
        RECT 2387.930 52.260 2388.250 52.320 ;
        RECT 1896.650 52.120 2388.250 52.260 ;
        RECT 1896.650 52.060 1896.970 52.120 ;
        RECT 2387.930 52.060 2388.250 52.120 ;
      LAYER via ;
        RECT 1896.680 52.060 1896.940 52.320 ;
        RECT 2387.960 52.060 2388.220 52.320 ;
      LAYER met2 ;
        RECT 1896.450 600.000 1896.730 604.000 ;
        RECT 1896.510 598.810 1896.650 600.000 ;
        RECT 1896.510 598.670 1896.880 598.810 ;
        RECT 1896.740 52.350 1896.880 598.670 ;
        RECT 1896.680 52.030 1896.940 52.350 ;
        RECT 2387.960 52.030 2388.220 52.350 ;
        RECT 2388.020 3.130 2388.160 52.030 ;
        RECT 2387.560 2.990 2388.160 3.130 ;
        RECT 2387.560 2.400 2387.700 2.990 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1907.230 586.740 1907.550 586.800 ;
        RECT 1910.910 586.740 1911.230 586.800 ;
        RECT 1907.230 586.600 1911.230 586.740 ;
        RECT 1907.230 586.540 1907.550 586.600 ;
        RECT 1910.910 586.540 1911.230 586.600 ;
        RECT 1910.910 52.600 1911.230 52.660 ;
        RECT 2401.270 52.600 2401.590 52.660 ;
        RECT 1910.910 52.460 2401.590 52.600 ;
        RECT 1910.910 52.400 1911.230 52.460 ;
        RECT 2401.270 52.400 2401.590 52.460 ;
      LAYER via ;
        RECT 1907.260 586.540 1907.520 586.800 ;
        RECT 1910.940 586.540 1911.200 586.800 ;
        RECT 1910.940 52.400 1911.200 52.660 ;
        RECT 2401.300 52.400 2401.560 52.660 ;
      LAYER met2 ;
        RECT 1905.650 600.170 1905.930 604.000 ;
        RECT 1905.650 600.030 1907.460 600.170 ;
        RECT 1905.650 600.000 1905.930 600.030 ;
        RECT 1907.320 586.830 1907.460 600.030 ;
        RECT 1907.260 586.510 1907.520 586.830 ;
        RECT 1910.940 586.510 1911.200 586.830 ;
        RECT 1911.000 52.690 1911.140 586.510 ;
        RECT 1910.940 52.370 1911.200 52.690 ;
        RECT 2401.300 52.370 2401.560 52.690 ;
        RECT 2401.360 18.090 2401.500 52.370 ;
        RECT 2401.360 17.950 2405.640 18.090 ;
        RECT 2405.500 2.400 2405.640 17.950 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1077.850 373.220 1078.170 373.280 ;
        RECT 1077.480 373.080 1078.170 373.220 ;
        RECT 1077.480 372.940 1077.620 373.080 ;
        RECT 1077.850 373.020 1078.170 373.080 ;
        RECT 1077.390 372.680 1077.710 372.940 ;
        RECT 1077.390 289.380 1077.710 289.640 ;
        RECT 1077.480 289.240 1077.620 289.380 ;
        RECT 1077.850 289.240 1078.170 289.300 ;
        RECT 1077.480 289.100 1078.170 289.240 ;
        RECT 1077.850 289.040 1078.170 289.100 ;
        RECT 1077.390 186.560 1077.710 186.620 ;
        RECT 1077.850 186.560 1078.170 186.620 ;
        RECT 1077.390 186.420 1078.170 186.560 ;
        RECT 1077.390 186.360 1077.710 186.420 ;
        RECT 1077.850 186.360 1078.170 186.420 ;
        RECT 1076.930 131.140 1077.250 131.200 ;
        RECT 1077.850 131.140 1078.170 131.200 ;
        RECT 1076.930 131.000 1078.170 131.140 ;
        RECT 1076.930 130.940 1077.250 131.000 ;
        RECT 1077.850 130.940 1078.170 131.000 ;
        RECT 1076.930 82.520 1077.250 82.580 ;
        RECT 1077.850 82.520 1078.170 82.580 ;
        RECT 1076.930 82.380 1078.170 82.520 ;
        RECT 1076.930 82.320 1077.250 82.380 ;
        RECT 1077.850 82.320 1078.170 82.380 ;
        RECT 1068.650 41.380 1068.970 41.440 ;
        RECT 1076.930 41.380 1077.250 41.440 ;
        RECT 1068.650 41.240 1077.250 41.380 ;
        RECT 1068.650 41.180 1068.970 41.240 ;
        RECT 1076.930 41.180 1077.250 41.240 ;
        RECT 959.170 33.900 959.490 33.960 ;
        RECT 1068.650 33.900 1068.970 33.960 ;
        RECT 959.170 33.760 1068.970 33.900 ;
        RECT 959.170 33.700 959.490 33.760 ;
        RECT 1068.650 33.700 1068.970 33.760 ;
        RECT 835.060 20.500 859.580 20.640 ;
        RECT 799.550 19.960 799.870 20.020 ;
        RECT 835.060 19.960 835.200 20.500 ;
        RECT 799.550 19.820 835.200 19.960 ;
        RECT 859.440 19.960 859.580 20.500 ;
        RECT 859.440 19.820 925.360 19.960 ;
        RECT 799.550 19.760 799.870 19.820 ;
        RECT 925.220 18.940 925.360 19.820 ;
        RECT 959.170 18.940 959.490 19.000 ;
        RECT 925.220 18.800 959.490 18.940 ;
        RECT 959.170 18.740 959.490 18.800 ;
      LAYER via ;
        RECT 1077.880 373.020 1078.140 373.280 ;
        RECT 1077.420 372.680 1077.680 372.940 ;
        RECT 1077.420 289.380 1077.680 289.640 ;
        RECT 1077.880 289.040 1078.140 289.300 ;
        RECT 1077.420 186.360 1077.680 186.620 ;
        RECT 1077.880 186.360 1078.140 186.620 ;
        RECT 1076.960 130.940 1077.220 131.200 ;
        RECT 1077.880 130.940 1078.140 131.200 ;
        RECT 1076.960 82.320 1077.220 82.580 ;
        RECT 1077.880 82.320 1078.140 82.580 ;
        RECT 1068.680 41.180 1068.940 41.440 ;
        RECT 1076.960 41.180 1077.220 41.440 ;
        RECT 959.200 33.700 959.460 33.960 ;
        RECT 1068.680 33.700 1068.940 33.960 ;
        RECT 799.580 19.760 799.840 20.020 ;
        RECT 959.200 18.740 959.460 19.000 ;
      LAYER met2 ;
        RECT 1080.410 600.170 1080.690 604.000 ;
        RECT 1078.400 600.030 1080.690 600.170 ;
        RECT 1078.400 498.850 1078.540 600.030 ;
        RECT 1080.410 600.000 1080.690 600.030 ;
        RECT 1077.940 498.710 1078.540 498.850 ;
        RECT 1077.940 373.310 1078.080 498.710 ;
        RECT 1077.880 372.990 1078.140 373.310 ;
        RECT 1077.420 372.650 1077.680 372.970 ;
        RECT 1077.480 289.670 1077.620 372.650 ;
        RECT 1077.420 289.350 1077.680 289.670 ;
        RECT 1077.880 289.010 1078.140 289.330 ;
        RECT 1077.940 186.650 1078.080 289.010 ;
        RECT 1077.420 186.330 1077.680 186.650 ;
        RECT 1077.880 186.330 1078.140 186.650 ;
        RECT 1077.480 158.850 1077.620 186.330 ;
        RECT 1077.480 158.710 1078.540 158.850 ;
        RECT 1078.400 158.170 1078.540 158.710 ;
        RECT 1077.940 158.030 1078.540 158.170 ;
        RECT 1077.940 131.230 1078.080 158.030 ;
        RECT 1076.960 130.910 1077.220 131.230 ;
        RECT 1077.880 130.910 1078.140 131.230 ;
        RECT 1077.020 124.285 1077.160 130.910 ;
        RECT 1076.950 123.915 1077.230 124.285 ;
        RECT 1077.870 123.915 1078.150 124.285 ;
        RECT 1077.940 82.610 1078.080 123.915 ;
        RECT 1076.960 82.290 1077.220 82.610 ;
        RECT 1077.880 82.290 1078.140 82.610 ;
        RECT 1077.020 41.470 1077.160 82.290 ;
        RECT 1068.680 41.150 1068.940 41.470 ;
        RECT 1076.960 41.150 1077.220 41.470 ;
        RECT 1068.740 33.990 1068.880 41.150 ;
        RECT 959.200 33.670 959.460 33.990 ;
        RECT 1068.680 33.670 1068.940 33.990 ;
        RECT 799.580 19.730 799.840 20.050 ;
        RECT 799.640 2.400 799.780 19.730 ;
        RECT 959.260 19.030 959.400 33.670 ;
        RECT 959.200 18.710 959.460 19.030 ;
        RECT 799.430 -4.800 799.990 2.400 ;
      LAYER via2 ;
        RECT 1076.950 123.960 1077.230 124.240 ;
        RECT 1077.870 123.960 1078.150 124.240 ;
      LAYER met3 ;
        RECT 1076.925 124.250 1077.255 124.265 ;
        RECT 1077.845 124.250 1078.175 124.265 ;
        RECT 1076.925 123.950 1078.175 124.250 ;
        RECT 1076.925 123.935 1077.255 123.950 ;
        RECT 1077.845 123.935 1078.175 123.950 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1001.490 579.940 1001.810 580.000 ;
        RECT 1001.950 579.940 1002.270 580.000 ;
        RECT 1001.490 579.800 1002.270 579.940 ;
        RECT 1001.490 579.740 1001.810 579.800 ;
        RECT 1001.950 579.740 1002.270 579.800 ;
        RECT 1001.030 483.040 1001.350 483.100 ;
        RECT 1001.950 483.040 1002.270 483.100 ;
        RECT 1001.030 482.900 1002.270 483.040 ;
        RECT 1001.030 482.840 1001.350 482.900 ;
        RECT 1001.950 482.840 1002.270 482.900 ;
        RECT 1001.030 317.800 1001.350 317.860 ;
        RECT 1002.410 317.800 1002.730 317.860 ;
        RECT 1001.030 317.660 1002.730 317.800 ;
        RECT 1001.030 317.600 1001.350 317.660 ;
        RECT 1002.410 317.600 1002.730 317.660 ;
        RECT 1002.410 241.780 1002.730 242.040 ;
        RECT 1002.500 241.360 1002.640 241.780 ;
        RECT 1002.410 241.100 1002.730 241.360 ;
        RECT 1001.030 186.560 1001.350 186.620 ;
        RECT 1002.410 186.560 1002.730 186.620 ;
        RECT 1001.030 186.420 1002.730 186.560 ;
        RECT 1001.030 186.360 1001.350 186.420 ;
        RECT 1002.410 186.360 1002.730 186.420 ;
        RECT 1001.030 96.460 1001.350 96.520 ;
        RECT 1001.950 96.460 1002.270 96.520 ;
        RECT 1001.030 96.320 1002.270 96.460 ;
        RECT 1001.030 96.260 1001.350 96.320 ;
        RECT 1001.950 96.260 1002.270 96.320 ;
        RECT 1001.030 62.120 1001.350 62.180 ;
        RECT 1001.950 62.120 1002.270 62.180 ;
        RECT 1001.030 61.980 1002.270 62.120 ;
        RECT 1001.030 61.920 1001.350 61.980 ;
        RECT 1001.950 61.920 1002.270 61.980 ;
        RECT 646.370 43.760 646.690 43.820 ;
        RECT 1001.030 43.760 1001.350 43.820 ;
        RECT 646.370 43.620 1001.350 43.760 ;
        RECT 646.370 43.560 646.690 43.620 ;
        RECT 1001.030 43.560 1001.350 43.620 ;
      LAYER via ;
        RECT 1001.520 579.740 1001.780 580.000 ;
        RECT 1001.980 579.740 1002.240 580.000 ;
        RECT 1001.060 482.840 1001.320 483.100 ;
        RECT 1001.980 482.840 1002.240 483.100 ;
        RECT 1001.060 317.600 1001.320 317.860 ;
        RECT 1002.440 317.600 1002.700 317.860 ;
        RECT 1002.440 241.780 1002.700 242.040 ;
        RECT 1002.440 241.100 1002.700 241.360 ;
        RECT 1001.060 186.360 1001.320 186.620 ;
        RECT 1002.440 186.360 1002.700 186.620 ;
        RECT 1001.060 96.260 1001.320 96.520 ;
        RECT 1001.980 96.260 1002.240 96.520 ;
        RECT 1001.060 61.920 1001.320 62.180 ;
        RECT 1001.980 61.920 1002.240 62.180 ;
        RECT 646.400 43.560 646.660 43.820 ;
        RECT 1001.060 43.560 1001.320 43.820 ;
      LAYER met2 ;
        RECT 1001.290 600.170 1001.570 604.000 ;
        RECT 1001.290 600.030 1002.180 600.170 ;
        RECT 1001.290 600.000 1001.570 600.030 ;
        RECT 1002.040 580.030 1002.180 600.030 ;
        RECT 1001.520 579.710 1001.780 580.030 ;
        RECT 1001.980 579.710 1002.240 580.030 ;
        RECT 1001.580 497.490 1001.720 579.710 ;
        RECT 1001.120 497.350 1001.720 497.490 ;
        RECT 1001.120 483.130 1001.260 497.350 ;
        RECT 1001.060 482.810 1001.320 483.130 ;
        RECT 1001.980 482.810 1002.240 483.130 ;
        RECT 1002.040 448.700 1002.180 482.810 ;
        RECT 1001.580 448.560 1002.180 448.700 ;
        RECT 1001.580 352.650 1001.720 448.560 ;
        RECT 1001.120 352.510 1001.720 352.650 ;
        RECT 1001.120 317.890 1001.260 352.510 ;
        RECT 1001.060 317.570 1001.320 317.890 ;
        RECT 1002.440 317.570 1002.700 317.890 ;
        RECT 1002.500 242.070 1002.640 317.570 ;
        RECT 1002.440 241.750 1002.700 242.070 ;
        RECT 1002.440 241.070 1002.700 241.390 ;
        RECT 1002.500 186.650 1002.640 241.070 ;
        RECT 1001.060 186.330 1001.320 186.650 ;
        RECT 1002.440 186.330 1002.700 186.650 ;
        RECT 1001.120 145.365 1001.260 186.330 ;
        RECT 1001.050 144.995 1001.330 145.365 ;
        RECT 1001.050 96.715 1001.330 97.085 ;
        RECT 1001.120 96.550 1001.260 96.715 ;
        RECT 1001.060 96.230 1001.320 96.550 ;
        RECT 1001.980 96.230 1002.240 96.550 ;
        RECT 1002.040 62.210 1002.180 96.230 ;
        RECT 1001.060 61.890 1001.320 62.210 ;
        RECT 1001.980 61.890 1002.240 62.210 ;
        RECT 1001.120 43.850 1001.260 61.890 ;
        RECT 646.400 43.530 646.660 43.850 ;
        RECT 1001.060 43.530 1001.320 43.850 ;
        RECT 646.460 3.130 646.600 43.530 ;
        RECT 645.080 2.990 646.600 3.130 ;
        RECT 645.080 2.400 645.220 2.990 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 1001.050 145.040 1001.330 145.320 ;
        RECT 1001.050 96.760 1001.330 97.040 ;
      LAYER met3 ;
        RECT 1001.025 145.330 1001.355 145.345 ;
        RECT 1001.025 145.030 1002.490 145.330 ;
        RECT 1001.025 145.015 1001.355 145.030 ;
        RECT 1001.230 143.970 1001.610 143.980 ;
        RECT 1002.190 143.970 1002.490 145.030 ;
        RECT 1001.230 143.670 1002.490 143.970 ;
        RECT 1001.230 143.660 1001.610 143.670 ;
        RECT 1001.025 97.060 1001.355 97.065 ;
        RECT 1001.025 97.050 1001.610 97.060 ;
        RECT 1000.800 96.750 1001.610 97.050 ;
        RECT 1001.025 96.740 1001.610 96.750 ;
        RECT 1001.025 96.735 1001.355 96.740 ;
      LAYER via3 ;
        RECT 1001.260 143.660 1001.580 143.980 ;
        RECT 1001.260 96.740 1001.580 97.060 ;
      LAYER met4 ;
        RECT 1001.255 143.655 1001.585 143.985 ;
        RECT 1001.270 97.065 1001.570 143.655 ;
        RECT 1001.255 96.735 1001.585 97.065 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1916.890 51.580 1917.210 51.640 ;
        RECT 2428.870 51.580 2429.190 51.640 ;
        RECT 1916.890 51.440 2429.190 51.580 ;
        RECT 1916.890 51.380 1917.210 51.440 ;
        RECT 2428.870 51.380 2429.190 51.440 ;
      LAYER via ;
        RECT 1916.920 51.380 1917.180 51.640 ;
        RECT 2428.900 51.380 2429.160 51.640 ;
      LAYER met2 ;
        RECT 1917.610 600.170 1917.890 604.000 ;
        RECT 1916.980 600.030 1917.890 600.170 ;
        RECT 1916.980 51.670 1917.120 600.030 ;
        RECT 1917.610 600.000 1917.890 600.030 ;
        RECT 1916.920 51.350 1917.180 51.670 ;
        RECT 2428.900 51.350 2429.160 51.670 ;
        RECT 2428.960 2.400 2429.100 51.350 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1928.390 586.740 1928.710 586.800 ;
        RECT 1931.150 586.740 1931.470 586.800 ;
        RECT 1928.390 586.600 1931.470 586.740 ;
        RECT 1928.390 586.540 1928.710 586.600 ;
        RECT 1931.150 586.540 1931.470 586.600 ;
        RECT 1931.150 51.920 1931.470 51.980 ;
        RECT 2442.670 51.920 2442.990 51.980 ;
        RECT 1931.150 51.780 2442.990 51.920 ;
        RECT 1931.150 51.720 1931.470 51.780 ;
        RECT 2442.670 51.720 2442.990 51.780 ;
      LAYER via ;
        RECT 1928.420 586.540 1928.680 586.800 ;
        RECT 1931.180 586.540 1931.440 586.800 ;
        RECT 1931.180 51.720 1931.440 51.980 ;
        RECT 2442.700 51.720 2442.960 51.980 ;
      LAYER met2 ;
        RECT 1926.810 600.170 1927.090 604.000 ;
        RECT 1926.810 600.030 1928.620 600.170 ;
        RECT 1926.810 600.000 1927.090 600.030 ;
        RECT 1928.480 586.830 1928.620 600.030 ;
        RECT 1928.420 586.510 1928.680 586.830 ;
        RECT 1931.180 586.510 1931.440 586.830 ;
        RECT 1931.240 52.010 1931.380 586.510 ;
        RECT 1931.180 51.690 1931.440 52.010 ;
        RECT 2442.700 51.690 2442.960 52.010 ;
        RECT 2442.760 18.090 2442.900 51.690 ;
        RECT 2442.760 17.950 2447.040 18.090 ;
        RECT 2446.900 2.400 2447.040 17.950 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.050 60.760 1938.370 60.820 ;
        RECT 2463.370 60.760 2463.690 60.820 ;
        RECT 1938.050 60.620 2463.690 60.760 ;
        RECT 1938.050 60.560 1938.370 60.620 ;
        RECT 2463.370 60.560 2463.690 60.620 ;
      LAYER via ;
        RECT 1938.080 60.560 1938.340 60.820 ;
        RECT 2463.400 60.560 2463.660 60.820 ;
      LAYER met2 ;
        RECT 1936.010 600.170 1936.290 604.000 ;
        RECT 1936.010 600.030 1938.280 600.170 ;
        RECT 1936.010 600.000 1936.290 600.030 ;
        RECT 1938.140 60.850 1938.280 600.030 ;
        RECT 1938.080 60.530 1938.340 60.850 ;
        RECT 2463.400 60.530 2463.660 60.850 ;
        RECT 2463.460 3.130 2463.600 60.530 ;
        RECT 2463.460 2.990 2464.520 3.130 ;
        RECT 2464.380 2.960 2464.520 2.990 ;
        RECT 2464.380 2.820 2464.980 2.960 ;
        RECT 2464.840 2.400 2464.980 2.820 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1944.490 60.420 1944.810 60.480 ;
        RECT 2477.170 60.420 2477.490 60.480 ;
        RECT 1944.490 60.280 2477.490 60.420 ;
        RECT 1944.490 60.220 1944.810 60.280 ;
        RECT 2477.170 60.220 2477.490 60.280 ;
        RECT 2477.170 2.960 2477.490 3.020 ;
        RECT 2482.690 2.960 2483.010 3.020 ;
        RECT 2477.170 2.820 2483.010 2.960 ;
        RECT 2477.170 2.760 2477.490 2.820 ;
        RECT 2482.690 2.760 2483.010 2.820 ;
      LAYER via ;
        RECT 1944.520 60.220 1944.780 60.480 ;
        RECT 2477.200 60.220 2477.460 60.480 ;
        RECT 2477.200 2.760 2477.460 3.020 ;
        RECT 2482.720 2.760 2482.980 3.020 ;
      LAYER met2 ;
        RECT 1945.210 600.170 1945.490 604.000 ;
        RECT 1944.580 600.030 1945.490 600.170 ;
        RECT 1944.580 60.510 1944.720 600.030 ;
        RECT 1945.210 600.000 1945.490 600.030 ;
        RECT 1944.520 60.190 1944.780 60.510 ;
        RECT 2477.200 60.190 2477.460 60.510 ;
        RECT 2477.260 3.050 2477.400 60.190 ;
        RECT 2477.200 2.730 2477.460 3.050 ;
        RECT 2482.720 2.730 2482.980 3.050 ;
        RECT 2482.780 2.400 2482.920 2.730 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1955.990 586.740 1956.310 586.800 ;
        RECT 1958.750 586.740 1959.070 586.800 ;
        RECT 1955.990 586.600 1959.070 586.740 ;
        RECT 1955.990 586.540 1956.310 586.600 ;
        RECT 1958.750 586.540 1959.070 586.600 ;
        RECT 1958.750 60.080 1959.070 60.140 ;
        RECT 2497.870 60.080 2498.190 60.140 ;
        RECT 1958.750 59.940 2498.190 60.080 ;
        RECT 1958.750 59.880 1959.070 59.940 ;
        RECT 2497.870 59.880 2498.190 59.940 ;
        RECT 2497.870 2.960 2498.190 3.020 ;
        RECT 2500.630 2.960 2500.950 3.020 ;
        RECT 2497.870 2.820 2500.950 2.960 ;
        RECT 2497.870 2.760 2498.190 2.820 ;
        RECT 2500.630 2.760 2500.950 2.820 ;
      LAYER via ;
        RECT 1956.020 586.540 1956.280 586.800 ;
        RECT 1958.780 586.540 1959.040 586.800 ;
        RECT 1958.780 59.880 1959.040 60.140 ;
        RECT 2497.900 59.880 2498.160 60.140 ;
        RECT 2497.900 2.760 2498.160 3.020 ;
        RECT 2500.660 2.760 2500.920 3.020 ;
      LAYER met2 ;
        RECT 1954.410 600.170 1954.690 604.000 ;
        RECT 1954.410 600.030 1956.220 600.170 ;
        RECT 1954.410 600.000 1954.690 600.030 ;
        RECT 1956.080 586.830 1956.220 600.030 ;
        RECT 1956.020 586.510 1956.280 586.830 ;
        RECT 1958.780 586.510 1959.040 586.830 ;
        RECT 1958.840 60.170 1958.980 586.510 ;
        RECT 1958.780 59.850 1959.040 60.170 ;
        RECT 2497.900 59.850 2498.160 60.170 ;
        RECT 2497.960 3.050 2498.100 59.850 ;
        RECT 2497.900 2.730 2498.160 3.050 ;
        RECT 2500.660 2.730 2500.920 3.050 ;
        RECT 2500.720 2.400 2500.860 2.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1965.650 59.740 1965.970 59.800 ;
        RECT 2511.670 59.740 2511.990 59.800 ;
        RECT 1965.650 59.600 2511.990 59.740 ;
        RECT 1965.650 59.540 1965.970 59.600 ;
        RECT 2511.670 59.540 2511.990 59.600 ;
        RECT 2511.670 14.180 2511.990 14.240 ;
        RECT 2518.110 14.180 2518.430 14.240 ;
        RECT 2511.670 14.040 2518.430 14.180 ;
        RECT 2511.670 13.980 2511.990 14.040 ;
        RECT 2518.110 13.980 2518.430 14.040 ;
      LAYER via ;
        RECT 1965.680 59.540 1965.940 59.800 ;
        RECT 2511.700 59.540 2511.960 59.800 ;
        RECT 2511.700 13.980 2511.960 14.240 ;
        RECT 2518.140 13.980 2518.400 14.240 ;
      LAYER met2 ;
        RECT 1963.610 600.170 1963.890 604.000 ;
        RECT 1963.610 600.030 1965.880 600.170 ;
        RECT 1963.610 600.000 1963.890 600.030 ;
        RECT 1965.740 59.830 1965.880 600.030 ;
        RECT 1965.680 59.510 1965.940 59.830 ;
        RECT 2511.700 59.510 2511.960 59.830 ;
        RECT 2511.760 14.270 2511.900 59.510 ;
        RECT 2511.700 13.950 2511.960 14.270 ;
        RECT 2518.140 13.950 2518.400 14.270 ;
        RECT 2518.200 2.400 2518.340 13.950 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1972.090 59.400 1972.410 59.460 ;
        RECT 2532.370 59.400 2532.690 59.460 ;
        RECT 1972.090 59.260 2532.690 59.400 ;
        RECT 1972.090 59.200 1972.410 59.260 ;
        RECT 2532.370 59.200 2532.690 59.260 ;
        RECT 2532.370 2.960 2532.690 3.020 ;
        RECT 2536.050 2.960 2536.370 3.020 ;
        RECT 2532.370 2.820 2536.370 2.960 ;
        RECT 2532.370 2.760 2532.690 2.820 ;
        RECT 2536.050 2.760 2536.370 2.820 ;
      LAYER via ;
        RECT 1972.120 59.200 1972.380 59.460 ;
        RECT 2532.400 59.200 2532.660 59.460 ;
        RECT 2532.400 2.760 2532.660 3.020 ;
        RECT 2536.080 2.760 2536.340 3.020 ;
      LAYER met2 ;
        RECT 1972.810 600.170 1973.090 604.000 ;
        RECT 1972.180 600.030 1973.090 600.170 ;
        RECT 1972.180 59.490 1972.320 600.030 ;
        RECT 1972.810 600.000 1973.090 600.030 ;
        RECT 1972.120 59.170 1972.380 59.490 ;
        RECT 2532.400 59.170 2532.660 59.490 ;
        RECT 2532.460 3.050 2532.600 59.170 ;
        RECT 2532.400 2.730 2532.660 3.050 ;
        RECT 2536.080 2.730 2536.340 3.050 ;
        RECT 2536.140 2.400 2536.280 2.730 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1983.590 586.740 1983.910 586.800 ;
        RECT 1986.350 586.740 1986.670 586.800 ;
        RECT 1983.590 586.600 1986.670 586.740 ;
        RECT 1983.590 586.540 1983.910 586.600 ;
        RECT 1986.350 586.540 1986.670 586.600 ;
        RECT 1986.350 59.060 1986.670 59.120 ;
        RECT 2553.070 59.060 2553.390 59.120 ;
        RECT 1986.350 58.920 2553.390 59.060 ;
        RECT 1986.350 58.860 1986.670 58.920 ;
        RECT 2553.070 58.860 2553.390 58.920 ;
        RECT 2553.070 2.960 2553.390 3.020 ;
        RECT 2553.990 2.960 2554.310 3.020 ;
        RECT 2553.070 2.820 2554.310 2.960 ;
        RECT 2553.070 2.760 2553.390 2.820 ;
        RECT 2553.990 2.760 2554.310 2.820 ;
      LAYER via ;
        RECT 1983.620 586.540 1983.880 586.800 ;
        RECT 1986.380 586.540 1986.640 586.800 ;
        RECT 1986.380 58.860 1986.640 59.120 ;
        RECT 2553.100 58.860 2553.360 59.120 ;
        RECT 2553.100 2.760 2553.360 3.020 ;
        RECT 2554.020 2.760 2554.280 3.020 ;
      LAYER met2 ;
        RECT 1982.010 600.170 1982.290 604.000 ;
        RECT 1982.010 600.030 1983.820 600.170 ;
        RECT 1982.010 600.000 1982.290 600.030 ;
        RECT 1983.680 586.830 1983.820 600.030 ;
        RECT 1983.620 586.510 1983.880 586.830 ;
        RECT 1986.380 586.510 1986.640 586.830 ;
        RECT 1986.440 59.150 1986.580 586.510 ;
        RECT 1986.380 58.830 1986.640 59.150 ;
        RECT 2553.100 58.830 2553.360 59.150 ;
        RECT 2553.160 3.050 2553.300 58.830 ;
        RECT 2553.100 2.730 2553.360 3.050 ;
        RECT 2554.020 2.730 2554.280 3.050 ;
        RECT 2554.080 2.400 2554.220 2.730 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.250 58.720 1993.570 58.780 ;
        RECT 2566.870 58.720 2567.190 58.780 ;
        RECT 1993.250 58.580 2567.190 58.720 ;
        RECT 1993.250 58.520 1993.570 58.580 ;
        RECT 2566.870 58.520 2567.190 58.580 ;
        RECT 2566.870 2.960 2567.190 3.020 ;
        RECT 2571.930 2.960 2572.250 3.020 ;
        RECT 2566.870 2.820 2572.250 2.960 ;
        RECT 2566.870 2.760 2567.190 2.820 ;
        RECT 2571.930 2.760 2572.250 2.820 ;
      LAYER via ;
        RECT 1993.280 58.520 1993.540 58.780 ;
        RECT 2566.900 58.520 2567.160 58.780 ;
        RECT 2566.900 2.760 2567.160 3.020 ;
        RECT 2571.960 2.760 2572.220 3.020 ;
      LAYER met2 ;
        RECT 1991.210 600.170 1991.490 604.000 ;
        RECT 1991.210 600.030 1993.480 600.170 ;
        RECT 1991.210 600.000 1991.490 600.030 ;
        RECT 1993.340 58.810 1993.480 600.030 ;
        RECT 1993.280 58.490 1993.540 58.810 ;
        RECT 2566.900 58.490 2567.160 58.810 ;
        RECT 2566.960 3.050 2567.100 58.490 ;
        RECT 2566.900 2.730 2567.160 3.050 ;
        RECT 2571.960 2.730 2572.220 3.050 ;
        RECT 2572.020 2.400 2572.160 2.730 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2000.150 587.760 2000.470 587.820 ;
        RECT 2004.290 587.760 2004.610 587.820 ;
        RECT 2000.150 587.620 2004.610 587.760 ;
        RECT 2000.150 587.560 2000.470 587.620 ;
        RECT 2004.290 587.560 2004.610 587.620 ;
        RECT 2004.290 20.300 2004.610 20.360 ;
        RECT 2589.410 20.300 2589.730 20.360 ;
        RECT 2004.290 20.160 2589.730 20.300 ;
        RECT 2004.290 20.100 2004.610 20.160 ;
        RECT 2589.410 20.100 2589.730 20.160 ;
      LAYER via ;
        RECT 2000.180 587.560 2000.440 587.820 ;
        RECT 2004.320 587.560 2004.580 587.820 ;
        RECT 2004.320 20.100 2004.580 20.360 ;
        RECT 2589.440 20.100 2589.700 20.360 ;
      LAYER met2 ;
        RECT 2000.410 600.000 2000.690 604.000 ;
        RECT 2000.470 598.810 2000.610 600.000 ;
        RECT 2000.240 598.670 2000.610 598.810 ;
        RECT 2000.240 587.850 2000.380 598.670 ;
        RECT 2000.180 587.530 2000.440 587.850 ;
        RECT 2004.320 587.530 2004.580 587.850 ;
        RECT 2004.380 20.390 2004.520 587.530 ;
        RECT 2004.320 20.070 2004.580 20.390 ;
        RECT 2589.440 20.070 2589.700 20.390 ;
        RECT 2589.500 2.400 2589.640 20.070 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 942.610 33.560 942.930 33.620 ;
        RECT 1090.730 33.560 1091.050 33.620 ;
        RECT 942.610 33.420 1091.050 33.560 ;
        RECT 942.610 33.360 942.930 33.420 ;
        RECT 1090.730 33.360 1091.050 33.420 ;
        RECT 823.470 15.200 823.790 15.260 ;
        RECT 823.470 15.060 907.420 15.200 ;
        RECT 823.470 15.000 823.790 15.060 ;
        RECT 907.280 14.860 907.420 15.060 ;
        RECT 942.610 14.860 942.930 14.920 ;
        RECT 907.280 14.720 942.930 14.860 ;
        RECT 942.610 14.660 942.930 14.720 ;
      LAYER via ;
        RECT 942.640 33.360 942.900 33.620 ;
        RECT 1090.760 33.360 1091.020 33.620 ;
        RECT 823.500 15.000 823.760 15.260 ;
        RECT 942.640 14.660 942.900 14.920 ;
      LAYER met2 ;
        RECT 1092.830 600.170 1093.110 604.000 ;
        RECT 1090.820 600.030 1093.110 600.170 ;
        RECT 1090.820 33.650 1090.960 600.030 ;
        RECT 1092.830 600.000 1093.110 600.030 ;
        RECT 942.640 33.330 942.900 33.650 ;
        RECT 1090.760 33.330 1091.020 33.650 ;
        RECT 823.500 14.970 823.760 15.290 ;
        RECT 823.560 2.400 823.700 14.970 ;
        RECT 942.700 14.950 942.840 33.330 ;
        RECT 942.640 14.630 942.900 14.950 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2010.730 593.200 2011.050 593.260 ;
        RECT 2349.290 593.200 2349.610 593.260 ;
        RECT 2010.730 593.060 2349.610 593.200 ;
        RECT 2010.730 593.000 2011.050 593.060 ;
        RECT 2349.290 593.000 2349.610 593.060 ;
        RECT 2349.290 14.520 2349.610 14.580 ;
        RECT 2607.350 14.520 2607.670 14.580 ;
        RECT 2349.290 14.380 2607.670 14.520 ;
        RECT 2349.290 14.320 2349.610 14.380 ;
        RECT 2607.350 14.320 2607.670 14.380 ;
      LAYER via ;
        RECT 2010.760 593.000 2011.020 593.260 ;
        RECT 2349.320 593.000 2349.580 593.260 ;
        RECT 2349.320 14.320 2349.580 14.580 ;
        RECT 2607.380 14.320 2607.640 14.580 ;
      LAYER met2 ;
        RECT 2009.150 600.170 2009.430 604.000 ;
        RECT 2009.150 600.030 2010.960 600.170 ;
        RECT 2009.150 600.000 2009.430 600.030 ;
        RECT 2010.820 593.290 2010.960 600.030 ;
        RECT 2010.760 592.970 2011.020 593.290 ;
        RECT 2349.320 592.970 2349.580 593.290 ;
        RECT 2349.380 14.610 2349.520 592.970 ;
        RECT 2349.320 14.290 2349.580 14.610 ;
        RECT 2607.380 14.290 2607.640 14.610 ;
        RECT 2607.440 2.400 2607.580 14.290 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2019.930 587.080 2020.250 587.140 ;
        RECT 2024.990 587.080 2025.310 587.140 ;
        RECT 2019.930 586.940 2025.310 587.080 ;
        RECT 2019.930 586.880 2020.250 586.940 ;
        RECT 2024.990 586.880 2025.310 586.940 ;
        RECT 2024.990 19.960 2025.310 20.020 ;
        RECT 2625.290 19.960 2625.610 20.020 ;
        RECT 2024.990 19.820 2625.610 19.960 ;
        RECT 2024.990 19.760 2025.310 19.820 ;
        RECT 2625.290 19.760 2625.610 19.820 ;
      LAYER via ;
        RECT 2019.960 586.880 2020.220 587.140 ;
        RECT 2025.020 586.880 2025.280 587.140 ;
        RECT 2025.020 19.760 2025.280 20.020 ;
        RECT 2625.320 19.760 2625.580 20.020 ;
      LAYER met2 ;
        RECT 2018.350 600.170 2018.630 604.000 ;
        RECT 2018.350 600.030 2020.160 600.170 ;
        RECT 2018.350 600.000 2018.630 600.030 ;
        RECT 2020.020 587.170 2020.160 600.030 ;
        RECT 2019.960 586.850 2020.220 587.170 ;
        RECT 2025.020 586.850 2025.280 587.170 ;
        RECT 2025.080 20.050 2025.220 586.850 ;
        RECT 2025.020 19.730 2025.280 20.050 ;
        RECT 2625.320 19.730 2625.580 20.050 ;
        RECT 2625.380 2.400 2625.520 19.730 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2028.210 589.460 2028.530 589.520 ;
        RECT 2356.190 589.460 2356.510 589.520 ;
        RECT 2028.210 589.320 2356.510 589.460 ;
        RECT 2028.210 589.260 2028.530 589.320 ;
        RECT 2356.190 589.260 2356.510 589.320 ;
        RECT 2356.190 14.860 2356.510 14.920 ;
        RECT 2643.230 14.860 2643.550 14.920 ;
        RECT 2356.190 14.720 2643.550 14.860 ;
        RECT 2356.190 14.660 2356.510 14.720 ;
        RECT 2643.230 14.660 2643.550 14.720 ;
      LAYER via ;
        RECT 2028.240 589.260 2028.500 589.520 ;
        RECT 2356.220 589.260 2356.480 589.520 ;
        RECT 2356.220 14.660 2356.480 14.920 ;
        RECT 2643.260 14.660 2643.520 14.920 ;
      LAYER met2 ;
        RECT 2027.550 600.170 2027.830 604.000 ;
        RECT 2027.550 600.030 2028.440 600.170 ;
        RECT 2027.550 600.000 2027.830 600.030 ;
        RECT 2028.300 589.550 2028.440 600.030 ;
        RECT 2028.240 589.230 2028.500 589.550 ;
        RECT 2356.220 589.230 2356.480 589.550 ;
        RECT 2356.280 14.950 2356.420 589.230 ;
        RECT 2356.220 14.630 2356.480 14.950 ;
        RECT 2643.260 14.630 2643.520 14.950 ;
        RECT 2643.320 2.400 2643.460 14.630 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2038.330 586.740 2038.650 586.800 ;
        RECT 2042.010 586.740 2042.330 586.800 ;
        RECT 2038.330 586.600 2042.330 586.740 ;
        RECT 2038.330 586.540 2038.650 586.600 ;
        RECT 2042.010 586.540 2042.330 586.600 ;
        RECT 2042.010 19.620 2042.330 19.680 ;
        RECT 2661.170 19.620 2661.490 19.680 ;
        RECT 2042.010 19.480 2661.490 19.620 ;
        RECT 2042.010 19.420 2042.330 19.480 ;
        RECT 2661.170 19.420 2661.490 19.480 ;
      LAYER via ;
        RECT 2038.360 586.540 2038.620 586.800 ;
        RECT 2042.040 586.540 2042.300 586.800 ;
        RECT 2042.040 19.420 2042.300 19.680 ;
        RECT 2661.200 19.420 2661.460 19.680 ;
      LAYER met2 ;
        RECT 2036.750 600.170 2037.030 604.000 ;
        RECT 2036.750 600.030 2038.560 600.170 ;
        RECT 2036.750 600.000 2037.030 600.030 ;
        RECT 2038.420 586.830 2038.560 600.030 ;
        RECT 2038.360 586.510 2038.620 586.830 ;
        RECT 2042.040 586.510 2042.300 586.830 ;
        RECT 2042.100 19.710 2042.240 586.510 ;
        RECT 2042.040 19.390 2042.300 19.710 ;
        RECT 2661.200 19.390 2661.460 19.710 ;
        RECT 2661.260 2.400 2661.400 19.390 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2066.850 589.120 2067.170 589.180 ;
        RECT 2369.990 589.120 2370.310 589.180 ;
        RECT 2066.850 588.980 2370.310 589.120 ;
        RECT 2066.850 588.920 2067.170 588.980 ;
        RECT 2369.990 588.920 2370.310 588.980 ;
        RECT 2047.530 588.100 2047.850 588.160 ;
        RECT 2066.850 588.100 2067.170 588.160 ;
        RECT 2047.530 587.960 2067.170 588.100 ;
        RECT 2047.530 587.900 2047.850 587.960 ;
        RECT 2066.850 587.900 2067.170 587.960 ;
        RECT 2369.990 15.200 2370.310 15.260 ;
        RECT 2678.650 15.200 2678.970 15.260 ;
        RECT 2369.990 15.060 2678.970 15.200 ;
        RECT 2369.990 15.000 2370.310 15.060 ;
        RECT 2678.650 15.000 2678.970 15.060 ;
      LAYER via ;
        RECT 2066.880 588.920 2067.140 589.180 ;
        RECT 2370.020 588.920 2370.280 589.180 ;
        RECT 2047.560 587.900 2047.820 588.160 ;
        RECT 2066.880 587.900 2067.140 588.160 ;
        RECT 2370.020 15.000 2370.280 15.260 ;
        RECT 2678.680 15.000 2678.940 15.260 ;
      LAYER met2 ;
        RECT 2045.950 600.170 2046.230 604.000 ;
        RECT 2045.950 600.030 2047.760 600.170 ;
        RECT 2045.950 600.000 2046.230 600.030 ;
        RECT 2047.620 588.190 2047.760 600.030 ;
        RECT 2066.880 588.890 2067.140 589.210 ;
        RECT 2370.020 588.890 2370.280 589.210 ;
        RECT 2066.940 588.190 2067.080 588.890 ;
        RECT 2047.560 587.870 2047.820 588.190 ;
        RECT 2066.880 587.870 2067.140 588.190 ;
        RECT 2370.080 15.290 2370.220 588.890 ;
        RECT 2370.020 14.970 2370.280 15.290 ;
        RECT 2678.680 14.970 2678.940 15.290 ;
        RECT 2678.740 2.400 2678.880 14.970 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 19.280 2090.630 19.340 ;
        RECT 2696.590 19.280 2696.910 19.340 ;
        RECT 2090.310 19.140 2696.910 19.280 ;
        RECT 2090.310 19.080 2090.630 19.140 ;
        RECT 2696.590 19.080 2696.910 19.140 ;
        RECT 2055.810 15.200 2056.130 15.260 ;
        RECT 2090.310 15.200 2090.630 15.260 ;
        RECT 2055.810 15.060 2090.630 15.200 ;
        RECT 2055.810 15.000 2056.130 15.060 ;
        RECT 2090.310 15.000 2090.630 15.060 ;
      LAYER via ;
        RECT 2090.340 19.080 2090.600 19.340 ;
        RECT 2696.620 19.080 2696.880 19.340 ;
        RECT 2055.840 15.000 2056.100 15.260 ;
        RECT 2090.340 15.000 2090.600 15.260 ;
      LAYER met2 ;
        RECT 2055.150 600.170 2055.430 604.000 ;
        RECT 2055.150 600.030 2056.040 600.170 ;
        RECT 2055.150 600.000 2055.430 600.030 ;
        RECT 2055.900 15.290 2056.040 600.030 ;
        RECT 2090.340 19.050 2090.600 19.370 ;
        RECT 2696.620 19.050 2696.880 19.370 ;
        RECT 2090.400 15.290 2090.540 19.050 ;
        RECT 2055.840 14.970 2056.100 15.290 ;
        RECT 2090.340 14.970 2090.600 15.290 ;
        RECT 2696.680 2.400 2696.820 19.050 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2065.930 588.780 2066.250 588.840 ;
        RECT 2390.690 588.780 2391.010 588.840 ;
        RECT 2065.930 588.640 2391.010 588.780 ;
        RECT 2065.930 588.580 2066.250 588.640 ;
        RECT 2390.690 588.580 2391.010 588.640 ;
        RECT 2390.690 15.540 2391.010 15.600 ;
        RECT 2714.530 15.540 2714.850 15.600 ;
        RECT 2390.690 15.400 2714.850 15.540 ;
        RECT 2390.690 15.340 2391.010 15.400 ;
        RECT 2714.530 15.340 2714.850 15.400 ;
      LAYER via ;
        RECT 2065.960 588.580 2066.220 588.840 ;
        RECT 2390.720 588.580 2390.980 588.840 ;
        RECT 2390.720 15.340 2390.980 15.600 ;
        RECT 2714.560 15.340 2714.820 15.600 ;
      LAYER met2 ;
        RECT 2064.350 600.170 2064.630 604.000 ;
        RECT 2064.350 600.030 2066.160 600.170 ;
        RECT 2064.350 600.000 2064.630 600.030 ;
        RECT 2066.020 588.870 2066.160 600.030 ;
        RECT 2065.960 588.550 2066.220 588.870 ;
        RECT 2390.720 588.550 2390.980 588.870 ;
        RECT 2390.780 15.630 2390.920 588.550 ;
        RECT 2390.720 15.310 2390.980 15.630 ;
        RECT 2714.560 15.310 2714.820 15.630 ;
        RECT 2714.620 2.400 2714.760 15.310 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2075.590 545.260 2075.910 545.320 ;
        RECT 2076.510 545.260 2076.830 545.320 ;
        RECT 2075.590 545.120 2076.830 545.260 ;
        RECT 2075.590 545.060 2075.910 545.120 ;
        RECT 2076.510 545.060 2076.830 545.120 ;
        RECT 2076.510 18.940 2076.830 19.000 ;
        RECT 2732.470 18.940 2732.790 19.000 ;
        RECT 2076.510 18.800 2732.790 18.940 ;
        RECT 2076.510 18.740 2076.830 18.800 ;
        RECT 2732.470 18.740 2732.790 18.800 ;
      LAYER via ;
        RECT 2075.620 545.060 2075.880 545.320 ;
        RECT 2076.540 545.060 2076.800 545.320 ;
        RECT 2076.540 18.740 2076.800 19.000 ;
        RECT 2732.500 18.740 2732.760 19.000 ;
      LAYER met2 ;
        RECT 2073.550 600.170 2073.830 604.000 ;
        RECT 2073.550 600.030 2076.280 600.170 ;
        RECT 2073.550 600.000 2073.830 600.030 ;
        RECT 2076.140 593.370 2076.280 600.030 ;
        RECT 2075.680 593.230 2076.280 593.370 ;
        RECT 2075.680 545.350 2075.820 593.230 ;
        RECT 2075.620 545.030 2075.880 545.350 ;
        RECT 2076.540 545.030 2076.800 545.350 ;
        RECT 2076.600 19.030 2076.740 545.030 ;
        RECT 2076.540 18.710 2076.800 19.030 ;
        RECT 2732.500 18.710 2732.760 19.030 ;
        RECT 2732.560 2.400 2732.700 18.710 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2082.720 598.980 2083.040 599.040 ;
        RECT 2122.050 598.980 2122.370 599.040 ;
        RECT 2082.720 598.840 2122.370 598.980 ;
        RECT 2082.720 598.780 2083.040 598.840 ;
        RECT 2122.050 598.780 2122.370 598.840 ;
        RECT 2122.050 587.420 2122.370 587.480 ;
        RECT 2391.150 587.420 2391.470 587.480 ;
        RECT 2122.050 587.280 2145.740 587.420 ;
        RECT 2122.050 587.220 2122.370 587.280 ;
        RECT 2145.600 587.080 2145.740 587.280 ;
        RECT 2338.800 587.280 2391.470 587.420 ;
        RECT 2145.970 587.080 2146.290 587.140 ;
        RECT 2145.600 586.940 2146.290 587.080 ;
        RECT 2145.970 586.880 2146.290 586.940 ;
        RECT 2187.370 587.080 2187.690 587.140 ;
        RECT 2242.570 587.080 2242.890 587.140 ;
        RECT 2187.370 586.940 2194.960 587.080 ;
        RECT 2187.370 586.880 2187.690 586.940 ;
        RECT 2194.820 586.740 2194.960 586.940 ;
        RECT 2236.220 586.940 2242.890 587.080 ;
        RECT 2236.220 586.740 2236.360 586.940 ;
        RECT 2242.570 586.880 2242.890 586.940 ;
        RECT 2290.410 587.080 2290.730 587.140 ;
        RECT 2304.210 587.080 2304.530 587.140 ;
        RECT 2290.410 586.940 2304.530 587.080 ;
        RECT 2290.410 586.880 2290.730 586.940 ;
        RECT 2304.210 586.880 2304.530 586.940 ;
        RECT 2304.670 587.080 2304.990 587.140 ;
        RECT 2338.800 587.080 2338.940 587.280 ;
        RECT 2391.150 587.220 2391.470 587.280 ;
        RECT 2304.670 586.940 2338.940 587.080 ;
        RECT 2304.670 586.880 2304.990 586.940 ;
        RECT 2194.820 586.600 2236.360 586.740 ;
        RECT 2145.970 586.060 2146.290 586.120 ;
        RECT 2187.370 586.060 2187.690 586.120 ;
        RECT 2145.970 585.920 2187.690 586.060 ;
        RECT 2145.970 585.860 2146.290 585.920 ;
        RECT 2187.370 585.860 2187.690 585.920 ;
        RECT 2391.150 15.880 2391.470 15.940 ;
        RECT 2750.410 15.880 2750.730 15.940 ;
        RECT 2391.150 15.740 2750.730 15.880 ;
        RECT 2391.150 15.680 2391.470 15.740 ;
        RECT 2750.410 15.680 2750.730 15.740 ;
      LAYER via ;
        RECT 2082.750 598.780 2083.010 599.040 ;
        RECT 2122.080 598.780 2122.340 599.040 ;
        RECT 2122.080 587.220 2122.340 587.480 ;
        RECT 2146.000 586.880 2146.260 587.140 ;
        RECT 2187.400 586.880 2187.660 587.140 ;
        RECT 2242.600 586.880 2242.860 587.140 ;
        RECT 2290.440 586.880 2290.700 587.140 ;
        RECT 2304.240 586.880 2304.500 587.140 ;
        RECT 2304.700 586.880 2304.960 587.140 ;
        RECT 2391.180 587.220 2391.440 587.480 ;
        RECT 2146.000 585.860 2146.260 586.120 ;
        RECT 2187.400 585.860 2187.660 586.120 ;
        RECT 2391.180 15.680 2391.440 15.940 ;
        RECT 2750.440 15.680 2750.700 15.940 ;
      LAYER met2 ;
        RECT 2082.750 600.000 2083.030 604.000 ;
        RECT 2082.810 599.070 2082.950 600.000 ;
        RECT 2082.750 598.750 2083.010 599.070 ;
        RECT 2122.080 598.750 2122.340 599.070 ;
        RECT 2122.140 587.510 2122.280 598.750 ;
        RECT 2122.080 587.190 2122.340 587.510 ;
        RECT 2146.000 586.850 2146.260 587.170 ;
        RECT 2187.400 586.850 2187.660 587.170 ;
        RECT 2242.590 586.995 2242.870 587.365 ;
        RECT 2304.300 587.170 2304.900 587.250 ;
        RECT 2391.180 587.190 2391.440 587.510 ;
        RECT 2242.600 586.850 2242.860 586.995 ;
        RECT 2290.440 586.850 2290.700 587.170 ;
        RECT 2304.240 587.110 2304.960 587.170 ;
        RECT 2304.240 586.850 2304.500 587.110 ;
        RECT 2304.700 586.850 2304.960 587.110 ;
        RECT 2146.060 586.150 2146.200 586.850 ;
        RECT 2187.460 586.150 2187.600 586.850 ;
        RECT 2290.500 586.685 2290.640 586.850 ;
        RECT 2290.430 586.315 2290.710 586.685 ;
        RECT 2146.000 585.830 2146.260 586.150 ;
        RECT 2187.400 585.830 2187.660 586.150 ;
        RECT 2391.240 15.970 2391.380 587.190 ;
        RECT 2391.180 15.650 2391.440 15.970 ;
        RECT 2750.440 15.650 2750.700 15.970 ;
        RECT 2750.500 2.400 2750.640 15.650 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
      LAYER via2 ;
        RECT 2242.590 587.040 2242.870 587.320 ;
        RECT 2290.430 586.360 2290.710 586.640 ;
      LAYER met3 ;
        RECT 2242.565 587.330 2242.895 587.345 ;
        RECT 2242.565 587.030 2243.570 587.330 ;
        RECT 2242.565 587.015 2242.895 587.030 ;
        RECT 2243.270 586.650 2243.570 587.030 ;
        RECT 2290.405 586.650 2290.735 586.665 ;
        RECT 2243.270 586.350 2290.735 586.650 ;
        RECT 2290.405 586.335 2290.735 586.350 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2093.530 586.740 2093.850 586.800 ;
        RECT 2097.210 586.740 2097.530 586.800 ;
        RECT 2093.530 586.600 2097.530 586.740 ;
        RECT 2093.530 586.540 2093.850 586.600 ;
        RECT 2097.210 586.540 2097.530 586.600 ;
        RECT 2126.190 18.600 2126.510 18.660 ;
        RECT 2767.890 18.600 2768.210 18.660 ;
        RECT 2126.190 18.460 2768.210 18.600 ;
        RECT 2126.190 18.400 2126.510 18.460 ;
        RECT 2767.890 18.400 2768.210 18.460 ;
        RECT 2097.210 17.580 2097.530 17.640 ;
        RECT 2126.190 17.580 2126.510 17.640 ;
        RECT 2097.210 17.440 2126.510 17.580 ;
        RECT 2097.210 17.380 2097.530 17.440 ;
        RECT 2126.190 17.380 2126.510 17.440 ;
      LAYER via ;
        RECT 2093.560 586.540 2093.820 586.800 ;
        RECT 2097.240 586.540 2097.500 586.800 ;
        RECT 2126.220 18.400 2126.480 18.660 ;
        RECT 2767.920 18.400 2768.180 18.660 ;
        RECT 2097.240 17.380 2097.500 17.640 ;
        RECT 2126.220 17.380 2126.480 17.640 ;
      LAYER met2 ;
        RECT 2091.950 600.170 2092.230 604.000 ;
        RECT 2091.950 600.030 2093.760 600.170 ;
        RECT 2091.950 600.000 2092.230 600.030 ;
        RECT 2093.620 586.830 2093.760 600.030 ;
        RECT 2093.560 586.510 2093.820 586.830 ;
        RECT 2097.240 586.510 2097.500 586.830 ;
        RECT 2097.300 17.670 2097.440 586.510 ;
        RECT 2126.220 18.370 2126.480 18.690 ;
        RECT 2767.920 18.370 2768.180 18.690 ;
        RECT 2126.280 17.670 2126.420 18.370 ;
        RECT 2097.240 17.350 2097.500 17.670 ;
        RECT 2126.220 17.350 2126.480 17.670 ;
        RECT 2767.980 2.400 2768.120 18.370 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1098.090 420.820 1098.410 420.880 ;
        RECT 1099.010 420.820 1099.330 420.880 ;
        RECT 1098.090 420.680 1099.330 420.820 ;
        RECT 1098.090 420.620 1098.410 420.680 ;
        RECT 1099.010 420.620 1099.330 420.680 ;
        RECT 1097.630 372.880 1097.950 372.940 ;
        RECT 1099.010 372.880 1099.330 372.940 ;
        RECT 1097.630 372.740 1099.330 372.880 ;
        RECT 1097.630 372.680 1097.950 372.740 ;
        RECT 1099.010 372.680 1099.330 372.740 ;
        RECT 1097.630 331.400 1097.950 331.460 ;
        RECT 1098.090 331.400 1098.410 331.460 ;
        RECT 1097.630 331.260 1098.410 331.400 ;
        RECT 1097.630 331.200 1097.950 331.260 ;
        RECT 1098.090 331.200 1098.410 331.260 ;
        RECT 1098.090 324.260 1098.410 324.320 ;
        RECT 1099.010 324.260 1099.330 324.320 ;
        RECT 1098.090 324.120 1099.330 324.260 ;
        RECT 1098.090 324.060 1098.410 324.120 ;
        RECT 1099.010 324.060 1099.330 324.120 ;
        RECT 1097.630 276.320 1097.950 276.380 ;
        RECT 1099.010 276.320 1099.330 276.380 ;
        RECT 1097.630 276.180 1099.330 276.320 ;
        RECT 1097.630 276.120 1097.950 276.180 ;
        RECT 1099.010 276.120 1099.330 276.180 ;
        RECT 1097.630 227.700 1097.950 227.760 ;
        RECT 1098.090 227.700 1098.410 227.760 ;
        RECT 1097.630 227.560 1098.410 227.700 ;
        RECT 1097.630 227.500 1097.950 227.560 ;
        RECT 1098.090 227.500 1098.410 227.560 ;
        RECT 1098.090 131.140 1098.410 131.200 ;
        RECT 1098.550 131.140 1098.870 131.200 ;
        RECT 1098.090 131.000 1098.870 131.140 ;
        RECT 1098.090 130.940 1098.410 131.000 ;
        RECT 1098.550 130.940 1098.870 131.000 ;
        RECT 1097.630 41.720 1097.950 41.780 ;
        RECT 1098.090 41.720 1098.410 41.780 ;
        RECT 1097.630 41.580 1098.410 41.720 ;
        RECT 1097.630 41.520 1097.950 41.580 ;
        RECT 1098.090 41.520 1098.410 41.580 ;
        RECT 931.110 33.220 931.430 33.280 ;
        RECT 1097.630 33.220 1097.950 33.280 ;
        RECT 931.110 33.080 1097.950 33.220 ;
        RECT 931.110 33.020 931.430 33.080 ;
        RECT 1097.630 33.020 1097.950 33.080 ;
        RECT 840.950 14.860 841.270 14.920 ;
        RECT 840.950 14.720 883.500 14.860 ;
        RECT 840.950 14.660 841.270 14.720 ;
        RECT 883.360 14.520 883.500 14.720 ;
        RECT 931.110 14.520 931.430 14.580 ;
        RECT 883.360 14.380 931.430 14.520 ;
        RECT 931.110 14.320 931.430 14.380 ;
      LAYER via ;
        RECT 1098.120 420.620 1098.380 420.880 ;
        RECT 1099.040 420.620 1099.300 420.880 ;
        RECT 1097.660 372.680 1097.920 372.940 ;
        RECT 1099.040 372.680 1099.300 372.940 ;
        RECT 1097.660 331.200 1097.920 331.460 ;
        RECT 1098.120 331.200 1098.380 331.460 ;
        RECT 1098.120 324.060 1098.380 324.320 ;
        RECT 1099.040 324.060 1099.300 324.320 ;
        RECT 1097.660 276.120 1097.920 276.380 ;
        RECT 1099.040 276.120 1099.300 276.380 ;
        RECT 1097.660 227.500 1097.920 227.760 ;
        RECT 1098.120 227.500 1098.380 227.760 ;
        RECT 1098.120 130.940 1098.380 131.200 ;
        RECT 1098.580 130.940 1098.840 131.200 ;
        RECT 1097.660 41.520 1097.920 41.780 ;
        RECT 1098.120 41.520 1098.380 41.780 ;
        RECT 931.140 33.020 931.400 33.280 ;
        RECT 1097.660 33.020 1097.920 33.280 ;
        RECT 840.980 14.660 841.240 14.920 ;
        RECT 931.140 14.320 931.400 14.580 ;
      LAYER met2 ;
        RECT 1102.030 600.170 1102.310 604.000 ;
        RECT 1100.940 600.030 1102.310 600.170 ;
        RECT 1100.940 579.885 1101.080 600.030 ;
        RECT 1102.030 600.000 1102.310 600.030 ;
        RECT 1099.490 579.515 1099.770 579.885 ;
        RECT 1100.870 579.515 1101.150 579.885 ;
        RECT 1099.560 476.410 1099.700 579.515 ;
        RECT 1098.180 476.270 1099.700 476.410 ;
        RECT 1098.180 420.910 1098.320 476.270 ;
        RECT 1098.120 420.590 1098.380 420.910 ;
        RECT 1099.040 420.590 1099.300 420.910 ;
        RECT 1099.100 372.970 1099.240 420.590 ;
        RECT 1097.660 372.650 1097.920 372.970 ;
        RECT 1099.040 372.650 1099.300 372.970 ;
        RECT 1097.720 331.490 1097.860 372.650 ;
        RECT 1097.660 331.170 1097.920 331.490 ;
        RECT 1098.120 331.170 1098.380 331.490 ;
        RECT 1098.180 324.350 1098.320 331.170 ;
        RECT 1098.120 324.030 1098.380 324.350 ;
        RECT 1099.040 324.030 1099.300 324.350 ;
        RECT 1099.100 276.410 1099.240 324.030 ;
        RECT 1097.660 276.090 1097.920 276.410 ;
        RECT 1099.040 276.090 1099.300 276.410 ;
        RECT 1097.720 227.790 1097.860 276.090 ;
        RECT 1097.660 227.470 1097.920 227.790 ;
        RECT 1098.120 227.470 1098.380 227.790 ;
        RECT 1098.180 220.845 1098.320 227.470 ;
        RECT 1098.110 220.475 1098.390 220.845 ;
        RECT 1099.030 220.475 1099.310 220.845 ;
        RECT 1099.100 154.770 1099.240 220.475 ;
        RECT 1098.180 154.630 1099.240 154.770 ;
        RECT 1098.180 131.230 1098.320 154.630 ;
        RECT 1098.120 130.910 1098.380 131.230 ;
        RECT 1098.580 130.910 1098.840 131.230 ;
        RECT 1098.640 110.400 1098.780 130.910 ;
        RECT 1098.180 110.260 1098.780 110.400 ;
        RECT 1098.180 41.810 1098.320 110.260 ;
        RECT 1097.660 41.490 1097.920 41.810 ;
        RECT 1098.120 41.490 1098.380 41.810 ;
        RECT 1097.720 33.310 1097.860 41.490 ;
        RECT 931.140 32.990 931.400 33.310 ;
        RECT 1097.660 32.990 1097.920 33.310 ;
        RECT 840.980 14.630 841.240 14.950 ;
        RECT 841.040 2.400 841.180 14.630 ;
        RECT 931.200 14.610 931.340 32.990 ;
        RECT 931.140 14.290 931.400 14.610 ;
        RECT 840.830 -4.800 841.390 2.400 ;
      LAYER via2 ;
        RECT 1099.490 579.560 1099.770 579.840 ;
        RECT 1100.870 579.560 1101.150 579.840 ;
        RECT 1098.110 220.520 1098.390 220.800 ;
        RECT 1099.030 220.520 1099.310 220.800 ;
      LAYER met3 ;
        RECT 1099.465 579.850 1099.795 579.865 ;
        RECT 1100.845 579.850 1101.175 579.865 ;
        RECT 1099.465 579.550 1101.175 579.850 ;
        RECT 1099.465 579.535 1099.795 579.550 ;
        RECT 1100.845 579.535 1101.175 579.550 ;
        RECT 1098.085 220.810 1098.415 220.825 ;
        RECT 1099.005 220.810 1099.335 220.825 ;
        RECT 1098.085 220.510 1099.335 220.810 ;
        RECT 1098.085 220.495 1098.415 220.510 ;
        RECT 1099.005 220.495 1099.335 220.510 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2102.730 588.440 2103.050 588.500 ;
        RECT 2102.730 588.300 2131.480 588.440 ;
        RECT 2102.730 588.240 2103.050 588.300 ;
        RECT 2131.340 588.100 2131.480 588.300 ;
        RECT 2404.490 588.100 2404.810 588.160 ;
        RECT 2131.340 587.960 2404.810 588.100 ;
        RECT 2404.490 587.900 2404.810 587.960 ;
        RECT 2404.490 20.640 2404.810 20.700 ;
        RECT 2406.330 20.640 2406.650 20.700 ;
        RECT 2404.490 20.500 2406.650 20.640 ;
        RECT 2404.490 20.440 2404.810 20.500 ;
        RECT 2406.330 20.440 2406.650 20.500 ;
        RECT 2406.330 16.220 2406.650 16.280 ;
        RECT 2785.830 16.220 2786.150 16.280 ;
        RECT 2406.330 16.080 2786.150 16.220 ;
        RECT 2406.330 16.020 2406.650 16.080 ;
        RECT 2785.830 16.020 2786.150 16.080 ;
      LAYER via ;
        RECT 2102.760 588.240 2103.020 588.500 ;
        RECT 2404.520 587.900 2404.780 588.160 ;
        RECT 2404.520 20.440 2404.780 20.700 ;
        RECT 2406.360 20.440 2406.620 20.700 ;
        RECT 2406.360 16.020 2406.620 16.280 ;
        RECT 2785.860 16.020 2786.120 16.280 ;
      LAYER met2 ;
        RECT 2101.150 600.170 2101.430 604.000 ;
        RECT 2101.150 600.030 2102.960 600.170 ;
        RECT 2101.150 600.000 2101.430 600.030 ;
        RECT 2102.820 588.530 2102.960 600.030 ;
        RECT 2102.760 588.210 2103.020 588.530 ;
        RECT 2404.520 587.870 2404.780 588.190 ;
        RECT 2404.580 20.730 2404.720 587.870 ;
        RECT 2404.520 20.410 2404.780 20.730 ;
        RECT 2406.360 20.410 2406.620 20.730 ;
        RECT 2406.420 16.310 2406.560 20.410 ;
        RECT 2406.360 15.990 2406.620 16.310 ;
        RECT 2785.860 15.990 2786.120 16.310 ;
        RECT 2785.920 2.400 2786.060 15.990 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2111.010 17.920 2111.330 17.980 ;
        RECT 2803.770 17.920 2804.090 17.980 ;
        RECT 2111.010 17.780 2804.090 17.920 ;
        RECT 2111.010 17.720 2111.330 17.780 ;
        RECT 2803.770 17.720 2804.090 17.780 ;
      LAYER via ;
        RECT 2111.040 17.720 2111.300 17.980 ;
        RECT 2803.800 17.720 2804.060 17.980 ;
      LAYER met2 ;
        RECT 2110.350 600.170 2110.630 604.000 ;
        RECT 2110.350 600.030 2111.240 600.170 ;
        RECT 2110.350 600.000 2110.630 600.030 ;
        RECT 2111.100 18.010 2111.240 600.030 ;
        RECT 2111.040 17.690 2111.300 18.010 ;
        RECT 2803.800 17.690 2804.060 18.010 ;
        RECT 2803.860 2.400 2804.000 17.690 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2121.130 592.860 2121.450 592.920 ;
        RECT 2432.090 592.860 2432.410 592.920 ;
        RECT 2121.130 592.720 2432.410 592.860 ;
        RECT 2121.130 592.660 2121.450 592.720 ;
        RECT 2432.090 592.660 2432.410 592.720 ;
        RECT 2432.090 16.560 2432.410 16.620 ;
        RECT 2821.710 16.560 2822.030 16.620 ;
        RECT 2432.090 16.420 2822.030 16.560 ;
        RECT 2432.090 16.360 2432.410 16.420 ;
        RECT 2821.710 16.360 2822.030 16.420 ;
      LAYER via ;
        RECT 2121.160 592.660 2121.420 592.920 ;
        RECT 2432.120 592.660 2432.380 592.920 ;
        RECT 2432.120 16.360 2432.380 16.620 ;
        RECT 2821.740 16.360 2822.000 16.620 ;
      LAYER met2 ;
        RECT 2119.550 600.170 2119.830 604.000 ;
        RECT 2119.550 600.030 2121.360 600.170 ;
        RECT 2119.550 600.000 2119.830 600.030 ;
        RECT 2121.220 592.950 2121.360 600.030 ;
        RECT 2121.160 592.630 2121.420 592.950 ;
        RECT 2432.120 592.630 2432.380 592.950 ;
        RECT 2432.180 16.650 2432.320 592.630 ;
        RECT 2432.120 16.330 2432.380 16.650 ;
        RECT 2821.740 16.330 2822.000 16.650 ;
        RECT 2821.800 2.400 2821.940 16.330 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2130.330 586.740 2130.650 586.800 ;
        RECT 2131.710 586.740 2132.030 586.800 ;
        RECT 2130.330 586.600 2132.030 586.740 ;
        RECT 2130.330 586.540 2130.650 586.600 ;
        RECT 2131.710 586.540 2132.030 586.600 ;
        RECT 2131.250 17.580 2131.570 17.640 ;
        RECT 2839.190 17.580 2839.510 17.640 ;
        RECT 2131.250 17.440 2839.510 17.580 ;
        RECT 2131.250 17.380 2131.570 17.440 ;
        RECT 2839.190 17.380 2839.510 17.440 ;
      LAYER via ;
        RECT 2130.360 586.540 2130.620 586.800 ;
        RECT 2131.740 586.540 2132.000 586.800 ;
        RECT 2131.280 17.380 2131.540 17.640 ;
        RECT 2839.220 17.380 2839.480 17.640 ;
      LAYER met2 ;
        RECT 2128.750 600.170 2129.030 604.000 ;
        RECT 2128.750 600.030 2130.560 600.170 ;
        RECT 2128.750 600.000 2129.030 600.030 ;
        RECT 2130.420 586.830 2130.560 600.030 ;
        RECT 2130.360 586.510 2130.620 586.830 ;
        RECT 2131.740 586.510 2132.000 586.830 ;
        RECT 2131.800 44.610 2131.940 586.510 ;
        RECT 2131.340 44.470 2131.940 44.610 ;
        RECT 2131.340 17.670 2131.480 44.470 ;
        RECT 2131.280 17.350 2131.540 17.670 ;
        RECT 2839.220 17.350 2839.480 17.670 ;
        RECT 2839.280 2.400 2839.420 17.350 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2138.610 592.520 2138.930 592.580 ;
        RECT 2445.890 592.520 2446.210 592.580 ;
        RECT 2138.610 592.380 2446.210 592.520 ;
        RECT 2138.610 592.320 2138.930 592.380 ;
        RECT 2445.890 592.320 2446.210 592.380 ;
        RECT 2447.270 16.900 2447.590 16.960 ;
        RECT 2857.130 16.900 2857.450 16.960 ;
        RECT 2447.270 16.760 2857.450 16.900 ;
        RECT 2447.270 16.700 2447.590 16.760 ;
        RECT 2857.130 16.700 2857.450 16.760 ;
      LAYER via ;
        RECT 2138.640 592.320 2138.900 592.580 ;
        RECT 2445.920 592.320 2446.180 592.580 ;
        RECT 2447.300 16.700 2447.560 16.960 ;
        RECT 2857.160 16.700 2857.420 16.960 ;
      LAYER met2 ;
        RECT 2137.490 600.170 2137.770 604.000 ;
        RECT 2137.490 600.030 2138.840 600.170 ;
        RECT 2137.490 600.000 2137.770 600.030 ;
        RECT 2138.700 592.610 2138.840 600.030 ;
        RECT 2138.640 592.290 2138.900 592.610 ;
        RECT 2445.920 592.290 2446.180 592.610 ;
        RECT 2445.980 25.570 2446.120 592.290 ;
        RECT 2445.980 25.430 2447.500 25.570 ;
        RECT 2447.360 16.990 2447.500 25.430 ;
        RECT 2447.300 16.670 2447.560 16.990 ;
        RECT 2857.160 16.670 2857.420 16.990 ;
        RECT 2857.220 2.400 2857.360 16.670 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2146.660 598.980 2146.980 599.040 ;
        RECT 2190.590 598.980 2190.910 599.040 ;
        RECT 2146.660 598.840 2190.910 598.980 ;
        RECT 2146.660 598.780 2146.980 598.840 ;
        RECT 2190.590 598.780 2190.910 598.840 ;
        RECT 2190.590 18.260 2190.910 18.320 ;
        RECT 2875.070 18.260 2875.390 18.320 ;
        RECT 2190.590 18.120 2875.390 18.260 ;
        RECT 2190.590 18.060 2190.910 18.120 ;
        RECT 2875.070 18.060 2875.390 18.120 ;
      LAYER via ;
        RECT 2146.690 598.780 2146.950 599.040 ;
        RECT 2190.620 598.780 2190.880 599.040 ;
        RECT 2190.620 18.060 2190.880 18.320 ;
        RECT 2875.100 18.060 2875.360 18.320 ;
      LAYER met2 ;
        RECT 2146.690 600.000 2146.970 604.000 ;
        RECT 2146.750 599.070 2146.890 600.000 ;
        RECT 2146.690 598.750 2146.950 599.070 ;
        RECT 2190.620 598.750 2190.880 599.070 ;
        RECT 2190.680 18.350 2190.820 598.750 ;
        RECT 2190.620 18.030 2190.880 18.350 ;
        RECT 2875.100 18.030 2875.360 18.350 ;
        RECT 2875.160 2.400 2875.300 18.030 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2157.470 592.180 2157.790 592.240 ;
        RECT 2466.590 592.180 2466.910 592.240 ;
        RECT 2157.470 592.040 2466.910 592.180 ;
        RECT 2157.470 591.980 2157.790 592.040 ;
        RECT 2466.590 591.980 2466.910 592.040 ;
        RECT 2466.590 20.640 2466.910 20.700 ;
        RECT 2893.010 20.640 2893.330 20.700 ;
        RECT 2466.590 20.500 2893.330 20.640 ;
        RECT 2466.590 20.440 2466.910 20.500 ;
        RECT 2893.010 20.440 2893.330 20.500 ;
      LAYER via ;
        RECT 2157.500 591.980 2157.760 592.240 ;
        RECT 2466.620 591.980 2466.880 592.240 ;
        RECT 2466.620 20.440 2466.880 20.700 ;
        RECT 2893.040 20.440 2893.300 20.700 ;
      LAYER met2 ;
        RECT 2155.890 600.170 2156.170 604.000 ;
        RECT 2155.890 600.030 2157.700 600.170 ;
        RECT 2155.890 600.000 2156.170 600.030 ;
        RECT 2157.560 592.270 2157.700 600.030 ;
        RECT 2157.500 591.950 2157.760 592.270 ;
        RECT 2466.620 591.950 2466.880 592.270 ;
        RECT 2466.680 20.730 2466.820 591.950 ;
        RECT 2466.620 20.410 2466.880 20.730 ;
        RECT 2893.040 20.410 2893.300 20.730 ;
        RECT 2893.100 2.400 2893.240 20.410 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2166.210 18.260 2166.530 18.320 ;
        RECT 2179.550 18.260 2179.870 18.320 ;
        RECT 2166.210 18.120 2179.870 18.260 ;
        RECT 2166.210 18.060 2166.530 18.120 ;
        RECT 2179.550 18.060 2179.870 18.120 ;
        RECT 2179.550 17.240 2179.870 17.300 ;
        RECT 2910.950 17.240 2911.270 17.300 ;
        RECT 2179.550 17.100 2911.270 17.240 ;
        RECT 2179.550 17.040 2179.870 17.100 ;
        RECT 2910.950 17.040 2911.270 17.100 ;
      LAYER via ;
        RECT 2166.240 18.060 2166.500 18.320 ;
        RECT 2179.580 18.060 2179.840 18.320 ;
        RECT 2179.580 17.040 2179.840 17.300 ;
        RECT 2910.980 17.040 2911.240 17.300 ;
      LAYER met2 ;
        RECT 2165.090 600.170 2165.370 604.000 ;
        RECT 2165.090 600.030 2166.440 600.170 ;
        RECT 2165.090 600.000 2165.370 600.030 ;
        RECT 2166.300 18.350 2166.440 600.030 ;
        RECT 2166.240 18.030 2166.500 18.350 ;
        RECT 2179.580 18.030 2179.840 18.350 ;
        RECT 2179.640 17.330 2179.780 18.030 ;
        RECT 2179.580 17.010 2179.840 17.330 ;
        RECT 2910.980 17.010 2911.240 17.330 ;
        RECT 2911.040 2.400 2911.180 17.010 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 955.030 32.880 955.350 32.940 ;
        RECT 1111.430 32.880 1111.750 32.940 ;
        RECT 955.030 32.740 1111.750 32.880 ;
        RECT 955.030 32.680 955.350 32.740 ;
        RECT 1111.430 32.680 1111.750 32.740 ;
        RECT 858.890 15.540 859.210 15.600 ;
        RECT 955.030 15.540 955.350 15.600 ;
        RECT 858.890 15.400 955.350 15.540 ;
        RECT 858.890 15.340 859.210 15.400 ;
        RECT 955.030 15.340 955.350 15.400 ;
      LAYER via ;
        RECT 955.060 32.680 955.320 32.940 ;
        RECT 1111.460 32.680 1111.720 32.940 ;
        RECT 858.920 15.340 859.180 15.600 ;
        RECT 955.060 15.340 955.320 15.600 ;
      LAYER met2 ;
        RECT 1111.230 600.000 1111.510 604.000 ;
        RECT 1111.290 598.810 1111.430 600.000 ;
        RECT 1111.290 598.670 1111.660 598.810 ;
        RECT 1111.520 32.970 1111.660 598.670 ;
        RECT 955.060 32.650 955.320 32.970 ;
        RECT 1111.460 32.650 1111.720 32.970 ;
        RECT 955.120 15.630 955.260 32.650 ;
        RECT 858.920 15.310 859.180 15.630 ;
        RECT 955.060 15.310 955.320 15.630 ;
        RECT 858.980 2.400 859.120 15.310 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 591.160 883.130 591.220 ;
        RECT 1118.790 591.160 1119.110 591.220 ;
        RECT 882.810 591.020 1119.110 591.160 ;
        RECT 882.810 590.960 883.130 591.020 ;
        RECT 1118.790 590.960 1119.110 591.020 ;
        RECT 876.830 18.940 877.150 19.000 ;
        RECT 882.810 18.940 883.130 19.000 ;
        RECT 876.830 18.800 883.130 18.940 ;
        RECT 876.830 18.740 877.150 18.800 ;
        RECT 882.810 18.740 883.130 18.800 ;
      LAYER via ;
        RECT 882.840 590.960 883.100 591.220 ;
        RECT 1118.820 590.960 1119.080 591.220 ;
        RECT 876.860 18.740 877.120 19.000 ;
        RECT 882.840 18.740 883.100 19.000 ;
      LAYER met2 ;
        RECT 1120.430 600.170 1120.710 604.000 ;
        RECT 1118.880 600.030 1120.710 600.170 ;
        RECT 1118.880 591.250 1119.020 600.030 ;
        RECT 1120.430 600.000 1120.710 600.030 ;
        RECT 882.840 590.930 883.100 591.250 ;
        RECT 1118.820 590.930 1119.080 591.250 ;
        RECT 882.900 19.030 883.040 590.930 ;
        RECT 876.860 18.710 877.120 19.030 ;
        RECT 882.840 18.710 883.100 19.030 ;
        RECT 876.920 2.400 877.060 18.710 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.610 590.820 896.930 590.880 ;
        RECT 1127.990 590.820 1128.310 590.880 ;
        RECT 896.610 590.680 1128.310 590.820 ;
        RECT 896.610 590.620 896.930 590.680 ;
        RECT 1127.990 590.620 1128.310 590.680 ;
        RECT 894.770 2.960 895.090 3.020 ;
        RECT 896.610 2.960 896.930 3.020 ;
        RECT 894.770 2.820 896.930 2.960 ;
        RECT 894.770 2.760 895.090 2.820 ;
        RECT 896.610 2.760 896.930 2.820 ;
      LAYER via ;
        RECT 896.640 590.620 896.900 590.880 ;
        RECT 1128.020 590.620 1128.280 590.880 ;
        RECT 894.800 2.760 895.060 3.020 ;
        RECT 896.640 2.760 896.900 3.020 ;
      LAYER met2 ;
        RECT 1129.630 600.170 1129.910 604.000 ;
        RECT 1128.080 600.030 1129.910 600.170 ;
        RECT 1128.080 590.910 1128.220 600.030 ;
        RECT 1129.630 600.000 1129.910 600.030 ;
        RECT 896.640 590.590 896.900 590.910 ;
        RECT 1128.020 590.590 1128.280 590.910 ;
        RECT 896.700 3.050 896.840 590.590 ;
        RECT 894.800 2.730 895.060 3.050 ;
        RECT 896.640 2.730 896.900 3.050 ;
        RECT 894.860 2.400 895.000 2.730 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 591.500 917.630 591.560 ;
        RECT 1139.030 591.500 1139.350 591.560 ;
        RECT 917.310 591.360 1139.350 591.500 ;
        RECT 917.310 591.300 917.630 591.360 ;
        RECT 1139.030 591.300 1139.350 591.360 ;
        RECT 912.710 20.640 913.030 20.700 ;
        RECT 917.310 20.640 917.630 20.700 ;
        RECT 912.710 20.500 917.630 20.640 ;
        RECT 912.710 20.440 913.030 20.500 ;
        RECT 917.310 20.440 917.630 20.500 ;
      LAYER via ;
        RECT 917.340 591.300 917.600 591.560 ;
        RECT 1139.060 591.300 1139.320 591.560 ;
        RECT 912.740 20.440 913.000 20.700 ;
        RECT 917.340 20.440 917.600 20.700 ;
      LAYER met2 ;
        RECT 1138.830 600.000 1139.110 604.000 ;
        RECT 1138.890 598.810 1139.030 600.000 ;
        RECT 1138.890 598.670 1139.260 598.810 ;
        RECT 1139.120 591.590 1139.260 598.670 ;
        RECT 917.340 591.270 917.600 591.590 ;
        RECT 1139.060 591.270 1139.320 591.590 ;
        RECT 917.400 20.730 917.540 591.270 ;
        RECT 912.740 20.410 913.000 20.730 ;
        RECT 917.340 20.410 917.600 20.730 ;
        RECT 912.800 2.400 912.940 20.410 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1128.450 586.740 1128.770 586.800 ;
        RECT 1146.390 586.740 1146.710 586.800 ;
        RECT 1128.450 586.600 1146.710 586.740 ;
        RECT 1128.450 586.540 1128.770 586.600 ;
        RECT 1146.390 586.540 1146.710 586.600 ;
        RECT 930.190 19.620 930.510 19.680 ;
        RECT 930.190 19.480 1082.220 19.620 ;
        RECT 930.190 19.420 930.510 19.480 ;
        RECT 1082.080 19.280 1082.220 19.480 ;
        RECT 1128.450 19.280 1128.770 19.340 ;
        RECT 1082.080 19.140 1128.770 19.280 ;
        RECT 1128.450 19.080 1128.770 19.140 ;
      LAYER via ;
        RECT 1128.480 586.540 1128.740 586.800 ;
        RECT 1146.420 586.540 1146.680 586.800 ;
        RECT 930.220 19.420 930.480 19.680 ;
        RECT 1128.480 19.080 1128.740 19.340 ;
      LAYER met2 ;
        RECT 1148.030 600.170 1148.310 604.000 ;
        RECT 1146.480 600.030 1148.310 600.170 ;
        RECT 1146.480 586.830 1146.620 600.030 ;
        RECT 1148.030 600.000 1148.310 600.030 ;
        RECT 1128.480 586.510 1128.740 586.830 ;
        RECT 1146.420 586.510 1146.680 586.830 ;
        RECT 930.220 19.390 930.480 19.710 ;
        RECT 930.280 2.400 930.420 19.390 ;
        RECT 1128.540 19.370 1128.680 586.510 ;
        RECT 1128.480 19.050 1128.740 19.370 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 593.200 952.130 593.260 ;
        RECT 1155.590 593.200 1155.910 593.260 ;
        RECT 951.810 593.060 1155.910 593.200 ;
        RECT 951.810 593.000 952.130 593.060 ;
        RECT 1155.590 593.000 1155.910 593.060 ;
        RECT 948.130 19.960 948.450 20.020 ;
        RECT 951.810 19.960 952.130 20.020 ;
        RECT 948.130 19.820 952.130 19.960 ;
        RECT 948.130 19.760 948.450 19.820 ;
        RECT 951.810 19.760 952.130 19.820 ;
      LAYER via ;
        RECT 951.840 593.000 952.100 593.260 ;
        RECT 1155.620 593.000 1155.880 593.260 ;
        RECT 948.160 19.760 948.420 20.020 ;
        RECT 951.840 19.760 952.100 20.020 ;
      LAYER met2 ;
        RECT 1157.230 600.170 1157.510 604.000 ;
        RECT 1155.680 600.030 1157.510 600.170 ;
        RECT 1155.680 593.290 1155.820 600.030 ;
        RECT 1157.230 600.000 1157.510 600.030 ;
        RECT 951.840 592.970 952.100 593.290 ;
        RECT 1155.620 592.970 1155.880 593.290 ;
        RECT 951.900 20.050 952.040 592.970 ;
        RECT 948.160 19.730 948.420 20.050 ;
        RECT 951.840 19.730 952.100 20.050 ;
        RECT 948.220 2.400 948.360 19.730 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.510 591.840 972.830 591.900 ;
        RECT 1166.170 591.840 1166.490 591.900 ;
        RECT 972.510 591.700 1166.490 591.840 ;
        RECT 972.510 591.640 972.830 591.700 ;
        RECT 1166.170 591.640 1166.490 591.700 ;
        RECT 966.070 11.800 966.390 11.860 ;
        RECT 972.510 11.800 972.830 11.860 ;
        RECT 966.070 11.660 972.830 11.800 ;
        RECT 966.070 11.600 966.390 11.660 ;
        RECT 972.510 11.600 972.830 11.660 ;
      LAYER via ;
        RECT 972.540 591.640 972.800 591.900 ;
        RECT 1166.200 591.640 1166.460 591.900 ;
        RECT 966.100 11.600 966.360 11.860 ;
        RECT 972.540 11.600 972.800 11.860 ;
      LAYER met2 ;
        RECT 1165.970 600.000 1166.250 604.000 ;
        RECT 1166.030 598.810 1166.170 600.000 ;
        RECT 1166.030 598.670 1166.400 598.810 ;
        RECT 1166.260 591.930 1166.400 598.670 ;
        RECT 972.540 591.610 972.800 591.930 ;
        RECT 1166.200 591.610 1166.460 591.930 ;
        RECT 972.600 11.890 972.740 591.610 ;
        RECT 966.100 11.570 966.360 11.890 ;
        RECT 972.540 11.570 972.800 11.890 ;
        RECT 966.160 2.400 966.300 11.570 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1114.190 588.100 1114.510 588.160 ;
        RECT 1173.530 588.100 1173.850 588.160 ;
        RECT 1114.190 587.960 1173.850 588.100 ;
        RECT 1114.190 587.900 1114.510 587.960 ;
        RECT 1173.530 587.900 1173.850 587.960 ;
        RECT 1080.610 17.580 1080.930 17.640 ;
        RECT 1114.190 17.580 1114.510 17.640 ;
        RECT 1080.610 17.440 1114.510 17.580 ;
        RECT 1080.610 17.380 1080.930 17.440 ;
        RECT 1114.190 17.380 1114.510 17.440 ;
        RECT 984.010 16.560 984.330 16.620 ;
        RECT 1080.610 16.560 1080.930 16.620 ;
        RECT 984.010 16.420 1080.930 16.560 ;
        RECT 984.010 16.360 984.330 16.420 ;
        RECT 1080.610 16.360 1080.930 16.420 ;
      LAYER via ;
        RECT 1114.220 587.900 1114.480 588.160 ;
        RECT 1173.560 587.900 1173.820 588.160 ;
        RECT 1080.640 17.380 1080.900 17.640 ;
        RECT 1114.220 17.380 1114.480 17.640 ;
        RECT 984.040 16.360 984.300 16.620 ;
        RECT 1080.640 16.360 1080.900 16.620 ;
      LAYER met2 ;
        RECT 1175.170 600.170 1175.450 604.000 ;
        RECT 1173.620 600.030 1175.450 600.170 ;
        RECT 1173.620 588.190 1173.760 600.030 ;
        RECT 1175.170 600.000 1175.450 600.030 ;
        RECT 1114.220 587.870 1114.480 588.190 ;
        RECT 1173.560 587.870 1173.820 588.190 ;
        RECT 1114.280 17.670 1114.420 587.870 ;
        RECT 1080.640 17.350 1080.900 17.670 ;
        RECT 1114.220 17.350 1114.480 17.670 ;
        RECT 1080.700 16.650 1080.840 17.350 ;
        RECT 984.040 16.330 984.300 16.650 ;
        RECT 1080.640 16.330 1080.900 16.650 ;
        RECT 984.100 2.400 984.240 16.330 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.450 45.460 668.770 45.520 ;
        RECT 1008.390 45.460 1008.710 45.520 ;
        RECT 668.450 45.320 1008.710 45.460 ;
        RECT 668.450 45.260 668.770 45.320 ;
        RECT 1008.390 45.260 1008.710 45.320 ;
        RECT 662.930 41.720 663.250 41.780 ;
        RECT 668.450 41.720 668.770 41.780 ;
        RECT 662.930 41.580 668.770 41.720 ;
        RECT 662.930 41.520 663.250 41.580 ;
        RECT 668.450 41.520 668.770 41.580 ;
      LAYER via ;
        RECT 668.480 45.260 668.740 45.520 ;
        RECT 1008.420 45.260 1008.680 45.520 ;
        RECT 662.960 41.520 663.220 41.780 ;
        RECT 668.480 41.520 668.740 41.780 ;
      LAYER met2 ;
        RECT 1010.490 600.170 1010.770 604.000 ;
        RECT 1008.480 600.030 1010.770 600.170 ;
        RECT 1008.480 45.550 1008.620 600.030 ;
        RECT 1010.490 600.000 1010.770 600.030 ;
        RECT 668.480 45.230 668.740 45.550 ;
        RECT 1008.420 45.230 1008.680 45.550 ;
        RECT 668.540 41.810 668.680 45.230 ;
        RECT 662.960 41.490 663.220 41.810 ;
        RECT 668.480 41.490 668.740 41.810 ;
        RECT 663.020 2.400 663.160 41.490 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1182.730 591.840 1183.050 591.900 ;
        RECT 1166.720 591.700 1183.050 591.840 ;
        RECT 1166.720 591.500 1166.860 591.700 ;
        RECT 1182.730 591.640 1183.050 591.700 ;
        RECT 1139.580 591.360 1166.860 591.500 ;
        RECT 1128.450 591.160 1128.770 591.220 ;
        RECT 1139.580 591.160 1139.720 591.360 ;
        RECT 1128.450 591.020 1139.720 591.160 ;
        RECT 1128.450 590.960 1128.770 591.020 ;
        RECT 1001.950 15.540 1002.270 15.600 ;
        RECT 1127.990 15.540 1128.310 15.600 ;
        RECT 1001.950 15.400 1128.310 15.540 ;
        RECT 1001.950 15.340 1002.270 15.400 ;
        RECT 1127.990 15.340 1128.310 15.400 ;
      LAYER via ;
        RECT 1182.760 591.640 1183.020 591.900 ;
        RECT 1128.480 590.960 1128.740 591.220 ;
        RECT 1001.980 15.340 1002.240 15.600 ;
        RECT 1128.020 15.340 1128.280 15.600 ;
      LAYER met2 ;
        RECT 1184.370 600.170 1184.650 604.000 ;
        RECT 1182.820 600.030 1184.650 600.170 ;
        RECT 1182.820 591.930 1182.960 600.030 ;
        RECT 1184.370 600.000 1184.650 600.030 ;
        RECT 1182.760 591.610 1183.020 591.930 ;
        RECT 1128.480 590.930 1128.740 591.250 ;
        RECT 1128.540 587.250 1128.680 590.930 ;
        RECT 1128.080 587.110 1128.680 587.250 ;
        RECT 1128.080 15.630 1128.220 587.110 ;
        RECT 1001.980 15.310 1002.240 15.630 ;
        RECT 1128.020 15.310 1128.280 15.630 ;
        RECT 1002.040 2.400 1002.180 15.310 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1148.230 587.420 1148.550 587.480 ;
        RECT 1193.770 587.420 1194.090 587.480 ;
        RECT 1148.230 587.280 1194.090 587.420 ;
        RECT 1148.230 587.220 1148.550 587.280 ;
        RECT 1193.770 587.220 1194.090 587.280 ;
        RECT 1148.690 531.320 1149.010 531.380 ;
        RECT 1149.150 531.320 1149.470 531.380 ;
        RECT 1148.690 531.180 1149.470 531.320 ;
        RECT 1148.690 531.120 1149.010 531.180 ;
        RECT 1149.150 531.120 1149.470 531.180 ;
        RECT 1149.150 496.980 1149.470 497.040 ;
        RECT 1148.780 496.840 1149.470 496.980 ;
        RECT 1148.780 496.700 1148.920 496.840 ;
        RECT 1149.150 496.780 1149.470 496.840 ;
        RECT 1148.690 496.440 1149.010 496.700 ;
        RECT 1148.230 448.700 1148.550 448.760 ;
        RECT 1149.150 448.700 1149.470 448.760 ;
        RECT 1148.230 448.560 1149.470 448.700 ;
        RECT 1148.230 448.500 1148.550 448.560 ;
        RECT 1149.150 448.500 1149.470 448.560 ;
        RECT 1148.690 145.080 1149.010 145.140 ;
        RECT 1149.150 145.080 1149.470 145.140 ;
        RECT 1148.690 144.940 1149.470 145.080 ;
        RECT 1148.690 144.880 1149.010 144.940 ;
        RECT 1149.150 144.880 1149.470 144.940 ;
        RECT 1019.430 16.220 1019.750 16.280 ;
        RECT 1148.230 16.220 1148.550 16.280 ;
        RECT 1019.430 16.080 1148.550 16.220 ;
        RECT 1019.430 16.020 1019.750 16.080 ;
        RECT 1148.230 16.020 1148.550 16.080 ;
      LAYER via ;
        RECT 1148.260 587.220 1148.520 587.480 ;
        RECT 1193.800 587.220 1194.060 587.480 ;
        RECT 1148.720 531.120 1148.980 531.380 ;
        RECT 1149.180 531.120 1149.440 531.380 ;
        RECT 1149.180 496.780 1149.440 497.040 ;
        RECT 1148.720 496.440 1148.980 496.700 ;
        RECT 1148.260 448.500 1148.520 448.760 ;
        RECT 1149.180 448.500 1149.440 448.760 ;
        RECT 1148.720 144.880 1148.980 145.140 ;
        RECT 1149.180 144.880 1149.440 145.140 ;
        RECT 1019.460 16.020 1019.720 16.280 ;
        RECT 1148.260 16.020 1148.520 16.280 ;
      LAYER met2 ;
        RECT 1193.570 600.000 1193.850 604.000 ;
        RECT 1193.630 598.810 1193.770 600.000 ;
        RECT 1193.630 598.670 1194.000 598.810 ;
        RECT 1193.860 587.510 1194.000 598.670 ;
        RECT 1148.260 587.190 1148.520 587.510 ;
        RECT 1193.800 587.190 1194.060 587.510 ;
        RECT 1148.320 545.090 1148.460 587.190 ;
        RECT 1148.320 544.950 1148.920 545.090 ;
        RECT 1148.780 531.410 1148.920 544.950 ;
        RECT 1148.720 531.090 1148.980 531.410 ;
        RECT 1149.180 531.090 1149.440 531.410 ;
        RECT 1149.240 497.070 1149.380 531.090 ;
        RECT 1149.180 496.750 1149.440 497.070 ;
        RECT 1148.720 496.410 1148.980 496.730 ;
        RECT 1148.780 483.210 1148.920 496.410 ;
        RECT 1148.780 483.070 1149.380 483.210 ;
        RECT 1149.240 448.790 1149.380 483.070 ;
        RECT 1148.260 448.530 1148.520 448.790 ;
        RECT 1148.260 448.470 1148.920 448.530 ;
        RECT 1149.180 448.470 1149.440 448.790 ;
        RECT 1148.320 448.390 1148.920 448.470 ;
        RECT 1148.780 447.850 1148.920 448.390 ;
        RECT 1148.780 447.710 1149.380 447.850 ;
        RECT 1149.240 351.290 1149.380 447.710 ;
        RECT 1148.780 351.150 1149.380 351.290 ;
        RECT 1148.780 303.690 1148.920 351.150 ;
        RECT 1148.780 303.550 1149.380 303.690 ;
        RECT 1149.240 145.170 1149.380 303.550 ;
        RECT 1148.720 144.850 1148.980 145.170 ;
        RECT 1149.180 144.850 1149.440 145.170 ;
        RECT 1148.780 110.570 1148.920 144.850 ;
        RECT 1148.780 110.430 1149.380 110.570 ;
        RECT 1149.240 62.290 1149.380 110.430 ;
        RECT 1148.320 62.150 1149.380 62.290 ;
        RECT 1148.320 16.310 1148.460 62.150 ;
        RECT 1019.460 15.990 1019.720 16.310 ;
        RECT 1148.260 15.990 1148.520 16.310 ;
        RECT 1019.520 2.400 1019.660 15.990 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.950 592.520 1163.270 592.580 ;
        RECT 1201.130 592.520 1201.450 592.580 ;
        RECT 1162.950 592.380 1201.450 592.520 ;
        RECT 1162.950 592.320 1163.270 592.380 ;
        RECT 1201.130 592.320 1201.450 592.380 ;
        RECT 1037.370 15.880 1037.690 15.940 ;
        RECT 1162.950 15.880 1163.270 15.940 ;
        RECT 1037.370 15.740 1163.270 15.880 ;
        RECT 1037.370 15.680 1037.690 15.740 ;
        RECT 1162.950 15.680 1163.270 15.740 ;
      LAYER via ;
        RECT 1162.980 592.320 1163.240 592.580 ;
        RECT 1201.160 592.320 1201.420 592.580 ;
        RECT 1037.400 15.680 1037.660 15.940 ;
        RECT 1162.980 15.680 1163.240 15.940 ;
      LAYER met2 ;
        RECT 1202.770 600.170 1203.050 604.000 ;
        RECT 1201.220 600.030 1203.050 600.170 ;
        RECT 1201.220 592.610 1201.360 600.030 ;
        RECT 1202.770 600.000 1203.050 600.030 ;
        RECT 1162.980 592.290 1163.240 592.610 ;
        RECT 1201.160 592.290 1201.420 592.610 ;
        RECT 1163.040 15.970 1163.180 592.290 ;
        RECT 1037.400 15.650 1037.660 15.970 ;
        RECT 1162.980 15.650 1163.240 15.970 ;
        RECT 1037.460 2.400 1037.600 15.650 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.990 586.740 1197.310 586.800 ;
        RECT 1210.330 586.740 1210.650 586.800 ;
        RECT 1196.990 586.600 1210.650 586.740 ;
        RECT 1196.990 586.540 1197.310 586.600 ;
        RECT 1210.330 586.540 1210.650 586.600 ;
        RECT 1163.410 22.680 1163.730 22.740 ;
        RECT 1196.990 22.680 1197.310 22.740 ;
        RECT 1163.410 22.540 1197.310 22.680 ;
        RECT 1163.410 22.480 1163.730 22.540 ;
        RECT 1196.990 22.480 1197.310 22.540 ;
        RECT 1055.310 16.900 1055.630 16.960 ;
        RECT 1163.410 16.900 1163.730 16.960 ;
        RECT 1055.310 16.760 1163.730 16.900 ;
        RECT 1055.310 16.700 1055.630 16.760 ;
        RECT 1163.410 16.700 1163.730 16.760 ;
      LAYER via ;
        RECT 1197.020 586.540 1197.280 586.800 ;
        RECT 1210.360 586.540 1210.620 586.800 ;
        RECT 1163.440 22.480 1163.700 22.740 ;
        RECT 1197.020 22.480 1197.280 22.740 ;
        RECT 1055.340 16.700 1055.600 16.960 ;
        RECT 1163.440 16.700 1163.700 16.960 ;
      LAYER met2 ;
        RECT 1211.970 600.170 1212.250 604.000 ;
        RECT 1210.420 600.030 1212.250 600.170 ;
        RECT 1210.420 586.830 1210.560 600.030 ;
        RECT 1211.970 600.000 1212.250 600.030 ;
        RECT 1197.020 586.510 1197.280 586.830 ;
        RECT 1210.360 586.510 1210.620 586.830 ;
        RECT 1197.080 22.770 1197.220 586.510 ;
        RECT 1163.440 22.450 1163.700 22.770 ;
        RECT 1197.020 22.450 1197.280 22.770 ;
        RECT 1163.500 16.990 1163.640 22.450 ;
        RECT 1055.340 16.670 1055.600 16.990 ;
        RECT 1163.440 16.670 1163.700 16.990 ;
        RECT 1055.400 2.400 1055.540 16.670 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 589.120 1076.330 589.180 ;
        RECT 1221.370 589.120 1221.690 589.180 ;
        RECT 1076.010 588.980 1221.690 589.120 ;
        RECT 1076.010 588.920 1076.330 588.980 ;
        RECT 1221.370 588.920 1221.690 588.980 ;
        RECT 1073.250 17.580 1073.570 17.640 ;
        RECT 1076.010 17.580 1076.330 17.640 ;
        RECT 1073.250 17.440 1076.330 17.580 ;
        RECT 1073.250 17.380 1073.570 17.440 ;
        RECT 1076.010 17.380 1076.330 17.440 ;
      LAYER via ;
        RECT 1076.040 588.920 1076.300 589.180 ;
        RECT 1221.400 588.920 1221.660 589.180 ;
        RECT 1073.280 17.380 1073.540 17.640 ;
        RECT 1076.040 17.380 1076.300 17.640 ;
      LAYER met2 ;
        RECT 1221.170 600.000 1221.450 604.000 ;
        RECT 1221.230 598.810 1221.370 600.000 ;
        RECT 1221.230 598.670 1221.600 598.810 ;
        RECT 1221.460 589.210 1221.600 598.670 ;
        RECT 1076.040 588.890 1076.300 589.210 ;
        RECT 1221.400 588.890 1221.660 589.210 ;
        RECT 1076.100 17.670 1076.240 588.890 ;
        RECT 1073.280 17.350 1073.540 17.670 ;
        RECT 1076.040 17.350 1076.300 17.670 ;
        RECT 1073.340 2.400 1073.480 17.350 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1111.430 17.240 1111.750 17.300 ;
        RECT 1172.610 17.240 1172.930 17.300 ;
        RECT 1111.430 17.100 1172.930 17.240 ;
        RECT 1111.430 17.040 1111.750 17.100 ;
        RECT 1172.610 17.040 1172.930 17.100 ;
        RECT 1173.070 16.900 1173.390 16.960 ;
        RECT 1229.190 16.900 1229.510 16.960 ;
        RECT 1173.070 16.760 1229.510 16.900 ;
        RECT 1173.070 16.700 1173.390 16.760 ;
        RECT 1229.190 16.700 1229.510 16.760 ;
        RECT 1090.730 5.000 1091.050 5.060 ;
        RECT 1110.050 5.000 1110.370 5.060 ;
        RECT 1090.730 4.860 1110.370 5.000 ;
        RECT 1090.730 4.800 1091.050 4.860 ;
        RECT 1110.050 4.800 1110.370 4.860 ;
      LAYER via ;
        RECT 1111.460 17.040 1111.720 17.300 ;
        RECT 1172.640 17.040 1172.900 17.300 ;
        RECT 1173.100 16.700 1173.360 16.960 ;
        RECT 1229.220 16.700 1229.480 16.960 ;
        RECT 1090.760 4.800 1091.020 5.060 ;
        RECT 1110.080 4.800 1110.340 5.060 ;
      LAYER met2 ;
        RECT 1230.370 600.170 1230.650 604.000 ;
        RECT 1229.280 600.030 1230.650 600.170 ;
        RECT 1172.700 17.330 1173.300 17.410 ;
        RECT 1111.460 17.240 1111.720 17.330 ;
        RECT 1110.140 17.100 1111.720 17.240 ;
        RECT 1110.140 5.090 1110.280 17.100 ;
        RECT 1111.460 17.010 1111.720 17.100 ;
        RECT 1172.640 17.270 1173.300 17.330 ;
        RECT 1172.640 17.010 1172.900 17.270 ;
        RECT 1173.160 16.990 1173.300 17.270 ;
        RECT 1229.280 16.990 1229.420 600.030 ;
        RECT 1230.370 600.000 1230.650 600.030 ;
        RECT 1173.100 16.670 1173.360 16.990 ;
        RECT 1229.220 16.670 1229.480 16.990 ;
        RECT 1090.760 4.770 1091.020 5.090 ;
        RECT 1110.080 4.770 1110.340 5.090 ;
        RECT 1090.820 2.400 1090.960 4.770 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1169.390 587.760 1169.710 587.820 ;
        RECT 1237.930 587.760 1238.250 587.820 ;
        RECT 1169.390 587.620 1238.250 587.760 ;
        RECT 1169.390 587.560 1169.710 587.620 ;
        RECT 1237.930 587.560 1238.250 587.620 ;
        RECT 1169.390 15.540 1169.710 15.600 ;
        RECT 1138.200 15.400 1169.710 15.540 ;
        RECT 1108.670 15.200 1108.990 15.260 ;
        RECT 1138.200 15.200 1138.340 15.400 ;
        RECT 1169.390 15.340 1169.710 15.400 ;
        RECT 1108.670 15.060 1138.340 15.200 ;
        RECT 1108.670 15.000 1108.990 15.060 ;
      LAYER via ;
        RECT 1169.420 587.560 1169.680 587.820 ;
        RECT 1237.960 587.560 1238.220 587.820 ;
        RECT 1108.700 15.000 1108.960 15.260 ;
        RECT 1169.420 15.340 1169.680 15.600 ;
      LAYER met2 ;
        RECT 1239.570 600.170 1239.850 604.000 ;
        RECT 1238.020 600.030 1239.850 600.170 ;
        RECT 1238.020 587.850 1238.160 600.030 ;
        RECT 1239.570 600.000 1239.850 600.030 ;
        RECT 1169.420 587.530 1169.680 587.850 ;
        RECT 1237.960 587.530 1238.220 587.850 ;
        RECT 1169.480 15.630 1169.620 587.530 ;
        RECT 1169.420 15.310 1169.680 15.630 ;
        RECT 1108.700 14.970 1108.960 15.290 ;
        RECT 1108.760 2.400 1108.900 14.970 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1126.610 17.920 1126.930 17.980 ;
        RECT 1249.890 17.920 1250.210 17.980 ;
        RECT 1126.610 17.780 1250.210 17.920 ;
        RECT 1126.610 17.720 1126.930 17.780 ;
        RECT 1249.890 17.720 1250.210 17.780 ;
      LAYER via ;
        RECT 1126.640 17.720 1126.900 17.980 ;
        RECT 1249.920 17.720 1250.180 17.980 ;
      LAYER met2 ;
        RECT 1248.770 600.170 1249.050 604.000 ;
        RECT 1248.770 600.030 1250.120 600.170 ;
        RECT 1248.770 600.000 1249.050 600.030 ;
        RECT 1249.980 18.010 1250.120 600.030 ;
        RECT 1126.640 17.690 1126.900 18.010 ;
        RECT 1249.920 17.690 1250.180 18.010 ;
        RECT 1126.700 2.400 1126.840 17.690 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.010 589.800 1145.330 589.860 ;
        RECT 1256.330 589.800 1256.650 589.860 ;
        RECT 1145.010 589.660 1256.650 589.800 ;
        RECT 1145.010 589.600 1145.330 589.660 ;
        RECT 1256.330 589.600 1256.650 589.660 ;
        RECT 1144.090 579.600 1144.410 579.660 ;
        RECT 1145.010 579.600 1145.330 579.660 ;
        RECT 1144.090 579.460 1145.330 579.600 ;
        RECT 1144.090 579.400 1144.410 579.460 ;
        RECT 1145.010 579.400 1145.330 579.460 ;
        RECT 1144.090 531.660 1144.410 531.720 ;
        RECT 1145.010 531.660 1145.330 531.720 ;
        RECT 1144.090 531.520 1145.330 531.660 ;
        RECT 1144.090 531.460 1144.410 531.520 ;
        RECT 1145.010 531.460 1145.330 531.520 ;
        RECT 1143.630 476.240 1143.950 476.300 ;
        RECT 1145.010 476.240 1145.330 476.300 ;
        RECT 1143.630 476.100 1145.330 476.240 ;
        RECT 1143.630 476.040 1143.950 476.100 ;
        RECT 1145.010 476.040 1145.330 476.100 ;
        RECT 1143.630 435.100 1143.950 435.160 ;
        RECT 1145.010 435.100 1145.330 435.160 ;
        RECT 1143.630 434.960 1145.330 435.100 ;
        RECT 1143.630 434.900 1143.950 434.960 ;
        RECT 1145.010 434.900 1145.330 434.960 ;
        RECT 1145.010 427.620 1145.330 427.680 ;
        RECT 1146.850 427.620 1147.170 427.680 ;
        RECT 1145.010 427.480 1147.170 427.620 ;
        RECT 1145.010 427.420 1145.330 427.480 ;
        RECT 1146.850 427.420 1147.170 427.480 ;
        RECT 1145.010 331.400 1145.330 331.460 ;
        RECT 1146.850 331.400 1147.170 331.460 ;
        RECT 1145.010 331.260 1147.170 331.400 ;
        RECT 1145.010 331.200 1145.330 331.260 ;
        RECT 1146.850 331.200 1147.170 331.260 ;
        RECT 1144.090 283.120 1144.410 283.180 ;
        RECT 1145.470 283.120 1145.790 283.180 ;
        RECT 1144.090 282.980 1145.790 283.120 ;
        RECT 1144.090 282.920 1144.410 282.980 ;
        RECT 1145.470 282.920 1145.790 282.980 ;
        RECT 1144.090 241.640 1144.410 241.700 ;
        RECT 1145.010 241.640 1145.330 241.700 ;
        RECT 1144.090 241.500 1145.330 241.640 ;
        RECT 1144.090 241.440 1144.410 241.500 ;
        RECT 1145.010 241.440 1145.330 241.500 ;
        RECT 1145.010 234.500 1145.330 234.560 ;
        RECT 1145.470 234.500 1145.790 234.560 ;
        RECT 1145.010 234.360 1145.790 234.500 ;
        RECT 1145.010 234.300 1145.330 234.360 ;
        RECT 1145.470 234.300 1145.790 234.360 ;
        RECT 1145.470 186.560 1145.790 186.620 ;
        RECT 1145.930 186.560 1146.250 186.620 ;
        RECT 1145.470 186.420 1146.250 186.560 ;
        RECT 1145.470 186.360 1145.790 186.420 ;
        RECT 1145.930 186.360 1146.250 186.420 ;
        RECT 1145.930 145.420 1146.250 145.480 ;
        RECT 1145.100 145.280 1146.250 145.420 ;
        RECT 1145.100 144.800 1145.240 145.280 ;
        RECT 1145.930 145.220 1146.250 145.280 ;
        RECT 1145.010 144.540 1145.330 144.800 ;
        RECT 1145.010 62.800 1145.330 62.860 ;
        RECT 1144.180 62.660 1145.330 62.800 ;
        RECT 1144.180 62.180 1144.320 62.660 ;
        RECT 1145.010 62.600 1145.330 62.660 ;
        RECT 1144.090 61.920 1144.410 62.180 ;
        RECT 1143.630 13.840 1143.950 13.900 ;
        RECT 1144.550 13.840 1144.870 13.900 ;
        RECT 1143.630 13.700 1144.870 13.840 ;
        RECT 1143.630 13.640 1143.950 13.700 ;
        RECT 1144.550 13.640 1144.870 13.700 ;
      LAYER via ;
        RECT 1145.040 589.600 1145.300 589.860 ;
        RECT 1256.360 589.600 1256.620 589.860 ;
        RECT 1144.120 579.400 1144.380 579.660 ;
        RECT 1145.040 579.400 1145.300 579.660 ;
        RECT 1144.120 531.460 1144.380 531.720 ;
        RECT 1145.040 531.460 1145.300 531.720 ;
        RECT 1143.660 476.040 1143.920 476.300 ;
        RECT 1145.040 476.040 1145.300 476.300 ;
        RECT 1143.660 434.900 1143.920 435.160 ;
        RECT 1145.040 434.900 1145.300 435.160 ;
        RECT 1145.040 427.420 1145.300 427.680 ;
        RECT 1146.880 427.420 1147.140 427.680 ;
        RECT 1145.040 331.200 1145.300 331.460 ;
        RECT 1146.880 331.200 1147.140 331.460 ;
        RECT 1144.120 282.920 1144.380 283.180 ;
        RECT 1145.500 282.920 1145.760 283.180 ;
        RECT 1144.120 241.440 1144.380 241.700 ;
        RECT 1145.040 241.440 1145.300 241.700 ;
        RECT 1145.040 234.300 1145.300 234.560 ;
        RECT 1145.500 234.300 1145.760 234.560 ;
        RECT 1145.500 186.360 1145.760 186.620 ;
        RECT 1145.960 186.360 1146.220 186.620 ;
        RECT 1145.960 145.220 1146.220 145.480 ;
        RECT 1145.040 144.540 1145.300 144.800 ;
        RECT 1145.040 62.600 1145.300 62.860 ;
        RECT 1144.120 61.920 1144.380 62.180 ;
        RECT 1143.660 13.640 1143.920 13.900 ;
        RECT 1144.580 13.640 1144.840 13.900 ;
      LAYER met2 ;
        RECT 1257.970 600.170 1258.250 604.000 ;
        RECT 1256.420 600.030 1258.250 600.170 ;
        RECT 1256.420 589.890 1256.560 600.030 ;
        RECT 1257.970 600.000 1258.250 600.030 ;
        RECT 1145.040 589.570 1145.300 589.890 ;
        RECT 1256.360 589.570 1256.620 589.890 ;
        RECT 1145.100 579.690 1145.240 589.570 ;
        RECT 1144.120 579.370 1144.380 579.690 ;
        RECT 1145.040 579.370 1145.300 579.690 ;
        RECT 1144.180 531.750 1144.320 579.370 ;
        RECT 1144.120 531.430 1144.380 531.750 ;
        RECT 1145.040 531.430 1145.300 531.750 ;
        RECT 1145.100 476.330 1145.240 531.430 ;
        RECT 1143.660 476.010 1143.920 476.330 ;
        RECT 1145.040 476.010 1145.300 476.330 ;
        RECT 1143.720 435.190 1143.860 476.010 ;
        RECT 1143.660 434.870 1143.920 435.190 ;
        RECT 1145.040 434.870 1145.300 435.190 ;
        RECT 1145.100 427.710 1145.240 434.870 ;
        RECT 1145.040 427.390 1145.300 427.710 ;
        RECT 1146.880 427.390 1147.140 427.710 ;
        RECT 1146.940 331.490 1147.080 427.390 ;
        RECT 1145.040 331.170 1145.300 331.490 ;
        RECT 1146.880 331.170 1147.140 331.490 ;
        RECT 1145.100 330.890 1145.240 331.170 ;
        RECT 1145.100 330.750 1145.700 330.890 ;
        RECT 1145.560 283.210 1145.700 330.750 ;
        RECT 1144.120 282.890 1144.380 283.210 ;
        RECT 1145.500 282.890 1145.760 283.210 ;
        RECT 1144.180 241.730 1144.320 282.890 ;
        RECT 1144.120 241.410 1144.380 241.730 ;
        RECT 1145.040 241.410 1145.300 241.730 ;
        RECT 1145.100 234.590 1145.240 241.410 ;
        RECT 1145.040 234.270 1145.300 234.590 ;
        RECT 1145.500 234.270 1145.760 234.590 ;
        RECT 1145.560 186.650 1145.700 234.270 ;
        RECT 1145.500 186.330 1145.760 186.650 ;
        RECT 1145.960 186.330 1146.220 186.650 ;
        RECT 1146.020 145.510 1146.160 186.330 ;
        RECT 1145.960 145.190 1146.220 145.510 ;
        RECT 1145.040 144.510 1145.300 144.830 ;
        RECT 1145.100 62.890 1145.240 144.510 ;
        RECT 1145.040 62.570 1145.300 62.890 ;
        RECT 1144.120 61.890 1144.380 62.210 ;
        RECT 1144.180 48.010 1144.320 61.890 ;
        RECT 1143.720 47.870 1144.320 48.010 ;
        RECT 1143.720 13.930 1143.860 47.870 ;
        RECT 1143.660 13.610 1143.920 13.930 ;
        RECT 1144.580 13.610 1144.840 13.930 ;
        RECT 1144.640 2.400 1144.780 13.610 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1197.450 591.500 1197.770 591.560 ;
        RECT 1265.530 591.500 1265.850 591.560 ;
        RECT 1197.450 591.360 1265.850 591.500 ;
        RECT 1197.450 591.300 1197.770 591.360 ;
        RECT 1265.530 591.300 1265.850 591.360 ;
        RECT 1197.450 587.080 1197.770 587.140 ;
        RECT 1196.620 586.940 1197.770 587.080 ;
        RECT 1165.710 586.740 1166.030 586.800 ;
        RECT 1196.620 586.740 1196.760 586.940 ;
        RECT 1197.450 586.880 1197.770 586.940 ;
        RECT 1165.710 586.600 1196.760 586.740 ;
        RECT 1165.710 586.540 1166.030 586.600 ;
        RECT 1162.490 19.960 1162.810 20.020 ;
        RECT 1165.710 19.960 1166.030 20.020 ;
        RECT 1162.490 19.820 1166.030 19.960 ;
        RECT 1162.490 19.760 1162.810 19.820 ;
        RECT 1165.710 19.760 1166.030 19.820 ;
      LAYER via ;
        RECT 1197.480 591.300 1197.740 591.560 ;
        RECT 1265.560 591.300 1265.820 591.560 ;
        RECT 1165.740 586.540 1166.000 586.800 ;
        RECT 1197.480 586.880 1197.740 587.140 ;
        RECT 1162.520 19.760 1162.780 20.020 ;
        RECT 1165.740 19.760 1166.000 20.020 ;
      LAYER met2 ;
        RECT 1267.170 600.170 1267.450 604.000 ;
        RECT 1265.620 600.030 1267.450 600.170 ;
        RECT 1265.620 591.590 1265.760 600.030 ;
        RECT 1267.170 600.000 1267.450 600.030 ;
        RECT 1197.480 591.270 1197.740 591.590 ;
        RECT 1265.560 591.270 1265.820 591.590 ;
        RECT 1197.540 587.170 1197.680 591.270 ;
        RECT 1197.480 586.850 1197.740 587.170 ;
        RECT 1165.740 586.510 1166.000 586.830 ;
        RECT 1165.800 20.050 1165.940 586.510 ;
        RECT 1162.520 19.730 1162.780 20.050 ;
        RECT 1165.740 19.730 1166.000 20.050 ;
        RECT 1162.580 2.400 1162.720 19.730 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1015.290 545.260 1015.610 545.320 ;
        RECT 1018.050 545.260 1018.370 545.320 ;
        RECT 1015.290 545.120 1018.370 545.260 ;
        RECT 1015.290 545.060 1015.610 545.120 ;
        RECT 1018.050 545.060 1018.370 545.120 ;
        RECT 1013.910 400.760 1014.230 400.820 ;
        RECT 1015.290 400.760 1015.610 400.820 ;
        RECT 1013.910 400.620 1015.610 400.760 ;
        RECT 1013.910 400.560 1014.230 400.620 ;
        RECT 1015.290 400.560 1015.610 400.620 ;
        RECT 1013.910 372.880 1014.230 372.940 ;
        RECT 1014.830 372.880 1015.150 372.940 ;
        RECT 1013.910 372.740 1015.150 372.880 ;
        RECT 1013.910 372.680 1014.230 372.740 ;
        RECT 1014.830 372.680 1015.150 372.740 ;
        RECT 1013.910 331.400 1014.230 331.460 ;
        RECT 1014.830 331.400 1015.150 331.460 ;
        RECT 1013.910 331.260 1015.150 331.400 ;
        RECT 1013.910 331.200 1014.230 331.260 ;
        RECT 1014.830 331.200 1015.150 331.260 ;
        RECT 1013.910 283.120 1014.230 283.180 ;
        RECT 1014.830 283.120 1015.150 283.180 ;
        RECT 1013.910 282.980 1015.150 283.120 ;
        RECT 1013.910 282.920 1014.230 282.980 ;
        RECT 1014.830 282.920 1015.150 282.980 ;
        RECT 1014.830 193.360 1015.150 193.420 ;
        RECT 1015.290 193.360 1015.610 193.420 ;
        RECT 1014.830 193.220 1015.610 193.360 ;
        RECT 1014.830 193.160 1015.150 193.220 ;
        RECT 1015.290 193.160 1015.610 193.220 ;
        RECT 1014.830 144.740 1015.150 144.800 ;
        RECT 1016.210 144.740 1016.530 144.800 ;
        RECT 1014.830 144.600 1016.530 144.740 ;
        RECT 1014.830 144.540 1015.150 144.600 ;
        RECT 1016.210 144.540 1016.530 144.600 ;
        RECT 1015.750 96.460 1016.070 96.520 ;
        RECT 1016.210 96.460 1016.530 96.520 ;
        RECT 1015.750 96.320 1016.530 96.460 ;
        RECT 1015.750 96.260 1016.070 96.320 ;
        RECT 1016.210 96.260 1016.530 96.320 ;
        RECT 680.410 42.740 680.730 42.800 ;
        RECT 1015.750 42.740 1016.070 42.800 ;
        RECT 680.410 42.600 1016.070 42.740 ;
        RECT 680.410 42.540 680.730 42.600 ;
        RECT 1015.750 42.540 1016.070 42.600 ;
      LAYER via ;
        RECT 1015.320 545.060 1015.580 545.320 ;
        RECT 1018.080 545.060 1018.340 545.320 ;
        RECT 1013.940 400.560 1014.200 400.820 ;
        RECT 1015.320 400.560 1015.580 400.820 ;
        RECT 1013.940 372.680 1014.200 372.940 ;
        RECT 1014.860 372.680 1015.120 372.940 ;
        RECT 1013.940 331.200 1014.200 331.460 ;
        RECT 1014.860 331.200 1015.120 331.460 ;
        RECT 1013.940 282.920 1014.200 283.180 ;
        RECT 1014.860 282.920 1015.120 283.180 ;
        RECT 1014.860 193.160 1015.120 193.420 ;
        RECT 1015.320 193.160 1015.580 193.420 ;
        RECT 1014.860 144.540 1015.120 144.800 ;
        RECT 1016.240 144.540 1016.500 144.800 ;
        RECT 1015.780 96.260 1016.040 96.520 ;
        RECT 1016.240 96.260 1016.500 96.520 ;
        RECT 680.440 42.540 680.700 42.800 ;
        RECT 1015.780 42.540 1016.040 42.800 ;
      LAYER met2 ;
        RECT 1019.690 600.170 1019.970 604.000 ;
        RECT 1018.140 600.030 1019.970 600.170 ;
        RECT 1018.140 545.350 1018.280 600.030 ;
        RECT 1019.690 600.000 1019.970 600.030 ;
        RECT 1015.320 545.030 1015.580 545.350 ;
        RECT 1018.080 545.030 1018.340 545.350 ;
        RECT 1015.380 400.850 1015.520 545.030 ;
        RECT 1013.940 400.530 1014.200 400.850 ;
        RECT 1015.320 400.530 1015.580 400.850 ;
        RECT 1014.000 372.970 1014.140 400.530 ;
        RECT 1013.940 372.650 1014.200 372.970 ;
        RECT 1014.860 372.650 1015.120 372.970 ;
        RECT 1014.920 331.490 1015.060 372.650 ;
        RECT 1013.940 331.170 1014.200 331.490 ;
        RECT 1014.860 331.170 1015.120 331.490 ;
        RECT 1014.000 283.210 1014.140 331.170 ;
        RECT 1013.940 282.890 1014.200 283.210 ;
        RECT 1014.860 282.890 1015.120 283.210 ;
        RECT 1014.920 241.925 1015.060 282.890 ;
        RECT 1014.850 241.555 1015.130 241.925 ;
        RECT 1015.310 240.195 1015.590 240.565 ;
        RECT 1015.380 193.450 1015.520 240.195 ;
        RECT 1014.860 193.130 1015.120 193.450 ;
        RECT 1015.320 193.130 1015.580 193.450 ;
        RECT 1014.920 144.830 1015.060 193.130 ;
        RECT 1014.860 144.510 1015.120 144.830 ;
        RECT 1016.240 144.510 1016.500 144.830 ;
        RECT 1016.300 96.550 1016.440 144.510 ;
        RECT 1015.780 96.230 1016.040 96.550 ;
        RECT 1016.240 96.230 1016.500 96.550 ;
        RECT 1015.840 42.830 1015.980 96.230 ;
        RECT 680.440 42.510 680.700 42.830 ;
        RECT 1015.780 42.510 1016.040 42.830 ;
        RECT 680.500 2.400 680.640 42.510 ;
        RECT 680.290 -4.800 680.850 2.400 ;
      LAYER via2 ;
        RECT 1014.850 241.600 1015.130 241.880 ;
        RECT 1015.310 240.240 1015.590 240.520 ;
      LAYER met3 ;
        RECT 1014.825 241.890 1015.155 241.905 ;
        RECT 1014.825 241.575 1015.370 241.890 ;
        RECT 1015.070 240.545 1015.370 241.575 ;
        RECT 1015.070 240.230 1015.615 240.545 ;
        RECT 1015.285 240.215 1015.615 240.230 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1185.950 591.840 1186.270 591.900 ;
        RECT 1276.570 591.840 1276.890 591.900 ;
        RECT 1185.950 591.700 1276.890 591.840 ;
        RECT 1185.950 591.640 1186.270 591.700 ;
        RECT 1276.570 591.640 1276.890 591.700 ;
        RECT 1185.950 62.260 1186.270 62.520 ;
        RECT 1186.040 61.840 1186.180 62.260 ;
        RECT 1185.950 61.580 1186.270 61.840 ;
        RECT 1179.970 23.360 1180.290 23.420 ;
        RECT 1185.950 23.360 1186.270 23.420 ;
        RECT 1179.970 23.220 1186.270 23.360 ;
        RECT 1179.970 23.160 1180.290 23.220 ;
        RECT 1185.950 23.160 1186.270 23.220 ;
      LAYER via ;
        RECT 1185.980 591.640 1186.240 591.900 ;
        RECT 1276.600 591.640 1276.860 591.900 ;
        RECT 1185.980 62.260 1186.240 62.520 ;
        RECT 1185.980 61.580 1186.240 61.840 ;
        RECT 1180.000 23.160 1180.260 23.420 ;
        RECT 1185.980 23.160 1186.240 23.420 ;
      LAYER met2 ;
        RECT 1276.370 600.000 1276.650 604.000 ;
        RECT 1276.430 598.810 1276.570 600.000 ;
        RECT 1276.430 598.670 1276.800 598.810 ;
        RECT 1276.660 591.930 1276.800 598.670 ;
        RECT 1185.980 591.610 1186.240 591.930 ;
        RECT 1276.600 591.610 1276.860 591.930 ;
        RECT 1186.040 62.550 1186.180 591.610 ;
        RECT 1185.980 62.230 1186.240 62.550 ;
        RECT 1185.980 61.550 1186.240 61.870 ;
        RECT 1186.040 23.450 1186.180 61.550 ;
        RECT 1180.000 23.130 1180.260 23.450 ;
        RECT 1185.980 23.130 1186.240 23.450 ;
        RECT 1180.060 2.400 1180.200 23.130 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 592.860 1200.530 592.920 ;
        RECT 1283.470 592.860 1283.790 592.920 ;
        RECT 1200.210 592.720 1283.790 592.860 ;
        RECT 1200.210 592.660 1200.530 592.720 ;
        RECT 1283.470 592.660 1283.790 592.720 ;
        RECT 1197.910 20.640 1198.230 20.700 ;
        RECT 1200.210 20.640 1200.530 20.700 ;
        RECT 1197.910 20.500 1200.530 20.640 ;
        RECT 1197.910 20.440 1198.230 20.500 ;
        RECT 1200.210 20.440 1200.530 20.500 ;
      LAYER via ;
        RECT 1200.240 592.660 1200.500 592.920 ;
        RECT 1283.500 592.660 1283.760 592.920 ;
        RECT 1197.940 20.440 1198.200 20.700 ;
        RECT 1200.240 20.440 1200.500 20.700 ;
      LAYER met2 ;
        RECT 1285.110 600.170 1285.390 604.000 ;
        RECT 1283.560 600.030 1285.390 600.170 ;
        RECT 1283.560 592.950 1283.700 600.030 ;
        RECT 1285.110 600.000 1285.390 600.030 ;
        RECT 1200.240 592.630 1200.500 592.950 ;
        RECT 1283.500 592.630 1283.760 592.950 ;
        RECT 1200.300 20.730 1200.440 592.630 ;
        RECT 1197.940 20.410 1198.200 20.730 ;
        RECT 1200.240 20.410 1200.500 20.730 ;
        RECT 1198.000 2.400 1198.140 20.410 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 587.420 1221.230 587.480 ;
        RECT 1292.670 587.420 1292.990 587.480 ;
        RECT 1220.910 587.280 1292.990 587.420 ;
        RECT 1220.910 587.220 1221.230 587.280 ;
        RECT 1292.670 587.220 1292.990 587.280 ;
        RECT 1215.850 16.560 1216.170 16.620 ;
        RECT 1220.910 16.560 1221.230 16.620 ;
        RECT 1215.850 16.420 1221.230 16.560 ;
        RECT 1215.850 16.360 1216.170 16.420 ;
        RECT 1220.910 16.360 1221.230 16.420 ;
      LAYER via ;
        RECT 1220.940 587.220 1221.200 587.480 ;
        RECT 1292.700 587.220 1292.960 587.480 ;
        RECT 1215.880 16.360 1216.140 16.620 ;
        RECT 1220.940 16.360 1221.200 16.620 ;
      LAYER met2 ;
        RECT 1294.310 600.170 1294.590 604.000 ;
        RECT 1292.760 600.030 1294.590 600.170 ;
        RECT 1292.760 587.510 1292.900 600.030 ;
        RECT 1294.310 600.000 1294.590 600.030 ;
        RECT 1220.940 587.190 1221.200 587.510 ;
        RECT 1292.700 587.190 1292.960 587.510 ;
        RECT 1221.000 16.650 1221.140 587.190 ;
        RECT 1215.880 16.330 1216.140 16.650 ;
        RECT 1220.940 16.330 1221.200 16.650 ;
        RECT 1215.940 2.400 1216.080 16.330 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.710 587.080 1235.030 587.140 ;
        RECT 1301.870 587.080 1302.190 587.140 ;
        RECT 1234.710 586.940 1302.190 587.080 ;
        RECT 1234.710 586.880 1235.030 586.940 ;
        RECT 1301.870 586.880 1302.190 586.940 ;
      LAYER via ;
        RECT 1234.740 586.880 1235.000 587.140 ;
        RECT 1301.900 586.880 1302.160 587.140 ;
      LAYER met2 ;
        RECT 1303.510 600.170 1303.790 604.000 ;
        RECT 1301.960 600.030 1303.790 600.170 ;
        RECT 1301.960 587.170 1302.100 600.030 ;
        RECT 1303.510 600.000 1303.790 600.030 ;
        RECT 1234.740 586.850 1235.000 587.170 ;
        RECT 1301.900 586.850 1302.160 587.170 ;
        RECT 1234.800 3.130 1234.940 586.850 ;
        RECT 1234.340 2.990 1234.940 3.130 ;
        RECT 1234.340 2.960 1234.480 2.990 ;
        RECT 1233.880 2.820 1234.480 2.960 ;
        RECT 1233.880 2.400 1234.020 2.820 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 590.140 1255.730 590.200 ;
        RECT 1311.070 590.140 1311.390 590.200 ;
        RECT 1255.410 590.000 1311.390 590.140 ;
        RECT 1255.410 589.940 1255.730 590.000 ;
        RECT 1311.070 589.940 1311.390 590.000 ;
        RECT 1251.730 16.900 1252.050 16.960 ;
        RECT 1255.410 16.900 1255.730 16.960 ;
        RECT 1251.730 16.760 1255.730 16.900 ;
        RECT 1251.730 16.700 1252.050 16.760 ;
        RECT 1255.410 16.700 1255.730 16.760 ;
      LAYER via ;
        RECT 1255.440 589.940 1255.700 590.200 ;
        RECT 1311.100 589.940 1311.360 590.200 ;
        RECT 1251.760 16.700 1252.020 16.960 ;
        RECT 1255.440 16.700 1255.700 16.960 ;
      LAYER met2 ;
        RECT 1312.710 600.170 1312.990 604.000 ;
        RECT 1311.160 600.030 1312.990 600.170 ;
        RECT 1311.160 590.230 1311.300 600.030 ;
        RECT 1312.710 600.000 1312.990 600.030 ;
        RECT 1255.440 589.910 1255.700 590.230 ;
        RECT 1311.100 589.910 1311.360 590.230 ;
        RECT 1255.500 16.990 1255.640 589.910 ;
        RECT 1251.760 16.670 1252.020 16.990 ;
        RECT 1255.440 16.670 1255.700 16.990 ;
        RECT 1251.820 2.400 1251.960 16.670 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1268.750 589.800 1269.070 589.860 ;
        RECT 1320.270 589.800 1320.590 589.860 ;
        RECT 1268.750 589.660 1320.590 589.800 ;
        RECT 1268.750 589.600 1269.070 589.660 ;
        RECT 1320.270 589.600 1320.590 589.660 ;
      LAYER via ;
        RECT 1268.780 589.600 1269.040 589.860 ;
        RECT 1320.300 589.600 1320.560 589.860 ;
      LAYER met2 ;
        RECT 1321.910 600.170 1322.190 604.000 ;
        RECT 1320.360 600.030 1322.190 600.170 ;
        RECT 1320.360 589.890 1320.500 600.030 ;
        RECT 1321.910 600.000 1322.190 600.030 ;
        RECT 1268.780 589.570 1269.040 589.890 ;
        RECT 1320.300 589.570 1320.560 589.890 ;
        RECT 1268.840 16.050 1268.980 589.570 ;
        RECT 1268.840 15.910 1269.440 16.050 ;
        RECT 1269.300 2.400 1269.440 15.910 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 592.520 1290.230 592.580 ;
        RECT 1329.470 592.520 1329.790 592.580 ;
        RECT 1289.910 592.380 1329.790 592.520 ;
        RECT 1289.910 592.320 1290.230 592.380 ;
        RECT 1329.470 592.320 1329.790 592.380 ;
        RECT 1287.150 17.580 1287.470 17.640 ;
        RECT 1289.910 17.580 1290.230 17.640 ;
        RECT 1287.150 17.440 1290.230 17.580 ;
        RECT 1287.150 17.380 1287.470 17.440 ;
        RECT 1289.910 17.380 1290.230 17.440 ;
      LAYER via ;
        RECT 1289.940 592.320 1290.200 592.580 ;
        RECT 1329.500 592.320 1329.760 592.580 ;
        RECT 1287.180 17.380 1287.440 17.640 ;
        RECT 1289.940 17.380 1290.200 17.640 ;
      LAYER met2 ;
        RECT 1331.110 600.170 1331.390 604.000 ;
        RECT 1329.560 600.030 1331.390 600.170 ;
        RECT 1329.560 592.610 1329.700 600.030 ;
        RECT 1331.110 600.000 1331.390 600.030 ;
        RECT 1289.940 592.290 1290.200 592.610 ;
        RECT 1329.500 592.290 1329.760 592.610 ;
        RECT 1290.000 17.670 1290.140 592.290 ;
        RECT 1287.180 17.350 1287.440 17.670 ;
        RECT 1289.940 17.350 1290.200 17.670 ;
        RECT 1287.240 2.400 1287.380 17.350 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 590.480 1310.930 590.540 ;
        RECT 1339.130 590.480 1339.450 590.540 ;
        RECT 1310.610 590.340 1339.450 590.480 ;
        RECT 1310.610 590.280 1310.930 590.340 ;
        RECT 1339.130 590.280 1339.450 590.340 ;
        RECT 1305.090 16.220 1305.410 16.280 ;
        RECT 1310.610 16.220 1310.930 16.280 ;
        RECT 1305.090 16.080 1310.930 16.220 ;
        RECT 1305.090 16.020 1305.410 16.080 ;
        RECT 1310.610 16.020 1310.930 16.080 ;
      LAYER via ;
        RECT 1310.640 590.280 1310.900 590.540 ;
        RECT 1339.160 590.280 1339.420 590.540 ;
        RECT 1305.120 16.020 1305.380 16.280 ;
        RECT 1310.640 16.020 1310.900 16.280 ;
      LAYER met2 ;
        RECT 1340.310 600.170 1340.590 604.000 ;
        RECT 1339.220 600.030 1340.590 600.170 ;
        RECT 1339.220 590.570 1339.360 600.030 ;
        RECT 1340.310 600.000 1340.590 600.030 ;
        RECT 1310.640 590.250 1310.900 590.570 ;
        RECT 1339.160 590.250 1339.420 590.570 ;
        RECT 1310.700 16.310 1310.840 590.250 ;
        RECT 1305.120 15.990 1305.380 16.310 ;
        RECT 1310.640 15.990 1310.900 16.310 ;
        RECT 1305.180 2.400 1305.320 15.990 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.410 589.120 1324.730 589.180 ;
        RECT 1347.870 589.120 1348.190 589.180 ;
        RECT 1324.410 588.980 1348.190 589.120 ;
        RECT 1324.410 588.920 1324.730 588.980 ;
        RECT 1347.870 588.920 1348.190 588.980 ;
      LAYER via ;
        RECT 1324.440 588.920 1324.700 589.180 ;
        RECT 1347.900 588.920 1348.160 589.180 ;
      LAYER met2 ;
        RECT 1349.510 600.170 1349.790 604.000 ;
        RECT 1347.960 600.030 1349.790 600.170 ;
        RECT 1347.960 589.210 1348.100 600.030 ;
        RECT 1349.510 600.000 1349.790 600.030 ;
        RECT 1324.440 588.890 1324.700 589.210 ;
        RECT 1347.900 588.890 1348.160 589.210 ;
        RECT 1324.500 17.410 1324.640 588.890 ;
        RECT 1323.120 17.270 1324.640 17.410 ;
        RECT 1323.120 2.400 1323.260 17.270 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1345.110 586.740 1345.430 586.800 ;
        RECT 1357.070 586.740 1357.390 586.800 ;
        RECT 1345.110 586.600 1357.390 586.740 ;
        RECT 1345.110 586.540 1345.430 586.600 ;
        RECT 1357.070 586.540 1357.390 586.600 ;
        RECT 1340.510 19.960 1340.830 20.020 ;
        RECT 1345.110 19.960 1345.430 20.020 ;
        RECT 1340.510 19.820 1345.430 19.960 ;
        RECT 1340.510 19.760 1340.830 19.820 ;
        RECT 1345.110 19.760 1345.430 19.820 ;
      LAYER via ;
        RECT 1345.140 586.540 1345.400 586.800 ;
        RECT 1357.100 586.540 1357.360 586.800 ;
        RECT 1340.540 19.760 1340.800 20.020 ;
        RECT 1345.140 19.760 1345.400 20.020 ;
      LAYER met2 ;
        RECT 1358.710 600.170 1358.990 604.000 ;
        RECT 1357.160 600.030 1358.990 600.170 ;
        RECT 1357.160 586.830 1357.300 600.030 ;
        RECT 1358.710 600.000 1358.990 600.030 ;
        RECT 1345.140 586.510 1345.400 586.830 ;
        RECT 1357.100 586.510 1357.360 586.830 ;
        RECT 1345.200 20.050 1345.340 586.510 ;
        RECT 1340.540 19.730 1340.800 20.050 ;
        RECT 1345.140 19.730 1345.400 20.050 ;
        RECT 1340.600 2.400 1340.740 19.730 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1029.090 579.940 1029.410 580.000 ;
        RECT 1029.550 579.940 1029.870 580.000 ;
        RECT 1029.090 579.800 1029.870 579.940 ;
        RECT 1029.090 579.740 1029.410 579.800 ;
        RECT 1029.550 579.740 1029.870 579.800 ;
        RECT 1028.630 448.840 1028.950 449.100 ;
        RECT 1028.720 448.420 1028.860 448.840 ;
        RECT 1028.630 448.160 1028.950 448.420 ;
        RECT 1028.630 283.460 1028.950 283.520 ;
        RECT 1028.630 283.320 1029.320 283.460 ;
        RECT 1028.630 283.260 1028.950 283.320 ;
        RECT 1029.180 283.180 1029.320 283.320 ;
        RECT 1029.090 282.920 1029.410 283.180 ;
        RECT 1028.630 241.300 1028.950 241.360 ;
        RECT 1029.090 241.300 1029.410 241.360 ;
        RECT 1028.630 241.160 1029.410 241.300 ;
        RECT 1028.630 241.100 1028.950 241.160 ;
        RECT 1029.090 241.100 1029.410 241.160 ;
        RECT 1027.250 186.220 1027.570 186.280 ;
        RECT 1028.630 186.220 1028.950 186.280 ;
        RECT 1027.250 186.080 1028.950 186.220 ;
        RECT 1027.250 186.020 1027.570 186.080 ;
        RECT 1028.630 186.020 1028.950 186.080 ;
        RECT 1027.250 138.280 1027.570 138.340 ;
        RECT 1028.630 138.280 1028.950 138.340 ;
        RECT 1027.250 138.140 1028.950 138.280 ;
        RECT 1027.250 138.080 1027.570 138.140 ;
        RECT 1028.630 138.080 1028.950 138.140 ;
        RECT 1020.350 48.180 1020.670 48.240 ;
        RECT 1029.090 48.180 1029.410 48.240 ;
        RECT 1020.350 48.040 1029.410 48.180 ;
        RECT 1020.350 47.980 1020.670 48.040 ;
        RECT 1029.090 47.980 1029.410 48.040 ;
        RECT 698.350 44.780 698.670 44.840 ;
        RECT 1020.350 44.780 1020.670 44.840 ;
        RECT 698.350 44.640 1020.670 44.780 ;
        RECT 698.350 44.580 698.670 44.640 ;
        RECT 1020.350 44.580 1020.670 44.640 ;
      LAYER via ;
        RECT 1029.120 579.740 1029.380 580.000 ;
        RECT 1029.580 579.740 1029.840 580.000 ;
        RECT 1028.660 448.840 1028.920 449.100 ;
        RECT 1028.660 448.160 1028.920 448.420 ;
        RECT 1028.660 283.260 1028.920 283.520 ;
        RECT 1029.120 282.920 1029.380 283.180 ;
        RECT 1028.660 241.100 1028.920 241.360 ;
        RECT 1029.120 241.100 1029.380 241.360 ;
        RECT 1027.280 186.020 1027.540 186.280 ;
        RECT 1028.660 186.020 1028.920 186.280 ;
        RECT 1027.280 138.080 1027.540 138.340 ;
        RECT 1028.660 138.080 1028.920 138.340 ;
        RECT 1020.380 47.980 1020.640 48.240 ;
        RECT 1029.120 47.980 1029.380 48.240 ;
        RECT 698.380 44.580 698.640 44.840 ;
        RECT 1020.380 44.580 1020.640 44.840 ;
      LAYER met2 ;
        RECT 1028.890 600.170 1029.170 604.000 ;
        RECT 1028.890 600.030 1029.780 600.170 ;
        RECT 1028.890 600.000 1029.170 600.030 ;
        RECT 1029.640 580.030 1029.780 600.030 ;
        RECT 1029.120 579.710 1029.380 580.030 ;
        RECT 1029.580 579.710 1029.840 580.030 ;
        RECT 1029.180 497.490 1029.320 579.710 ;
        RECT 1028.720 497.350 1029.320 497.490 ;
        RECT 1028.720 449.130 1028.860 497.350 ;
        RECT 1028.660 448.810 1028.920 449.130 ;
        RECT 1028.660 448.130 1028.920 448.450 ;
        RECT 1028.720 283.550 1028.860 448.130 ;
        RECT 1028.660 283.230 1028.920 283.550 ;
        RECT 1029.120 282.890 1029.380 283.210 ;
        RECT 1029.180 241.390 1029.320 282.890 ;
        RECT 1028.660 241.070 1028.920 241.390 ;
        RECT 1029.120 241.070 1029.380 241.390 ;
        RECT 1028.720 186.310 1028.860 241.070 ;
        RECT 1027.280 185.990 1027.540 186.310 ;
        RECT 1028.660 185.990 1028.920 186.310 ;
        RECT 1027.340 138.370 1027.480 185.990 ;
        RECT 1027.280 138.050 1027.540 138.370 ;
        RECT 1028.660 138.050 1028.920 138.370 ;
        RECT 1028.720 137.885 1028.860 138.050 ;
        RECT 1028.650 137.515 1028.930 137.885 ;
        RECT 1029.110 136.835 1029.390 137.205 ;
        RECT 1029.180 48.270 1029.320 136.835 ;
        RECT 1020.380 47.950 1020.640 48.270 ;
        RECT 1029.120 47.950 1029.380 48.270 ;
        RECT 1020.440 44.870 1020.580 47.950 ;
        RECT 698.380 44.550 698.640 44.870 ;
        RECT 1020.380 44.550 1020.640 44.870 ;
        RECT 698.440 2.400 698.580 44.550 ;
        RECT 698.230 -4.800 698.790 2.400 ;
      LAYER via2 ;
        RECT 1028.650 137.560 1028.930 137.840 ;
        RECT 1029.110 136.880 1029.390 137.160 ;
      LAYER met3 ;
        RECT 1028.625 137.850 1028.955 137.865 ;
        RECT 1027.950 137.550 1028.955 137.850 ;
        RECT 1027.950 137.170 1028.250 137.550 ;
        RECT 1028.625 137.535 1028.955 137.550 ;
        RECT 1029.085 137.170 1029.415 137.185 ;
        RECT 1027.950 136.870 1029.415 137.170 ;
        RECT 1029.085 136.855 1029.415 136.870 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1358.910 587.080 1359.230 587.140 ;
        RECT 1366.270 587.080 1366.590 587.140 ;
        RECT 1358.910 586.940 1366.590 587.080 ;
        RECT 1358.910 586.880 1359.230 586.940 ;
        RECT 1366.270 586.880 1366.590 586.940 ;
      LAYER via ;
        RECT 1358.940 586.880 1359.200 587.140 ;
        RECT 1366.300 586.880 1366.560 587.140 ;
      LAYER met2 ;
        RECT 1367.910 600.170 1368.190 604.000 ;
        RECT 1366.360 600.030 1368.190 600.170 ;
        RECT 1366.360 587.170 1366.500 600.030 ;
        RECT 1367.910 600.000 1368.190 600.030 ;
        RECT 1358.940 586.850 1359.200 587.170 ;
        RECT 1366.300 586.850 1366.560 587.170 ;
        RECT 1359.000 24.210 1359.140 586.850 ;
        RECT 1358.540 24.070 1359.140 24.210 ;
        RECT 1358.540 2.400 1358.680 24.070 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1373.170 569.400 1373.490 569.460 ;
        RECT 1375.470 569.400 1375.790 569.460 ;
        RECT 1373.170 569.260 1375.790 569.400 ;
        RECT 1373.170 569.200 1373.490 569.260 ;
        RECT 1375.470 569.200 1375.790 569.260 ;
        RECT 1373.170 20.300 1373.490 20.360 ;
        RECT 1376.390 20.300 1376.710 20.360 ;
        RECT 1373.170 20.160 1376.710 20.300 ;
        RECT 1373.170 20.100 1373.490 20.160 ;
        RECT 1376.390 20.100 1376.710 20.160 ;
      LAYER via ;
        RECT 1373.200 569.200 1373.460 569.460 ;
        RECT 1375.500 569.200 1375.760 569.460 ;
        RECT 1373.200 20.100 1373.460 20.360 ;
        RECT 1376.420 20.100 1376.680 20.360 ;
      LAYER met2 ;
        RECT 1377.110 600.170 1377.390 604.000 ;
        RECT 1375.560 600.030 1377.390 600.170 ;
        RECT 1375.560 569.490 1375.700 600.030 ;
        RECT 1377.110 600.000 1377.390 600.030 ;
        RECT 1373.200 569.170 1373.460 569.490 ;
        RECT 1375.500 569.170 1375.760 569.490 ;
        RECT 1373.260 20.390 1373.400 569.170 ;
        RECT 1373.200 20.070 1373.460 20.390 ;
        RECT 1376.420 20.070 1376.680 20.390 ;
        RECT 1376.480 2.400 1376.620 20.070 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.050 587.420 1386.370 587.480 ;
        RECT 1390.190 587.420 1390.510 587.480 ;
        RECT 1386.050 587.280 1390.510 587.420 ;
        RECT 1386.050 587.220 1386.370 587.280 ;
        RECT 1390.190 587.220 1390.510 587.280 ;
        RECT 1390.190 20.640 1390.510 20.700 ;
        RECT 1394.330 20.640 1394.650 20.700 ;
        RECT 1390.190 20.500 1394.650 20.640 ;
        RECT 1390.190 20.440 1390.510 20.500 ;
        RECT 1394.330 20.440 1394.650 20.500 ;
      LAYER via ;
        RECT 1386.080 587.220 1386.340 587.480 ;
        RECT 1390.220 587.220 1390.480 587.480 ;
        RECT 1390.220 20.440 1390.480 20.700 ;
        RECT 1394.360 20.440 1394.620 20.700 ;
      LAYER met2 ;
        RECT 1386.310 600.000 1386.590 604.000 ;
        RECT 1386.370 598.810 1386.510 600.000 ;
        RECT 1386.140 598.670 1386.510 598.810 ;
        RECT 1386.140 587.510 1386.280 598.670 ;
        RECT 1386.080 587.190 1386.340 587.510 ;
        RECT 1390.220 587.190 1390.480 587.510 ;
        RECT 1390.280 20.730 1390.420 587.190 ;
        RECT 1390.220 20.410 1390.480 20.730 ;
        RECT 1394.360 20.410 1394.620 20.730 ;
        RECT 1394.420 2.400 1394.560 20.410 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1397.090 586.740 1397.410 586.800 ;
        RECT 1400.310 586.740 1400.630 586.800 ;
        RECT 1397.090 586.600 1400.630 586.740 ;
        RECT 1397.090 586.540 1397.410 586.600 ;
        RECT 1400.310 586.540 1400.630 586.600 ;
        RECT 1400.310 20.780 1400.630 21.040 ;
        RECT 1400.400 20.640 1400.540 20.780 ;
        RECT 1412.270 20.640 1412.590 20.700 ;
        RECT 1400.400 20.500 1412.590 20.640 ;
        RECT 1412.270 20.440 1412.590 20.500 ;
      LAYER via ;
        RECT 1397.120 586.540 1397.380 586.800 ;
        RECT 1400.340 586.540 1400.600 586.800 ;
        RECT 1400.340 20.780 1400.600 21.040 ;
        RECT 1412.300 20.440 1412.560 20.700 ;
      LAYER met2 ;
        RECT 1395.510 600.170 1395.790 604.000 ;
        RECT 1395.510 600.030 1397.320 600.170 ;
        RECT 1395.510 600.000 1395.790 600.030 ;
        RECT 1397.180 586.830 1397.320 600.030 ;
        RECT 1397.120 586.510 1397.380 586.830 ;
        RECT 1400.340 586.510 1400.600 586.830 ;
        RECT 1400.400 21.070 1400.540 586.510 ;
        RECT 1400.340 20.750 1400.600 21.070 ;
        RECT 1412.300 20.410 1412.560 20.730 ;
        RECT 1412.360 2.400 1412.500 20.410 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1407.210 17.240 1407.530 17.300 ;
        RECT 1429.750 17.240 1430.070 17.300 ;
        RECT 1407.210 17.100 1430.070 17.240 ;
        RECT 1407.210 17.040 1407.530 17.100 ;
        RECT 1429.750 17.040 1430.070 17.100 ;
      LAYER via ;
        RECT 1407.240 17.040 1407.500 17.300 ;
        RECT 1429.780 17.040 1430.040 17.300 ;
      LAYER met2 ;
        RECT 1404.250 600.170 1404.530 604.000 ;
        RECT 1404.250 600.030 1406.980 600.170 ;
        RECT 1404.250 600.000 1404.530 600.030 ;
        RECT 1406.840 587.930 1406.980 600.030 ;
        RECT 1406.840 587.790 1407.440 587.930 ;
        RECT 1407.300 17.330 1407.440 587.790 ;
        RECT 1407.240 17.010 1407.500 17.330 ;
        RECT 1429.780 17.010 1430.040 17.330 ;
        RECT 1429.840 2.400 1429.980 17.010 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1414.110 18.260 1414.430 18.320 ;
        RECT 1447.690 18.260 1448.010 18.320 ;
        RECT 1414.110 18.120 1448.010 18.260 ;
        RECT 1414.110 18.060 1414.430 18.120 ;
        RECT 1447.690 18.060 1448.010 18.120 ;
      LAYER via ;
        RECT 1414.140 18.060 1414.400 18.320 ;
        RECT 1447.720 18.060 1447.980 18.320 ;
      LAYER met2 ;
        RECT 1413.450 600.170 1413.730 604.000 ;
        RECT 1413.450 600.030 1414.340 600.170 ;
        RECT 1413.450 600.000 1413.730 600.030 ;
        RECT 1414.200 18.350 1414.340 600.030 ;
        RECT 1414.140 18.030 1414.400 18.350 ;
        RECT 1447.720 18.030 1447.980 18.350 ;
        RECT 1447.780 2.400 1447.920 18.030 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1424.230 586.740 1424.550 586.800 ;
        RECT 1427.910 586.740 1428.230 586.800 ;
        RECT 1424.230 586.600 1428.230 586.740 ;
        RECT 1424.230 586.540 1424.550 586.600 ;
        RECT 1427.910 586.540 1428.230 586.600 ;
        RECT 1427.910 17.920 1428.230 17.980 ;
        RECT 1465.630 17.920 1465.950 17.980 ;
        RECT 1427.910 17.780 1465.950 17.920 ;
        RECT 1427.910 17.720 1428.230 17.780 ;
        RECT 1465.630 17.720 1465.950 17.780 ;
      LAYER via ;
        RECT 1424.260 586.540 1424.520 586.800 ;
        RECT 1427.940 586.540 1428.200 586.800 ;
        RECT 1427.940 17.720 1428.200 17.980 ;
        RECT 1465.660 17.720 1465.920 17.980 ;
      LAYER met2 ;
        RECT 1422.650 600.170 1422.930 604.000 ;
        RECT 1422.650 600.030 1424.460 600.170 ;
        RECT 1422.650 600.000 1422.930 600.030 ;
        RECT 1424.320 586.830 1424.460 600.030 ;
        RECT 1424.260 586.510 1424.520 586.830 ;
        RECT 1427.940 586.510 1428.200 586.830 ;
        RECT 1428.000 18.010 1428.140 586.510 ;
        RECT 1427.940 17.690 1428.200 18.010 ;
        RECT 1465.660 17.690 1465.920 18.010 ;
        RECT 1465.720 2.400 1465.860 17.690 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.350 19.960 1434.670 20.020 ;
        RECT 1483.570 19.960 1483.890 20.020 ;
        RECT 1434.350 19.820 1483.890 19.960 ;
        RECT 1434.350 19.760 1434.670 19.820 ;
        RECT 1483.570 19.760 1483.890 19.820 ;
      LAYER via ;
        RECT 1434.380 19.760 1434.640 20.020 ;
        RECT 1483.600 19.760 1483.860 20.020 ;
      LAYER met2 ;
        RECT 1431.850 600.170 1432.130 604.000 ;
        RECT 1431.850 600.030 1434.580 600.170 ;
        RECT 1431.850 600.000 1432.130 600.030 ;
        RECT 1434.440 20.050 1434.580 600.030 ;
        RECT 1434.380 19.730 1434.640 20.050 ;
        RECT 1483.600 19.730 1483.860 20.050 ;
        RECT 1483.660 2.400 1483.800 19.730 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1441.710 19.620 1442.030 19.680 ;
        RECT 1501.510 19.620 1501.830 19.680 ;
        RECT 1441.710 19.480 1501.830 19.620 ;
        RECT 1441.710 19.420 1442.030 19.480 ;
        RECT 1501.510 19.420 1501.830 19.480 ;
      LAYER via ;
        RECT 1441.740 19.420 1442.000 19.680 ;
        RECT 1501.540 19.420 1501.800 19.680 ;
      LAYER met2 ;
        RECT 1441.050 600.170 1441.330 604.000 ;
        RECT 1441.050 600.030 1441.940 600.170 ;
        RECT 1441.050 600.000 1441.330 600.030 ;
        RECT 1441.800 19.710 1441.940 600.030 ;
        RECT 1441.740 19.390 1442.000 19.710 ;
        RECT 1501.540 19.390 1501.800 19.710 ;
        RECT 1501.600 2.400 1501.740 19.390 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1451.830 586.740 1452.150 586.800 ;
        RECT 1455.510 586.740 1455.830 586.800 ;
        RECT 1451.830 586.600 1455.830 586.740 ;
        RECT 1451.830 586.540 1452.150 586.600 ;
        RECT 1455.510 586.540 1455.830 586.600 ;
        RECT 1455.510 18.600 1455.830 18.660 ;
        RECT 1518.990 18.600 1519.310 18.660 ;
        RECT 1455.510 18.460 1519.310 18.600 ;
        RECT 1455.510 18.400 1455.830 18.460 ;
        RECT 1518.990 18.400 1519.310 18.460 ;
      LAYER via ;
        RECT 1451.860 586.540 1452.120 586.800 ;
        RECT 1455.540 586.540 1455.800 586.800 ;
        RECT 1455.540 18.400 1455.800 18.660 ;
        RECT 1519.020 18.400 1519.280 18.660 ;
      LAYER met2 ;
        RECT 1450.250 600.170 1450.530 604.000 ;
        RECT 1450.250 600.030 1452.060 600.170 ;
        RECT 1450.250 600.000 1450.530 600.030 ;
        RECT 1451.920 586.830 1452.060 600.030 ;
        RECT 1451.860 586.510 1452.120 586.830 ;
        RECT 1455.540 586.510 1455.800 586.830 ;
        RECT 1455.600 18.690 1455.740 586.510 ;
        RECT 1455.540 18.370 1455.800 18.690 ;
        RECT 1519.020 18.370 1519.280 18.690 ;
        RECT 1519.080 2.400 1519.220 18.370 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 716.290 45.120 716.610 45.180 ;
        RECT 1035.990 45.120 1036.310 45.180 ;
        RECT 716.290 44.980 1036.310 45.120 ;
        RECT 716.290 44.920 716.610 44.980 ;
        RECT 1035.990 44.920 1036.310 44.980 ;
      LAYER via ;
        RECT 716.320 44.920 716.580 45.180 ;
        RECT 1036.020 44.920 1036.280 45.180 ;
      LAYER met2 ;
        RECT 1037.630 600.170 1037.910 604.000 ;
        RECT 1036.080 600.030 1037.910 600.170 ;
        RECT 1036.080 45.210 1036.220 600.030 ;
        RECT 1037.630 600.000 1037.910 600.030 ;
        RECT 716.320 44.890 716.580 45.210 ;
        RECT 1036.020 44.890 1036.280 45.210 ;
        RECT 716.380 2.400 716.520 44.890 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1461.950 18.260 1462.270 18.320 ;
        RECT 1536.930 18.260 1537.250 18.320 ;
        RECT 1461.950 18.120 1537.250 18.260 ;
        RECT 1461.950 18.060 1462.270 18.120 ;
        RECT 1536.930 18.060 1537.250 18.120 ;
      LAYER via ;
        RECT 1461.980 18.060 1462.240 18.320 ;
        RECT 1536.960 18.060 1537.220 18.320 ;
      LAYER met2 ;
        RECT 1459.450 600.170 1459.730 604.000 ;
        RECT 1459.450 600.030 1462.180 600.170 ;
        RECT 1459.450 600.000 1459.730 600.030 ;
        RECT 1462.040 18.350 1462.180 600.030 ;
        RECT 1461.980 18.030 1462.240 18.350 ;
        RECT 1536.960 18.030 1537.220 18.350 ;
        RECT 1537.020 2.400 1537.160 18.030 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.310 17.580 1469.630 17.640 ;
        RECT 1554.870 17.580 1555.190 17.640 ;
        RECT 1469.310 17.440 1555.190 17.580 ;
        RECT 1469.310 17.380 1469.630 17.440 ;
        RECT 1554.870 17.380 1555.190 17.440 ;
      LAYER via ;
        RECT 1469.340 17.380 1469.600 17.640 ;
        RECT 1554.900 17.380 1555.160 17.640 ;
      LAYER met2 ;
        RECT 1468.650 600.170 1468.930 604.000 ;
        RECT 1468.650 600.030 1469.540 600.170 ;
        RECT 1468.650 600.000 1468.930 600.030 ;
        RECT 1469.400 17.670 1469.540 600.030 ;
        RECT 1469.340 17.350 1469.600 17.670 ;
        RECT 1554.900 17.350 1555.160 17.670 ;
        RECT 1554.960 2.400 1555.100 17.350 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1479.430 586.740 1479.750 586.800 ;
        RECT 1483.110 586.740 1483.430 586.800 ;
        RECT 1479.430 586.600 1483.430 586.740 ;
        RECT 1479.430 586.540 1479.750 586.600 ;
        RECT 1483.110 586.540 1483.430 586.600 ;
        RECT 1483.110 20.300 1483.430 20.360 ;
        RECT 1572.810 20.300 1573.130 20.360 ;
        RECT 1483.110 20.160 1573.130 20.300 ;
        RECT 1483.110 20.100 1483.430 20.160 ;
        RECT 1572.810 20.100 1573.130 20.160 ;
      LAYER via ;
        RECT 1479.460 586.540 1479.720 586.800 ;
        RECT 1483.140 586.540 1483.400 586.800 ;
        RECT 1483.140 20.100 1483.400 20.360 ;
        RECT 1572.840 20.100 1573.100 20.360 ;
      LAYER met2 ;
        RECT 1477.850 600.170 1478.130 604.000 ;
        RECT 1477.850 600.030 1479.660 600.170 ;
        RECT 1477.850 600.000 1478.130 600.030 ;
        RECT 1479.520 586.830 1479.660 600.030 ;
        RECT 1479.460 586.510 1479.720 586.830 ;
        RECT 1483.140 586.510 1483.400 586.830 ;
        RECT 1483.200 20.390 1483.340 586.510 ;
        RECT 1483.140 20.070 1483.400 20.390 ;
        RECT 1572.840 20.070 1573.100 20.390 ;
        RECT 1572.900 2.400 1573.040 20.070 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1488.170 559.200 1488.490 559.260 ;
        RECT 1489.550 559.200 1489.870 559.260 ;
        RECT 1488.170 559.060 1489.870 559.200 ;
        RECT 1488.170 559.000 1488.490 559.060 ;
        RECT 1489.550 559.000 1489.870 559.060 ;
        RECT 1489.550 510.580 1489.870 510.640 ;
        RECT 1490.470 510.580 1490.790 510.640 ;
        RECT 1489.550 510.440 1490.790 510.580 ;
        RECT 1489.550 510.380 1489.870 510.440 ;
        RECT 1490.470 510.380 1490.790 510.440 ;
        RECT 1489.550 462.640 1489.870 462.700 ;
        RECT 1490.470 462.640 1490.790 462.700 ;
        RECT 1489.550 462.500 1490.790 462.640 ;
        RECT 1489.550 462.440 1489.870 462.500 ;
        RECT 1490.470 462.440 1490.790 462.500 ;
        RECT 1489.550 427.760 1489.870 428.020 ;
        RECT 1489.640 427.280 1489.780 427.760 ;
        RECT 1490.010 427.280 1490.330 427.340 ;
        RECT 1489.640 427.140 1490.330 427.280 ;
        RECT 1490.010 427.080 1490.330 427.140 ;
        RECT 1489.090 414.020 1489.410 414.080 ;
        RECT 1490.010 414.020 1490.330 414.080 ;
        RECT 1489.090 413.880 1490.330 414.020 ;
        RECT 1489.090 413.820 1489.410 413.880 ;
        RECT 1490.010 413.820 1490.330 413.880 ;
        RECT 1489.090 366.080 1489.410 366.140 ;
        RECT 1490.010 366.080 1490.330 366.140 ;
        RECT 1489.090 365.940 1490.330 366.080 ;
        RECT 1489.090 365.880 1489.410 365.940 ;
        RECT 1490.010 365.880 1490.330 365.940 ;
        RECT 1489.090 317.460 1489.410 317.520 ;
        RECT 1490.010 317.460 1490.330 317.520 ;
        RECT 1489.090 317.320 1490.330 317.460 ;
        RECT 1489.090 317.260 1489.410 317.320 ;
        RECT 1490.010 317.260 1490.330 317.320 ;
        RECT 1489.090 269.180 1489.410 269.240 ;
        RECT 1490.010 269.180 1490.330 269.240 ;
        RECT 1489.090 269.040 1490.330 269.180 ;
        RECT 1489.090 268.980 1489.410 269.040 ;
        RECT 1490.010 268.980 1490.330 269.040 ;
        RECT 1490.010 255.580 1490.330 255.640 ;
        RECT 1489.180 255.440 1490.330 255.580 ;
        RECT 1489.180 255.300 1489.320 255.440 ;
        RECT 1490.010 255.380 1490.330 255.440 ;
        RECT 1489.090 255.040 1489.410 255.300 ;
        RECT 1489.090 138.280 1489.410 138.340 ;
        RECT 1488.720 138.140 1489.410 138.280 ;
        RECT 1488.720 137.660 1488.860 138.140 ;
        RECT 1489.090 138.080 1489.410 138.140 ;
        RECT 1488.630 137.400 1488.950 137.660 ;
        RECT 1488.170 131.140 1488.490 131.200 ;
        RECT 1488.630 131.140 1488.950 131.200 ;
        RECT 1488.170 131.000 1488.950 131.140 ;
        RECT 1488.170 130.940 1488.490 131.000 ;
        RECT 1488.630 130.940 1488.950 131.000 ;
        RECT 1488.170 107.000 1488.490 107.060 ;
        RECT 1489.550 107.000 1489.870 107.060 ;
        RECT 1488.170 106.860 1489.870 107.000 ;
        RECT 1488.170 106.800 1488.490 106.860 ;
        RECT 1489.550 106.800 1489.870 106.860 ;
        RECT 1490.010 19.960 1490.330 20.020 ;
        RECT 1590.290 19.960 1590.610 20.020 ;
        RECT 1490.010 19.820 1590.610 19.960 ;
        RECT 1490.010 19.760 1490.330 19.820 ;
        RECT 1590.290 19.760 1590.610 19.820 ;
      LAYER via ;
        RECT 1488.200 559.000 1488.460 559.260 ;
        RECT 1489.580 559.000 1489.840 559.260 ;
        RECT 1489.580 510.380 1489.840 510.640 ;
        RECT 1490.500 510.380 1490.760 510.640 ;
        RECT 1489.580 462.440 1489.840 462.700 ;
        RECT 1490.500 462.440 1490.760 462.700 ;
        RECT 1489.580 427.760 1489.840 428.020 ;
        RECT 1490.040 427.080 1490.300 427.340 ;
        RECT 1489.120 413.820 1489.380 414.080 ;
        RECT 1490.040 413.820 1490.300 414.080 ;
        RECT 1489.120 365.880 1489.380 366.140 ;
        RECT 1490.040 365.880 1490.300 366.140 ;
        RECT 1489.120 317.260 1489.380 317.520 ;
        RECT 1490.040 317.260 1490.300 317.520 ;
        RECT 1489.120 268.980 1489.380 269.240 ;
        RECT 1490.040 268.980 1490.300 269.240 ;
        RECT 1490.040 255.380 1490.300 255.640 ;
        RECT 1489.120 255.040 1489.380 255.300 ;
        RECT 1489.120 138.080 1489.380 138.340 ;
        RECT 1488.660 137.400 1488.920 137.660 ;
        RECT 1488.200 130.940 1488.460 131.200 ;
        RECT 1488.660 130.940 1488.920 131.200 ;
        RECT 1488.200 106.800 1488.460 107.060 ;
        RECT 1489.580 106.800 1489.840 107.060 ;
        RECT 1490.040 19.760 1490.300 20.020 ;
        RECT 1590.320 19.760 1590.580 20.020 ;
      LAYER met2 ;
        RECT 1487.050 600.170 1487.330 604.000 ;
        RECT 1487.050 600.030 1488.400 600.170 ;
        RECT 1487.050 600.000 1487.330 600.030 ;
        RECT 1488.260 559.290 1488.400 600.030 ;
        RECT 1488.200 558.970 1488.460 559.290 ;
        RECT 1489.580 558.970 1489.840 559.290 ;
        RECT 1489.640 510.670 1489.780 558.970 ;
        RECT 1489.580 510.350 1489.840 510.670 ;
        RECT 1490.500 510.350 1490.760 510.670 ;
        RECT 1490.560 462.730 1490.700 510.350 ;
        RECT 1489.580 462.410 1489.840 462.730 ;
        RECT 1490.500 462.410 1490.760 462.730 ;
        RECT 1489.640 428.050 1489.780 462.410 ;
        RECT 1489.580 427.730 1489.840 428.050 ;
        RECT 1490.040 427.050 1490.300 427.370 ;
        RECT 1490.100 414.110 1490.240 427.050 ;
        RECT 1489.120 413.790 1489.380 414.110 ;
        RECT 1490.040 413.790 1490.300 414.110 ;
        RECT 1489.180 366.170 1489.320 413.790 ;
        RECT 1489.120 365.850 1489.380 366.170 ;
        RECT 1490.040 365.850 1490.300 366.170 ;
        RECT 1490.100 317.550 1490.240 365.850 ;
        RECT 1489.120 317.230 1489.380 317.550 ;
        RECT 1490.040 317.230 1490.300 317.550 ;
        RECT 1489.180 269.270 1489.320 317.230 ;
        RECT 1489.120 268.950 1489.380 269.270 ;
        RECT 1490.040 268.950 1490.300 269.270 ;
        RECT 1490.100 255.670 1490.240 268.950 ;
        RECT 1490.040 255.350 1490.300 255.670 ;
        RECT 1489.120 255.010 1489.380 255.330 ;
        RECT 1489.180 211.325 1489.320 255.010 ;
        RECT 1489.110 210.955 1489.390 211.325 ;
        RECT 1488.650 179.675 1488.930 180.045 ;
        RECT 1488.720 179.250 1488.860 179.675 ;
        RECT 1488.720 179.110 1489.320 179.250 ;
        RECT 1489.180 138.370 1489.320 179.110 ;
        RECT 1489.120 138.050 1489.380 138.370 ;
        RECT 1488.660 137.370 1488.920 137.690 ;
        RECT 1488.720 131.230 1488.860 137.370 ;
        RECT 1488.200 130.910 1488.460 131.230 ;
        RECT 1488.660 130.910 1488.920 131.230 ;
        RECT 1488.260 107.090 1488.400 130.910 ;
        RECT 1488.200 106.770 1488.460 107.090 ;
        RECT 1489.580 106.770 1489.840 107.090 ;
        RECT 1489.640 62.290 1489.780 106.770 ;
        RECT 1489.640 62.150 1490.240 62.290 ;
        RECT 1490.100 20.050 1490.240 62.150 ;
        RECT 1490.040 19.730 1490.300 20.050 ;
        RECT 1590.320 19.730 1590.580 20.050 ;
        RECT 1590.380 2.400 1590.520 19.730 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
      LAYER via2 ;
        RECT 1489.110 211.000 1489.390 211.280 ;
        RECT 1488.650 179.720 1488.930 180.000 ;
      LAYER met3 ;
        RECT 1489.085 211.300 1489.415 211.305 ;
        RECT 1488.830 211.290 1489.415 211.300 ;
        RECT 1488.630 210.990 1489.415 211.290 ;
        RECT 1488.830 210.980 1489.415 210.990 ;
        RECT 1489.085 210.975 1489.415 210.980 ;
        RECT 1488.625 180.020 1488.955 180.025 ;
        RECT 1488.625 180.010 1489.210 180.020 ;
        RECT 1488.625 179.710 1489.410 180.010 ;
        RECT 1488.625 179.700 1489.210 179.710 ;
        RECT 1488.625 179.695 1488.955 179.700 ;
      LAYER via3 ;
        RECT 1488.860 210.980 1489.180 211.300 ;
        RECT 1488.860 179.700 1489.180 180.020 ;
      LAYER met4 ;
        RECT 1488.855 210.975 1489.185 211.305 ;
        RECT 1488.870 180.025 1489.170 210.975 ;
        RECT 1488.855 179.695 1489.185 180.025 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1496.910 19.280 1497.230 19.340 ;
        RECT 1608.230 19.280 1608.550 19.340 ;
        RECT 1496.910 19.140 1608.550 19.280 ;
        RECT 1496.910 19.080 1497.230 19.140 ;
        RECT 1608.230 19.080 1608.550 19.140 ;
      LAYER via ;
        RECT 1496.940 19.080 1497.200 19.340 ;
        RECT 1608.260 19.080 1608.520 19.340 ;
      LAYER met2 ;
        RECT 1496.250 600.170 1496.530 604.000 ;
        RECT 1496.250 600.030 1497.140 600.170 ;
        RECT 1496.250 600.000 1496.530 600.030 ;
        RECT 1497.000 19.370 1497.140 600.030 ;
        RECT 1496.940 19.050 1497.200 19.370 ;
        RECT 1608.260 19.050 1608.520 19.370 ;
        RECT 1608.320 2.400 1608.460 19.050 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1507.030 586.740 1507.350 586.800 ;
        RECT 1510.710 586.740 1511.030 586.800 ;
        RECT 1507.030 586.600 1511.030 586.740 ;
        RECT 1507.030 586.540 1507.350 586.600 ;
        RECT 1510.710 586.540 1511.030 586.600 ;
        RECT 1510.710 19.620 1511.030 19.680 ;
        RECT 1626.170 19.620 1626.490 19.680 ;
        RECT 1510.710 19.480 1626.490 19.620 ;
        RECT 1510.710 19.420 1511.030 19.480 ;
        RECT 1626.170 19.420 1626.490 19.480 ;
      LAYER via ;
        RECT 1507.060 586.540 1507.320 586.800 ;
        RECT 1510.740 586.540 1511.000 586.800 ;
        RECT 1510.740 19.420 1511.000 19.680 ;
        RECT 1626.200 19.420 1626.460 19.680 ;
      LAYER met2 ;
        RECT 1505.450 600.170 1505.730 604.000 ;
        RECT 1505.450 600.030 1507.260 600.170 ;
        RECT 1505.450 600.000 1505.730 600.030 ;
        RECT 1507.120 586.830 1507.260 600.030 ;
        RECT 1507.060 586.510 1507.320 586.830 ;
        RECT 1510.740 586.510 1511.000 586.830 ;
        RECT 1510.800 19.710 1510.940 586.510 ;
        RECT 1510.740 19.390 1511.000 19.710 ;
        RECT 1626.200 19.390 1626.460 19.710 ;
        RECT 1626.260 2.400 1626.400 19.390 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1516.230 586.740 1516.550 586.800 ;
        RECT 1521.290 586.740 1521.610 586.800 ;
        RECT 1516.230 586.600 1521.610 586.740 ;
        RECT 1516.230 586.540 1516.550 586.600 ;
        RECT 1521.290 586.540 1521.610 586.600 ;
        RECT 1521.290 18.940 1521.610 19.000 ;
        RECT 1644.110 18.940 1644.430 19.000 ;
        RECT 1521.290 18.800 1644.430 18.940 ;
        RECT 1521.290 18.740 1521.610 18.800 ;
        RECT 1644.110 18.740 1644.430 18.800 ;
      LAYER via ;
        RECT 1516.260 586.540 1516.520 586.800 ;
        RECT 1521.320 586.540 1521.580 586.800 ;
        RECT 1521.320 18.740 1521.580 19.000 ;
        RECT 1644.140 18.740 1644.400 19.000 ;
      LAYER met2 ;
        RECT 1514.650 600.170 1514.930 604.000 ;
        RECT 1514.650 600.030 1516.460 600.170 ;
        RECT 1514.650 600.000 1514.930 600.030 ;
        RECT 1516.320 586.830 1516.460 600.030 ;
        RECT 1516.260 586.510 1516.520 586.830 ;
        RECT 1521.320 586.510 1521.580 586.830 ;
        RECT 1521.380 19.030 1521.520 586.510 ;
        RECT 1521.320 18.710 1521.580 19.030 ;
        RECT 1644.140 18.710 1644.400 19.030 ;
        RECT 1644.200 2.400 1644.340 18.710 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.510 588.780 1524.830 588.840 ;
        RECT 1562.690 588.780 1563.010 588.840 ;
        RECT 1524.510 588.640 1563.010 588.780 ;
        RECT 1524.510 588.580 1524.830 588.640 ;
        RECT 1562.690 588.580 1563.010 588.640 ;
        RECT 1562.690 16.900 1563.010 16.960 ;
        RECT 1662.050 16.900 1662.370 16.960 ;
        RECT 1562.690 16.760 1662.370 16.900 ;
        RECT 1562.690 16.700 1563.010 16.760 ;
        RECT 1662.050 16.700 1662.370 16.760 ;
      LAYER via ;
        RECT 1524.540 588.580 1524.800 588.840 ;
        RECT 1562.720 588.580 1562.980 588.840 ;
        RECT 1562.720 16.700 1562.980 16.960 ;
        RECT 1662.080 16.700 1662.340 16.960 ;
      LAYER met2 ;
        RECT 1523.390 600.170 1523.670 604.000 ;
        RECT 1523.390 600.030 1524.740 600.170 ;
        RECT 1523.390 600.000 1523.670 600.030 ;
        RECT 1524.600 588.870 1524.740 600.030 ;
        RECT 1524.540 588.550 1524.800 588.870 ;
        RECT 1562.720 588.550 1562.980 588.870 ;
        RECT 1562.780 16.990 1562.920 588.550 ;
        RECT 1562.720 16.670 1562.980 16.990 ;
        RECT 1662.080 16.670 1662.340 16.990 ;
        RECT 1662.140 2.400 1662.280 16.670 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1534.170 590.140 1534.490 590.200 ;
        RECT 1538.310 590.140 1538.630 590.200 ;
        RECT 1534.170 590.000 1538.630 590.140 ;
        RECT 1534.170 589.940 1534.490 590.000 ;
        RECT 1538.310 589.940 1538.630 590.000 ;
        RECT 1538.310 18.600 1538.630 18.660 ;
        RECT 1679.530 18.600 1679.850 18.660 ;
        RECT 1538.310 18.460 1679.850 18.600 ;
        RECT 1538.310 18.400 1538.630 18.460 ;
        RECT 1679.530 18.400 1679.850 18.460 ;
      LAYER via ;
        RECT 1534.200 589.940 1534.460 590.200 ;
        RECT 1538.340 589.940 1538.600 590.200 ;
        RECT 1538.340 18.400 1538.600 18.660 ;
        RECT 1679.560 18.400 1679.820 18.660 ;
      LAYER met2 ;
        RECT 1532.590 600.170 1532.870 604.000 ;
        RECT 1532.590 600.030 1534.400 600.170 ;
        RECT 1532.590 600.000 1532.870 600.030 ;
        RECT 1534.260 590.230 1534.400 600.030 ;
        RECT 1534.200 589.910 1534.460 590.230 ;
        RECT 1538.340 589.910 1538.600 590.230 ;
        RECT 1538.400 18.690 1538.540 589.910 ;
        RECT 1538.340 18.370 1538.600 18.690 ;
        RECT 1679.560 18.370 1679.820 18.690 ;
        RECT 1679.620 2.400 1679.760 18.370 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1543.370 581.640 1543.690 581.700 ;
        RECT 1545.210 581.640 1545.530 581.700 ;
        RECT 1543.370 581.500 1545.530 581.640 ;
        RECT 1543.370 581.440 1543.690 581.500 ;
        RECT 1545.210 581.440 1545.530 581.500 ;
        RECT 1545.210 18.260 1545.530 18.320 ;
        RECT 1697.470 18.260 1697.790 18.320 ;
        RECT 1545.210 18.120 1697.790 18.260 ;
        RECT 1545.210 18.060 1545.530 18.120 ;
        RECT 1697.470 18.060 1697.790 18.120 ;
      LAYER via ;
        RECT 1543.400 581.440 1543.660 581.700 ;
        RECT 1545.240 581.440 1545.500 581.700 ;
        RECT 1545.240 18.060 1545.500 18.320 ;
        RECT 1697.500 18.060 1697.760 18.320 ;
      LAYER met2 ;
        RECT 1541.790 600.170 1542.070 604.000 ;
        RECT 1541.790 600.030 1543.600 600.170 ;
        RECT 1541.790 600.000 1542.070 600.030 ;
        RECT 1543.460 581.730 1543.600 600.030 ;
        RECT 1543.400 581.410 1543.660 581.730 ;
        RECT 1545.240 581.410 1545.500 581.730 ;
        RECT 1545.300 18.350 1545.440 581.410 ;
        RECT 1545.240 18.030 1545.500 18.350 ;
        RECT 1697.500 18.030 1697.760 18.350 ;
        RECT 1697.560 2.400 1697.700 18.030 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.510 461.960 1041.830 462.020 ;
        RECT 1045.190 461.960 1045.510 462.020 ;
        RECT 1041.510 461.820 1045.510 461.960 ;
        RECT 1041.510 461.760 1041.830 461.820 ;
        RECT 1045.190 461.760 1045.510 461.820 ;
        RECT 1041.510 444.960 1041.830 445.020 ;
        RECT 1043.350 444.960 1043.670 445.020 ;
        RECT 1041.510 444.820 1043.670 444.960 ;
        RECT 1041.510 444.760 1041.830 444.820 ;
        RECT 1043.350 444.760 1043.670 444.820 ;
        RECT 1042.890 372.880 1043.210 372.940 ;
        RECT 1043.350 372.880 1043.670 372.940 ;
        RECT 1042.890 372.740 1043.670 372.880 ;
        RECT 1042.890 372.680 1043.210 372.740 ;
        RECT 1043.350 372.680 1043.670 372.740 ;
        RECT 1043.350 110.880 1043.670 111.140 ;
        RECT 1043.440 110.460 1043.580 110.880 ;
        RECT 1043.350 110.200 1043.670 110.460 ;
        RECT 1042.430 96.800 1042.750 96.860 ;
        RECT 1043.350 96.800 1043.670 96.860 ;
        RECT 1042.430 96.660 1043.670 96.800 ;
        RECT 1042.430 96.600 1042.750 96.660 ;
        RECT 1043.350 96.600 1043.670 96.660 ;
        RECT 1041.050 72.660 1041.370 72.720 ;
        RECT 1042.430 72.660 1042.750 72.720 ;
        RECT 1041.050 72.520 1042.750 72.660 ;
        RECT 1041.050 72.460 1041.370 72.520 ;
        RECT 1042.430 72.460 1042.750 72.520 ;
        RECT 821.170 22.340 821.490 22.400 ;
        RECT 1041.050 22.340 1041.370 22.400 ;
        RECT 821.170 22.200 1041.370 22.340 ;
        RECT 821.170 22.140 821.490 22.200 ;
        RECT 1041.050 22.140 1041.370 22.200 ;
        RECT 734.230 17.580 734.550 17.640 ;
        RECT 821.170 17.580 821.490 17.640 ;
        RECT 734.230 17.440 821.490 17.580 ;
        RECT 734.230 17.380 734.550 17.440 ;
        RECT 821.170 17.380 821.490 17.440 ;
      LAYER via ;
        RECT 1041.540 461.760 1041.800 462.020 ;
        RECT 1045.220 461.760 1045.480 462.020 ;
        RECT 1041.540 444.760 1041.800 445.020 ;
        RECT 1043.380 444.760 1043.640 445.020 ;
        RECT 1042.920 372.680 1043.180 372.940 ;
        RECT 1043.380 372.680 1043.640 372.940 ;
        RECT 1043.380 110.880 1043.640 111.140 ;
        RECT 1043.380 110.200 1043.640 110.460 ;
        RECT 1042.460 96.600 1042.720 96.860 ;
        RECT 1043.380 96.600 1043.640 96.860 ;
        RECT 1041.080 72.460 1041.340 72.720 ;
        RECT 1042.460 72.460 1042.720 72.720 ;
        RECT 821.200 22.140 821.460 22.400 ;
        RECT 1041.080 22.140 1041.340 22.400 ;
        RECT 734.260 17.380 734.520 17.640 ;
        RECT 821.200 17.380 821.460 17.640 ;
      LAYER met2 ;
        RECT 1046.830 600.000 1047.110 604.000 ;
        RECT 1046.890 598.810 1047.030 600.000 ;
        RECT 1046.660 598.670 1047.030 598.810 ;
        RECT 1046.660 579.885 1046.800 598.670 ;
        RECT 1045.210 579.515 1045.490 579.885 ;
        RECT 1046.590 579.515 1046.870 579.885 ;
        RECT 1045.280 462.050 1045.420 579.515 ;
        RECT 1041.540 461.730 1041.800 462.050 ;
        RECT 1045.220 461.730 1045.480 462.050 ;
        RECT 1041.600 445.050 1041.740 461.730 ;
        RECT 1041.540 444.730 1041.800 445.050 ;
        RECT 1043.380 444.730 1043.640 445.050 ;
        RECT 1043.440 372.970 1043.580 444.730 ;
        RECT 1042.920 372.650 1043.180 372.970 ;
        RECT 1043.380 372.650 1043.640 372.970 ;
        RECT 1042.980 351.970 1043.120 372.650 ;
        RECT 1042.980 351.830 1043.580 351.970 ;
        RECT 1043.440 316.610 1043.580 351.830 ;
        RECT 1042.980 316.470 1043.580 316.610 ;
        RECT 1042.980 255.410 1043.120 316.470 ;
        RECT 1042.980 255.270 1043.580 255.410 ;
        RECT 1043.440 207.130 1043.580 255.270 ;
        RECT 1042.980 206.990 1043.580 207.130 ;
        RECT 1042.980 158.850 1043.120 206.990 ;
        RECT 1042.980 158.710 1043.580 158.850 ;
        RECT 1043.440 111.170 1043.580 158.710 ;
        RECT 1043.380 110.850 1043.640 111.170 ;
        RECT 1043.380 110.170 1043.640 110.490 ;
        RECT 1043.440 96.890 1043.580 110.170 ;
        RECT 1042.460 96.570 1042.720 96.890 ;
        RECT 1043.380 96.570 1043.640 96.890 ;
        RECT 1042.520 72.750 1042.660 96.570 ;
        RECT 1041.080 72.430 1041.340 72.750 ;
        RECT 1042.460 72.430 1042.720 72.750 ;
        RECT 1041.140 22.430 1041.280 72.430 ;
        RECT 821.200 22.110 821.460 22.430 ;
        RECT 1041.080 22.110 1041.340 22.430 ;
        RECT 821.260 17.670 821.400 22.110 ;
        RECT 734.260 17.350 734.520 17.670 ;
        RECT 821.200 17.350 821.460 17.670 ;
        RECT 734.320 2.400 734.460 17.350 ;
        RECT 734.110 -4.800 734.670 2.400 ;
      LAYER via2 ;
        RECT 1045.210 579.560 1045.490 579.840 ;
        RECT 1046.590 579.560 1046.870 579.840 ;
      LAYER met3 ;
        RECT 1045.185 579.850 1045.515 579.865 ;
        RECT 1046.565 579.850 1046.895 579.865 ;
        RECT 1045.185 579.550 1046.895 579.850 ;
        RECT 1045.185 579.535 1045.515 579.550 ;
        RECT 1046.565 579.535 1046.895 579.550 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1552.110 17.920 1552.430 17.980 ;
        RECT 1715.410 17.920 1715.730 17.980 ;
        RECT 1552.110 17.780 1715.730 17.920 ;
        RECT 1552.110 17.720 1552.430 17.780 ;
        RECT 1715.410 17.720 1715.730 17.780 ;
      LAYER via ;
        RECT 1552.140 17.720 1552.400 17.980 ;
        RECT 1715.440 17.720 1715.700 17.980 ;
      LAYER met2 ;
        RECT 1550.990 600.170 1551.270 604.000 ;
        RECT 1550.990 600.030 1552.340 600.170 ;
        RECT 1550.990 600.000 1551.270 600.030 ;
        RECT 1552.200 18.010 1552.340 600.030 ;
        RECT 1552.140 17.690 1552.400 18.010 ;
        RECT 1715.440 17.690 1715.700 18.010 ;
        RECT 1715.500 2.400 1715.640 17.690 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1561.770 586.740 1562.090 586.800 ;
        RECT 1565.910 586.740 1566.230 586.800 ;
        RECT 1561.770 586.600 1566.230 586.740 ;
        RECT 1561.770 586.540 1562.090 586.600 ;
        RECT 1565.910 586.540 1566.230 586.600 ;
        RECT 1565.910 17.580 1566.230 17.640 ;
        RECT 1733.350 17.580 1733.670 17.640 ;
        RECT 1565.910 17.440 1733.670 17.580 ;
        RECT 1565.910 17.380 1566.230 17.440 ;
        RECT 1733.350 17.380 1733.670 17.440 ;
      LAYER via ;
        RECT 1561.800 586.540 1562.060 586.800 ;
        RECT 1565.940 586.540 1566.200 586.800 ;
        RECT 1565.940 17.380 1566.200 17.640 ;
        RECT 1733.380 17.380 1733.640 17.640 ;
      LAYER met2 ;
        RECT 1560.190 600.170 1560.470 604.000 ;
        RECT 1560.190 600.030 1562.000 600.170 ;
        RECT 1560.190 600.000 1560.470 600.030 ;
        RECT 1561.860 586.830 1562.000 600.030 ;
        RECT 1561.800 586.510 1562.060 586.830 ;
        RECT 1565.940 586.510 1566.200 586.830 ;
        RECT 1566.000 17.670 1566.140 586.510 ;
        RECT 1565.940 17.350 1566.200 17.670 ;
        RECT 1733.380 17.350 1733.640 17.670 ;
        RECT 1733.440 2.400 1733.580 17.350 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1610.990 589.460 1611.310 589.520 ;
        RECT 1581.640 589.320 1611.310 589.460 ;
        RECT 1570.970 588.440 1571.290 588.500 ;
        RECT 1581.640 588.440 1581.780 589.320 ;
        RECT 1610.990 589.260 1611.310 589.320 ;
        RECT 1570.970 588.300 1581.780 588.440 ;
        RECT 1570.970 588.240 1571.290 588.300 ;
        RECT 1610.990 15.880 1611.310 15.940 ;
        RECT 1751.290 15.880 1751.610 15.940 ;
        RECT 1610.990 15.740 1751.610 15.880 ;
        RECT 1610.990 15.680 1611.310 15.740 ;
        RECT 1751.290 15.680 1751.610 15.740 ;
      LAYER via ;
        RECT 1571.000 588.240 1571.260 588.500 ;
        RECT 1611.020 589.260 1611.280 589.520 ;
        RECT 1611.020 15.680 1611.280 15.940 ;
        RECT 1751.320 15.680 1751.580 15.940 ;
      LAYER met2 ;
        RECT 1569.390 600.170 1569.670 604.000 ;
        RECT 1569.390 600.030 1571.200 600.170 ;
        RECT 1569.390 600.000 1569.670 600.030 ;
        RECT 1571.060 588.530 1571.200 600.030 ;
        RECT 1611.020 589.230 1611.280 589.550 ;
        RECT 1571.000 588.210 1571.260 588.530 ;
        RECT 1611.080 15.970 1611.220 589.230 ;
        RECT 1611.020 15.650 1611.280 15.970 ;
        RECT 1751.320 15.650 1751.580 15.970 ;
        RECT 1751.380 2.400 1751.520 15.650 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.710 17.240 1580.030 17.300 ;
        RECT 1768.770 17.240 1769.090 17.300 ;
        RECT 1579.710 17.100 1769.090 17.240 ;
        RECT 1579.710 17.040 1580.030 17.100 ;
        RECT 1768.770 17.040 1769.090 17.100 ;
      LAYER via ;
        RECT 1579.740 17.040 1580.000 17.300 ;
        RECT 1768.800 17.040 1769.060 17.300 ;
      LAYER met2 ;
        RECT 1578.590 600.170 1578.870 604.000 ;
        RECT 1578.590 600.030 1579.940 600.170 ;
        RECT 1578.590 600.000 1578.870 600.030 ;
        RECT 1579.800 17.330 1579.940 600.030 ;
        RECT 1579.740 17.010 1580.000 17.330 ;
        RECT 1768.800 17.010 1769.060 17.330 ;
        RECT 1768.860 2.400 1769.000 17.010 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1589.370 589.120 1589.690 589.180 ;
        RECT 1652.390 589.120 1652.710 589.180 ;
        RECT 1589.370 588.980 1652.710 589.120 ;
        RECT 1589.370 588.920 1589.690 588.980 ;
        RECT 1652.390 588.920 1652.710 588.980 ;
        RECT 1652.390 15.540 1652.710 15.600 ;
        RECT 1786.710 15.540 1787.030 15.600 ;
        RECT 1652.390 15.400 1787.030 15.540 ;
        RECT 1652.390 15.340 1652.710 15.400 ;
        RECT 1786.710 15.340 1787.030 15.400 ;
      LAYER via ;
        RECT 1589.400 588.920 1589.660 589.180 ;
        RECT 1652.420 588.920 1652.680 589.180 ;
        RECT 1652.420 15.340 1652.680 15.600 ;
        RECT 1786.740 15.340 1787.000 15.600 ;
      LAYER met2 ;
        RECT 1587.790 600.170 1588.070 604.000 ;
        RECT 1587.790 600.030 1589.600 600.170 ;
        RECT 1587.790 600.000 1588.070 600.030 ;
        RECT 1589.460 589.210 1589.600 600.030 ;
        RECT 1589.400 588.890 1589.660 589.210 ;
        RECT 1652.420 588.890 1652.680 589.210 ;
        RECT 1652.480 15.630 1652.620 588.890 ;
        RECT 1652.420 15.310 1652.680 15.630 ;
        RECT 1786.740 15.310 1787.000 15.630 ;
        RECT 1786.800 2.400 1786.940 15.310 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1598.570 592.860 1598.890 592.920 ;
        RECT 1659.290 592.860 1659.610 592.920 ;
        RECT 1598.570 592.720 1659.610 592.860 ;
        RECT 1598.570 592.660 1598.890 592.720 ;
        RECT 1659.290 592.660 1659.610 592.720 ;
        RECT 1659.290 16.220 1659.610 16.280 ;
        RECT 1804.650 16.220 1804.970 16.280 ;
        RECT 1659.290 16.080 1804.970 16.220 ;
        RECT 1659.290 16.020 1659.610 16.080 ;
        RECT 1804.650 16.020 1804.970 16.080 ;
      LAYER via ;
        RECT 1598.600 592.660 1598.860 592.920 ;
        RECT 1659.320 592.660 1659.580 592.920 ;
        RECT 1659.320 16.020 1659.580 16.280 ;
        RECT 1804.680 16.020 1804.940 16.280 ;
      LAYER met2 ;
        RECT 1596.990 600.170 1597.270 604.000 ;
        RECT 1596.990 600.030 1598.800 600.170 ;
        RECT 1596.990 600.000 1597.270 600.030 ;
        RECT 1598.660 592.950 1598.800 600.030 ;
        RECT 1598.600 592.630 1598.860 592.950 ;
        RECT 1659.320 592.630 1659.580 592.950 ;
        RECT 1659.380 16.310 1659.520 592.630 ;
        RECT 1659.320 15.990 1659.580 16.310 ;
        RECT 1804.680 15.990 1804.940 16.310 ;
        RECT 1804.740 2.400 1804.880 15.990 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1607.310 20.640 1607.630 20.700 ;
        RECT 1822.590 20.640 1822.910 20.700 ;
        RECT 1607.310 20.500 1822.910 20.640 ;
        RECT 1607.310 20.440 1607.630 20.500 ;
        RECT 1822.590 20.440 1822.910 20.500 ;
      LAYER via ;
        RECT 1607.340 20.440 1607.600 20.700 ;
        RECT 1822.620 20.440 1822.880 20.700 ;
      LAYER met2 ;
        RECT 1606.190 600.170 1606.470 604.000 ;
        RECT 1606.190 600.030 1607.540 600.170 ;
        RECT 1606.190 600.000 1606.470 600.030 ;
        RECT 1607.400 20.730 1607.540 600.030 ;
        RECT 1607.340 20.410 1607.600 20.730 ;
        RECT 1822.620 20.410 1822.880 20.730 ;
        RECT 1822.680 2.400 1822.820 20.410 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1616.970 593.200 1617.290 593.260 ;
        RECT 1666.190 593.200 1666.510 593.260 ;
        RECT 1616.970 593.060 1666.510 593.200 ;
        RECT 1616.970 593.000 1617.290 593.060 ;
        RECT 1666.190 593.000 1666.510 593.060 ;
        RECT 1666.190 16.560 1666.510 16.620 ;
        RECT 1840.070 16.560 1840.390 16.620 ;
        RECT 1666.190 16.420 1840.390 16.560 ;
        RECT 1666.190 16.360 1666.510 16.420 ;
        RECT 1840.070 16.360 1840.390 16.420 ;
      LAYER via ;
        RECT 1617.000 593.000 1617.260 593.260 ;
        RECT 1666.220 593.000 1666.480 593.260 ;
        RECT 1666.220 16.360 1666.480 16.620 ;
        RECT 1840.100 16.360 1840.360 16.620 ;
      LAYER met2 ;
        RECT 1615.390 600.170 1615.670 604.000 ;
        RECT 1615.390 600.030 1617.200 600.170 ;
        RECT 1615.390 600.000 1615.670 600.030 ;
        RECT 1617.060 593.290 1617.200 600.030 ;
        RECT 1617.000 592.970 1617.260 593.290 ;
        RECT 1666.220 592.970 1666.480 593.290 ;
        RECT 1666.280 16.650 1666.420 592.970 ;
        RECT 1666.220 16.330 1666.480 16.650 ;
        RECT 1840.100 16.330 1840.360 16.650 ;
        RECT 1840.160 2.400 1840.300 16.330 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1626.170 587.080 1626.490 587.140 ;
        RECT 1628.010 587.080 1628.330 587.140 ;
        RECT 1626.170 586.940 1628.330 587.080 ;
        RECT 1626.170 586.880 1626.490 586.940 ;
        RECT 1628.010 586.880 1628.330 586.940 ;
        RECT 1628.010 20.300 1628.330 20.360 ;
        RECT 1858.010 20.300 1858.330 20.360 ;
        RECT 1628.010 20.160 1858.330 20.300 ;
        RECT 1628.010 20.100 1628.330 20.160 ;
        RECT 1858.010 20.100 1858.330 20.160 ;
      LAYER via ;
        RECT 1626.200 586.880 1626.460 587.140 ;
        RECT 1628.040 586.880 1628.300 587.140 ;
        RECT 1628.040 20.100 1628.300 20.360 ;
        RECT 1858.040 20.100 1858.300 20.360 ;
      LAYER met2 ;
        RECT 1624.590 600.170 1624.870 604.000 ;
        RECT 1624.590 600.030 1626.400 600.170 ;
        RECT 1624.590 600.000 1624.870 600.030 ;
        RECT 1626.260 587.170 1626.400 600.030 ;
        RECT 1626.200 586.850 1626.460 587.170 ;
        RECT 1628.040 586.850 1628.300 587.170 ;
        RECT 1628.100 20.390 1628.240 586.850 ;
        RECT 1628.040 20.070 1628.300 20.390 ;
        RECT 1858.040 20.070 1858.300 20.390 ;
        RECT 1858.100 2.400 1858.240 20.070 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1634.450 587.080 1634.770 587.140 ;
        RECT 1673.090 587.080 1673.410 587.140 ;
        RECT 1634.450 586.940 1673.410 587.080 ;
        RECT 1634.450 586.880 1634.770 586.940 ;
        RECT 1673.090 586.880 1673.410 586.940 ;
        RECT 1673.090 16.900 1673.410 16.960 ;
        RECT 1875.950 16.900 1876.270 16.960 ;
        RECT 1673.090 16.760 1876.270 16.900 ;
        RECT 1673.090 16.700 1673.410 16.760 ;
        RECT 1875.950 16.700 1876.270 16.760 ;
      LAYER via ;
        RECT 1634.480 586.880 1634.740 587.140 ;
        RECT 1673.120 586.880 1673.380 587.140 ;
        RECT 1673.120 16.700 1673.380 16.960 ;
        RECT 1875.980 16.700 1876.240 16.960 ;
      LAYER met2 ;
        RECT 1633.790 600.170 1634.070 604.000 ;
        RECT 1633.790 600.030 1634.680 600.170 ;
        RECT 1633.790 600.000 1634.070 600.030 ;
        RECT 1634.540 587.170 1634.680 600.030 ;
        RECT 1634.480 586.850 1634.740 587.170 ;
        RECT 1673.120 586.850 1673.380 587.170 ;
        RECT 1673.180 16.990 1673.320 586.850 ;
        RECT 1673.120 16.670 1673.380 16.990 ;
        RECT 1875.980 16.670 1876.240 16.990 ;
        RECT 1876.040 2.400 1876.180 16.670 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 894.310 32.540 894.630 32.600 ;
        RECT 1056.230 32.540 1056.550 32.600 ;
        RECT 894.310 32.400 1056.550 32.540 ;
        RECT 894.310 32.340 894.630 32.400 ;
        RECT 1056.230 32.340 1056.550 32.400 ;
        RECT 752.170 19.280 752.490 19.340 ;
        RECT 765.970 19.280 766.290 19.340 ;
        RECT 752.170 19.140 766.290 19.280 ;
        RECT 752.170 19.080 752.490 19.140 ;
        RECT 765.970 19.080 766.290 19.140 ;
        RECT 811.510 19.280 811.830 19.340 ;
        RECT 894.310 19.280 894.630 19.340 ;
        RECT 811.510 19.140 894.630 19.280 ;
        RECT 811.510 19.080 811.830 19.140 ;
        RECT 894.310 19.080 894.630 19.140 ;
      LAYER via ;
        RECT 894.340 32.340 894.600 32.600 ;
        RECT 1056.260 32.340 1056.520 32.600 ;
        RECT 752.200 19.080 752.460 19.340 ;
        RECT 766.000 19.080 766.260 19.340 ;
        RECT 811.540 19.080 811.800 19.340 ;
        RECT 894.340 19.080 894.600 19.340 ;
      LAYER met2 ;
        RECT 1056.030 600.000 1056.310 604.000 ;
        RECT 1056.090 598.810 1056.230 600.000 ;
        RECT 1056.090 598.670 1056.460 598.810 ;
        RECT 1056.320 32.630 1056.460 598.670 ;
        RECT 894.340 32.310 894.600 32.630 ;
        RECT 1056.260 32.310 1056.520 32.630 ;
        RECT 894.400 19.370 894.540 32.310 ;
        RECT 752.200 19.050 752.460 19.370 ;
        RECT 766.000 19.050 766.260 19.370 ;
        RECT 811.540 19.050 811.800 19.370 ;
        RECT 894.340 19.050 894.600 19.370 ;
        RECT 752.260 2.400 752.400 19.050 ;
        RECT 766.060 18.885 766.200 19.050 ;
        RECT 811.600 18.885 811.740 19.050 ;
        RECT 765.990 18.515 766.270 18.885 ;
        RECT 811.530 18.515 811.810 18.885 ;
        RECT 752.050 -4.800 752.610 2.400 ;
      LAYER via2 ;
        RECT 765.990 18.560 766.270 18.840 ;
        RECT 811.530 18.560 811.810 18.840 ;
      LAYER met3 ;
        RECT 765.965 18.850 766.295 18.865 ;
        RECT 811.505 18.850 811.835 18.865 ;
        RECT 765.965 18.550 811.835 18.850 ;
        RECT 765.965 18.535 766.295 18.550 ;
        RECT 811.505 18.535 811.835 18.550 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1644.570 586.740 1644.890 586.800 ;
        RECT 1648.710 586.740 1649.030 586.800 ;
        RECT 1644.570 586.600 1649.030 586.740 ;
        RECT 1644.570 586.540 1644.890 586.600 ;
        RECT 1648.710 586.540 1649.030 586.600 ;
        RECT 1648.710 19.620 1649.030 19.680 ;
        RECT 1893.890 19.620 1894.210 19.680 ;
        RECT 1648.710 19.480 1894.210 19.620 ;
        RECT 1648.710 19.420 1649.030 19.480 ;
        RECT 1893.890 19.420 1894.210 19.480 ;
      LAYER via ;
        RECT 1644.600 586.540 1644.860 586.800 ;
        RECT 1648.740 586.540 1649.000 586.800 ;
        RECT 1648.740 19.420 1649.000 19.680 ;
        RECT 1893.920 19.420 1894.180 19.680 ;
      LAYER met2 ;
        RECT 1642.990 600.170 1643.270 604.000 ;
        RECT 1642.990 600.030 1644.800 600.170 ;
        RECT 1642.990 600.000 1643.270 600.030 ;
        RECT 1644.660 586.830 1644.800 600.030 ;
        RECT 1644.600 586.510 1644.860 586.830 ;
        RECT 1648.740 586.510 1649.000 586.830 ;
        RECT 1648.800 19.710 1648.940 586.510 ;
        RECT 1648.740 19.390 1649.000 19.710 ;
        RECT 1893.920 19.390 1894.180 19.710 ;
        RECT 1893.980 2.400 1894.120 19.390 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1653.310 588.440 1653.630 588.500 ;
        RECT 1907.690 588.440 1908.010 588.500 ;
        RECT 1653.310 588.300 1908.010 588.440 ;
        RECT 1653.310 588.240 1653.630 588.300 ;
        RECT 1907.690 588.240 1908.010 588.300 ;
        RECT 1907.690 20.640 1908.010 20.700 ;
        RECT 1911.830 20.640 1912.150 20.700 ;
        RECT 1907.690 20.500 1912.150 20.640 ;
        RECT 1907.690 20.440 1908.010 20.500 ;
        RECT 1911.830 20.440 1912.150 20.500 ;
      LAYER via ;
        RECT 1653.340 588.240 1653.600 588.500 ;
        RECT 1907.720 588.240 1907.980 588.500 ;
        RECT 1907.720 20.440 1907.980 20.700 ;
        RECT 1911.860 20.440 1912.120 20.700 ;
      LAYER met2 ;
        RECT 1651.730 600.170 1652.010 604.000 ;
        RECT 1651.730 600.030 1653.540 600.170 ;
        RECT 1651.730 600.000 1652.010 600.030 ;
        RECT 1653.400 588.530 1653.540 600.030 ;
        RECT 1653.340 588.210 1653.600 588.530 ;
        RECT 1907.720 588.210 1907.980 588.530 ;
        RECT 1907.780 20.730 1907.920 588.210 ;
        RECT 1907.720 20.410 1907.980 20.730 ;
        RECT 1911.860 20.410 1912.120 20.730 ;
        RECT 1911.920 2.400 1912.060 20.410 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.510 587.420 1662.830 587.480 ;
        RECT 1686.890 587.420 1687.210 587.480 ;
        RECT 1662.510 587.280 1687.210 587.420 ;
        RECT 1662.510 587.220 1662.830 587.280 ;
        RECT 1686.890 587.220 1687.210 587.280 ;
        RECT 1686.890 19.960 1687.210 20.020 ;
        RECT 1929.310 19.960 1929.630 20.020 ;
        RECT 1686.890 19.820 1929.630 19.960 ;
        RECT 1686.890 19.760 1687.210 19.820 ;
        RECT 1929.310 19.760 1929.630 19.820 ;
      LAYER via ;
        RECT 1662.540 587.220 1662.800 587.480 ;
        RECT 1686.920 587.220 1687.180 587.480 ;
        RECT 1686.920 19.760 1687.180 20.020 ;
        RECT 1929.340 19.760 1929.600 20.020 ;
      LAYER met2 ;
        RECT 1660.930 600.170 1661.210 604.000 ;
        RECT 1660.930 600.030 1662.740 600.170 ;
        RECT 1660.930 600.000 1661.210 600.030 ;
        RECT 1662.600 587.510 1662.740 600.030 ;
        RECT 1662.540 587.190 1662.800 587.510 ;
        RECT 1686.920 587.190 1687.180 587.510 ;
        RECT 1686.980 20.050 1687.120 587.190 ;
        RECT 1686.920 19.730 1687.180 20.050 ;
        RECT 1929.340 19.730 1929.600 20.050 ;
        RECT 1929.400 2.400 1929.540 19.730 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1690.110 589.120 1690.430 589.180 ;
        RECT 1787.630 589.120 1787.950 589.180 ;
        RECT 1690.110 588.980 1787.950 589.120 ;
        RECT 1690.110 588.920 1690.430 588.980 ;
        RECT 1787.630 588.920 1787.950 588.980 ;
        RECT 1788.550 589.120 1788.870 589.180 ;
        RECT 1935.290 589.120 1935.610 589.180 ;
        RECT 1788.550 588.980 1935.610 589.120 ;
        RECT 1788.550 588.920 1788.870 588.980 ;
        RECT 1935.290 588.920 1935.610 588.980 ;
        RECT 1934.830 15.200 1935.150 15.260 ;
        RECT 1947.250 15.200 1947.570 15.260 ;
        RECT 1934.830 15.060 1947.570 15.200 ;
        RECT 1934.830 15.000 1935.150 15.060 ;
        RECT 1947.250 15.000 1947.570 15.060 ;
      LAYER via ;
        RECT 1690.140 588.920 1690.400 589.180 ;
        RECT 1787.660 588.920 1787.920 589.180 ;
        RECT 1788.580 588.920 1788.840 589.180 ;
        RECT 1935.320 588.920 1935.580 589.180 ;
        RECT 1934.860 15.000 1935.120 15.260 ;
        RECT 1947.280 15.000 1947.540 15.260 ;
      LAYER met2 ;
        RECT 1670.130 600.170 1670.410 604.000 ;
        RECT 1670.130 600.030 1671.940 600.170 ;
        RECT 1670.130 600.000 1670.410 600.030 ;
        RECT 1671.800 589.405 1671.940 600.030 ;
        RECT 1671.730 589.035 1672.010 589.405 ;
        RECT 1690.130 589.035 1690.410 589.405 ;
        RECT 1787.720 589.210 1788.780 589.290 ;
        RECT 1787.660 589.150 1788.840 589.210 ;
        RECT 1690.140 588.890 1690.400 589.035 ;
        RECT 1787.660 588.890 1787.920 589.150 ;
        RECT 1788.580 588.890 1788.840 589.150 ;
        RECT 1935.320 588.890 1935.580 589.210 ;
        RECT 1935.380 38.490 1935.520 588.890 ;
        RECT 1934.920 38.350 1935.520 38.490 ;
        RECT 1934.920 15.290 1935.060 38.350 ;
        RECT 1934.860 14.970 1935.120 15.290 ;
        RECT 1947.280 14.970 1947.540 15.290 ;
        RECT 1947.340 2.400 1947.480 14.970 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER via2 ;
        RECT 1671.730 589.080 1672.010 589.360 ;
        RECT 1690.130 589.080 1690.410 589.360 ;
      LAYER met3 ;
        RECT 1671.705 589.370 1672.035 589.385 ;
        RECT 1690.105 589.370 1690.435 589.385 ;
        RECT 1671.705 589.070 1690.435 589.370 ;
        RECT 1671.705 589.055 1672.035 589.070 ;
        RECT 1690.105 589.055 1690.435 589.070 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1680.910 587.080 1681.230 587.140 ;
        RECT 1693.790 587.080 1694.110 587.140 ;
        RECT 1680.910 586.940 1694.110 587.080 ;
        RECT 1680.910 586.880 1681.230 586.940 ;
        RECT 1693.790 586.880 1694.110 586.940 ;
        RECT 1965.190 19.960 1965.510 20.020 ;
        RECT 1945.040 19.820 1965.510 19.960 ;
        RECT 1693.790 19.280 1694.110 19.340 ;
        RECT 1945.040 19.280 1945.180 19.820 ;
        RECT 1965.190 19.760 1965.510 19.820 ;
        RECT 1693.790 19.140 1945.180 19.280 ;
        RECT 1693.790 19.080 1694.110 19.140 ;
      LAYER via ;
        RECT 1680.940 586.880 1681.200 587.140 ;
        RECT 1693.820 586.880 1694.080 587.140 ;
        RECT 1693.820 19.080 1694.080 19.340 ;
        RECT 1965.220 19.760 1965.480 20.020 ;
      LAYER met2 ;
        RECT 1679.330 600.170 1679.610 604.000 ;
        RECT 1679.330 600.030 1681.140 600.170 ;
        RECT 1679.330 600.000 1679.610 600.030 ;
        RECT 1681.000 587.170 1681.140 600.030 ;
        RECT 1680.940 586.850 1681.200 587.170 ;
        RECT 1693.820 586.850 1694.080 587.170 ;
        RECT 1693.880 19.370 1694.020 586.850 ;
        RECT 1965.220 19.730 1965.480 20.050 ;
        RECT 1693.820 19.050 1694.080 19.370 ;
        RECT 1965.280 2.400 1965.420 19.730 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1690.110 593.200 1690.430 593.260 ;
        RECT 1969.330 593.200 1969.650 593.260 ;
        RECT 1690.110 593.060 1969.650 593.200 ;
        RECT 1690.110 593.000 1690.430 593.060 ;
        RECT 1969.330 593.000 1969.650 593.060 ;
        RECT 1969.790 20.300 1970.110 20.360 ;
        RECT 1983.130 20.300 1983.450 20.360 ;
        RECT 1969.790 20.160 1983.450 20.300 ;
        RECT 1969.790 20.100 1970.110 20.160 ;
        RECT 1983.130 20.100 1983.450 20.160 ;
      LAYER via ;
        RECT 1690.140 593.000 1690.400 593.260 ;
        RECT 1969.360 593.000 1969.620 593.260 ;
        RECT 1969.820 20.100 1970.080 20.360 ;
        RECT 1983.160 20.100 1983.420 20.360 ;
      LAYER met2 ;
        RECT 1688.530 600.170 1688.810 604.000 ;
        RECT 1688.530 600.030 1690.340 600.170 ;
        RECT 1688.530 600.000 1688.810 600.030 ;
        RECT 1690.200 593.290 1690.340 600.030 ;
        RECT 1690.140 592.970 1690.400 593.290 ;
        RECT 1969.360 592.970 1969.620 593.290 ;
        RECT 1969.420 586.570 1969.560 592.970 ;
        RECT 1969.420 586.430 1970.020 586.570 ;
        RECT 1969.880 20.390 1970.020 586.430 ;
        RECT 1969.820 20.070 1970.080 20.390 ;
        RECT 1983.160 20.070 1983.420 20.390 ;
        RECT 1983.220 2.400 1983.360 20.070 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1699.310 587.080 1699.630 587.140 ;
        RECT 1714.490 587.080 1714.810 587.140 ;
        RECT 1699.310 586.940 1714.810 587.080 ;
        RECT 1699.310 586.880 1699.630 586.940 ;
        RECT 1714.490 586.880 1714.810 586.940 ;
        RECT 1973.010 19.620 1973.330 19.680 ;
        RECT 1980.370 19.620 1980.690 19.680 ;
        RECT 1973.010 19.480 1980.690 19.620 ;
        RECT 1973.010 19.420 1973.330 19.480 ;
        RECT 1980.370 19.420 1980.690 19.480 ;
        RECT 1714.490 18.940 1714.810 19.000 ;
        RECT 1925.170 18.940 1925.490 19.000 ;
        RECT 1714.490 18.800 1925.490 18.940 ;
        RECT 1714.490 18.740 1714.810 18.800 ;
        RECT 1925.170 18.740 1925.490 18.800 ;
        RECT 1980.370 18.940 1980.690 19.000 ;
        RECT 2001.070 18.940 2001.390 19.000 ;
        RECT 1980.370 18.800 2001.390 18.940 ;
        RECT 1980.370 18.740 1980.690 18.800 ;
        RECT 2001.070 18.740 2001.390 18.800 ;
      LAYER via ;
        RECT 1699.340 586.880 1699.600 587.140 ;
        RECT 1714.520 586.880 1714.780 587.140 ;
        RECT 1973.040 19.420 1973.300 19.680 ;
        RECT 1980.400 19.420 1980.660 19.680 ;
        RECT 1714.520 18.740 1714.780 19.000 ;
        RECT 1925.200 18.740 1925.460 19.000 ;
        RECT 1980.400 18.740 1980.660 19.000 ;
        RECT 2001.100 18.740 2001.360 19.000 ;
      LAYER met2 ;
        RECT 1697.730 600.170 1698.010 604.000 ;
        RECT 1697.730 600.030 1699.540 600.170 ;
        RECT 1697.730 600.000 1698.010 600.030 ;
        RECT 1699.400 587.170 1699.540 600.030 ;
        RECT 1699.340 586.850 1699.600 587.170 ;
        RECT 1714.520 586.850 1714.780 587.170 ;
        RECT 1714.580 19.030 1714.720 586.850 ;
        RECT 1972.180 19.990 1973.240 20.130 ;
        RECT 1714.520 18.710 1714.780 19.030 ;
        RECT 1925.200 18.885 1925.460 19.030 ;
        RECT 1972.180 18.885 1972.320 19.990 ;
        RECT 1973.100 19.710 1973.240 19.990 ;
        RECT 1973.040 19.390 1973.300 19.710 ;
        RECT 1980.400 19.390 1980.660 19.710 ;
        RECT 1980.460 19.030 1980.600 19.390 ;
        RECT 1925.190 18.515 1925.470 18.885 ;
        RECT 1972.110 18.515 1972.390 18.885 ;
        RECT 1980.400 18.710 1980.660 19.030 ;
        RECT 2001.100 18.710 2001.360 19.030 ;
        RECT 2001.160 2.400 2001.300 18.710 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
      LAYER via2 ;
        RECT 1925.190 18.560 1925.470 18.840 ;
        RECT 1972.110 18.560 1972.390 18.840 ;
      LAYER met3 ;
        RECT 1925.165 18.850 1925.495 18.865 ;
        RECT 1972.085 18.850 1972.415 18.865 ;
        RECT 1925.165 18.550 1972.415 18.850 ;
        RECT 1925.165 18.535 1925.495 18.550 ;
        RECT 1972.085 18.535 1972.415 18.550 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1787.260 590.000 1801.200 590.140 ;
        RECT 1708.510 589.460 1708.830 589.520 ;
        RECT 1738.870 589.460 1739.190 589.520 ;
        RECT 1708.510 589.320 1739.190 589.460 ;
        RECT 1708.510 589.260 1708.830 589.320 ;
        RECT 1738.870 589.260 1739.190 589.320 ;
        RECT 1786.710 589.460 1787.030 589.520 ;
        RECT 1787.260 589.460 1787.400 590.000 ;
        RECT 1801.060 589.800 1801.200 590.000 ;
        RECT 1909.530 589.800 1909.850 589.860 ;
        RECT 1801.060 589.660 1909.850 589.800 ;
        RECT 1909.530 589.600 1909.850 589.660 ;
        RECT 1786.710 589.320 1787.400 589.460 ;
        RECT 1786.710 589.260 1787.030 589.320 ;
        RECT 1945.870 589.120 1946.190 589.180 ;
        RECT 2014.870 589.120 2015.190 589.180 ;
        RECT 1945.870 588.980 2015.190 589.120 ;
        RECT 1945.870 588.920 1946.190 588.980 ;
        RECT 2014.870 588.920 2015.190 588.980 ;
        RECT 1909.530 588.440 1909.850 588.500 ;
        RECT 1945.870 588.440 1946.190 588.500 ;
        RECT 1909.530 588.300 1946.190 588.440 ;
        RECT 1909.530 588.240 1909.850 588.300 ;
        RECT 1945.870 588.240 1946.190 588.300 ;
        RECT 2014.870 2.960 2015.190 3.020 ;
        RECT 2018.550 2.960 2018.870 3.020 ;
        RECT 2014.870 2.820 2018.870 2.960 ;
        RECT 2014.870 2.760 2015.190 2.820 ;
        RECT 2018.550 2.760 2018.870 2.820 ;
      LAYER via ;
        RECT 1708.540 589.260 1708.800 589.520 ;
        RECT 1738.900 589.260 1739.160 589.520 ;
        RECT 1786.740 589.260 1787.000 589.520 ;
        RECT 1909.560 589.600 1909.820 589.860 ;
        RECT 1945.900 588.920 1946.160 589.180 ;
        RECT 2014.900 588.920 2015.160 589.180 ;
        RECT 1909.560 588.240 1909.820 588.500 ;
        RECT 1945.900 588.240 1946.160 588.500 ;
        RECT 2014.900 2.760 2015.160 3.020 ;
        RECT 2018.580 2.760 2018.840 3.020 ;
      LAYER met2 ;
        RECT 1706.930 600.170 1707.210 604.000 ;
        RECT 1706.930 600.030 1708.740 600.170 ;
        RECT 1706.930 600.000 1707.210 600.030 ;
        RECT 1708.600 589.550 1708.740 600.030 ;
        RECT 1909.560 589.570 1909.820 589.890 ;
        RECT 1708.540 589.230 1708.800 589.550 ;
        RECT 1738.900 589.405 1739.160 589.550 ;
        RECT 1786.740 589.405 1787.000 589.550 ;
        RECT 1738.890 589.035 1739.170 589.405 ;
        RECT 1786.730 589.035 1787.010 589.405 ;
        RECT 1909.620 588.530 1909.760 589.570 ;
        RECT 1945.900 588.890 1946.160 589.210 ;
        RECT 2014.900 588.890 2015.160 589.210 ;
        RECT 1945.960 588.530 1946.100 588.890 ;
        RECT 1909.560 588.210 1909.820 588.530 ;
        RECT 1945.900 588.210 1946.160 588.530 ;
        RECT 2014.960 3.050 2015.100 588.890 ;
        RECT 2014.900 2.730 2015.160 3.050 ;
        RECT 2018.580 2.730 2018.840 3.050 ;
        RECT 2018.640 2.400 2018.780 2.730 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
      LAYER via2 ;
        RECT 1738.890 589.080 1739.170 589.360 ;
        RECT 1786.730 589.080 1787.010 589.360 ;
      LAYER met3 ;
        RECT 1738.865 589.370 1739.195 589.385 ;
        RECT 1786.705 589.370 1787.035 589.385 ;
        RECT 1738.865 589.070 1787.035 589.370 ;
        RECT 1738.865 589.055 1739.195 589.070 ;
        RECT 1786.705 589.055 1787.035 589.070 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1717.710 592.180 1718.030 592.240 ;
        RECT 1728.290 592.180 1728.610 592.240 ;
        RECT 1717.710 592.040 1728.610 592.180 ;
        RECT 1717.710 591.980 1718.030 592.040 ;
        RECT 1728.290 591.980 1728.610 592.040 ;
        RECT 1728.290 18.600 1728.610 18.660 ;
        RECT 2036.490 18.600 2036.810 18.660 ;
        RECT 1728.290 18.460 2036.810 18.600 ;
        RECT 1728.290 18.400 1728.610 18.460 ;
        RECT 2036.490 18.400 2036.810 18.460 ;
      LAYER via ;
        RECT 1717.740 591.980 1718.000 592.240 ;
        RECT 1728.320 591.980 1728.580 592.240 ;
        RECT 1728.320 18.400 1728.580 18.660 ;
        RECT 2036.520 18.400 2036.780 18.660 ;
      LAYER met2 ;
        RECT 1716.130 600.170 1716.410 604.000 ;
        RECT 1716.130 600.030 1717.940 600.170 ;
        RECT 1716.130 600.000 1716.410 600.030 ;
        RECT 1717.800 592.270 1717.940 600.030 ;
        RECT 1717.740 591.950 1718.000 592.270 ;
        RECT 1728.320 591.950 1728.580 592.270 ;
        RECT 1728.380 18.690 1728.520 591.950 ;
        RECT 1728.320 18.370 1728.580 18.690 ;
        RECT 2036.520 18.370 2036.780 18.690 ;
        RECT 2036.580 2.400 2036.720 18.370 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1726.910 588.780 1727.230 588.840 ;
        RECT 2045.690 588.780 2046.010 588.840 ;
        RECT 1726.910 588.640 2046.010 588.780 ;
        RECT 1726.910 588.580 1727.230 588.640 ;
        RECT 2045.690 588.580 2046.010 588.640 ;
        RECT 2045.690 19.280 2046.010 19.340 ;
        RECT 2054.430 19.280 2054.750 19.340 ;
        RECT 2045.690 19.140 2054.750 19.280 ;
        RECT 2045.690 19.080 2046.010 19.140 ;
        RECT 2054.430 19.080 2054.750 19.140 ;
      LAYER via ;
        RECT 1726.940 588.580 1727.200 588.840 ;
        RECT 2045.720 588.580 2045.980 588.840 ;
        RECT 2045.720 19.080 2045.980 19.340 ;
        RECT 2054.460 19.080 2054.720 19.340 ;
      LAYER met2 ;
        RECT 1725.330 600.170 1725.610 604.000 ;
        RECT 1725.330 600.030 1727.140 600.170 ;
        RECT 1725.330 600.000 1725.610 600.030 ;
        RECT 1727.000 588.870 1727.140 600.030 ;
        RECT 1726.940 588.550 1727.200 588.870 ;
        RECT 2045.720 588.550 2045.980 588.870 ;
        RECT 2045.780 19.370 2045.920 588.550 ;
        RECT 2045.720 19.050 2045.980 19.370 ;
        RECT 2054.460 19.050 2054.720 19.370 ;
        RECT 2054.520 2.400 2054.660 19.050 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 769.650 30.840 769.970 30.900 ;
        RECT 1063.590 30.840 1063.910 30.900 ;
        RECT 769.650 30.700 1063.910 30.840 ;
        RECT 769.650 30.640 769.970 30.700 ;
        RECT 1063.590 30.640 1063.910 30.700 ;
      LAYER via ;
        RECT 769.680 30.640 769.940 30.900 ;
        RECT 1063.620 30.640 1063.880 30.900 ;
      LAYER met2 ;
        RECT 1065.230 600.170 1065.510 604.000 ;
        RECT 1063.680 600.030 1065.510 600.170 ;
        RECT 1063.680 30.930 1063.820 600.030 ;
        RECT 1065.230 600.000 1065.510 600.030 ;
        RECT 769.680 30.610 769.940 30.930 ;
        RECT 1063.620 30.610 1063.880 30.930 ;
        RECT 769.740 2.400 769.880 30.610 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1736.110 586.740 1736.430 586.800 ;
        RECT 1741.170 586.740 1741.490 586.800 ;
        RECT 1736.110 586.600 1741.490 586.740 ;
        RECT 1736.110 586.540 1736.430 586.600 ;
        RECT 1741.170 586.540 1741.490 586.600 ;
        RECT 1740.250 572.460 1740.570 572.520 ;
        RECT 1741.170 572.460 1741.490 572.520 ;
        RECT 1740.250 572.320 1741.490 572.460 ;
        RECT 1740.250 572.260 1740.570 572.320 ;
        RECT 1741.170 572.260 1741.490 572.320 ;
        RECT 1740.250 524.520 1740.570 524.580 ;
        RECT 1742.090 524.520 1742.410 524.580 ;
        RECT 1740.250 524.380 1742.410 524.520 ;
        RECT 1740.250 524.320 1740.570 524.380 ;
        RECT 1742.090 524.320 1742.410 524.380 ;
        RECT 1740.710 476.580 1741.030 476.640 ;
        RECT 1743.470 476.580 1743.790 476.640 ;
        RECT 1740.710 476.440 1743.790 476.580 ;
        RECT 1740.710 476.380 1741.030 476.440 ;
        RECT 1743.470 476.380 1743.790 476.440 ;
        RECT 1740.710 475.900 1741.030 475.960 ;
        RECT 1741.170 475.900 1741.490 475.960 ;
        RECT 1740.710 475.760 1741.490 475.900 ;
        RECT 1740.710 475.700 1741.030 475.760 ;
        RECT 1741.170 475.700 1741.490 475.760 ;
        RECT 1740.710 434.760 1741.030 434.820 ;
        RECT 1741.170 434.760 1741.490 434.820 ;
        RECT 1740.710 434.620 1741.490 434.760 ;
        RECT 1740.710 434.560 1741.030 434.620 ;
        RECT 1741.170 434.560 1741.490 434.620 ;
        RECT 1741.170 427.420 1741.490 427.680 ;
        RECT 1740.710 427.280 1741.030 427.340 ;
        RECT 1741.260 427.280 1741.400 427.420 ;
        RECT 1740.710 427.140 1741.400 427.280 ;
        RECT 1740.710 427.080 1741.030 427.140 ;
        RECT 1740.710 399.400 1741.030 399.460 ;
        RECT 1742.090 399.400 1742.410 399.460 ;
        RECT 1740.710 399.260 1742.410 399.400 ;
        RECT 1740.710 399.200 1741.030 399.260 ;
        RECT 1742.090 399.200 1742.410 399.260 ;
        RECT 1740.710 379.340 1741.030 379.400 ;
        RECT 1742.090 379.340 1742.410 379.400 ;
        RECT 1740.710 379.200 1742.410 379.340 ;
        RECT 1740.710 379.140 1741.030 379.200 ;
        RECT 1742.090 379.140 1742.410 379.200 ;
        RECT 1740.710 331.400 1741.030 331.460 ;
        RECT 1741.170 331.400 1741.490 331.460 ;
        RECT 1740.710 331.260 1741.490 331.400 ;
        RECT 1740.710 331.200 1741.030 331.260 ;
        RECT 1741.170 331.200 1741.490 331.260 ;
        RECT 1740.710 289.580 1741.030 289.640 ;
        RECT 1742.090 289.580 1742.410 289.640 ;
        RECT 1740.710 289.440 1742.410 289.580 ;
        RECT 1740.710 289.380 1741.030 289.440 ;
        RECT 1742.090 289.380 1742.410 289.440 ;
        RECT 1740.710 241.640 1741.030 241.700 ;
        RECT 1741.170 241.640 1741.490 241.700 ;
        RECT 1740.710 241.500 1741.490 241.640 ;
        RECT 1740.710 241.440 1741.030 241.500 ;
        RECT 1741.170 241.440 1741.490 241.500 ;
        RECT 1740.710 193.020 1741.030 193.080 ;
        RECT 1742.090 193.020 1742.410 193.080 ;
        RECT 1740.710 192.880 1742.410 193.020 ;
        RECT 1740.710 192.820 1741.030 192.880 ;
        RECT 1742.090 192.820 1742.410 192.880 ;
        RECT 1740.710 145.080 1741.030 145.140 ;
        RECT 1741.170 145.080 1741.490 145.140 ;
        RECT 1740.710 144.940 1741.490 145.080 ;
        RECT 1740.710 144.880 1741.030 144.940 ;
        RECT 1741.170 144.880 1741.490 144.940 ;
        RECT 1742.090 96.460 1742.410 96.520 ;
        RECT 1743.010 96.460 1743.330 96.520 ;
        RECT 1742.090 96.320 1743.330 96.460 ;
        RECT 1742.090 96.260 1742.410 96.320 ;
        RECT 1743.010 96.260 1743.330 96.320 ;
        RECT 1743.010 17.920 1743.330 17.980 ;
        RECT 2031.430 17.920 2031.750 17.980 ;
        RECT 1743.010 17.780 2031.750 17.920 ;
        RECT 1743.010 17.720 1743.330 17.780 ;
        RECT 2031.430 17.720 2031.750 17.780 ;
        RECT 2031.430 10.780 2031.750 10.840 ;
        RECT 2072.370 10.780 2072.690 10.840 ;
        RECT 2031.430 10.640 2072.690 10.780 ;
        RECT 2031.430 10.580 2031.750 10.640 ;
        RECT 2072.370 10.580 2072.690 10.640 ;
      LAYER via ;
        RECT 1736.140 586.540 1736.400 586.800 ;
        RECT 1741.200 586.540 1741.460 586.800 ;
        RECT 1740.280 572.260 1740.540 572.520 ;
        RECT 1741.200 572.260 1741.460 572.520 ;
        RECT 1740.280 524.320 1740.540 524.580 ;
        RECT 1742.120 524.320 1742.380 524.580 ;
        RECT 1740.740 476.380 1741.000 476.640 ;
        RECT 1743.500 476.380 1743.760 476.640 ;
        RECT 1740.740 475.700 1741.000 475.960 ;
        RECT 1741.200 475.700 1741.460 475.960 ;
        RECT 1740.740 434.560 1741.000 434.820 ;
        RECT 1741.200 434.560 1741.460 434.820 ;
        RECT 1741.200 427.420 1741.460 427.680 ;
        RECT 1740.740 427.080 1741.000 427.340 ;
        RECT 1740.740 399.200 1741.000 399.460 ;
        RECT 1742.120 399.200 1742.380 399.460 ;
        RECT 1740.740 379.140 1741.000 379.400 ;
        RECT 1742.120 379.140 1742.380 379.400 ;
        RECT 1740.740 331.200 1741.000 331.460 ;
        RECT 1741.200 331.200 1741.460 331.460 ;
        RECT 1740.740 289.380 1741.000 289.640 ;
        RECT 1742.120 289.380 1742.380 289.640 ;
        RECT 1740.740 241.440 1741.000 241.700 ;
        RECT 1741.200 241.440 1741.460 241.700 ;
        RECT 1740.740 192.820 1741.000 193.080 ;
        RECT 1742.120 192.820 1742.380 193.080 ;
        RECT 1740.740 144.880 1741.000 145.140 ;
        RECT 1741.200 144.880 1741.460 145.140 ;
        RECT 1742.120 96.260 1742.380 96.520 ;
        RECT 1743.040 96.260 1743.300 96.520 ;
        RECT 1743.040 17.720 1743.300 17.980 ;
        RECT 2031.460 17.720 2031.720 17.980 ;
        RECT 2031.460 10.580 2031.720 10.840 ;
        RECT 2072.400 10.580 2072.660 10.840 ;
      LAYER met2 ;
        RECT 1734.530 600.170 1734.810 604.000 ;
        RECT 1734.530 600.030 1736.340 600.170 ;
        RECT 1734.530 600.000 1734.810 600.030 ;
        RECT 1736.200 586.830 1736.340 600.030 ;
        RECT 1736.140 586.510 1736.400 586.830 ;
        RECT 1741.200 586.510 1741.460 586.830 ;
        RECT 1741.260 572.550 1741.400 586.510 ;
        RECT 1740.280 572.230 1740.540 572.550 ;
        RECT 1741.200 572.230 1741.460 572.550 ;
        RECT 1740.340 524.610 1740.480 572.230 ;
        RECT 1740.280 524.290 1740.540 524.610 ;
        RECT 1742.120 524.290 1742.380 524.610 ;
        RECT 1742.180 524.125 1742.320 524.290 ;
        RECT 1742.110 523.755 1742.390 524.125 ;
        RECT 1743.490 523.755 1743.770 524.125 ;
        RECT 1743.560 476.670 1743.700 523.755 ;
        RECT 1740.740 476.350 1741.000 476.670 ;
        RECT 1743.500 476.350 1743.760 476.670 ;
        RECT 1740.800 475.990 1740.940 476.350 ;
        RECT 1740.740 475.670 1741.000 475.990 ;
        RECT 1741.200 475.670 1741.460 475.990 ;
        RECT 1741.260 434.850 1741.400 475.670 ;
        RECT 1740.740 434.530 1741.000 434.850 ;
        RECT 1741.200 434.530 1741.460 434.850 ;
        RECT 1740.800 428.130 1740.940 434.530 ;
        RECT 1740.800 427.990 1741.400 428.130 ;
        RECT 1741.260 427.710 1741.400 427.990 ;
        RECT 1741.200 427.390 1741.460 427.710 ;
        RECT 1740.740 427.050 1741.000 427.370 ;
        RECT 1740.800 399.490 1740.940 427.050 ;
        RECT 1740.740 399.170 1741.000 399.490 ;
        RECT 1742.120 399.170 1742.380 399.490 ;
        RECT 1742.180 379.430 1742.320 399.170 ;
        RECT 1740.740 379.110 1741.000 379.430 ;
        RECT 1742.120 379.110 1742.380 379.430 ;
        RECT 1740.800 331.490 1740.940 379.110 ;
        RECT 1740.740 331.170 1741.000 331.490 ;
        RECT 1741.200 331.170 1741.460 331.490 ;
        RECT 1741.260 303.690 1741.400 331.170 ;
        RECT 1741.260 303.550 1742.320 303.690 ;
        RECT 1742.180 289.670 1742.320 303.550 ;
        RECT 1740.740 289.350 1741.000 289.670 ;
        RECT 1742.120 289.350 1742.380 289.670 ;
        RECT 1740.800 241.730 1740.940 289.350 ;
        RECT 1740.740 241.410 1741.000 241.730 ;
        RECT 1741.200 241.410 1741.460 241.730 ;
        RECT 1741.260 207.130 1741.400 241.410 ;
        RECT 1741.260 206.990 1742.320 207.130 ;
        RECT 1742.180 193.110 1742.320 206.990 ;
        RECT 1740.740 192.790 1741.000 193.110 ;
        RECT 1742.120 192.790 1742.380 193.110 ;
        RECT 1740.800 145.170 1740.940 192.790 ;
        RECT 1740.740 144.850 1741.000 145.170 ;
        RECT 1741.200 144.850 1741.460 145.170 ;
        RECT 1741.260 110.570 1741.400 144.850 ;
        RECT 1741.260 110.430 1742.320 110.570 ;
        RECT 1742.180 96.550 1742.320 110.430 ;
        RECT 1742.120 96.230 1742.380 96.550 ;
        RECT 1743.040 96.230 1743.300 96.550 ;
        RECT 1743.100 18.010 1743.240 96.230 ;
        RECT 1743.040 17.690 1743.300 18.010 ;
        RECT 2031.460 17.690 2031.720 18.010 ;
        RECT 2031.520 10.870 2031.660 17.690 ;
        RECT 2031.460 10.550 2031.720 10.870 ;
        RECT 2072.400 10.550 2072.660 10.870 ;
        RECT 2072.460 2.400 2072.600 10.550 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
      LAYER via2 ;
        RECT 1742.110 523.800 1742.390 524.080 ;
        RECT 1743.490 523.800 1743.770 524.080 ;
      LAYER met3 ;
        RECT 1742.085 524.090 1742.415 524.105 ;
        RECT 1743.465 524.090 1743.795 524.105 ;
        RECT 1742.085 523.790 1743.795 524.090 ;
        RECT 1742.085 523.775 1742.415 523.790 ;
        RECT 1743.465 523.775 1743.795 523.790 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1745.310 592.860 1745.630 592.920 ;
        RECT 2080.190 592.860 2080.510 592.920 ;
        RECT 1745.310 592.720 2080.510 592.860 ;
        RECT 1745.310 592.660 1745.630 592.720 ;
        RECT 2080.190 592.660 2080.510 592.720 ;
        RECT 2080.190 19.280 2080.510 19.340 ;
        RECT 2089.850 19.280 2090.170 19.340 ;
        RECT 2080.190 19.140 2090.170 19.280 ;
        RECT 2080.190 19.080 2080.510 19.140 ;
        RECT 2089.850 19.080 2090.170 19.140 ;
      LAYER via ;
        RECT 1745.340 592.660 1745.600 592.920 ;
        RECT 2080.220 592.660 2080.480 592.920 ;
        RECT 2080.220 19.080 2080.480 19.340 ;
        RECT 2089.880 19.080 2090.140 19.340 ;
      LAYER met2 ;
        RECT 1743.730 600.170 1744.010 604.000 ;
        RECT 1743.730 600.030 1745.540 600.170 ;
        RECT 1743.730 600.000 1744.010 600.030 ;
        RECT 1745.400 592.950 1745.540 600.030 ;
        RECT 1745.340 592.630 1745.600 592.950 ;
        RECT 2080.220 592.630 2080.480 592.950 ;
        RECT 2080.280 19.370 2080.420 592.630 ;
        RECT 2080.220 19.050 2080.480 19.370 ;
        RECT 2089.880 19.050 2090.140 19.370 ;
        RECT 2089.940 2.400 2090.080 19.050 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1754.510 587.080 1754.830 587.140 ;
        RECT 1762.790 587.080 1763.110 587.140 ;
        RECT 1754.510 586.940 1763.110 587.080 ;
        RECT 1754.510 586.880 1754.830 586.940 ;
        RECT 1762.790 586.880 1763.110 586.940 ;
        RECT 2042.930 17.920 2043.250 17.980 ;
        RECT 2107.790 17.920 2108.110 17.980 ;
        RECT 2042.930 17.780 2108.110 17.920 ;
        RECT 2042.930 17.720 2043.250 17.780 ;
        RECT 2107.790 17.720 2108.110 17.780 ;
        RECT 1762.330 17.580 1762.650 17.640 ;
        RECT 2028.670 17.580 2028.990 17.640 ;
        RECT 1762.330 17.440 2028.990 17.580 ;
        RECT 1762.330 17.380 1762.650 17.440 ;
        RECT 2028.670 17.380 2028.990 17.440 ;
      LAYER via ;
        RECT 1754.540 586.880 1754.800 587.140 ;
        RECT 1762.820 586.880 1763.080 587.140 ;
        RECT 2042.960 17.720 2043.220 17.980 ;
        RECT 2107.820 17.720 2108.080 17.980 ;
        RECT 1762.360 17.380 1762.620 17.640 ;
        RECT 2028.700 17.380 2028.960 17.640 ;
      LAYER met2 ;
        RECT 1752.930 600.170 1753.210 604.000 ;
        RECT 1752.930 600.030 1754.740 600.170 ;
        RECT 1752.930 600.000 1753.210 600.030 ;
        RECT 1754.600 587.170 1754.740 600.030 ;
        RECT 1754.540 586.850 1754.800 587.170 ;
        RECT 1762.820 586.850 1763.080 587.170 ;
        RECT 1762.880 39.850 1763.020 586.850 ;
        RECT 1762.420 39.710 1763.020 39.850 ;
        RECT 1762.420 17.670 1762.560 39.710 ;
        RECT 2028.690 17.835 2028.970 18.205 ;
        RECT 2042.950 17.835 2043.230 18.205 ;
        RECT 2028.760 17.670 2028.900 17.835 ;
        RECT 2042.960 17.690 2043.220 17.835 ;
        RECT 2107.820 17.690 2108.080 18.010 ;
        RECT 1762.360 17.350 1762.620 17.670 ;
        RECT 2028.700 17.350 2028.960 17.670 ;
        RECT 2107.880 2.400 2108.020 17.690 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
      LAYER via2 ;
        RECT 2028.690 17.880 2028.970 18.160 ;
        RECT 2042.950 17.880 2043.230 18.160 ;
      LAYER met3 ;
        RECT 2028.665 18.170 2028.995 18.185 ;
        RECT 2042.925 18.170 2043.255 18.185 ;
        RECT 2028.665 17.870 2043.255 18.170 ;
        RECT 2028.665 17.855 2028.995 17.870 ;
        RECT 2042.925 17.855 2043.255 17.870 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1763.710 592.520 1764.030 592.580 ;
        RECT 2121.590 592.520 2121.910 592.580 ;
        RECT 1763.710 592.380 2121.910 592.520 ;
        RECT 1763.710 592.320 1764.030 592.380 ;
        RECT 2121.590 592.320 2121.910 592.380 ;
        RECT 2121.590 18.600 2121.910 18.660 ;
        RECT 2125.730 18.600 2126.050 18.660 ;
        RECT 2121.590 18.460 2126.050 18.600 ;
        RECT 2121.590 18.400 2121.910 18.460 ;
        RECT 2125.730 18.400 2126.050 18.460 ;
      LAYER via ;
        RECT 1763.740 592.320 1764.000 592.580 ;
        RECT 2121.620 592.320 2121.880 592.580 ;
        RECT 2121.620 18.400 2121.880 18.660 ;
        RECT 2125.760 18.400 2126.020 18.660 ;
      LAYER met2 ;
        RECT 1762.130 600.170 1762.410 604.000 ;
        RECT 1762.130 600.030 1763.940 600.170 ;
        RECT 1762.130 600.000 1762.410 600.030 ;
        RECT 1763.800 592.610 1763.940 600.030 ;
        RECT 1763.740 592.290 1764.000 592.610 ;
        RECT 2121.620 592.290 2121.880 592.610 ;
        RECT 2121.680 18.690 2121.820 592.290 ;
        RECT 2121.620 18.370 2121.880 18.690 ;
        RECT 2125.760 18.370 2126.020 18.690 ;
        RECT 2125.820 2.400 2125.960 18.370 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.450 586.740 1772.770 586.800 ;
        RECT 1783.490 586.740 1783.810 586.800 ;
        RECT 1772.450 586.600 1783.810 586.740 ;
        RECT 1772.450 586.540 1772.770 586.600 ;
        RECT 1783.490 586.540 1783.810 586.600 ;
        RECT 1783.490 17.240 1783.810 17.300 ;
        RECT 2143.670 17.240 2143.990 17.300 ;
        RECT 1783.490 17.100 2143.990 17.240 ;
        RECT 1783.490 17.040 1783.810 17.100 ;
        RECT 2143.670 17.040 2143.990 17.100 ;
      LAYER via ;
        RECT 1772.480 586.540 1772.740 586.800 ;
        RECT 1783.520 586.540 1783.780 586.800 ;
        RECT 1783.520 17.040 1783.780 17.300 ;
        RECT 2143.700 17.040 2143.960 17.300 ;
      LAYER met2 ;
        RECT 1770.870 600.170 1771.150 604.000 ;
        RECT 1770.870 600.030 1772.680 600.170 ;
        RECT 1770.870 600.000 1771.150 600.030 ;
        RECT 1772.540 586.830 1772.680 600.030 ;
        RECT 1772.480 586.510 1772.740 586.830 ;
        RECT 1783.520 586.510 1783.780 586.830 ;
        RECT 1783.580 17.330 1783.720 586.510 ;
        RECT 1783.520 17.010 1783.780 17.330 ;
        RECT 2143.700 17.010 2143.960 17.330 ;
        RECT 2143.760 2.400 2143.900 17.010 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1781.650 592.180 1781.970 592.240 ;
        RECT 1921.030 592.180 1921.350 592.240 ;
        RECT 1781.650 592.040 1921.350 592.180 ;
        RECT 1781.650 591.980 1781.970 592.040 ;
        RECT 1921.030 591.980 1921.350 592.040 ;
        RECT 1969.790 592.180 1970.110 592.240 ;
        RECT 2018.090 592.180 2018.410 592.240 ;
        RECT 1969.790 592.040 2018.410 592.180 ;
        RECT 1969.790 591.980 1970.110 592.040 ;
        RECT 2018.090 591.980 2018.410 592.040 ;
        RECT 2066.390 592.180 2066.710 592.240 ;
        RECT 2149.190 592.180 2149.510 592.240 ;
        RECT 2066.390 592.040 2149.510 592.180 ;
        RECT 2066.390 591.980 2066.710 592.040 ;
        RECT 2149.190 591.980 2149.510 592.040 ;
        RECT 2018.090 589.120 2018.410 589.180 ;
        RECT 2066.390 589.120 2066.710 589.180 ;
        RECT 2018.090 588.980 2066.710 589.120 ;
        RECT 2018.090 588.920 2018.410 588.980 ;
        RECT 2066.390 588.920 2066.710 588.980 ;
        RECT 1921.030 587.760 1921.350 587.820 ;
        RECT 1969.790 587.760 1970.110 587.820 ;
        RECT 1921.030 587.620 1970.110 587.760 ;
        RECT 1921.030 587.560 1921.350 587.620 ;
        RECT 1969.790 587.560 1970.110 587.620 ;
        RECT 2149.190 18.260 2149.510 18.320 ;
        RECT 2161.610 18.260 2161.930 18.320 ;
        RECT 2149.190 18.120 2161.930 18.260 ;
        RECT 2149.190 18.060 2149.510 18.120 ;
        RECT 2161.610 18.060 2161.930 18.120 ;
      LAYER via ;
        RECT 1781.680 591.980 1781.940 592.240 ;
        RECT 1921.060 591.980 1921.320 592.240 ;
        RECT 1969.820 591.980 1970.080 592.240 ;
        RECT 2018.120 591.980 2018.380 592.240 ;
        RECT 2066.420 591.980 2066.680 592.240 ;
        RECT 2149.220 591.980 2149.480 592.240 ;
        RECT 2018.120 588.920 2018.380 589.180 ;
        RECT 2066.420 588.920 2066.680 589.180 ;
        RECT 1921.060 587.560 1921.320 587.820 ;
        RECT 1969.820 587.560 1970.080 587.820 ;
        RECT 2149.220 18.060 2149.480 18.320 ;
        RECT 2161.640 18.060 2161.900 18.320 ;
      LAYER met2 ;
        RECT 1780.070 600.170 1780.350 604.000 ;
        RECT 1780.070 600.030 1781.880 600.170 ;
        RECT 1780.070 600.000 1780.350 600.030 ;
        RECT 1781.740 592.270 1781.880 600.030 ;
        RECT 1781.680 591.950 1781.940 592.270 ;
        RECT 1921.060 591.950 1921.320 592.270 ;
        RECT 1969.820 591.950 1970.080 592.270 ;
        RECT 2018.120 591.950 2018.380 592.270 ;
        RECT 2066.420 591.950 2066.680 592.270 ;
        RECT 2149.220 591.950 2149.480 592.270 ;
        RECT 1921.120 587.850 1921.260 591.950 ;
        RECT 1969.880 587.850 1970.020 591.950 ;
        RECT 2018.180 589.210 2018.320 591.950 ;
        RECT 2066.480 589.210 2066.620 591.950 ;
        RECT 2018.120 588.890 2018.380 589.210 ;
        RECT 2066.420 588.890 2066.680 589.210 ;
        RECT 1921.060 587.530 1921.320 587.850 ;
        RECT 1969.820 587.530 1970.080 587.850 ;
        RECT 2149.280 18.350 2149.420 591.950 ;
        RECT 2149.220 18.030 2149.480 18.350 ;
        RECT 2161.640 18.030 2161.900 18.350 ;
        RECT 2161.700 2.400 2161.840 18.030 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1790.850 587.080 1791.170 587.140 ;
        RECT 1804.190 587.080 1804.510 587.140 ;
        RECT 1790.850 586.940 1804.510 587.080 ;
        RECT 1790.850 586.880 1791.170 586.940 ;
        RECT 1804.190 586.880 1804.510 586.940 ;
        RECT 2044.770 19.280 2045.090 19.340 ;
        RECT 2041.640 19.140 2045.090 19.280 ;
        RECT 1804.190 18.260 1804.510 18.320 ;
        RECT 2041.640 18.260 2041.780 19.140 ;
        RECT 2044.770 19.080 2045.090 19.140 ;
        RECT 1804.190 18.120 2041.780 18.260 ;
        RECT 2044.770 18.260 2045.090 18.320 ;
        RECT 2148.730 18.260 2149.050 18.320 ;
        RECT 2044.770 18.120 2149.050 18.260 ;
        RECT 1804.190 18.060 1804.510 18.120 ;
        RECT 2044.770 18.060 2045.090 18.120 ;
        RECT 2148.730 18.060 2149.050 18.120 ;
        RECT 2148.730 17.240 2149.050 17.300 ;
        RECT 2179.090 17.240 2179.410 17.300 ;
        RECT 2148.730 17.100 2179.410 17.240 ;
        RECT 2148.730 17.040 2149.050 17.100 ;
        RECT 2179.090 17.040 2179.410 17.100 ;
      LAYER via ;
        RECT 1790.880 586.880 1791.140 587.140 ;
        RECT 1804.220 586.880 1804.480 587.140 ;
        RECT 1804.220 18.060 1804.480 18.320 ;
        RECT 2044.800 19.080 2045.060 19.340 ;
        RECT 2044.800 18.060 2045.060 18.320 ;
        RECT 2148.760 18.060 2149.020 18.320 ;
        RECT 2148.760 17.040 2149.020 17.300 ;
        RECT 2179.120 17.040 2179.380 17.300 ;
      LAYER met2 ;
        RECT 1789.270 600.170 1789.550 604.000 ;
        RECT 1789.270 600.030 1791.080 600.170 ;
        RECT 1789.270 600.000 1789.550 600.030 ;
        RECT 1790.940 587.170 1791.080 600.030 ;
        RECT 1790.880 586.850 1791.140 587.170 ;
        RECT 1804.220 586.850 1804.480 587.170 ;
        RECT 1804.280 18.350 1804.420 586.850 ;
        RECT 2044.800 19.050 2045.060 19.370 ;
        RECT 2044.860 18.350 2045.000 19.050 ;
        RECT 1804.220 18.030 1804.480 18.350 ;
        RECT 2044.800 18.030 2045.060 18.350 ;
        RECT 2148.760 18.030 2149.020 18.350 ;
        RECT 2148.820 17.330 2148.960 18.030 ;
        RECT 2148.760 17.010 2149.020 17.330 ;
        RECT 2179.120 17.010 2179.380 17.330 ;
        RECT 2179.180 2.400 2179.320 17.010 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.050 591.840 1800.370 591.900 ;
        RECT 2194.270 591.840 2194.590 591.900 ;
        RECT 1800.050 591.700 2194.590 591.840 ;
        RECT 1800.050 591.640 1800.370 591.700 ;
        RECT 2194.270 591.640 2194.590 591.700 ;
      LAYER via ;
        RECT 1800.080 591.640 1800.340 591.900 ;
        RECT 2194.300 591.640 2194.560 591.900 ;
      LAYER met2 ;
        RECT 1798.470 600.170 1798.750 604.000 ;
        RECT 1798.470 600.030 1800.280 600.170 ;
        RECT 1798.470 600.000 1798.750 600.030 ;
        RECT 1800.140 591.930 1800.280 600.030 ;
        RECT 1800.080 591.610 1800.340 591.930 ;
        RECT 2194.300 591.610 2194.560 591.930 ;
        RECT 2194.360 17.410 2194.500 591.610 ;
        RECT 2194.360 17.270 2197.260 17.410 ;
        RECT 2197.120 2.400 2197.260 17.270 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1809.250 589.460 1809.570 589.520 ;
        RECT 1861.230 589.460 1861.550 589.520 ;
        RECT 1809.250 589.320 1861.550 589.460 ;
        RECT 1809.250 589.260 1809.570 589.320 ;
        RECT 1861.230 589.260 1861.550 589.320 ;
        RECT 1861.230 588.100 1861.550 588.160 ;
        RECT 1873.190 588.100 1873.510 588.160 ;
        RECT 1861.230 587.960 1873.510 588.100 ;
        RECT 1861.230 587.900 1861.550 587.960 ;
        RECT 1873.190 587.900 1873.510 587.960 ;
        RECT 1873.190 15.540 1873.510 15.600 ;
        RECT 2214.970 15.540 2215.290 15.600 ;
        RECT 1873.190 15.400 2215.290 15.540 ;
        RECT 1873.190 15.340 1873.510 15.400 ;
        RECT 2214.970 15.340 2215.290 15.400 ;
      LAYER via ;
        RECT 1809.280 589.260 1809.540 589.520 ;
        RECT 1861.260 589.260 1861.520 589.520 ;
        RECT 1861.260 587.900 1861.520 588.160 ;
        RECT 1873.220 587.900 1873.480 588.160 ;
        RECT 1873.220 15.340 1873.480 15.600 ;
        RECT 2215.000 15.340 2215.260 15.600 ;
      LAYER met2 ;
        RECT 1807.670 600.170 1807.950 604.000 ;
        RECT 1807.670 600.030 1809.480 600.170 ;
        RECT 1807.670 600.000 1807.950 600.030 ;
        RECT 1809.340 589.550 1809.480 600.030 ;
        RECT 1809.280 589.230 1809.540 589.550 ;
        RECT 1861.260 589.230 1861.520 589.550 ;
        RECT 1861.320 588.190 1861.460 589.230 ;
        RECT 1861.260 587.870 1861.520 588.190 ;
        RECT 1873.220 587.870 1873.480 588.190 ;
        RECT 1873.280 15.630 1873.420 587.870 ;
        RECT 1873.220 15.310 1873.480 15.630 ;
        RECT 2215.000 15.310 2215.260 15.630 ;
        RECT 2215.060 2.400 2215.200 15.310 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1818.450 591.500 1818.770 591.560 ;
        RECT 2228.770 591.500 2229.090 591.560 ;
        RECT 1818.450 591.360 2229.090 591.500 ;
        RECT 1818.450 591.300 1818.770 591.360 ;
        RECT 2228.770 591.300 2229.090 591.360 ;
      LAYER via ;
        RECT 1818.480 591.300 1818.740 591.560 ;
        RECT 2228.800 591.300 2229.060 591.560 ;
      LAYER met2 ;
        RECT 1816.870 600.170 1817.150 604.000 ;
        RECT 1816.870 600.030 1818.680 600.170 ;
        RECT 1816.870 600.000 1817.150 600.030 ;
        RECT 1818.540 591.590 1818.680 600.030 ;
        RECT 1818.480 591.270 1818.740 591.590 ;
        RECT 2228.800 591.270 2229.060 591.590 ;
        RECT 2228.860 17.410 2229.000 591.270 ;
        RECT 2228.860 17.270 2233.140 17.410 ;
        RECT 2233.000 2.400 2233.140 17.270 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1069.110 469.100 1069.430 469.160 ;
        RECT 1070.030 469.100 1070.350 469.160 ;
        RECT 1069.110 468.960 1070.350 469.100 ;
        RECT 1069.110 468.900 1069.430 468.960 ;
        RECT 1070.030 468.900 1070.350 468.960 ;
        RECT 1069.110 421.160 1069.430 421.220 ;
        RECT 1070.490 421.160 1070.810 421.220 ;
        RECT 1069.110 421.020 1070.810 421.160 ;
        RECT 1069.110 420.960 1069.430 421.020 ;
        RECT 1070.490 420.960 1070.810 421.020 ;
        RECT 1070.950 373.220 1071.270 373.280 ;
        RECT 1070.120 373.080 1071.270 373.220 ;
        RECT 1070.120 372.940 1070.260 373.080 ;
        RECT 1070.950 373.020 1071.270 373.080 ;
        RECT 1070.030 372.680 1070.350 372.940 ;
        RECT 787.590 31.520 787.910 31.580 ;
        RECT 1070.490 31.520 1070.810 31.580 ;
        RECT 787.590 31.380 1070.810 31.520 ;
        RECT 787.590 31.320 787.910 31.380 ;
        RECT 1070.490 31.320 1070.810 31.380 ;
      LAYER via ;
        RECT 1069.140 468.900 1069.400 469.160 ;
        RECT 1070.060 468.900 1070.320 469.160 ;
        RECT 1069.140 420.960 1069.400 421.220 ;
        RECT 1070.520 420.960 1070.780 421.220 ;
        RECT 1070.980 373.020 1071.240 373.280 ;
        RECT 1070.060 372.680 1070.320 372.940 ;
        RECT 787.620 31.320 787.880 31.580 ;
        RECT 1070.520 31.320 1070.780 31.580 ;
      LAYER met2 ;
        RECT 1074.430 601.530 1074.710 604.000 ;
        RECT 1072.880 601.390 1074.710 601.530 ;
        RECT 1072.880 579.770 1073.020 601.390 ;
        RECT 1074.430 600.000 1074.710 601.390 ;
        RECT 1072.420 579.630 1073.020 579.770 ;
        RECT 1072.420 470.405 1072.560 579.630 ;
        RECT 1072.350 470.035 1072.630 470.405 ;
        RECT 1070.050 469.355 1070.330 469.725 ;
        RECT 1070.120 469.190 1070.260 469.355 ;
        RECT 1069.140 468.870 1069.400 469.190 ;
        RECT 1070.060 468.870 1070.320 469.190 ;
        RECT 1069.200 421.250 1069.340 468.870 ;
        RECT 1069.140 420.930 1069.400 421.250 ;
        RECT 1070.520 420.930 1070.780 421.250 ;
        RECT 1070.580 420.650 1070.720 420.930 ;
        RECT 1070.580 420.510 1071.180 420.650 ;
        RECT 1071.040 373.310 1071.180 420.510 ;
        RECT 1070.980 372.990 1071.240 373.310 ;
        RECT 1070.060 372.650 1070.320 372.970 ;
        RECT 1070.120 109.890 1070.260 372.650 ;
        RECT 1070.120 109.750 1070.720 109.890 ;
        RECT 1070.580 31.610 1070.720 109.750 ;
        RECT 787.620 31.290 787.880 31.610 ;
        RECT 1070.520 31.290 1070.780 31.610 ;
        RECT 787.680 2.400 787.820 31.290 ;
        RECT 787.470 -4.800 788.030 2.400 ;
      LAYER via2 ;
        RECT 1072.350 470.080 1072.630 470.360 ;
        RECT 1070.050 469.400 1070.330 469.680 ;
      LAYER met3 ;
        RECT 1072.325 470.370 1072.655 470.385 ;
        RECT 1069.350 470.070 1072.655 470.370 ;
        RECT 1069.350 469.690 1069.650 470.070 ;
        RECT 1072.325 470.055 1072.655 470.070 ;
        RECT 1070.025 469.690 1070.355 469.705 ;
        RECT 1069.350 469.390 1070.355 469.690 ;
        RECT 1070.025 469.375 1070.355 469.390 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1827.650 587.080 1827.970 587.140 ;
        RECT 1838.690 587.080 1839.010 587.140 ;
        RECT 1827.650 586.940 1839.010 587.080 ;
        RECT 1827.650 586.880 1827.970 586.940 ;
        RECT 1838.690 586.880 1839.010 586.940 ;
        RECT 1838.690 15.880 1839.010 15.940 ;
        RECT 2250.850 15.880 2251.170 15.940 ;
        RECT 1838.690 15.740 2251.170 15.880 ;
        RECT 1838.690 15.680 1839.010 15.740 ;
        RECT 2250.850 15.680 2251.170 15.740 ;
      LAYER via ;
        RECT 1827.680 586.880 1827.940 587.140 ;
        RECT 1838.720 586.880 1838.980 587.140 ;
        RECT 1838.720 15.680 1838.980 15.940 ;
        RECT 2250.880 15.680 2251.140 15.940 ;
      LAYER met2 ;
        RECT 1826.070 600.170 1826.350 604.000 ;
        RECT 1826.070 600.030 1827.880 600.170 ;
        RECT 1826.070 600.000 1826.350 600.030 ;
        RECT 1827.740 587.170 1827.880 600.030 ;
        RECT 1827.680 586.850 1827.940 587.170 ;
        RECT 1838.720 586.850 1838.980 587.170 ;
        RECT 1838.780 15.970 1838.920 586.850 ;
        RECT 1838.720 15.650 1838.980 15.970 ;
        RECT 2250.880 15.650 2251.140 15.970 ;
        RECT 2250.940 2.400 2251.080 15.650 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1836.850 591.160 1837.170 591.220 ;
        RECT 2264.650 591.160 2264.970 591.220 ;
        RECT 1836.850 591.020 2264.970 591.160 ;
        RECT 1836.850 590.960 1837.170 591.020 ;
        RECT 2264.650 590.960 2264.970 591.020 ;
        RECT 2263.270 586.060 2263.590 586.120 ;
        RECT 2264.650 586.060 2264.970 586.120 ;
        RECT 2263.270 585.920 2264.970 586.060 ;
        RECT 2263.270 585.860 2263.590 585.920 ;
        RECT 2264.650 585.860 2264.970 585.920 ;
        RECT 2263.270 2.960 2263.590 3.020 ;
        RECT 2268.330 2.960 2268.650 3.020 ;
        RECT 2263.270 2.820 2268.650 2.960 ;
        RECT 2263.270 2.760 2263.590 2.820 ;
        RECT 2268.330 2.760 2268.650 2.820 ;
      LAYER via ;
        RECT 1836.880 590.960 1837.140 591.220 ;
        RECT 2264.680 590.960 2264.940 591.220 ;
        RECT 2263.300 585.860 2263.560 586.120 ;
        RECT 2264.680 585.860 2264.940 586.120 ;
        RECT 2263.300 2.760 2263.560 3.020 ;
        RECT 2268.360 2.760 2268.620 3.020 ;
      LAYER met2 ;
        RECT 1835.270 600.170 1835.550 604.000 ;
        RECT 1835.270 600.030 1837.080 600.170 ;
        RECT 1835.270 600.000 1835.550 600.030 ;
        RECT 1836.940 591.250 1837.080 600.030 ;
        RECT 1836.880 590.930 1837.140 591.250 ;
        RECT 2264.680 590.930 2264.940 591.250 ;
        RECT 2264.740 586.150 2264.880 590.930 ;
        RECT 2263.300 585.830 2263.560 586.150 ;
        RECT 2264.680 585.830 2264.940 586.150 ;
        RECT 2263.360 3.050 2263.500 585.830 ;
        RECT 2263.300 2.730 2263.560 3.050 ;
        RECT 2268.360 2.730 2268.620 3.050 ;
        RECT 2268.420 2.400 2268.560 2.730 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1846.050 586.740 1846.370 586.800 ;
        RECT 1848.810 586.740 1849.130 586.800 ;
        RECT 1846.050 586.600 1849.130 586.740 ;
        RECT 1846.050 586.540 1846.370 586.600 ;
        RECT 1848.810 586.540 1849.130 586.600 ;
        RECT 1848.810 16.220 1849.130 16.280 ;
        RECT 2286.270 16.220 2286.590 16.280 ;
        RECT 1848.810 16.080 2286.590 16.220 ;
        RECT 1848.810 16.020 1849.130 16.080 ;
        RECT 2286.270 16.020 2286.590 16.080 ;
      LAYER via ;
        RECT 1846.080 586.540 1846.340 586.800 ;
        RECT 1848.840 586.540 1849.100 586.800 ;
        RECT 1848.840 16.020 1849.100 16.280 ;
        RECT 2286.300 16.020 2286.560 16.280 ;
      LAYER met2 ;
        RECT 1844.470 600.170 1844.750 604.000 ;
        RECT 1844.470 600.030 1846.280 600.170 ;
        RECT 1844.470 600.000 1844.750 600.030 ;
        RECT 1846.140 586.830 1846.280 600.030 ;
        RECT 1846.080 586.510 1846.340 586.830 ;
        RECT 1848.840 586.510 1849.100 586.830 ;
        RECT 1848.900 16.310 1849.040 586.510 ;
        RECT 1848.840 15.990 1849.100 16.310 ;
        RECT 2286.300 15.990 2286.560 16.310 ;
        RECT 2286.360 2.400 2286.500 15.990 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1855.250 590.820 1855.570 590.880 ;
        RECT 2297.770 590.820 2298.090 590.880 ;
        RECT 1855.250 590.680 2298.090 590.820 ;
        RECT 1855.250 590.620 1855.570 590.680 ;
        RECT 2297.770 590.620 2298.090 590.680 ;
        RECT 2297.770 16.220 2298.090 16.280 ;
        RECT 2304.210 16.220 2304.530 16.280 ;
        RECT 2297.770 16.080 2304.530 16.220 ;
        RECT 2297.770 16.020 2298.090 16.080 ;
        RECT 2304.210 16.020 2304.530 16.080 ;
      LAYER via ;
        RECT 1855.280 590.620 1855.540 590.880 ;
        RECT 2297.800 590.620 2298.060 590.880 ;
        RECT 2297.800 16.020 2298.060 16.280 ;
        RECT 2304.240 16.020 2304.500 16.280 ;
      LAYER met2 ;
        RECT 1853.670 600.170 1853.950 604.000 ;
        RECT 1853.670 600.030 1855.480 600.170 ;
        RECT 1853.670 600.000 1853.950 600.030 ;
        RECT 1855.340 590.910 1855.480 600.030 ;
        RECT 1855.280 590.590 1855.540 590.910 ;
        RECT 2297.800 590.590 2298.060 590.910 ;
        RECT 2297.860 16.310 2298.000 590.590 ;
        RECT 2297.800 15.990 2298.060 16.310 ;
        RECT 2304.240 15.990 2304.500 16.310 ;
        RECT 2304.300 2.400 2304.440 15.990 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1864.450 589.460 1864.770 589.520 ;
        RECT 1869.510 589.460 1869.830 589.520 ;
        RECT 1864.450 589.320 1869.830 589.460 ;
        RECT 1864.450 589.260 1864.770 589.320 ;
        RECT 1869.510 589.260 1869.830 589.320 ;
        RECT 1869.510 16.560 1869.830 16.620 ;
        RECT 2322.150 16.560 2322.470 16.620 ;
        RECT 1869.510 16.420 2322.470 16.560 ;
        RECT 1869.510 16.360 1869.830 16.420 ;
        RECT 2322.150 16.360 2322.470 16.420 ;
      LAYER via ;
        RECT 1864.480 589.260 1864.740 589.520 ;
        RECT 1869.540 589.260 1869.800 589.520 ;
        RECT 1869.540 16.360 1869.800 16.620 ;
        RECT 2322.180 16.360 2322.440 16.620 ;
      LAYER met2 ;
        RECT 1862.870 600.170 1863.150 604.000 ;
        RECT 1862.870 600.030 1864.680 600.170 ;
        RECT 1862.870 600.000 1863.150 600.030 ;
        RECT 1864.540 589.550 1864.680 600.030 ;
        RECT 1864.480 589.230 1864.740 589.550 ;
        RECT 1869.540 589.230 1869.800 589.550 ;
        RECT 1869.600 16.650 1869.740 589.230 ;
        RECT 1869.540 16.330 1869.800 16.650 ;
        RECT 2322.180 16.330 2322.440 16.650 ;
        RECT 2322.240 2.400 2322.380 16.330 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1873.650 590.480 1873.970 590.540 ;
        RECT 2339.170 590.480 2339.490 590.540 ;
        RECT 1873.650 590.340 2339.490 590.480 ;
        RECT 1873.650 590.280 1873.970 590.340 ;
        RECT 2339.170 590.280 2339.490 590.340 ;
      LAYER via ;
        RECT 1873.680 590.280 1873.940 590.540 ;
        RECT 2339.200 590.280 2339.460 590.540 ;
      LAYER met2 ;
        RECT 1872.070 600.170 1872.350 604.000 ;
        RECT 1872.070 600.030 1873.880 600.170 ;
        RECT 1872.070 600.000 1872.350 600.030 ;
        RECT 1873.740 590.570 1873.880 600.030 ;
        RECT 1873.680 590.250 1873.940 590.570 ;
        RECT 2339.200 590.250 2339.460 590.570 ;
        RECT 2339.260 17.410 2339.400 590.250 ;
        RECT 2339.260 17.270 2339.860 17.410 ;
        RECT 2339.720 2.400 2339.860 17.270 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1883.310 20.300 1883.630 20.360 ;
        RECT 1921.490 20.300 1921.810 20.360 ;
        RECT 1883.310 20.160 1921.810 20.300 ;
        RECT 1883.310 20.100 1883.630 20.160 ;
        RECT 1921.490 20.100 1921.810 20.160 ;
        RECT 1921.490 16.900 1921.810 16.960 ;
        RECT 2357.570 16.900 2357.890 16.960 ;
        RECT 1921.490 16.760 2357.890 16.900 ;
        RECT 1921.490 16.700 1921.810 16.760 ;
        RECT 2357.570 16.700 2357.890 16.760 ;
      LAYER via ;
        RECT 1883.340 20.100 1883.600 20.360 ;
        RECT 1921.520 20.100 1921.780 20.360 ;
        RECT 1921.520 16.700 1921.780 16.960 ;
        RECT 2357.600 16.700 2357.860 16.960 ;
      LAYER met2 ;
        RECT 1881.270 600.170 1881.550 604.000 ;
        RECT 1881.270 600.030 1883.540 600.170 ;
        RECT 1881.270 600.000 1881.550 600.030 ;
        RECT 1883.400 20.390 1883.540 600.030 ;
        RECT 1883.340 20.070 1883.600 20.390 ;
        RECT 1921.520 20.070 1921.780 20.390 ;
        RECT 1921.580 16.990 1921.720 20.070 ;
        RECT 1921.520 16.670 1921.780 16.990 ;
        RECT 2357.600 16.670 2357.860 16.990 ;
        RECT 2357.660 2.400 2357.800 16.670 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1921.490 590.140 1921.810 590.200 ;
        RECT 2373.670 590.140 2373.990 590.200 ;
        RECT 1921.490 590.000 2373.990 590.140 ;
        RECT 1921.490 589.940 1921.810 590.000 ;
        RECT 2373.670 589.940 2373.990 590.000 ;
        RECT 1890.210 588.100 1890.530 588.160 ;
        RECT 1921.490 588.100 1921.810 588.160 ;
        RECT 1890.210 587.960 1921.810 588.100 ;
        RECT 1890.210 587.900 1890.530 587.960 ;
        RECT 1921.490 587.900 1921.810 587.960 ;
        RECT 2373.670 2.960 2373.990 3.020 ;
        RECT 2375.510 2.960 2375.830 3.020 ;
        RECT 2373.670 2.820 2375.830 2.960 ;
        RECT 2373.670 2.760 2373.990 2.820 ;
        RECT 2375.510 2.760 2375.830 2.820 ;
      LAYER via ;
        RECT 1921.520 589.940 1921.780 590.200 ;
        RECT 2373.700 589.940 2373.960 590.200 ;
        RECT 1890.240 587.900 1890.500 588.160 ;
        RECT 1921.520 587.900 1921.780 588.160 ;
        RECT 2373.700 2.760 2373.960 3.020 ;
        RECT 2375.540 2.760 2375.800 3.020 ;
      LAYER met2 ;
        RECT 1890.010 600.000 1890.290 604.000 ;
        RECT 1890.070 598.810 1890.210 600.000 ;
        RECT 1890.070 598.670 1890.440 598.810 ;
        RECT 1890.300 588.190 1890.440 598.670 ;
        RECT 1921.520 589.910 1921.780 590.230 ;
        RECT 2373.700 589.910 2373.960 590.230 ;
        RECT 1921.580 588.190 1921.720 589.910 ;
        RECT 1890.240 587.870 1890.500 588.190 ;
        RECT 1921.520 587.870 1921.780 588.190 ;
        RECT 2373.760 3.050 2373.900 589.910 ;
        RECT 2373.700 2.730 2373.960 3.050 ;
        RECT 2375.540 2.730 2375.800 3.050 ;
        RECT 2375.600 2.400 2375.740 2.730 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1900.790 586.740 1901.110 586.800 ;
        RECT 1904.010 586.740 1904.330 586.800 ;
        RECT 1900.790 586.600 1904.330 586.740 ;
        RECT 1900.790 586.540 1901.110 586.600 ;
        RECT 1904.010 586.540 1904.330 586.600 ;
        RECT 1907.320 20.840 1912.520 20.980 ;
        RECT 1904.010 20.640 1904.330 20.700 ;
        RECT 1907.320 20.640 1907.460 20.840 ;
        RECT 1904.010 20.500 1907.460 20.640 ;
        RECT 1912.380 20.640 1912.520 20.840 ;
        RECT 2393.450 20.640 2393.770 20.700 ;
        RECT 1912.380 20.500 2393.770 20.640 ;
        RECT 1904.010 20.440 1904.330 20.500 ;
        RECT 2393.450 20.440 2393.770 20.500 ;
      LAYER via ;
        RECT 1900.820 586.540 1901.080 586.800 ;
        RECT 1904.040 586.540 1904.300 586.800 ;
        RECT 1904.040 20.440 1904.300 20.700 ;
        RECT 2393.480 20.440 2393.740 20.700 ;
      LAYER met2 ;
        RECT 1899.210 600.170 1899.490 604.000 ;
        RECT 1899.210 600.030 1901.020 600.170 ;
        RECT 1899.210 600.000 1899.490 600.030 ;
        RECT 1900.880 586.830 1901.020 600.030 ;
        RECT 1900.820 586.510 1901.080 586.830 ;
        RECT 1904.040 586.510 1904.300 586.830 ;
        RECT 1904.100 20.730 1904.240 586.510 ;
        RECT 1904.040 20.410 1904.300 20.730 ;
        RECT 2393.480 20.410 2393.740 20.730 ;
        RECT 2393.540 2.400 2393.680 20.410 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1909.990 589.800 1910.310 589.860 ;
        RECT 2408.170 589.800 2408.490 589.860 ;
        RECT 1909.990 589.660 2408.490 589.800 ;
        RECT 1909.990 589.600 1910.310 589.660 ;
        RECT 2408.170 589.600 2408.490 589.660 ;
      LAYER via ;
        RECT 1910.020 589.600 1910.280 589.860 ;
        RECT 2408.200 589.600 2408.460 589.860 ;
      LAYER met2 ;
        RECT 1908.410 600.170 1908.690 604.000 ;
        RECT 1908.410 600.030 1910.220 600.170 ;
        RECT 1908.410 600.000 1908.690 600.030 ;
        RECT 1910.080 589.890 1910.220 600.030 ;
        RECT 1910.020 589.570 1910.280 589.890 ;
        RECT 2408.200 589.570 2408.460 589.890 ;
        RECT 2408.260 17.410 2408.400 589.570 ;
        RECT 2408.260 17.270 2411.620 17.410 ;
        RECT 2411.480 2.400 2411.620 17.270 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 805.530 31.180 805.850 31.240 ;
        RECT 1084.290 31.180 1084.610 31.240 ;
        RECT 805.530 31.040 1084.610 31.180 ;
        RECT 805.530 30.980 805.850 31.040 ;
        RECT 1084.290 30.980 1084.610 31.040 ;
      LAYER via ;
        RECT 805.560 30.980 805.820 31.240 ;
        RECT 1084.320 30.980 1084.580 31.240 ;
      LAYER met2 ;
        RECT 1083.630 600.170 1083.910 604.000 ;
        RECT 1083.630 600.030 1084.520 600.170 ;
        RECT 1083.630 600.000 1083.910 600.030 ;
        RECT 1084.380 31.270 1084.520 600.030 ;
        RECT 805.560 30.950 805.820 31.270 ;
        RECT 1084.320 30.950 1084.580 31.270 ;
        RECT 805.620 2.400 805.760 30.950 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 37.980 3.150 38.040 ;
        RECT 669.830 37.980 670.150 38.040 ;
        RECT 2.830 37.840 670.150 37.980 ;
        RECT 2.830 37.780 3.150 37.840 ;
        RECT 669.830 37.780 670.150 37.840 ;
      LAYER via ;
        RECT 2.860 37.780 3.120 38.040 ;
        RECT 669.860 37.780 670.120 38.040 ;
      LAYER met2 ;
        RECT 671.470 600.170 671.750 604.000 ;
        RECT 669.920 600.030 671.750 600.170 ;
        RECT 669.920 38.070 670.060 600.030 ;
        RECT 671.470 600.000 671.750 600.030 ;
        RECT 2.860 37.750 3.120 38.070 ;
        RECT 669.860 37.750 670.120 38.070 ;
        RECT 2.920 2.400 3.060 37.750 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 669.370 569.400 669.690 569.460 ;
        RECT 672.590 569.400 672.910 569.460 ;
        RECT 669.370 569.260 672.910 569.400 ;
        RECT 669.370 569.200 669.690 569.260 ;
        RECT 672.590 569.200 672.910 569.260 ;
        RECT 8.350 38.660 8.670 38.720 ;
        RECT 669.370 38.660 669.690 38.720 ;
        RECT 8.350 38.520 669.690 38.660 ;
        RECT 8.350 38.460 8.670 38.520 ;
        RECT 669.370 38.460 669.690 38.520 ;
      LAYER via ;
        RECT 669.400 569.200 669.660 569.460 ;
        RECT 672.620 569.200 672.880 569.460 ;
        RECT 8.380 38.460 8.640 38.720 ;
        RECT 669.400 38.460 669.660 38.720 ;
      LAYER met2 ;
        RECT 674.230 600.170 674.510 604.000 ;
        RECT 672.680 600.030 674.510 600.170 ;
        RECT 672.680 569.490 672.820 600.030 ;
        RECT 674.230 600.000 674.510 600.030 ;
        RECT 669.400 569.170 669.660 569.490 ;
        RECT 672.620 569.170 672.880 569.490 ;
        RECT 669.460 38.750 669.600 569.170 ;
        RECT 8.380 38.430 8.640 38.750 ;
        RECT 669.400 38.430 669.660 38.750 ;
        RECT 8.440 2.400 8.580 38.430 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 38.320 14.650 38.380 ;
        RECT 676.730 38.320 677.050 38.380 ;
        RECT 14.330 38.180 677.050 38.320 ;
        RECT 14.330 38.120 14.650 38.180 ;
        RECT 676.730 38.120 677.050 38.180 ;
      LAYER via ;
        RECT 14.360 38.120 14.620 38.380 ;
        RECT 676.760 38.120 677.020 38.380 ;
      LAYER met2 ;
        RECT 677.450 600.170 677.730 604.000 ;
        RECT 676.820 600.030 677.730 600.170 ;
        RECT 676.820 38.410 676.960 600.030 ;
        RECT 677.450 600.000 677.730 600.030 ;
        RECT 14.360 38.090 14.620 38.410 ;
        RECT 676.760 38.090 677.020 38.410 ;
        RECT 14.420 2.400 14.560 38.090 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 683.630 569.400 683.950 569.460 ;
        RECT 687.770 569.400 688.090 569.460 ;
        RECT 683.630 569.260 688.090 569.400 ;
        RECT 683.630 569.200 683.950 569.260 ;
        RECT 687.770 569.200 688.090 569.260 ;
        RECT 683.630 62.260 683.950 62.520 ;
        RECT 683.720 61.840 683.860 62.260 ;
        RECT 683.630 61.580 683.950 61.840 ;
        RECT 38.250 39.000 38.570 39.060 ;
        RECT 683.630 39.000 683.950 39.060 ;
        RECT 38.250 38.860 683.950 39.000 ;
        RECT 38.250 38.800 38.570 38.860 ;
        RECT 683.630 38.800 683.950 38.860 ;
      LAYER via ;
        RECT 683.660 569.200 683.920 569.460 ;
        RECT 687.800 569.200 688.060 569.460 ;
        RECT 683.660 62.260 683.920 62.520 ;
        RECT 683.660 61.580 683.920 61.840 ;
        RECT 38.280 38.800 38.540 39.060 ;
        RECT 683.660 38.800 683.920 39.060 ;
      LAYER met2 ;
        RECT 689.410 600.170 689.690 604.000 ;
        RECT 687.860 600.030 689.690 600.170 ;
        RECT 687.860 569.490 688.000 600.030 ;
        RECT 689.410 600.000 689.690 600.030 ;
        RECT 683.660 569.170 683.920 569.490 ;
        RECT 687.800 569.170 688.060 569.490 ;
        RECT 683.720 62.550 683.860 569.170 ;
        RECT 683.660 62.230 683.920 62.550 ;
        RECT 683.660 61.550 683.920 61.870 ;
        RECT 683.720 39.090 683.860 61.550 ;
        RECT 38.280 38.770 38.540 39.090 ;
        RECT 683.660 38.770 683.920 39.090 ;
        RECT 38.340 2.400 38.480 38.770 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 794.490 589.800 794.810 589.860 ;
        RECT 795.870 589.800 796.190 589.860 ;
        RECT 794.490 589.660 796.190 589.800 ;
        RECT 794.490 589.600 794.810 589.660 ;
        RECT 795.870 589.600 796.190 589.660 ;
        RECT 794.030 552.400 794.350 552.460 ;
        RECT 795.870 552.400 796.190 552.460 ;
        RECT 794.030 552.260 796.190 552.400 ;
        RECT 794.030 552.200 794.350 552.260 ;
        RECT 795.870 552.200 796.190 552.260 ;
        RECT 240.650 39.340 240.970 39.400 ;
        RECT 794.030 39.340 794.350 39.400 ;
        RECT 240.650 39.200 794.350 39.340 ;
        RECT 240.650 39.140 240.970 39.200 ;
        RECT 794.030 39.140 794.350 39.200 ;
      LAYER via ;
        RECT 794.520 589.600 794.780 589.860 ;
        RECT 795.900 589.600 796.160 589.860 ;
        RECT 794.060 552.200 794.320 552.460 ;
        RECT 795.900 552.200 796.160 552.460 ;
        RECT 240.680 39.140 240.940 39.400 ;
        RECT 794.060 39.140 794.320 39.400 ;
      LAYER met2 ;
        RECT 793.370 600.170 793.650 604.000 ;
        RECT 793.370 600.030 794.720 600.170 ;
        RECT 793.370 600.000 793.650 600.030 ;
        RECT 794.580 589.890 794.720 600.030 ;
        RECT 794.520 589.570 794.780 589.890 ;
        RECT 795.900 589.570 796.160 589.890 ;
        RECT 795.960 552.490 796.100 589.570 ;
        RECT 794.060 552.170 794.320 552.490 ;
        RECT 795.900 552.170 796.160 552.490 ;
        RECT 794.120 39.430 794.260 552.170 ;
        RECT 240.680 39.110 240.940 39.430 ;
        RECT 794.060 39.110 794.320 39.430 ;
        RECT 240.740 2.400 240.880 39.110 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 46.480 258.450 46.540 ;
        RECT 800.930 46.480 801.250 46.540 ;
        RECT 258.130 46.340 801.250 46.480 ;
        RECT 258.130 46.280 258.450 46.340 ;
        RECT 800.930 46.280 801.250 46.340 ;
      LAYER via ;
        RECT 258.160 46.280 258.420 46.540 ;
        RECT 800.960 46.280 801.220 46.540 ;
      LAYER met2 ;
        RECT 802.570 600.170 802.850 604.000 ;
        RECT 801.020 600.030 802.850 600.170 ;
        RECT 801.020 46.570 801.160 600.030 ;
        RECT 802.570 600.000 802.850 600.030 ;
        RECT 258.160 46.250 258.420 46.570 ;
        RECT 800.960 46.250 801.220 46.570 ;
        RECT 258.220 2.400 258.360 46.250 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 808.290 565.660 808.610 565.720 ;
        RECT 809.210 565.660 809.530 565.720 ;
        RECT 808.290 565.520 809.530 565.660 ;
        RECT 808.290 565.460 808.610 565.520 ;
        RECT 809.210 565.460 809.530 565.520 ;
        RECT 808.290 517.380 808.610 517.440 ;
        RECT 809.670 517.380 809.990 517.440 ;
        RECT 808.290 517.240 809.990 517.380 ;
        RECT 808.290 517.180 808.610 517.240 ;
        RECT 809.670 517.180 809.990 517.240 ;
        RECT 808.750 475.560 809.070 475.620 ;
        RECT 809.670 475.560 809.990 475.620 ;
        RECT 808.750 475.420 809.990 475.560 ;
        RECT 808.750 475.360 809.070 475.420 ;
        RECT 809.670 475.360 809.990 475.420 ;
        RECT 807.830 427.960 808.150 428.020 ;
        RECT 808.750 427.960 809.070 428.020 ;
        RECT 807.830 427.820 809.070 427.960 ;
        RECT 807.830 427.760 808.150 427.820 ;
        RECT 808.750 427.760 809.070 427.820 ;
        RECT 807.830 331.400 808.150 331.460 ;
        RECT 808.290 331.400 808.610 331.460 ;
        RECT 807.830 331.260 808.610 331.400 ;
        RECT 807.830 331.200 808.150 331.260 ;
        RECT 808.290 331.200 808.610 331.260 ;
        RECT 807.830 241.640 808.150 241.700 ;
        RECT 808.750 241.640 809.070 241.700 ;
        RECT 807.830 241.500 809.070 241.640 ;
        RECT 807.830 241.440 808.150 241.500 ;
        RECT 808.750 241.440 809.070 241.500 ;
        RECT 807.830 193.500 808.150 193.760 ;
        RECT 807.920 193.080 808.060 193.500 ;
        RECT 807.830 192.820 808.150 193.080 ;
        RECT 807.830 137.940 808.150 138.000 ;
        RECT 809.210 137.940 809.530 138.000 ;
        RECT 807.830 137.800 809.530 137.940 ;
        RECT 807.830 137.740 808.150 137.800 ;
        RECT 809.210 137.740 809.530 137.800 ;
        RECT 807.830 72.660 808.150 72.720 ;
        RECT 808.750 72.660 809.070 72.720 ;
        RECT 807.830 72.520 809.070 72.660 ;
        RECT 807.830 72.460 808.150 72.520 ;
        RECT 808.750 72.460 809.070 72.520 ;
        RECT 276.070 46.820 276.390 46.880 ;
        RECT 807.830 46.820 808.150 46.880 ;
        RECT 276.070 46.680 808.150 46.820 ;
        RECT 276.070 46.620 276.390 46.680 ;
        RECT 807.830 46.620 808.150 46.680 ;
      LAYER via ;
        RECT 808.320 565.460 808.580 565.720 ;
        RECT 809.240 565.460 809.500 565.720 ;
        RECT 808.320 517.180 808.580 517.440 ;
        RECT 809.700 517.180 809.960 517.440 ;
        RECT 808.780 475.360 809.040 475.620 ;
        RECT 809.700 475.360 809.960 475.620 ;
        RECT 807.860 427.760 808.120 428.020 ;
        RECT 808.780 427.760 809.040 428.020 ;
        RECT 807.860 331.200 808.120 331.460 ;
        RECT 808.320 331.200 808.580 331.460 ;
        RECT 807.860 241.440 808.120 241.700 ;
        RECT 808.780 241.440 809.040 241.700 ;
        RECT 807.860 193.500 808.120 193.760 ;
        RECT 807.860 192.820 808.120 193.080 ;
        RECT 807.860 137.740 808.120 138.000 ;
        RECT 809.240 137.740 809.500 138.000 ;
        RECT 807.860 72.460 808.120 72.720 ;
        RECT 808.780 72.460 809.040 72.720 ;
        RECT 276.100 46.620 276.360 46.880 ;
        RECT 807.860 46.620 808.120 46.880 ;
      LAYER met2 ;
        RECT 811.770 600.850 812.050 604.000 ;
        RECT 809.300 600.710 812.050 600.850 ;
        RECT 809.300 596.770 809.440 600.710 ;
        RECT 811.770 600.000 812.050 600.710 ;
        RECT 808.380 596.630 809.440 596.770 ;
        RECT 808.380 565.750 808.520 596.630 ;
        RECT 808.320 565.430 808.580 565.750 ;
        RECT 809.240 565.430 809.500 565.750 ;
        RECT 809.300 541.010 809.440 565.430 ;
        RECT 808.380 540.870 809.440 541.010 ;
        RECT 808.380 517.470 808.520 540.870 ;
        RECT 808.320 517.150 808.580 517.470 ;
        RECT 809.700 517.150 809.960 517.470 ;
        RECT 809.760 475.650 809.900 517.150 ;
        RECT 808.780 475.330 809.040 475.650 ;
        RECT 809.700 475.330 809.960 475.650 ;
        RECT 808.840 428.050 808.980 475.330 ;
        RECT 807.860 427.730 808.120 428.050 ;
        RECT 808.780 427.730 809.040 428.050 ;
        RECT 807.920 379.170 808.060 427.730 ;
        RECT 807.920 379.030 808.520 379.170 ;
        RECT 808.380 331.490 808.520 379.030 ;
        RECT 807.860 331.170 808.120 331.490 ;
        RECT 808.320 331.170 808.580 331.490 ;
        RECT 807.920 330.890 808.060 331.170 ;
        RECT 807.920 330.750 808.520 330.890 ;
        RECT 808.380 266.290 808.520 330.750 ;
        RECT 808.380 266.150 808.980 266.290 ;
        RECT 808.840 241.730 808.980 266.150 ;
        RECT 807.860 241.410 808.120 241.730 ;
        RECT 808.780 241.410 809.040 241.730 ;
        RECT 807.920 193.790 808.060 241.410 ;
        RECT 807.860 193.470 808.120 193.790 ;
        RECT 807.860 192.790 808.120 193.110 ;
        RECT 807.920 138.030 808.060 192.790 ;
        RECT 807.860 137.710 808.120 138.030 ;
        RECT 809.240 137.710 809.500 138.030 ;
        RECT 809.300 96.290 809.440 137.710 ;
        RECT 808.840 96.150 809.440 96.290 ;
        RECT 808.840 72.750 808.980 96.150 ;
        RECT 807.860 72.430 808.120 72.750 ;
        RECT 808.780 72.430 809.040 72.750 ;
        RECT 807.920 46.910 808.060 72.430 ;
        RECT 276.100 46.590 276.360 46.910 ;
        RECT 807.860 46.590 808.120 46.910 ;
        RECT 276.160 2.400 276.300 46.590 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 47.160 294.330 47.220 ;
        RECT 821.630 47.160 821.950 47.220 ;
        RECT 294.010 47.020 821.950 47.160 ;
        RECT 294.010 46.960 294.330 47.020 ;
        RECT 821.630 46.960 821.950 47.020 ;
      LAYER via ;
        RECT 294.040 46.960 294.300 47.220 ;
        RECT 821.660 46.960 821.920 47.220 ;
      LAYER met2 ;
        RECT 820.970 600.170 821.250 604.000 ;
        RECT 820.970 600.030 821.860 600.170 ;
        RECT 820.970 600.000 821.250 600.030 ;
        RECT 821.720 47.250 821.860 600.030 ;
        RECT 294.040 46.930 294.300 47.250 ;
        RECT 821.660 46.930 821.920 47.250 ;
        RECT 294.100 2.400 294.240 46.930 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 47.500 312.270 47.560 ;
        RECT 828.530 47.500 828.850 47.560 ;
        RECT 311.950 47.360 828.850 47.500 ;
        RECT 311.950 47.300 312.270 47.360 ;
        RECT 828.530 47.300 828.850 47.360 ;
      LAYER via ;
        RECT 311.980 47.300 312.240 47.560 ;
        RECT 828.560 47.300 828.820 47.560 ;
      LAYER met2 ;
        RECT 830.170 600.170 830.450 604.000 ;
        RECT 828.620 600.030 830.450 600.170 ;
        RECT 828.620 47.590 828.760 600.030 ;
        RECT 830.170 600.000 830.450 600.030 ;
        RECT 311.980 47.270 312.240 47.590 ;
        RECT 828.560 47.270 828.820 47.590 ;
        RECT 312.040 2.400 312.180 47.270 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.970 583.000 835.290 583.060 ;
        RECT 837.730 583.000 838.050 583.060 ;
        RECT 834.970 582.860 838.050 583.000 ;
        RECT 834.970 582.800 835.290 582.860 ;
        RECT 837.730 582.800 838.050 582.860 ;
        RECT 329.890 26.760 330.210 26.820 ;
        RECT 834.970 26.760 835.290 26.820 ;
        RECT 329.890 26.620 835.290 26.760 ;
        RECT 329.890 26.560 330.210 26.620 ;
        RECT 834.970 26.560 835.290 26.620 ;
      LAYER via ;
        RECT 835.000 582.800 835.260 583.060 ;
        RECT 837.760 582.800 838.020 583.060 ;
        RECT 329.920 26.560 330.180 26.820 ;
        RECT 835.000 26.560 835.260 26.820 ;
      LAYER met2 ;
        RECT 839.370 600.170 839.650 604.000 ;
        RECT 837.820 600.030 839.650 600.170 ;
        RECT 837.820 583.090 837.960 600.030 ;
        RECT 839.370 600.000 839.650 600.030 ;
        RECT 835.000 582.770 835.260 583.090 ;
        RECT 837.760 582.770 838.020 583.090 ;
        RECT 835.060 26.850 835.200 582.770 ;
        RECT 329.920 26.530 330.180 26.850 ;
        RECT 835.000 26.530 835.260 26.850 ;
        RECT 329.980 2.400 330.120 26.530 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 27.100 347.690 27.160 ;
        RECT 849.690 27.100 850.010 27.160 ;
        RECT 347.370 26.960 850.010 27.100 ;
        RECT 347.370 26.900 347.690 26.960 ;
        RECT 849.690 26.900 850.010 26.960 ;
      LAYER via ;
        RECT 347.400 26.900 347.660 27.160 ;
        RECT 849.720 26.900 849.980 27.160 ;
      LAYER met2 ;
        RECT 848.570 600.170 848.850 604.000 ;
        RECT 848.570 600.030 849.920 600.170 ;
        RECT 848.570 600.000 848.850 600.030 ;
        RECT 849.780 27.190 849.920 600.030 ;
        RECT 347.400 26.870 347.660 27.190 ;
        RECT 849.720 26.870 849.980 27.190 ;
        RECT 347.460 2.400 347.600 26.870 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 27.440 365.630 27.500 ;
        RECT 856.130 27.440 856.450 27.500 ;
        RECT 365.310 27.300 856.450 27.440 ;
        RECT 365.310 27.240 365.630 27.300 ;
        RECT 856.130 27.240 856.450 27.300 ;
      LAYER via ;
        RECT 365.340 27.240 365.600 27.500 ;
        RECT 856.160 27.240 856.420 27.500 ;
      LAYER met2 ;
        RECT 857.770 600.170 858.050 604.000 ;
        RECT 856.220 600.030 858.050 600.170 ;
        RECT 856.220 27.530 856.360 600.030 ;
        RECT 857.770 600.000 858.050 600.030 ;
        RECT 365.340 27.210 365.600 27.530 ;
        RECT 856.160 27.210 856.420 27.530 ;
        RECT 365.400 2.400 365.540 27.210 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.570 573.480 862.890 573.540 ;
        RECT 865.330 573.480 865.650 573.540 ;
        RECT 862.570 573.340 865.650 573.480 ;
        RECT 862.570 573.280 862.890 573.340 ;
        RECT 865.330 573.280 865.650 573.340 ;
        RECT 383.250 23.700 383.570 23.760 ;
        RECT 862.570 23.700 862.890 23.760 ;
        RECT 383.250 23.560 862.890 23.700 ;
        RECT 383.250 23.500 383.570 23.560 ;
        RECT 862.570 23.500 862.890 23.560 ;
      LAYER via ;
        RECT 862.600 573.280 862.860 573.540 ;
        RECT 865.360 573.280 865.620 573.540 ;
        RECT 383.280 23.500 383.540 23.760 ;
        RECT 862.600 23.500 862.860 23.760 ;
      LAYER met2 ;
        RECT 866.970 600.170 867.250 604.000 ;
        RECT 865.420 600.030 867.250 600.170 ;
        RECT 865.420 573.570 865.560 600.030 ;
        RECT 866.970 600.000 867.250 600.030 ;
        RECT 862.600 573.250 862.860 573.570 ;
        RECT 865.360 573.250 865.620 573.570 ;
        RECT 862.660 23.790 862.800 573.250 ;
        RECT 383.280 23.470 383.540 23.790 ;
        RECT 862.600 23.470 862.860 23.790 ;
        RECT 383.340 2.400 383.480 23.470 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 870.390 565.660 870.710 565.720 ;
        RECT 871.310 565.660 871.630 565.720 ;
        RECT 870.390 565.520 871.630 565.660 ;
        RECT 870.390 565.460 870.710 565.520 ;
        RECT 871.310 565.460 871.630 565.520 ;
        RECT 870.850 497.320 871.170 497.380 ;
        RECT 870.480 497.180 871.170 497.320 ;
        RECT 870.480 496.700 870.620 497.180 ;
        RECT 870.850 497.120 871.170 497.180 ;
        RECT 870.390 496.440 870.710 496.700 ;
        RECT 869.470 483.040 869.790 483.100 ;
        RECT 870.390 483.040 870.710 483.100 ;
        RECT 869.470 482.900 870.710 483.040 ;
        RECT 869.470 482.840 869.790 482.900 ;
        RECT 870.390 482.840 870.710 482.900 ;
        RECT 870.850 434.760 871.170 434.820 ;
        RECT 871.770 434.760 872.090 434.820 ;
        RECT 870.850 434.620 872.090 434.760 ;
        RECT 870.850 434.560 871.170 434.620 ;
        RECT 871.770 434.560 872.090 434.620 ;
        RECT 870.390 303.520 870.710 303.580 ;
        RECT 871.310 303.520 871.630 303.580 ;
        RECT 870.390 303.380 871.630 303.520 ;
        RECT 870.390 303.320 870.710 303.380 ;
        RECT 871.310 303.320 871.630 303.380 ;
        RECT 870.390 289.580 870.710 289.640 ;
        RECT 871.310 289.580 871.630 289.640 ;
        RECT 870.390 289.440 871.630 289.580 ;
        RECT 870.390 289.380 870.710 289.440 ;
        RECT 871.310 289.380 871.630 289.440 ;
        RECT 870.390 241.640 870.710 241.700 ;
        RECT 871.770 241.640 872.090 241.700 ;
        RECT 870.390 241.500 872.090 241.640 ;
        RECT 870.390 241.440 870.710 241.500 ;
        RECT 871.770 241.440 872.090 241.500 ;
        RECT 871.310 193.020 871.630 193.080 ;
        RECT 872.230 193.020 872.550 193.080 ;
        RECT 871.310 192.880 872.550 193.020 ;
        RECT 871.310 192.820 871.630 192.880 ;
        RECT 872.230 192.820 872.550 192.880 ;
        RECT 870.850 145.080 871.170 145.140 ;
        RECT 872.230 145.080 872.550 145.140 ;
        RECT 870.850 144.940 872.550 145.080 ;
        RECT 870.850 144.880 871.170 144.940 ;
        RECT 872.230 144.880 872.550 144.940 ;
        RECT 870.390 110.400 870.710 110.460 ;
        RECT 871.310 110.400 871.630 110.460 ;
        RECT 870.390 110.260 871.630 110.400 ;
        RECT 870.390 110.200 870.710 110.260 ;
        RECT 871.310 110.200 871.630 110.260 ;
        RECT 871.310 96.460 871.630 96.520 ;
        RECT 872.230 96.460 872.550 96.520 ;
        RECT 871.310 96.320 872.550 96.460 ;
        RECT 871.310 96.260 871.630 96.320 ;
        RECT 872.230 96.260 872.550 96.320 ;
        RECT 401.190 23.360 401.510 23.420 ;
        RECT 871.310 23.360 871.630 23.420 ;
        RECT 401.190 23.220 871.630 23.360 ;
        RECT 401.190 23.160 401.510 23.220 ;
        RECT 871.310 23.160 871.630 23.220 ;
      LAYER via ;
        RECT 870.420 565.460 870.680 565.720 ;
        RECT 871.340 565.460 871.600 565.720 ;
        RECT 870.880 497.120 871.140 497.380 ;
        RECT 870.420 496.440 870.680 496.700 ;
        RECT 869.500 482.840 869.760 483.100 ;
        RECT 870.420 482.840 870.680 483.100 ;
        RECT 870.880 434.560 871.140 434.820 ;
        RECT 871.800 434.560 872.060 434.820 ;
        RECT 870.420 303.320 870.680 303.580 ;
        RECT 871.340 303.320 871.600 303.580 ;
        RECT 870.420 289.380 870.680 289.640 ;
        RECT 871.340 289.380 871.600 289.640 ;
        RECT 870.420 241.440 870.680 241.700 ;
        RECT 871.800 241.440 872.060 241.700 ;
        RECT 871.340 192.820 871.600 193.080 ;
        RECT 872.260 192.820 872.520 193.080 ;
        RECT 870.880 144.880 871.140 145.140 ;
        RECT 872.260 144.880 872.520 145.140 ;
        RECT 870.420 110.200 870.680 110.460 ;
        RECT 871.340 110.200 871.600 110.460 ;
        RECT 871.340 96.260 871.600 96.520 ;
        RECT 872.260 96.260 872.520 96.520 ;
        RECT 401.220 23.160 401.480 23.420 ;
        RECT 871.340 23.160 871.600 23.420 ;
      LAYER met2 ;
        RECT 875.710 600.170 875.990 604.000 ;
        RECT 873.700 600.030 875.990 600.170 ;
        RECT 873.700 582.490 873.840 600.030 ;
        RECT 875.710 600.000 875.990 600.030 ;
        RECT 870.480 582.350 873.840 582.490 ;
        RECT 870.480 565.750 870.620 582.350 ;
        RECT 870.420 565.430 870.680 565.750 ;
        RECT 871.340 565.430 871.600 565.750 ;
        RECT 871.400 545.090 871.540 565.430 ;
        RECT 870.940 544.950 871.540 545.090 ;
        RECT 870.940 497.410 871.080 544.950 ;
        RECT 870.880 497.090 871.140 497.410 ;
        RECT 870.420 496.410 870.680 496.730 ;
        RECT 870.480 483.130 870.620 496.410 ;
        RECT 869.500 482.810 869.760 483.130 ;
        RECT 870.420 482.810 870.680 483.130 ;
        RECT 869.560 435.045 869.700 482.810 ;
        RECT 869.490 434.675 869.770 435.045 ;
        RECT 870.870 434.675 871.150 435.045 ;
        RECT 870.880 434.530 871.140 434.675 ;
        RECT 871.800 434.530 872.060 434.850 ;
        RECT 871.860 386.650 872.000 434.530 ;
        RECT 871.400 386.510 872.000 386.650 ;
        RECT 871.400 362.170 871.540 386.510 ;
        RECT 870.940 362.030 871.540 362.170 ;
        RECT 870.940 303.690 871.080 362.030 ;
        RECT 870.480 303.610 871.080 303.690 ;
        RECT 870.420 303.550 871.080 303.610 ;
        RECT 870.420 303.290 870.680 303.550 ;
        RECT 871.340 303.290 871.600 303.610 ;
        RECT 871.400 289.670 871.540 303.290 ;
        RECT 870.420 289.350 870.680 289.670 ;
        RECT 871.340 289.350 871.600 289.670 ;
        RECT 870.480 241.730 870.620 289.350 ;
        RECT 870.420 241.410 870.680 241.730 ;
        RECT 871.800 241.410 872.060 241.730 ;
        RECT 871.860 207.925 872.000 241.410 ;
        RECT 871.790 207.555 872.070 207.925 ;
        RECT 871.330 193.275 871.610 193.645 ;
        RECT 871.400 193.110 871.540 193.275 ;
        RECT 871.340 192.790 871.600 193.110 ;
        RECT 872.260 192.790 872.520 193.110 ;
        RECT 872.320 145.170 872.460 192.790 ;
        RECT 870.880 144.850 871.140 145.170 ;
        RECT 872.260 144.850 872.520 145.170 ;
        RECT 870.940 110.570 871.080 144.850 ;
        RECT 870.480 110.490 871.080 110.570 ;
        RECT 870.420 110.430 871.080 110.490 ;
        RECT 870.420 110.170 870.680 110.430 ;
        RECT 871.340 110.170 871.600 110.490 ;
        RECT 871.400 96.550 871.540 110.170 ;
        RECT 871.340 96.230 871.600 96.550 ;
        RECT 872.260 96.230 872.520 96.550 ;
        RECT 872.320 60.930 872.460 96.230 ;
        RECT 871.400 60.790 872.460 60.930 ;
        RECT 871.400 23.450 871.540 60.790 ;
        RECT 401.220 23.130 401.480 23.450 ;
        RECT 871.340 23.130 871.600 23.450 ;
        RECT 401.280 2.400 401.420 23.130 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 869.490 434.720 869.770 435.000 ;
        RECT 870.870 434.720 871.150 435.000 ;
        RECT 871.790 207.600 872.070 207.880 ;
        RECT 871.330 193.320 871.610 193.600 ;
      LAYER met3 ;
        RECT 869.465 435.010 869.795 435.025 ;
        RECT 870.845 435.010 871.175 435.025 ;
        RECT 869.465 434.710 871.175 435.010 ;
        RECT 869.465 434.695 869.795 434.710 ;
        RECT 870.845 434.695 871.175 434.710 ;
        RECT 871.765 207.900 872.095 207.905 ;
        RECT 871.510 207.890 872.095 207.900 ;
        RECT 871.310 207.590 872.095 207.890 ;
        RECT 871.510 207.580 872.095 207.590 ;
        RECT 871.765 207.575 872.095 207.580 ;
        RECT 871.305 193.620 871.635 193.625 ;
        RECT 871.305 193.610 871.890 193.620 ;
        RECT 871.305 193.310 872.090 193.610 ;
        RECT 871.305 193.300 871.890 193.310 ;
        RECT 871.305 193.295 871.635 193.300 ;
      LAYER via3 ;
        RECT 871.540 207.580 871.860 207.900 ;
        RECT 871.540 193.300 871.860 193.620 ;
      LAYER met4 ;
        RECT 871.535 207.575 871.865 207.905 ;
        RECT 871.550 193.625 871.850 207.575 ;
        RECT 871.535 193.295 871.865 193.625 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 697.430 569.400 697.750 569.460 ;
        RECT 700.190 569.400 700.510 569.460 ;
        RECT 697.430 569.260 700.510 569.400 ;
        RECT 697.430 569.200 697.750 569.260 ;
        RECT 700.190 569.200 700.510 569.260 ;
        RECT 62.170 24.380 62.490 24.440 ;
        RECT 697.430 24.380 697.750 24.440 ;
        RECT 62.170 24.240 697.750 24.380 ;
        RECT 62.170 24.180 62.490 24.240 ;
        RECT 697.430 24.180 697.750 24.240 ;
      LAYER via ;
        RECT 697.460 569.200 697.720 569.460 ;
        RECT 700.220 569.200 700.480 569.460 ;
        RECT 62.200 24.180 62.460 24.440 ;
        RECT 697.460 24.180 697.720 24.440 ;
      LAYER met2 ;
        RECT 701.830 600.170 702.110 604.000 ;
        RECT 700.280 600.030 702.110 600.170 ;
        RECT 700.280 569.490 700.420 600.030 ;
        RECT 701.830 600.000 702.110 600.030 ;
        RECT 697.460 569.170 697.720 569.490 ;
        RECT 700.220 569.170 700.480 569.490 ;
        RECT 697.520 24.470 697.660 569.170 ;
        RECT 62.200 24.150 62.460 24.470 ;
        RECT 697.460 24.150 697.720 24.470 ;
        RECT 62.260 2.400 62.400 24.150 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 23.020 419.450 23.080 ;
        RECT 883.730 23.020 884.050 23.080 ;
        RECT 419.130 22.880 884.050 23.020 ;
        RECT 419.130 22.820 419.450 22.880 ;
        RECT 883.730 22.820 884.050 22.880 ;
      LAYER via ;
        RECT 419.160 22.820 419.420 23.080 ;
        RECT 883.760 22.820 884.020 23.080 ;
      LAYER met2 ;
        RECT 884.910 600.170 885.190 604.000 ;
        RECT 883.820 600.030 885.190 600.170 ;
        RECT 883.820 23.110 883.960 600.030 ;
        RECT 884.910 600.000 885.190 600.030 ;
        RECT 419.160 22.790 419.420 23.110 ;
        RECT 883.760 22.790 884.020 23.110 ;
        RECT 419.220 2.400 419.360 22.790 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 890.170 569.400 890.490 569.460 ;
        RECT 892.470 569.400 892.790 569.460 ;
        RECT 890.170 569.260 892.790 569.400 ;
        RECT 890.170 569.200 890.490 569.260 ;
        RECT 892.470 569.200 892.790 569.260 ;
        RECT 436.610 48.180 436.930 48.240 ;
        RECT 890.170 48.180 890.490 48.240 ;
        RECT 436.610 48.040 890.490 48.180 ;
        RECT 436.610 47.980 436.930 48.040 ;
        RECT 890.170 47.980 890.490 48.040 ;
      LAYER via ;
        RECT 890.200 569.200 890.460 569.460 ;
        RECT 892.500 569.200 892.760 569.460 ;
        RECT 436.640 47.980 436.900 48.240 ;
        RECT 890.200 47.980 890.460 48.240 ;
      LAYER met2 ;
        RECT 894.110 600.170 894.390 604.000 ;
        RECT 892.560 600.030 894.390 600.170 ;
        RECT 892.560 569.490 892.700 600.030 ;
        RECT 894.110 600.000 894.390 600.030 ;
        RECT 890.200 569.170 890.460 569.490 ;
        RECT 892.500 569.170 892.760 569.490 ;
        RECT 890.260 48.270 890.400 569.170 ;
        RECT 436.640 47.950 436.900 48.270 ;
        RECT 890.200 47.950 890.460 48.270 ;
        RECT 436.700 2.400 436.840 47.950 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 897.530 569.400 897.850 569.460 ;
        RECT 901.670 569.400 901.990 569.460 ;
        RECT 897.530 569.260 901.990 569.400 ;
        RECT 897.530 569.200 897.850 569.260 ;
        RECT 901.670 569.200 901.990 569.260 ;
        RECT 454.550 44.440 454.870 44.500 ;
        RECT 897.530 44.440 897.850 44.500 ;
        RECT 454.550 44.300 897.850 44.440 ;
        RECT 454.550 44.240 454.870 44.300 ;
        RECT 897.530 44.240 897.850 44.300 ;
      LAYER via ;
        RECT 897.560 569.200 897.820 569.460 ;
        RECT 901.700 569.200 901.960 569.460 ;
        RECT 454.580 44.240 454.840 44.500 ;
        RECT 897.560 44.240 897.820 44.500 ;
      LAYER met2 ;
        RECT 903.310 600.170 903.590 604.000 ;
        RECT 901.760 600.030 903.590 600.170 ;
        RECT 901.760 569.490 901.900 600.030 ;
        RECT 903.310 600.000 903.590 600.030 ;
        RECT 897.560 569.170 897.820 569.490 ;
        RECT 901.700 569.170 901.960 569.490 ;
        RECT 897.620 44.530 897.760 569.170 ;
        RECT 454.580 44.210 454.840 44.530 ;
        RECT 897.560 44.210 897.820 44.530 ;
        RECT 454.640 2.400 454.780 44.210 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 33.560 472.810 33.620 ;
        RECT 911.330 33.560 911.650 33.620 ;
        RECT 472.490 33.420 911.650 33.560 ;
        RECT 472.490 33.360 472.810 33.420 ;
        RECT 911.330 33.360 911.650 33.420 ;
      LAYER via ;
        RECT 472.520 33.360 472.780 33.620 ;
        RECT 911.360 33.360 911.620 33.620 ;
      LAYER met2 ;
        RECT 912.510 600.170 912.790 604.000 ;
        RECT 911.420 600.030 912.790 600.170 ;
        RECT 911.420 33.650 911.560 600.030 ;
        RECT 912.510 600.000 912.790 600.030 ;
        RECT 472.520 33.330 472.780 33.650 ;
        RECT 911.360 33.330 911.620 33.650 ;
        RECT 472.580 2.400 472.720 33.330 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.770 569.400 918.090 569.460 ;
        RECT 920.070 569.400 920.390 569.460 ;
        RECT 917.770 569.260 920.390 569.400 ;
        RECT 917.770 569.200 918.090 569.260 ;
        RECT 920.070 569.200 920.390 569.260 ;
        RECT 490.430 33.900 490.750 33.960 ;
        RECT 917.770 33.900 918.090 33.960 ;
        RECT 490.430 33.760 918.090 33.900 ;
        RECT 490.430 33.700 490.750 33.760 ;
        RECT 917.770 33.700 918.090 33.760 ;
      LAYER via ;
        RECT 917.800 569.200 918.060 569.460 ;
        RECT 920.100 569.200 920.360 569.460 ;
        RECT 490.460 33.700 490.720 33.960 ;
        RECT 917.800 33.700 918.060 33.960 ;
      LAYER met2 ;
        RECT 921.710 600.170 921.990 604.000 ;
        RECT 920.160 600.030 921.990 600.170 ;
        RECT 920.160 569.490 920.300 600.030 ;
        RECT 921.710 600.000 921.990 600.030 ;
        RECT 917.800 569.170 918.060 569.490 ;
        RECT 920.100 569.170 920.360 569.490 ;
        RECT 917.860 33.990 918.000 569.170 ;
        RECT 490.460 33.670 490.720 33.990 ;
        RECT 917.800 33.670 918.060 33.990 ;
        RECT 490.520 2.400 490.660 33.670 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 926.510 524.180 926.830 524.240 ;
        RECT 927.430 524.180 927.750 524.240 ;
        RECT 926.510 524.040 927.750 524.180 ;
        RECT 926.510 523.980 926.830 524.040 ;
        RECT 927.430 523.980 927.750 524.040 ;
        RECT 925.590 476.240 925.910 476.300 ;
        RECT 927.430 476.240 927.750 476.300 ;
        RECT 925.590 476.100 927.750 476.240 ;
        RECT 925.590 476.040 925.910 476.100 ;
        RECT 927.430 476.040 927.750 476.100 ;
        RECT 925.590 427.620 925.910 427.680 ;
        RECT 926.510 427.620 926.830 427.680 ;
        RECT 925.590 427.480 926.830 427.620 ;
        RECT 925.590 427.420 925.910 427.480 ;
        RECT 926.510 427.420 926.830 427.480 ;
        RECT 925.590 352.140 925.910 352.200 ;
        RECT 925.590 352.000 926.280 352.140 ;
        RECT 925.590 351.940 925.910 352.000 ;
        RECT 926.140 351.860 926.280 352.000 ;
        RECT 926.050 351.600 926.370 351.860 ;
        RECT 925.590 338.200 925.910 338.260 ;
        RECT 926.050 338.200 926.370 338.260 ;
        RECT 925.590 338.060 926.370 338.200 ;
        RECT 925.590 338.000 925.910 338.060 ;
        RECT 926.050 338.000 926.370 338.060 ;
        RECT 925.590 326.980 925.910 327.040 ;
        RECT 926.510 326.980 926.830 327.040 ;
        RECT 925.590 326.840 926.830 326.980 ;
        RECT 925.590 326.780 925.910 326.840 ;
        RECT 926.510 326.780 926.830 326.840 ;
        RECT 926.050 241.640 926.370 241.700 ;
        RECT 926.510 241.640 926.830 241.700 ;
        RECT 926.050 241.500 926.830 241.640 ;
        RECT 926.050 241.440 926.370 241.500 ;
        RECT 926.510 241.440 926.830 241.500 ;
        RECT 926.050 131.140 926.370 131.200 ;
        RECT 927.430 131.140 927.750 131.200 ;
        RECT 926.050 131.000 927.750 131.140 ;
        RECT 926.050 130.940 926.370 131.000 ;
        RECT 927.430 130.940 927.750 131.000 ;
        RECT 507.910 30.500 508.230 30.560 ;
        RECT 925.130 30.500 925.450 30.560 ;
        RECT 507.910 30.360 925.450 30.500 ;
        RECT 507.910 30.300 508.230 30.360 ;
        RECT 925.130 30.300 925.450 30.360 ;
      LAYER via ;
        RECT 926.540 523.980 926.800 524.240 ;
        RECT 927.460 523.980 927.720 524.240 ;
        RECT 925.620 476.040 925.880 476.300 ;
        RECT 927.460 476.040 927.720 476.300 ;
        RECT 925.620 427.420 925.880 427.680 ;
        RECT 926.540 427.420 926.800 427.680 ;
        RECT 925.620 351.940 925.880 352.200 ;
        RECT 926.080 351.600 926.340 351.860 ;
        RECT 925.620 338.000 925.880 338.260 ;
        RECT 926.080 338.000 926.340 338.260 ;
        RECT 925.620 326.780 925.880 327.040 ;
        RECT 926.540 326.780 926.800 327.040 ;
        RECT 926.080 241.440 926.340 241.700 ;
        RECT 926.540 241.440 926.800 241.700 ;
        RECT 926.080 130.940 926.340 131.200 ;
        RECT 927.460 130.940 927.720 131.200 ;
        RECT 507.940 30.300 508.200 30.560 ;
        RECT 925.160 30.300 925.420 30.560 ;
      LAYER met2 ;
        RECT 930.910 600.850 931.190 604.000 ;
        RECT 928.440 600.710 931.190 600.850 ;
        RECT 928.440 596.770 928.580 600.710 ;
        RECT 930.910 600.000 931.190 600.710 ;
        RECT 926.140 596.630 928.580 596.770 ;
        RECT 926.140 568.890 926.280 596.630 ;
        RECT 925.680 568.750 926.280 568.890 ;
        RECT 925.680 545.090 925.820 568.750 ;
        RECT 925.680 544.950 926.740 545.090 ;
        RECT 926.600 524.270 926.740 544.950 ;
        RECT 926.540 523.950 926.800 524.270 ;
        RECT 927.460 523.950 927.720 524.270 ;
        RECT 927.520 476.330 927.660 523.950 ;
        RECT 925.620 476.010 925.880 476.330 ;
        RECT 927.460 476.010 927.720 476.330 ;
        RECT 925.680 434.930 925.820 476.010 ;
        RECT 925.680 434.790 926.280 434.930 ;
        RECT 926.140 434.250 926.280 434.790 ;
        RECT 925.680 434.110 926.280 434.250 ;
        RECT 925.680 427.710 925.820 434.110 ;
        RECT 925.620 427.390 925.880 427.710 ;
        RECT 926.540 427.390 926.800 427.710 ;
        RECT 926.600 385.290 926.740 427.390 ;
        RECT 925.680 385.150 926.740 385.290 ;
        RECT 925.680 352.230 925.820 385.150 ;
        RECT 925.620 351.910 925.880 352.230 ;
        RECT 926.080 351.570 926.340 351.890 ;
        RECT 926.140 338.290 926.280 351.570 ;
        RECT 925.620 337.970 925.880 338.290 ;
        RECT 926.080 337.970 926.340 338.290 ;
        RECT 925.680 327.070 925.820 337.970 ;
        RECT 925.620 326.750 925.880 327.070 ;
        RECT 926.540 326.750 926.800 327.070 ;
        RECT 926.600 241.730 926.740 326.750 ;
        RECT 926.080 241.410 926.340 241.730 ;
        RECT 926.540 241.410 926.800 241.730 ;
        RECT 926.140 207.130 926.280 241.410 ;
        RECT 925.680 206.990 926.280 207.130 ;
        RECT 925.680 138.280 925.820 206.990 ;
        RECT 925.680 138.140 926.280 138.280 ;
        RECT 926.140 131.230 926.280 138.140 ;
        RECT 926.080 130.910 926.340 131.230 ;
        RECT 927.460 130.910 927.720 131.230 ;
        RECT 927.520 88.810 927.660 130.910 ;
        RECT 926.140 88.670 927.660 88.810 ;
        RECT 926.140 48.690 926.280 88.670 ;
        RECT 926.140 48.550 926.740 48.690 ;
        RECT 926.600 48.010 926.740 48.550 ;
        RECT 925.680 47.870 926.740 48.010 ;
        RECT 925.680 41.210 925.820 47.870 ;
        RECT 925.220 41.070 925.820 41.210 ;
        RECT 925.220 30.590 925.360 41.070 ;
        RECT 507.940 30.270 508.200 30.590 ;
        RECT 925.160 30.270 925.420 30.590 ;
        RECT 508.000 2.400 508.140 30.270 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 30.160 526.170 30.220 ;
        RECT 938.930 30.160 939.250 30.220 ;
        RECT 525.850 30.020 939.250 30.160 ;
        RECT 525.850 29.960 526.170 30.020 ;
        RECT 938.930 29.960 939.250 30.020 ;
      LAYER via ;
        RECT 525.880 29.960 526.140 30.220 ;
        RECT 938.960 29.960 939.220 30.220 ;
      LAYER met2 ;
        RECT 940.110 600.170 940.390 604.000 ;
        RECT 939.020 600.030 940.390 600.170 ;
        RECT 939.020 30.250 939.160 600.030 ;
        RECT 940.110 600.000 940.390 600.030 ;
        RECT 525.880 29.930 526.140 30.250 ;
        RECT 938.960 29.930 939.220 30.250 ;
        RECT 525.940 2.400 526.080 29.930 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 945.830 556.820 946.150 556.880 ;
        RECT 947.670 556.820 947.990 556.880 ;
        RECT 945.830 556.680 947.990 556.820 ;
        RECT 945.830 556.620 946.150 556.680 ;
        RECT 947.670 556.620 947.990 556.680 ;
        RECT 543.790 29.820 544.110 29.880 ;
        RECT 945.830 29.820 946.150 29.880 ;
        RECT 543.790 29.680 946.150 29.820 ;
        RECT 543.790 29.620 544.110 29.680 ;
        RECT 945.830 29.620 946.150 29.680 ;
      LAYER via ;
        RECT 945.860 556.620 946.120 556.880 ;
        RECT 947.700 556.620 947.960 556.880 ;
        RECT 543.820 29.620 544.080 29.880 ;
        RECT 945.860 29.620 946.120 29.880 ;
      LAYER met2 ;
        RECT 949.310 600.170 949.590 604.000 ;
        RECT 947.760 600.030 949.590 600.170 ;
        RECT 947.760 556.910 947.900 600.030 ;
        RECT 949.310 600.000 949.590 600.030 ;
        RECT 945.860 556.590 946.120 556.910 ;
        RECT 947.700 556.590 947.960 556.910 ;
        RECT 945.920 29.910 946.060 556.590 ;
        RECT 543.820 29.590 544.080 29.910 ;
        RECT 945.860 29.590 946.120 29.910 ;
        RECT 543.880 2.400 544.020 29.590 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 954.110 497.320 954.430 497.380 ;
        RECT 953.740 497.180 954.430 497.320 ;
        RECT 953.740 497.040 953.880 497.180 ;
        RECT 954.110 497.120 954.430 497.180 ;
        RECT 953.650 496.780 953.970 497.040 ;
        RECT 561.730 29.140 562.050 29.200 ;
        RECT 953.650 29.140 953.970 29.200 ;
        RECT 561.730 29.000 953.970 29.140 ;
        RECT 561.730 28.940 562.050 29.000 ;
        RECT 953.650 28.940 953.970 29.000 ;
      LAYER via ;
        RECT 954.140 497.120 954.400 497.380 ;
        RECT 953.680 496.780 953.940 497.040 ;
        RECT 561.760 28.940 562.020 29.200 ;
        RECT 953.680 28.940 953.940 29.200 ;
      LAYER met2 ;
        RECT 958.510 600.170 958.790 604.000 ;
        RECT 956.040 600.030 958.790 600.170 ;
        RECT 956.040 589.290 956.180 600.030 ;
        RECT 958.510 600.000 958.790 600.030 ;
        RECT 954.200 589.150 956.180 589.290 ;
        RECT 954.200 497.410 954.340 589.150 ;
        RECT 954.140 497.090 954.400 497.410 ;
        RECT 953.680 496.750 953.940 497.070 ;
        RECT 953.740 207.130 953.880 496.750 ;
        RECT 953.280 206.990 953.880 207.130 ;
        RECT 953.280 206.450 953.420 206.990 ;
        RECT 953.280 206.310 953.880 206.450 ;
        RECT 953.740 110.570 953.880 206.310 ;
        RECT 953.280 110.430 953.880 110.570 ;
        RECT 953.280 109.890 953.420 110.430 ;
        RECT 953.280 109.750 953.880 109.890 ;
        RECT 953.740 29.230 953.880 109.750 ;
        RECT 561.760 28.910 562.020 29.230 ;
        RECT 953.680 28.910 953.940 29.230 ;
        RECT 561.820 2.400 561.960 28.910 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 580.130 28.800 580.450 28.860 ;
        RECT 966.070 28.800 966.390 28.860 ;
        RECT 580.130 28.660 966.390 28.800 ;
        RECT 580.130 28.600 580.450 28.660 ;
        RECT 966.070 28.600 966.390 28.660 ;
      LAYER via ;
        RECT 580.160 28.600 580.420 28.860 ;
        RECT 966.100 28.600 966.360 28.860 ;
      LAYER met2 ;
        RECT 967.710 600.170 967.990 604.000 ;
        RECT 966.160 600.030 967.990 600.170 ;
        RECT 966.160 28.890 966.300 600.030 ;
        RECT 967.710 600.000 967.990 600.030 ;
        RECT 580.160 28.570 580.420 28.890 ;
        RECT 966.100 28.570 966.360 28.890 ;
        RECT 580.220 14.690 580.360 28.570 ;
        RECT 579.760 14.550 580.360 14.690 ;
        RECT 579.760 2.400 579.900 14.550 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1901.710 2533.240 1902.030 2533.300 ;
        RECT 1903.090 2533.240 1903.410 2533.300 ;
        RECT 1901.710 2533.100 1903.410 2533.240 ;
        RECT 1901.710 2533.040 1902.030 2533.100 ;
        RECT 1903.090 2533.040 1903.410 2533.100 ;
        RECT 653.730 2501.960 654.050 2502.020 ;
        RECT 1903.090 2501.960 1903.410 2502.020 ;
        RECT 653.730 2501.820 1903.410 2501.960 ;
        RECT 653.730 2501.760 654.050 2501.820 ;
        RECT 1903.090 2501.760 1903.410 2501.820 ;
        RECT 653.730 594.900 654.050 594.960 ;
        RECT 711.230 594.900 711.550 594.960 ;
        RECT 712.150 594.900 712.470 594.960 ;
        RECT 653.730 594.760 712.470 594.900 ;
        RECT 653.730 594.700 654.050 594.760 ;
        RECT 711.230 594.700 711.550 594.760 ;
        RECT 712.150 594.700 712.470 594.760 ;
        RECT 86.090 24.720 86.410 24.780 ;
        RECT 711.230 24.720 711.550 24.780 ;
        RECT 86.090 24.580 711.550 24.720 ;
        RECT 86.090 24.520 86.410 24.580 ;
        RECT 711.230 24.520 711.550 24.580 ;
      LAYER via ;
        RECT 1901.740 2533.040 1902.000 2533.300 ;
        RECT 1903.120 2533.040 1903.380 2533.300 ;
        RECT 653.760 2501.760 654.020 2502.020 ;
        RECT 1903.120 2501.760 1903.380 2502.020 ;
        RECT 653.760 594.700 654.020 594.960 ;
        RECT 711.260 594.700 711.520 594.960 ;
        RECT 712.180 594.700 712.440 594.960 ;
        RECT 86.120 24.520 86.380 24.780 ;
        RECT 711.260 24.520 711.520 24.780 ;
      LAYER met2 ;
        RECT 1901.730 2705.195 1902.010 2705.565 ;
        RECT 1901.800 2533.330 1901.940 2705.195 ;
        RECT 1901.740 2533.010 1902.000 2533.330 ;
        RECT 1903.120 2533.010 1903.380 2533.330 ;
        RECT 1903.180 2502.050 1903.320 2533.010 ;
        RECT 653.760 2501.730 654.020 2502.050 ;
        RECT 1903.120 2501.730 1903.380 2502.050 ;
        RECT 653.820 594.990 653.960 2501.730 ;
        RECT 713.790 600.170 714.070 604.000 ;
        RECT 712.240 600.030 714.070 600.170 ;
        RECT 712.240 594.990 712.380 600.030 ;
        RECT 713.790 600.000 714.070 600.030 ;
        RECT 653.760 594.670 654.020 594.990 ;
        RECT 711.260 594.670 711.520 594.990 ;
        RECT 712.180 594.670 712.440 594.990 ;
        RECT 711.320 24.810 711.460 594.670 ;
        RECT 86.120 24.490 86.380 24.810 ;
        RECT 711.260 24.490 711.520 24.810 ;
        RECT 86.180 2.400 86.320 24.490 ;
        RECT 85.970 -4.800 86.530 2.400 ;
      LAYER via2 ;
        RECT 1901.730 2705.240 1902.010 2705.520 ;
      LAYER met3 ;
        RECT 1885.335 2707.080 1889.335 2707.360 ;
        RECT 1885.335 2706.760 1889.370 2707.080 ;
        RECT 1889.070 2705.530 1889.370 2706.760 ;
        RECT 1901.705 2705.530 1902.035 2705.545 ;
        RECT 1889.070 2705.230 1902.035 2705.530 ;
        RECT 1901.705 2705.215 1902.035 2705.230 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.970 569.400 973.290 569.460 ;
        RECT 975.270 569.400 975.590 569.460 ;
        RECT 972.970 569.260 975.590 569.400 ;
        RECT 972.970 569.200 973.290 569.260 ;
        RECT 975.270 569.200 975.590 569.260 ;
        RECT 597.150 28.460 597.470 28.520 ;
        RECT 972.970 28.460 973.290 28.520 ;
        RECT 597.150 28.320 973.290 28.460 ;
        RECT 597.150 28.260 597.470 28.320 ;
        RECT 972.970 28.260 973.290 28.320 ;
      LAYER via ;
        RECT 973.000 569.200 973.260 569.460 ;
        RECT 975.300 569.200 975.560 569.460 ;
        RECT 597.180 28.260 597.440 28.520 ;
        RECT 973.000 28.260 973.260 28.520 ;
      LAYER met2 ;
        RECT 976.910 600.170 977.190 604.000 ;
        RECT 975.360 600.030 977.190 600.170 ;
        RECT 975.360 569.490 975.500 600.030 ;
        RECT 976.910 600.000 977.190 600.030 ;
        RECT 973.000 569.170 973.260 569.490 ;
        RECT 975.300 569.170 975.560 569.490 ;
        RECT 973.060 28.550 973.200 569.170 ;
        RECT 597.180 28.230 597.440 28.550 ;
        RECT 973.000 28.230 973.260 28.550 ;
        RECT 597.240 2.400 597.380 28.230 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 979.870 561.240 980.190 561.300 ;
        RECT 984.470 561.240 984.790 561.300 ;
        RECT 979.870 561.100 984.790 561.240 ;
        RECT 979.870 561.040 980.190 561.100 ;
        RECT 984.470 561.040 984.790 561.100 ;
        RECT 615.090 28.120 615.410 28.180 ;
        RECT 979.870 28.120 980.190 28.180 ;
        RECT 615.090 27.980 980.190 28.120 ;
        RECT 615.090 27.920 615.410 27.980 ;
        RECT 979.870 27.920 980.190 27.980 ;
      LAYER via ;
        RECT 979.900 561.040 980.160 561.300 ;
        RECT 984.500 561.040 984.760 561.300 ;
        RECT 615.120 27.920 615.380 28.180 ;
        RECT 979.900 27.920 980.160 28.180 ;
      LAYER met2 ;
        RECT 986.110 600.170 986.390 604.000 ;
        RECT 984.560 600.030 986.390 600.170 ;
        RECT 984.560 561.330 984.700 600.030 ;
        RECT 986.110 600.000 986.390 600.030 ;
        RECT 979.900 561.010 980.160 561.330 ;
        RECT 984.500 561.010 984.760 561.330 ;
        RECT 979.960 28.210 980.100 561.010 ;
        RECT 615.120 27.890 615.380 28.210 ;
        RECT 979.900 27.890 980.160 28.210 ;
        RECT 615.180 2.400 615.320 27.890 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 654.190 2815.440 654.510 2815.500 ;
        RECT 1490.010 2815.440 1490.330 2815.500 ;
        RECT 654.190 2815.300 1490.330 2815.440 ;
        RECT 654.190 2815.240 654.510 2815.300 ;
        RECT 1490.010 2815.240 1490.330 2815.300 ;
        RECT 654.190 594.560 654.510 594.620 ;
        RECT 725.950 594.560 726.270 594.620 ;
        RECT 654.190 594.420 726.270 594.560 ;
        RECT 654.190 594.360 654.510 594.420 ;
        RECT 725.950 594.360 726.270 594.420 ;
        RECT 724.570 517.720 724.890 517.780 ;
        RECT 725.950 517.720 726.270 517.780 ;
        RECT 724.570 517.580 726.270 517.720 ;
        RECT 724.570 517.520 724.890 517.580 ;
        RECT 725.950 517.520 726.270 517.580 ;
        RECT 724.570 483.380 724.890 483.440 ;
        RECT 725.490 483.380 725.810 483.440 ;
        RECT 724.570 483.240 725.810 483.380 ;
        RECT 724.570 483.180 724.890 483.240 ;
        RECT 725.490 483.180 725.810 483.240 ;
        RECT 725.030 352.280 725.350 352.540 ;
        RECT 725.120 351.180 725.260 352.280 ;
        RECT 725.030 350.920 725.350 351.180 ;
        RECT 725.030 303.660 725.350 303.920 ;
        RECT 725.120 303.240 725.260 303.660 ;
        RECT 725.030 302.980 725.350 303.240 ;
        RECT 725.030 289.580 725.350 289.640 ;
        RECT 726.410 289.580 726.730 289.640 ;
        RECT 725.030 289.440 726.730 289.580 ;
        RECT 725.030 289.380 725.350 289.440 ;
        RECT 726.410 289.380 726.730 289.440 ;
        RECT 725.030 254.560 725.350 254.620 ;
        RECT 726.410 254.560 726.730 254.620 ;
        RECT 725.030 254.420 726.730 254.560 ;
        RECT 725.030 254.360 725.350 254.420 ;
        RECT 726.410 254.360 726.730 254.420 ;
        RECT 725.030 241.100 725.350 241.360 ;
        RECT 725.120 240.960 725.260 241.100 ;
        RECT 725.490 240.960 725.810 241.020 ;
        RECT 725.120 240.820 725.810 240.960 ;
        RECT 725.490 240.760 725.810 240.820 ;
        RECT 725.030 193.360 725.350 193.420 ;
        RECT 725.490 193.360 725.810 193.420 ;
        RECT 725.030 193.220 725.810 193.360 ;
        RECT 725.030 193.160 725.350 193.220 ;
        RECT 725.490 193.160 725.810 193.220 ;
        RECT 725.490 159.020 725.810 159.080 ;
        RECT 725.120 158.880 725.810 159.020 ;
        RECT 725.120 158.740 725.260 158.880 ;
        RECT 725.490 158.820 725.810 158.880 ;
        RECT 725.030 158.480 725.350 158.740 ;
        RECT 724.570 145.080 724.890 145.140 ;
        RECT 725.030 145.080 725.350 145.140 ;
        RECT 724.570 144.940 725.350 145.080 ;
        RECT 724.570 144.880 724.890 144.940 ;
        RECT 725.030 144.880 725.350 144.940 ;
        RECT 724.570 144.060 724.890 144.120 ;
        RECT 725.490 144.060 725.810 144.120 ;
        RECT 724.570 143.920 725.810 144.060 ;
        RECT 724.570 143.860 724.890 143.920 ;
        RECT 725.490 143.860 725.810 143.920 ;
        RECT 725.030 96.800 725.350 96.860 ;
        RECT 725.490 96.800 725.810 96.860 ;
        RECT 725.030 96.660 725.810 96.800 ;
        RECT 725.030 96.600 725.350 96.660 ;
        RECT 725.490 96.600 725.810 96.660 ;
        RECT 724.570 48.520 724.890 48.580 ;
        RECT 725.490 48.520 725.810 48.580 ;
        RECT 724.570 48.380 725.810 48.520 ;
        RECT 724.570 48.320 724.890 48.380 ;
        RECT 725.490 48.320 725.810 48.380 ;
        RECT 109.550 25.060 109.870 25.120 ;
        RECT 724.570 25.060 724.890 25.120 ;
        RECT 109.550 24.920 724.890 25.060 ;
        RECT 109.550 24.860 109.870 24.920 ;
        RECT 724.570 24.860 724.890 24.920 ;
      LAYER via ;
        RECT 654.220 2815.240 654.480 2815.500 ;
        RECT 1490.040 2815.240 1490.300 2815.500 ;
        RECT 654.220 594.360 654.480 594.620 ;
        RECT 725.980 594.360 726.240 594.620 ;
        RECT 724.600 517.520 724.860 517.780 ;
        RECT 725.980 517.520 726.240 517.780 ;
        RECT 724.600 483.180 724.860 483.440 ;
        RECT 725.520 483.180 725.780 483.440 ;
        RECT 725.060 352.280 725.320 352.540 ;
        RECT 725.060 350.920 725.320 351.180 ;
        RECT 725.060 303.660 725.320 303.920 ;
        RECT 725.060 302.980 725.320 303.240 ;
        RECT 725.060 289.380 725.320 289.640 ;
        RECT 726.440 289.380 726.700 289.640 ;
        RECT 725.060 254.360 725.320 254.620 ;
        RECT 726.440 254.360 726.700 254.620 ;
        RECT 725.060 241.100 725.320 241.360 ;
        RECT 725.520 240.760 725.780 241.020 ;
        RECT 725.060 193.160 725.320 193.420 ;
        RECT 725.520 193.160 725.780 193.420 ;
        RECT 725.520 158.820 725.780 159.080 ;
        RECT 725.060 158.480 725.320 158.740 ;
        RECT 724.600 144.880 724.860 145.140 ;
        RECT 725.060 144.880 725.320 145.140 ;
        RECT 724.600 143.860 724.860 144.120 ;
        RECT 725.520 143.860 725.780 144.120 ;
        RECT 725.060 96.600 725.320 96.860 ;
        RECT 725.520 96.600 725.780 96.860 ;
        RECT 724.600 48.320 724.860 48.580 ;
        RECT 725.520 48.320 725.780 48.580 ;
        RECT 109.580 24.860 109.840 25.120 ;
        RECT 724.600 24.860 724.860 25.120 ;
      LAYER met2 ;
        RECT 1490.030 2816.035 1490.310 2816.405 ;
        RECT 1490.100 2815.530 1490.240 2816.035 ;
        RECT 654.220 2815.210 654.480 2815.530 ;
        RECT 1490.040 2815.210 1490.300 2815.530 ;
        RECT 654.280 594.650 654.420 2815.210 ;
        RECT 726.210 600.000 726.490 604.000 ;
        RECT 726.270 598.810 726.410 600.000 ;
        RECT 726.040 598.670 726.410 598.810 ;
        RECT 726.040 594.650 726.180 598.670 ;
        RECT 654.220 594.330 654.480 594.650 ;
        RECT 725.980 594.330 726.240 594.650 ;
        RECT 726.040 517.810 726.180 594.330 ;
        RECT 724.600 517.490 724.860 517.810 ;
        RECT 725.980 517.490 726.240 517.810 ;
        RECT 724.660 483.470 724.800 517.490 ;
        RECT 724.600 483.150 724.860 483.470 ;
        RECT 725.520 483.150 725.780 483.470 ;
        RECT 725.580 400.930 725.720 483.150 ;
        RECT 725.120 400.790 725.720 400.930 ;
        RECT 725.120 352.570 725.260 400.790 ;
        RECT 725.060 352.250 725.320 352.570 ;
        RECT 725.060 350.890 725.320 351.210 ;
        RECT 725.120 303.950 725.260 350.890 ;
        RECT 725.060 303.630 725.320 303.950 ;
        RECT 725.060 302.950 725.320 303.270 ;
        RECT 725.120 289.670 725.260 302.950 ;
        RECT 725.060 289.350 725.320 289.670 ;
        RECT 726.440 289.350 726.700 289.670 ;
        RECT 726.500 254.650 726.640 289.350 ;
        RECT 725.060 254.330 725.320 254.650 ;
        RECT 726.440 254.330 726.700 254.650 ;
        RECT 725.120 241.390 725.260 254.330 ;
        RECT 725.060 241.070 725.320 241.390 ;
        RECT 725.520 240.730 725.780 241.050 ;
        RECT 725.580 193.450 725.720 240.730 ;
        RECT 725.060 193.130 725.320 193.450 ;
        RECT 725.520 193.130 725.780 193.450 ;
        RECT 725.120 192.850 725.260 193.130 ;
        RECT 725.120 192.710 725.720 192.850 ;
        RECT 725.580 159.110 725.720 192.710 ;
        RECT 725.520 158.790 725.780 159.110 ;
        RECT 725.060 158.450 725.320 158.770 ;
        RECT 725.120 145.170 725.260 158.450 ;
        RECT 724.600 144.850 724.860 145.170 ;
        RECT 725.060 144.850 725.320 145.170 ;
        RECT 724.660 144.150 724.800 144.850 ;
        RECT 724.600 143.830 724.860 144.150 ;
        RECT 725.520 143.830 725.780 144.150 ;
        RECT 725.580 96.890 725.720 143.830 ;
        RECT 725.060 96.570 725.320 96.890 ;
        RECT 725.520 96.570 725.780 96.890 ;
        RECT 725.120 96.290 725.260 96.570 ;
        RECT 725.120 96.150 725.720 96.290 ;
        RECT 725.580 48.610 725.720 96.150 ;
        RECT 724.600 48.290 724.860 48.610 ;
        RECT 725.520 48.290 725.780 48.610 ;
        RECT 724.660 25.150 724.800 48.290 ;
        RECT 109.580 24.830 109.840 25.150 ;
        RECT 724.600 24.830 724.860 25.150 ;
        RECT 109.640 2.400 109.780 24.830 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 1490.030 2816.080 1490.310 2816.360 ;
      LAYER met3 ;
        RECT 1500.000 2818.600 1504.000 2818.880 ;
        RECT 1499.910 2818.280 1504.000 2818.600 ;
        RECT 1490.005 2816.370 1490.335 2816.385 ;
        RECT 1499.910 2816.370 1500.210 2818.280 ;
        RECT 1490.005 2816.070 1500.210 2816.370 ;
        RECT 1490.005 2816.055 1490.335 2816.070 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 647.290 2916.760 647.610 2916.820 ;
        RECT 1747.610 2916.760 1747.930 2916.820 ;
        RECT 647.290 2916.620 1747.930 2916.760 ;
        RECT 647.290 2916.560 647.610 2916.620 ;
        RECT 1747.610 2916.560 1747.930 2916.620 ;
        RECT 647.290 594.220 647.610 594.280 ;
        RECT 738.830 594.220 739.150 594.280 ;
        RECT 647.290 594.080 739.150 594.220 ;
        RECT 647.290 594.020 647.610 594.080 ;
        RECT 738.830 594.020 739.150 594.080 ;
        RECT 133.470 25.400 133.790 25.460 ;
        RECT 738.830 25.400 739.150 25.460 ;
        RECT 133.470 25.260 739.150 25.400 ;
        RECT 133.470 25.200 133.790 25.260 ;
        RECT 738.830 25.200 739.150 25.260 ;
      LAYER via ;
        RECT 647.320 2916.560 647.580 2916.820 ;
        RECT 1747.640 2916.560 1747.900 2916.820 ;
        RECT 647.320 594.020 647.580 594.280 ;
        RECT 738.860 594.020 739.120 594.280 ;
        RECT 133.500 25.200 133.760 25.460 ;
        RECT 738.860 25.200 739.120 25.460 ;
      LAYER met2 ;
        RECT 647.320 2916.530 647.580 2916.850 ;
        RECT 1747.640 2916.530 1747.900 2916.850 ;
        RECT 647.380 594.310 647.520 2916.530 ;
        RECT 1747.700 2900.055 1747.840 2916.530 ;
        RECT 1747.570 2896.055 1747.850 2900.055 ;
        RECT 738.630 600.000 738.910 604.000 ;
        RECT 738.690 598.810 738.830 600.000 ;
        RECT 738.690 598.670 739.060 598.810 ;
        RECT 738.920 594.310 739.060 598.670 ;
        RECT 647.320 593.990 647.580 594.310 ;
        RECT 738.860 593.990 739.120 594.310 ;
        RECT 738.920 25.490 739.060 593.990 ;
        RECT 133.500 25.170 133.760 25.490 ;
        RECT 738.860 25.170 739.120 25.490 ;
        RECT 133.560 2.400 133.700 25.170 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 646.830 2502.300 647.150 2502.360 ;
        RECT 1886.990 2502.300 1887.310 2502.360 ;
        RECT 646.830 2502.160 1887.310 2502.300 ;
        RECT 646.830 2502.100 647.150 2502.160 ;
        RECT 1886.990 2502.100 1887.310 2502.160 ;
        RECT 646.830 593.880 647.150 593.940 ;
        RECT 745.270 593.880 745.590 593.940 ;
        RECT 646.830 593.740 745.590 593.880 ;
        RECT 646.830 593.680 647.150 593.740 ;
        RECT 745.270 593.680 745.590 593.740 ;
        RECT 151.410 25.740 151.730 25.800 ;
        RECT 745.270 25.740 745.590 25.800 ;
        RECT 151.410 25.600 745.590 25.740 ;
        RECT 151.410 25.540 151.730 25.600 ;
        RECT 745.270 25.540 745.590 25.600 ;
      LAYER via ;
        RECT 646.860 2502.100 647.120 2502.360 ;
        RECT 1887.020 2502.100 1887.280 2502.360 ;
        RECT 646.860 593.680 647.120 593.940 ;
        RECT 745.300 593.680 745.560 593.940 ;
        RECT 151.440 25.540 151.700 25.800 ;
        RECT 745.300 25.540 745.560 25.800 ;
      LAYER met2 ;
        RECT 1887.010 2860.235 1887.290 2860.605 ;
        RECT 1887.080 2502.390 1887.220 2860.235 ;
        RECT 646.860 2502.070 647.120 2502.390 ;
        RECT 1887.020 2502.070 1887.280 2502.390 ;
        RECT 646.920 593.970 647.060 2502.070 ;
        RECT 747.830 600.170 748.110 604.000 ;
        RECT 745.360 600.030 748.110 600.170 ;
        RECT 745.360 593.970 745.500 600.030 ;
        RECT 747.830 600.000 748.110 600.030 ;
        RECT 646.860 593.650 647.120 593.970 ;
        RECT 745.300 593.650 745.560 593.970 ;
        RECT 745.360 25.830 745.500 593.650 ;
        RECT 151.440 25.510 151.700 25.830 ;
        RECT 745.300 25.510 745.560 25.830 ;
        RECT 151.500 2.400 151.640 25.510 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 1887.010 2860.280 1887.290 2860.560 ;
      LAYER met3 ;
        RECT 1885.335 2863.160 1889.335 2863.760 ;
        RECT 1887.230 2860.585 1887.530 2863.160 ;
        RECT 1886.985 2860.270 1887.530 2860.585 ;
        RECT 1886.985 2860.255 1887.315 2860.270 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 752.170 569.400 752.490 569.460 ;
        RECT 754.930 569.400 755.250 569.460 ;
        RECT 752.170 569.260 755.250 569.400 ;
        RECT 752.170 569.200 752.490 569.260 ;
        RECT 754.930 569.200 755.250 569.260 ;
        RECT 169.350 26.080 169.670 26.140 ;
        RECT 752.170 26.080 752.490 26.140 ;
        RECT 169.350 25.940 752.490 26.080 ;
        RECT 169.350 25.880 169.670 25.940 ;
        RECT 752.170 25.880 752.490 25.940 ;
      LAYER via ;
        RECT 752.200 569.200 752.460 569.460 ;
        RECT 754.960 569.200 755.220 569.460 ;
        RECT 169.380 25.880 169.640 26.140 ;
        RECT 752.200 25.880 752.460 26.140 ;
      LAYER met2 ;
        RECT 756.570 600.170 756.850 604.000 ;
        RECT 755.020 600.030 756.850 600.170 ;
        RECT 755.020 569.490 755.160 600.030 ;
        RECT 756.570 600.000 756.850 600.030 ;
        RECT 752.200 569.170 752.460 569.490 ;
        RECT 754.960 569.170 755.220 569.490 ;
        RECT 752.260 26.170 752.400 569.170 ;
        RECT 169.380 25.850 169.640 26.170 ;
        RECT 752.200 25.850 752.460 26.170 ;
        RECT 169.440 2.400 169.580 25.850 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 26.420 187.150 26.480 ;
        RECT 766.890 26.420 767.210 26.480 ;
        RECT 186.830 26.280 767.210 26.420 ;
        RECT 186.830 26.220 187.150 26.280 ;
        RECT 766.890 26.220 767.210 26.280 ;
      LAYER via ;
        RECT 186.860 26.220 187.120 26.480 ;
        RECT 766.920 26.220 767.180 26.480 ;
      LAYER met2 ;
        RECT 765.770 600.170 766.050 604.000 ;
        RECT 765.770 600.030 767.120 600.170 ;
        RECT 765.770 600.000 766.050 600.030 ;
        RECT 766.980 26.510 767.120 600.030 ;
        RECT 186.860 26.190 187.120 26.510 ;
        RECT 766.920 26.190 767.180 26.510 ;
        RECT 186.920 2.400 187.060 26.190 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 45.800 205.090 45.860 ;
        RECT 772.870 45.800 773.190 45.860 ;
        RECT 204.770 45.660 773.190 45.800 ;
        RECT 204.770 45.600 205.090 45.660 ;
        RECT 772.870 45.600 773.190 45.660 ;
      LAYER via ;
        RECT 204.800 45.600 205.060 45.860 ;
        RECT 772.900 45.600 773.160 45.860 ;
      LAYER met2 ;
        RECT 774.970 600.170 775.250 604.000 ;
        RECT 772.960 600.030 775.250 600.170 ;
        RECT 772.960 45.890 773.100 600.030 ;
        RECT 774.970 600.000 775.250 600.030 ;
        RECT 204.800 45.570 205.060 45.890 ;
        RECT 772.900 45.570 773.160 45.890 ;
        RECT 204.860 2.400 205.000 45.570 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 782.070 600.340 782.390 600.400 ;
        RECT 782.990 600.340 783.310 600.400 ;
        RECT 782.070 600.200 783.310 600.340 ;
        RECT 782.070 600.140 782.390 600.200 ;
        RECT 782.990 600.140 783.310 600.200 ;
        RECT 782.530 517.720 782.850 517.780 ;
        RECT 782.990 517.720 783.310 517.780 ;
        RECT 782.530 517.580 783.310 517.720 ;
        RECT 782.530 517.520 782.850 517.580 ;
        RECT 782.990 517.520 783.310 517.580 ;
        RECT 780.230 469.440 780.550 469.500 ;
        RECT 782.530 469.440 782.850 469.500 ;
        RECT 780.230 469.300 782.850 469.440 ;
        RECT 780.230 469.240 780.550 469.300 ;
        RECT 782.530 469.240 782.850 469.300 ;
        RECT 780.230 338.200 780.550 338.260 ;
        RECT 780.690 338.200 781.010 338.260 ;
        RECT 780.230 338.060 781.010 338.200 ;
        RECT 780.230 338.000 780.550 338.060 ;
        RECT 780.690 338.000 781.010 338.060 ;
        RECT 780.230 331.060 780.550 331.120 ;
        RECT 781.150 331.060 781.470 331.120 ;
        RECT 780.230 330.920 781.470 331.060 ;
        RECT 780.230 330.860 780.550 330.920 ;
        RECT 781.150 330.860 781.470 330.920 ;
        RECT 781.150 283.460 781.470 283.520 ;
        RECT 781.150 283.320 781.840 283.460 ;
        RECT 781.150 283.260 781.470 283.320 ;
        RECT 781.700 283.180 781.840 283.320 ;
        RECT 781.610 282.920 781.930 283.180 ;
        RECT 780.690 234.500 781.010 234.560 ;
        RECT 780.690 234.360 781.380 234.500 ;
        RECT 780.690 234.300 781.010 234.360 ;
        RECT 781.240 234.220 781.380 234.360 ;
        RECT 781.150 233.960 781.470 234.220 ;
        RECT 780.690 96.800 781.010 96.860 ;
        RECT 781.150 96.800 781.470 96.860 ;
        RECT 780.690 96.660 781.470 96.800 ;
        RECT 780.690 96.600 781.010 96.660 ;
        RECT 781.150 96.600 781.470 96.660 ;
        RECT 780.690 48.860 781.010 48.920 ;
        RECT 780.320 48.720 781.010 48.860 ;
        RECT 780.320 48.580 780.460 48.720 ;
        RECT 780.690 48.660 781.010 48.720 ;
        RECT 780.230 48.320 780.550 48.580 ;
        RECT 222.710 31.860 223.030 31.920 ;
        RECT 780.230 31.860 780.550 31.920 ;
        RECT 222.710 31.720 780.550 31.860 ;
        RECT 222.710 31.660 223.030 31.720 ;
        RECT 780.230 31.660 780.550 31.720 ;
      LAYER via ;
        RECT 782.100 600.140 782.360 600.400 ;
        RECT 783.020 600.140 783.280 600.400 ;
        RECT 782.560 517.520 782.820 517.780 ;
        RECT 783.020 517.520 783.280 517.780 ;
        RECT 780.260 469.240 780.520 469.500 ;
        RECT 782.560 469.240 782.820 469.500 ;
        RECT 780.260 338.000 780.520 338.260 ;
        RECT 780.720 338.000 780.980 338.260 ;
        RECT 780.260 330.860 780.520 331.120 ;
        RECT 781.180 330.860 781.440 331.120 ;
        RECT 781.180 283.260 781.440 283.520 ;
        RECT 781.640 282.920 781.900 283.180 ;
        RECT 780.720 234.300 780.980 234.560 ;
        RECT 781.180 233.960 781.440 234.220 ;
        RECT 780.720 96.600 780.980 96.860 ;
        RECT 781.180 96.600 781.440 96.860 ;
        RECT 780.720 48.660 780.980 48.920 ;
        RECT 780.260 48.320 780.520 48.580 ;
        RECT 222.740 31.660 223.000 31.920 ;
        RECT 780.260 31.660 780.520 31.920 ;
      LAYER met2 ;
        RECT 784.170 600.850 784.450 604.000 ;
        RECT 782.160 600.710 784.450 600.850 ;
        RECT 782.160 600.430 782.300 600.710 ;
        RECT 782.100 600.110 782.360 600.430 ;
        RECT 783.020 600.110 783.280 600.430 ;
        RECT 783.080 517.810 783.220 600.110 ;
        RECT 784.170 600.000 784.450 600.710 ;
        RECT 782.560 517.490 782.820 517.810 ;
        RECT 783.020 517.490 783.280 517.810 ;
        RECT 782.620 469.530 782.760 517.490 ;
        RECT 780.260 469.210 780.520 469.530 ;
        RECT 782.560 469.210 782.820 469.530 ;
        RECT 780.320 428.245 780.460 469.210 ;
        RECT 780.250 427.875 780.530 428.245 ;
        RECT 780.710 426.515 780.990 426.885 ;
        RECT 780.780 338.290 780.920 426.515 ;
        RECT 780.260 337.970 780.520 338.290 ;
        RECT 780.720 337.970 780.980 338.290 ;
        RECT 780.320 331.150 780.460 337.970 ;
        RECT 780.260 330.830 780.520 331.150 ;
        RECT 781.180 330.830 781.440 331.150 ;
        RECT 781.240 283.550 781.380 330.830 ;
        RECT 781.180 283.230 781.440 283.550 ;
        RECT 781.640 282.890 781.900 283.210 ;
        RECT 781.700 258.810 781.840 282.890 ;
        RECT 780.780 258.670 781.840 258.810 ;
        RECT 780.780 234.590 780.920 258.670 ;
        RECT 780.720 234.270 780.980 234.590 ;
        RECT 781.180 233.930 781.440 234.250 ;
        RECT 781.240 96.890 781.380 233.930 ;
        RECT 780.720 96.570 780.980 96.890 ;
        RECT 781.180 96.570 781.440 96.890 ;
        RECT 780.780 48.950 780.920 96.570 ;
        RECT 780.720 48.630 780.980 48.950 ;
        RECT 780.260 48.290 780.520 48.610 ;
        RECT 780.320 31.950 780.460 48.290 ;
        RECT 222.740 31.630 223.000 31.950 ;
        RECT 780.260 31.630 780.520 31.950 ;
        RECT 222.800 2.400 222.940 31.630 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 780.250 427.920 780.530 428.200 ;
        RECT 780.710 426.560 780.990 426.840 ;
      LAYER met3 ;
        RECT 780.225 428.210 780.555 428.225 ;
        RECT 779.550 427.910 780.555 428.210 ;
        RECT 779.550 426.850 779.850 427.910 ;
        RECT 780.225 427.895 780.555 427.910 ;
        RECT 780.685 426.850 781.015 426.865 ;
        RECT 779.550 426.550 781.015 426.850 ;
        RECT 780.685 426.535 781.015 426.550 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 676.270 569.400 676.590 569.460 ;
        RECT 678.570 569.400 678.890 569.460 ;
        RECT 676.270 569.260 678.890 569.400 ;
        RECT 676.270 569.200 676.590 569.260 ;
        RECT 678.570 569.200 678.890 569.260 ;
        RECT 20.310 24.040 20.630 24.100 ;
        RECT 676.270 24.040 676.590 24.100 ;
        RECT 20.310 23.900 676.590 24.040 ;
        RECT 20.310 23.840 20.630 23.900 ;
        RECT 676.270 23.840 676.590 23.900 ;
      LAYER via ;
        RECT 676.300 569.200 676.560 569.460 ;
        RECT 678.600 569.200 678.860 569.460 ;
        RECT 20.340 23.840 20.600 24.100 ;
        RECT 676.300 23.840 676.560 24.100 ;
      LAYER met2 ;
        RECT 680.210 600.170 680.490 604.000 ;
        RECT 678.660 600.030 680.490 600.170 ;
        RECT 678.660 569.490 678.800 600.030 ;
        RECT 680.210 600.000 680.490 600.030 ;
        RECT 676.300 569.170 676.560 569.490 ;
        RECT 678.600 569.170 678.860 569.490 ;
        RECT 676.360 24.130 676.500 569.170 ;
        RECT 20.340 23.810 20.600 24.130 ;
        RECT 676.300 23.810 676.560 24.130 ;
        RECT 20.400 2.400 20.540 23.810 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.570 2504.680 517.890 2504.740 ;
        RECT 524.010 2504.680 524.330 2504.740 ;
        RECT 517.570 2504.540 524.330 2504.680 ;
        RECT 517.570 2504.480 517.890 2504.540 ;
        RECT 524.010 2504.480 524.330 2504.540 ;
        RECT 524.010 2503.660 524.330 2503.720 ;
        RECT 1888.370 2503.660 1888.690 2503.720 ;
        RECT 524.010 2503.520 1888.690 2503.660 ;
        RECT 524.010 2503.460 524.330 2503.520 ;
        RECT 1888.370 2503.460 1888.690 2503.520 ;
        RECT 350.590 2038.880 350.910 2038.940 ;
        RECT 524.010 2038.880 524.330 2038.940 ;
        RECT 2083.870 2038.880 2084.190 2038.940 ;
        RECT 350.590 2038.740 2084.190 2038.880 ;
        RECT 350.590 2038.680 350.910 2038.740 ;
        RECT 524.010 2038.680 524.330 2038.740 ;
        RECT 2083.870 2038.680 2084.190 2038.740 ;
        RECT 349.210 593.200 349.530 593.260 ;
        RECT 351.510 593.200 351.830 593.260 ;
        RECT 690.990 593.200 691.310 593.260 ;
        RECT 349.210 593.060 691.310 593.200 ;
        RECT 349.210 593.000 349.530 593.060 ;
        RECT 351.510 593.000 351.830 593.060 ;
        RECT 690.990 593.000 691.310 593.060 ;
        RECT 47.910 589.800 48.230 589.860 ;
        RECT 349.210 589.800 349.530 589.860 ;
        RECT 47.910 589.660 349.530 589.800 ;
        RECT 47.910 589.600 48.230 589.660 ;
        RECT 349.210 589.600 349.530 589.660 ;
        RECT 44.230 17.580 44.550 17.640 ;
        RECT 47.910 17.580 48.230 17.640 ;
        RECT 44.230 17.440 48.230 17.580 ;
        RECT 44.230 17.380 44.550 17.440 ;
        RECT 47.910 17.380 48.230 17.440 ;
      LAYER via ;
        RECT 517.600 2504.480 517.860 2504.740 ;
        RECT 524.040 2504.480 524.300 2504.740 ;
        RECT 524.040 2503.460 524.300 2503.720 ;
        RECT 1888.400 2503.460 1888.660 2503.720 ;
        RECT 350.620 2038.680 350.880 2038.940 ;
        RECT 524.040 2038.680 524.300 2038.940 ;
        RECT 2083.900 2038.680 2084.160 2038.940 ;
        RECT 349.240 593.000 349.500 593.260 ;
        RECT 351.540 593.000 351.800 593.260 ;
        RECT 691.020 593.000 691.280 593.260 ;
        RECT 47.940 589.600 48.200 589.860 ;
        RECT 349.240 589.600 349.500 589.860 ;
        RECT 44.260 17.380 44.520 17.640 ;
        RECT 47.940 17.380 48.200 17.640 ;
      LAYER met2 ;
        RECT 519.330 2600.730 519.610 2604.000 ;
        RECT 517.660 2600.590 519.610 2600.730 ;
        RECT 517.660 2504.770 517.800 2600.590 ;
        RECT 519.330 2600.000 519.610 2600.590 ;
        RECT 1888.390 2595.715 1888.670 2596.085 ;
        RECT 517.600 2504.450 517.860 2504.770 ;
        RECT 524.040 2504.450 524.300 2504.770 ;
        RECT 524.100 2503.750 524.240 2504.450 ;
        RECT 1888.460 2503.750 1888.600 2595.715 ;
        RECT 524.040 2503.430 524.300 2503.750 ;
        RECT 1888.400 2503.430 1888.660 2503.750 ;
        RECT 524.100 2038.970 524.240 2503.430 ;
        RECT 350.620 2038.650 350.880 2038.970 ;
        RECT 524.040 2038.650 524.300 2038.970 ;
        RECT 2083.900 2038.650 2084.160 2038.970 ;
        RECT 350.680 1851.485 350.820 2038.650 ;
        RECT 2083.960 1873.245 2084.100 2038.650 ;
        RECT 2083.890 1872.875 2084.170 1873.245 ;
        RECT 350.610 1851.115 350.890 1851.485 ;
        RECT 351.530 1851.115 351.810 1851.485 ;
        RECT 351.600 593.290 351.740 1851.115 ;
        RECT 692.630 600.170 692.910 604.000 ;
        RECT 691.080 600.030 692.910 600.170 ;
        RECT 691.080 593.290 691.220 600.030 ;
        RECT 692.630 600.000 692.910 600.030 ;
        RECT 349.240 592.970 349.500 593.290 ;
        RECT 351.540 592.970 351.800 593.290 ;
        RECT 691.020 592.970 691.280 593.290 ;
        RECT 349.300 589.890 349.440 592.970 ;
        RECT 47.940 589.570 48.200 589.890 ;
        RECT 349.240 589.570 349.500 589.890 ;
        RECT 48.000 17.670 48.140 589.570 ;
        RECT 44.260 17.350 44.520 17.670 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 44.320 2.400 44.460 17.350 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 1888.390 2595.760 1888.670 2596.040 ;
        RECT 2083.890 1872.920 2084.170 1873.200 ;
        RECT 350.610 1851.160 350.890 1851.440 ;
        RECT 351.530 1851.160 351.810 1851.440 ;
      LAYER met3 ;
        RECT 1885.335 2596.600 1889.335 2597.200 ;
        RECT 1888.150 2596.065 1888.450 2596.600 ;
        RECT 1888.150 2595.750 1888.695 2596.065 ;
        RECT 1888.365 2595.735 1888.695 2595.750 ;
        RECT 2083.865 1873.210 2084.195 1873.225 ;
        RECT 2075.830 1872.910 2084.195 1873.210 ;
        RECT 2075.830 1870.320 2076.130 1872.910 ;
        RECT 2083.865 1872.895 2084.195 1872.910 ;
        RECT 2072.375 1869.720 2076.375 1870.320 ;
        RECT 350.585 1851.450 350.915 1851.465 ;
        RECT 351.505 1851.450 351.835 1851.465 ;
        RECT 360.000 1851.450 364.000 1851.600 ;
        RECT 350.585 1851.150 364.000 1851.450 ;
        RECT 350.585 1851.135 350.915 1851.150 ;
        RECT 351.505 1851.135 351.835 1851.150 ;
        RECT 360.000 1851.000 364.000 1851.150 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1554.870 2896.500 1555.190 2896.760 ;
        RECT 787.130 2892.620 787.450 2892.680 ;
        RECT 883.730 2892.620 884.050 2892.680 ;
        RECT 980.330 2892.620 980.650 2892.680 ;
        RECT 1076.930 2892.620 1077.250 2892.680 ;
        RECT 1173.530 2892.620 1173.850 2892.680 ;
        RECT 1270.130 2892.620 1270.450 2892.680 ;
        RECT 1317.510 2892.620 1317.830 2892.680 ;
        RECT 787.130 2892.480 821.400 2892.620 ;
        RECT 787.130 2892.420 787.450 2892.480 ;
        RECT 821.260 2892.340 821.400 2892.480 ;
        RECT 883.730 2892.480 918.000 2892.620 ;
        RECT 883.730 2892.420 884.050 2892.480 ;
        RECT 917.860 2892.340 918.000 2892.480 ;
        RECT 980.330 2892.480 1014.600 2892.620 ;
        RECT 980.330 2892.420 980.650 2892.480 ;
        RECT 1014.460 2892.340 1014.600 2892.480 ;
        RECT 1076.930 2892.480 1111.200 2892.620 ;
        RECT 1076.930 2892.420 1077.250 2892.480 ;
        RECT 1111.060 2892.340 1111.200 2892.480 ;
        RECT 1173.530 2892.480 1207.800 2892.620 ;
        RECT 1173.530 2892.420 1173.850 2892.480 ;
        RECT 1207.660 2892.340 1207.800 2892.480 ;
        RECT 1270.130 2892.480 1317.830 2892.620 ;
        RECT 1270.130 2892.420 1270.450 2892.480 ;
        RECT 1317.510 2892.420 1317.830 2892.480 ;
        RECT 1366.730 2892.620 1367.050 2892.680 ;
        RECT 1366.730 2892.480 1401.000 2892.620 ;
        RECT 1366.730 2892.420 1367.050 2892.480 ;
        RECT 1400.860 2892.340 1401.000 2892.480 ;
        RECT 772.410 2892.280 772.730 2892.340 ;
        RECT 786.210 2892.280 786.530 2892.340 ;
        RECT 772.410 2892.140 786.530 2892.280 ;
        RECT 772.410 2892.080 772.730 2892.140 ;
        RECT 786.210 2892.080 786.530 2892.140 ;
        RECT 821.170 2892.080 821.490 2892.340 ;
        RECT 869.010 2892.280 869.330 2892.340 ;
        RECT 882.810 2892.280 883.130 2892.340 ;
        RECT 869.010 2892.140 883.130 2892.280 ;
        RECT 869.010 2892.080 869.330 2892.140 ;
        RECT 882.810 2892.080 883.130 2892.140 ;
        RECT 917.770 2892.080 918.090 2892.340 ;
        RECT 965.610 2892.280 965.930 2892.340 ;
        RECT 979.410 2892.280 979.730 2892.340 ;
        RECT 965.610 2892.140 979.730 2892.280 ;
        RECT 965.610 2892.080 965.930 2892.140 ;
        RECT 979.410 2892.080 979.730 2892.140 ;
        RECT 1014.370 2892.080 1014.690 2892.340 ;
        RECT 1062.210 2892.280 1062.530 2892.340 ;
        RECT 1076.010 2892.280 1076.330 2892.340 ;
        RECT 1062.210 2892.140 1076.330 2892.280 ;
        RECT 1062.210 2892.080 1062.530 2892.140 ;
        RECT 1076.010 2892.080 1076.330 2892.140 ;
        RECT 1110.970 2892.080 1111.290 2892.340 ;
        RECT 1158.810 2892.280 1159.130 2892.340 ;
        RECT 1172.610 2892.280 1172.930 2892.340 ;
        RECT 1158.810 2892.140 1172.930 2892.280 ;
        RECT 1158.810 2892.080 1159.130 2892.140 ;
        RECT 1172.610 2892.080 1172.930 2892.140 ;
        RECT 1207.570 2892.080 1207.890 2892.340 ;
        RECT 1255.410 2892.280 1255.730 2892.340 ;
        RECT 1269.210 2892.280 1269.530 2892.340 ;
        RECT 1255.410 2892.140 1269.530 2892.280 ;
        RECT 1255.410 2892.080 1255.730 2892.140 ;
        RECT 1269.210 2892.080 1269.530 2892.140 ;
        RECT 1317.970 2892.280 1318.290 2892.340 ;
        RECT 1365.810 2892.280 1366.130 2892.340 ;
        RECT 1317.970 2892.140 1366.130 2892.280 ;
        RECT 1317.970 2892.080 1318.290 2892.140 ;
        RECT 1365.810 2892.080 1366.130 2892.140 ;
        RECT 1400.770 2892.080 1401.090 2892.340 ;
        RECT 1448.610 2892.280 1448.930 2892.340 ;
        RECT 1462.410 2892.280 1462.730 2892.340 ;
        RECT 1448.610 2892.140 1462.730 2892.280 ;
        RECT 1448.610 2892.080 1448.930 2892.140 ;
        RECT 1462.410 2892.080 1462.730 2892.140 ;
        RECT 1462.870 2892.280 1463.190 2892.340 ;
        RECT 1462.870 2892.140 1497.140 2892.280 ;
        RECT 1462.870 2892.080 1463.190 2892.140 ;
        RECT 651.890 2891.940 652.210 2892.000 ;
        RECT 689.610 2891.940 689.930 2892.000 ;
        RECT 651.890 2891.800 689.930 2891.940 ;
        RECT 651.890 2891.740 652.210 2891.800 ;
        RECT 689.610 2891.740 689.930 2891.800 ;
        RECT 690.530 2891.600 690.850 2891.660 ;
        RECT 724.570 2891.600 724.890 2891.660 ;
        RECT 690.530 2891.460 724.890 2891.600 ;
        RECT 690.530 2891.400 690.850 2891.460 ;
        RECT 724.570 2891.400 724.890 2891.460 ;
        RECT 821.170 2891.600 821.490 2891.660 ;
        RECT 869.010 2891.600 869.330 2891.660 ;
        RECT 821.170 2891.460 869.330 2891.600 ;
        RECT 821.170 2891.400 821.490 2891.460 ;
        RECT 869.010 2891.400 869.330 2891.460 ;
        RECT 917.770 2891.600 918.090 2891.660 ;
        RECT 965.610 2891.600 965.930 2891.660 ;
        RECT 917.770 2891.460 965.930 2891.600 ;
        RECT 917.770 2891.400 918.090 2891.460 ;
        RECT 965.610 2891.400 965.930 2891.460 ;
        RECT 1014.370 2891.600 1014.690 2891.660 ;
        RECT 1062.210 2891.600 1062.530 2891.660 ;
        RECT 1014.370 2891.460 1062.530 2891.600 ;
        RECT 1014.370 2891.400 1014.690 2891.460 ;
        RECT 1062.210 2891.400 1062.530 2891.460 ;
        RECT 1110.970 2891.600 1111.290 2891.660 ;
        RECT 1158.810 2891.600 1159.130 2891.660 ;
        RECT 1110.970 2891.460 1159.130 2891.600 ;
        RECT 1110.970 2891.400 1111.290 2891.460 ;
        RECT 1158.810 2891.400 1159.130 2891.460 ;
        RECT 1207.570 2891.600 1207.890 2891.660 ;
        RECT 1255.410 2891.600 1255.730 2891.660 ;
        RECT 1207.570 2891.460 1255.730 2891.600 ;
        RECT 1207.570 2891.400 1207.890 2891.460 ;
        RECT 1255.410 2891.400 1255.730 2891.460 ;
        RECT 1400.770 2891.600 1401.090 2891.660 ;
        RECT 1448.610 2891.600 1448.930 2891.660 ;
        RECT 1400.770 2891.460 1448.930 2891.600 ;
        RECT 1497.000 2891.600 1497.140 2892.140 ;
        RECT 1554.960 2891.600 1555.100 2896.500 ;
        RECT 1497.000 2891.460 1555.100 2891.600 ;
        RECT 1400.770 2891.400 1401.090 2891.460 ;
        RECT 1448.610 2891.400 1448.930 2891.460 ;
        RECT 724.570 2890.920 724.890 2890.980 ;
        RECT 772.410 2890.920 772.730 2890.980 ;
        RECT 724.570 2890.780 772.730 2890.920 ;
        RECT 724.570 2890.720 724.890 2890.780 ;
        RECT 772.410 2890.720 772.730 2890.780 ;
        RECT 446.730 2594.440 447.050 2594.500 ;
        RECT 612.790 2594.440 613.110 2594.500 ;
        RECT 446.730 2594.300 613.110 2594.440 ;
        RECT 446.730 2594.240 447.050 2594.300 ;
        RECT 612.790 2594.240 613.110 2594.300 ;
        RECT 614.170 2594.440 614.490 2594.500 ;
        RECT 648.670 2594.440 648.990 2594.500 ;
        RECT 614.170 2594.300 648.990 2594.440 ;
        RECT 614.170 2594.240 614.490 2594.300 ;
        RECT 648.670 2594.240 648.990 2594.300 ;
        RECT 648.670 2592.740 648.990 2592.800 ;
        RECT 651.890 2592.740 652.210 2592.800 ;
        RECT 648.670 2592.600 652.210 2592.740 ;
        RECT 648.670 2592.540 648.990 2592.600 ;
        RECT 651.890 2592.540 652.210 2592.600 ;
        RECT 644.070 1758.720 644.390 1758.780 ;
        RECT 648.670 1758.720 648.990 1758.780 ;
        RECT 651.890 1758.720 652.210 1758.780 ;
        RECT 644.070 1758.580 652.210 1758.720 ;
        RECT 644.070 1758.520 644.390 1758.580 ;
        RECT 648.670 1758.520 648.990 1758.580 ;
        RECT 651.890 1758.520 652.210 1758.580 ;
        RECT 651.890 1703.300 652.210 1703.360 ;
        RECT 1401.230 1703.300 1401.550 1703.360 ;
        RECT 651.890 1703.160 1401.550 1703.300 ;
        RECT 651.890 1703.100 652.210 1703.160 ;
        RECT 1401.230 1703.100 1401.550 1703.160 ;
        RECT 1403.070 1703.300 1403.390 1703.360 ;
        RECT 1642.730 1703.300 1643.050 1703.360 ;
        RECT 1403.070 1703.160 1643.050 1703.300 ;
        RECT 1403.070 1703.100 1403.390 1703.160 ;
        RECT 1642.730 1703.100 1643.050 1703.160 ;
        RECT 1644.570 1703.300 1644.890 1703.360 ;
        RECT 1907.690 1703.300 1908.010 1703.360 ;
        RECT 1644.570 1703.160 1908.010 1703.300 ;
        RECT 1644.570 1703.100 1644.890 1703.160 ;
        RECT 1907.690 1703.100 1908.010 1703.160 ;
        RECT 651.890 588.440 652.210 588.500 ;
        RECT 651.890 588.300 666.380 588.440 ;
        RECT 651.890 588.240 652.210 588.300 ;
        RECT 666.240 588.100 666.380 588.300 ;
        RECT 794.950 588.100 795.270 588.160 ;
        RECT 666.240 587.960 795.270 588.100 ;
        RECT 794.950 587.900 795.270 587.960 ;
        RECT 246.630 22.680 246.950 22.740 ;
        RECT 651.890 22.680 652.210 22.740 ;
        RECT 246.630 22.540 652.210 22.680 ;
        RECT 246.630 22.480 246.950 22.540 ;
        RECT 651.890 22.480 652.210 22.540 ;
      LAYER via ;
        RECT 1554.900 2896.500 1555.160 2896.760 ;
        RECT 787.160 2892.420 787.420 2892.680 ;
        RECT 883.760 2892.420 884.020 2892.680 ;
        RECT 980.360 2892.420 980.620 2892.680 ;
        RECT 1076.960 2892.420 1077.220 2892.680 ;
        RECT 1173.560 2892.420 1173.820 2892.680 ;
        RECT 1270.160 2892.420 1270.420 2892.680 ;
        RECT 1317.540 2892.420 1317.800 2892.680 ;
        RECT 1366.760 2892.420 1367.020 2892.680 ;
        RECT 772.440 2892.080 772.700 2892.340 ;
        RECT 786.240 2892.080 786.500 2892.340 ;
        RECT 821.200 2892.080 821.460 2892.340 ;
        RECT 869.040 2892.080 869.300 2892.340 ;
        RECT 882.840 2892.080 883.100 2892.340 ;
        RECT 917.800 2892.080 918.060 2892.340 ;
        RECT 965.640 2892.080 965.900 2892.340 ;
        RECT 979.440 2892.080 979.700 2892.340 ;
        RECT 1014.400 2892.080 1014.660 2892.340 ;
        RECT 1062.240 2892.080 1062.500 2892.340 ;
        RECT 1076.040 2892.080 1076.300 2892.340 ;
        RECT 1111.000 2892.080 1111.260 2892.340 ;
        RECT 1158.840 2892.080 1159.100 2892.340 ;
        RECT 1172.640 2892.080 1172.900 2892.340 ;
        RECT 1207.600 2892.080 1207.860 2892.340 ;
        RECT 1255.440 2892.080 1255.700 2892.340 ;
        RECT 1269.240 2892.080 1269.500 2892.340 ;
        RECT 1318.000 2892.080 1318.260 2892.340 ;
        RECT 1365.840 2892.080 1366.100 2892.340 ;
        RECT 1400.800 2892.080 1401.060 2892.340 ;
        RECT 1448.640 2892.080 1448.900 2892.340 ;
        RECT 1462.440 2892.080 1462.700 2892.340 ;
        RECT 1462.900 2892.080 1463.160 2892.340 ;
        RECT 651.920 2891.740 652.180 2892.000 ;
        RECT 689.640 2891.740 689.900 2892.000 ;
        RECT 690.560 2891.400 690.820 2891.660 ;
        RECT 724.600 2891.400 724.860 2891.660 ;
        RECT 821.200 2891.400 821.460 2891.660 ;
        RECT 869.040 2891.400 869.300 2891.660 ;
        RECT 917.800 2891.400 918.060 2891.660 ;
        RECT 965.640 2891.400 965.900 2891.660 ;
        RECT 1014.400 2891.400 1014.660 2891.660 ;
        RECT 1062.240 2891.400 1062.500 2891.660 ;
        RECT 1111.000 2891.400 1111.260 2891.660 ;
        RECT 1158.840 2891.400 1159.100 2891.660 ;
        RECT 1207.600 2891.400 1207.860 2891.660 ;
        RECT 1255.440 2891.400 1255.700 2891.660 ;
        RECT 1400.800 2891.400 1401.060 2891.660 ;
        RECT 1448.640 2891.400 1448.900 2891.660 ;
        RECT 724.600 2890.720 724.860 2890.980 ;
        RECT 772.440 2890.720 772.700 2890.980 ;
        RECT 446.760 2594.240 447.020 2594.500 ;
        RECT 612.820 2594.240 613.080 2594.500 ;
        RECT 614.200 2594.240 614.460 2594.500 ;
        RECT 648.700 2594.240 648.960 2594.500 ;
        RECT 648.700 2592.540 648.960 2592.800 ;
        RECT 651.920 2592.540 652.180 2592.800 ;
        RECT 644.100 1758.520 644.360 1758.780 ;
        RECT 648.700 1758.520 648.960 1758.780 ;
        RECT 651.920 1758.520 652.180 1758.780 ;
        RECT 651.920 1703.100 652.180 1703.360 ;
        RECT 1401.260 1703.100 1401.520 1703.360 ;
        RECT 1403.100 1703.100 1403.360 1703.360 ;
        RECT 1642.760 1703.100 1643.020 1703.360 ;
        RECT 1644.600 1703.100 1644.860 1703.360 ;
        RECT 1907.720 1703.100 1907.980 1703.360 ;
        RECT 651.920 588.240 652.180 588.500 ;
        RECT 794.980 587.900 795.240 588.160 ;
        RECT 246.660 22.480 246.920 22.740 ;
        RECT 651.920 22.480 652.180 22.740 ;
      LAYER met2 ;
        RECT 1554.900 2896.530 1555.160 2896.790 ;
        RECT 1556.210 2896.530 1556.490 2900.055 ;
        RECT 1554.900 2896.470 1556.490 2896.530 ;
        RECT 1554.960 2896.390 1556.490 2896.470 ;
        RECT 1556.210 2896.055 1556.490 2896.390 ;
        RECT 787.160 2892.450 787.420 2892.710 ;
        RECT 883.760 2892.450 884.020 2892.710 ;
        RECT 980.360 2892.450 980.620 2892.710 ;
        RECT 1076.960 2892.450 1077.220 2892.710 ;
        RECT 1173.560 2892.450 1173.820 2892.710 ;
        RECT 1270.160 2892.450 1270.420 2892.710 ;
        RECT 786.300 2892.390 787.420 2892.450 ;
        RECT 882.900 2892.390 884.020 2892.450 ;
        RECT 979.500 2892.390 980.620 2892.450 ;
        RECT 1076.100 2892.390 1077.220 2892.450 ;
        RECT 1172.700 2892.390 1173.820 2892.450 ;
        RECT 1269.300 2892.390 1270.420 2892.450 ;
        RECT 1317.540 2892.450 1317.800 2892.710 ;
        RECT 1366.760 2892.450 1367.020 2892.710 ;
        RECT 1317.540 2892.390 1318.200 2892.450 ;
        RECT 786.300 2892.370 787.360 2892.390 ;
        RECT 882.900 2892.370 883.960 2892.390 ;
        RECT 979.500 2892.370 980.560 2892.390 ;
        RECT 1076.100 2892.370 1077.160 2892.390 ;
        RECT 1172.700 2892.370 1173.760 2892.390 ;
        RECT 1269.300 2892.370 1270.360 2892.390 ;
        RECT 772.440 2892.050 772.700 2892.370 ;
        RECT 786.240 2892.310 787.360 2892.370 ;
        RECT 786.240 2892.050 786.500 2892.310 ;
        RECT 821.200 2892.050 821.460 2892.370 ;
        RECT 869.040 2892.050 869.300 2892.370 ;
        RECT 882.840 2892.310 883.960 2892.370 ;
        RECT 882.840 2892.050 883.100 2892.310 ;
        RECT 917.800 2892.050 918.060 2892.370 ;
        RECT 965.640 2892.050 965.900 2892.370 ;
        RECT 979.440 2892.310 980.560 2892.370 ;
        RECT 979.440 2892.050 979.700 2892.310 ;
        RECT 1014.400 2892.050 1014.660 2892.370 ;
        RECT 1062.240 2892.050 1062.500 2892.370 ;
        RECT 1076.040 2892.310 1077.160 2892.370 ;
        RECT 1076.040 2892.050 1076.300 2892.310 ;
        RECT 1111.000 2892.050 1111.260 2892.370 ;
        RECT 1158.840 2892.050 1159.100 2892.370 ;
        RECT 1172.640 2892.310 1173.760 2892.370 ;
        RECT 1172.640 2892.050 1172.900 2892.310 ;
        RECT 1207.600 2892.050 1207.860 2892.370 ;
        RECT 1255.440 2892.050 1255.700 2892.370 ;
        RECT 1269.240 2892.310 1270.360 2892.370 ;
        RECT 1317.600 2892.370 1318.200 2892.390 ;
        RECT 1365.900 2892.390 1367.020 2892.450 ;
        RECT 1365.900 2892.370 1366.960 2892.390 ;
        RECT 1462.500 2892.370 1463.100 2892.450 ;
        RECT 1317.600 2892.310 1318.260 2892.370 ;
        RECT 1269.240 2892.050 1269.500 2892.310 ;
        RECT 1318.000 2892.050 1318.260 2892.310 ;
        RECT 1365.840 2892.310 1366.960 2892.370 ;
        RECT 1365.840 2892.050 1366.100 2892.310 ;
        RECT 1400.800 2892.050 1401.060 2892.370 ;
        RECT 1448.640 2892.050 1448.900 2892.370 ;
        RECT 1462.440 2892.310 1463.160 2892.370 ;
        RECT 1462.440 2892.050 1462.700 2892.310 ;
        RECT 1462.900 2892.050 1463.160 2892.310 ;
        RECT 651.920 2891.710 652.180 2892.030 ;
        RECT 689.640 2891.770 689.900 2892.030 ;
        RECT 689.640 2891.710 690.760 2891.770 ;
        RECT 446.650 2600.660 446.930 2604.000 ;
        RECT 446.650 2600.000 446.960 2600.660 ;
        RECT 446.820 2594.530 446.960 2600.000 ;
        RECT 446.760 2594.210 447.020 2594.530 ;
        RECT 612.820 2594.210 613.080 2594.530 ;
        RECT 614.200 2594.210 614.460 2594.530 ;
        RECT 648.700 2594.210 648.960 2594.530 ;
        RECT 612.880 2593.930 613.020 2594.210 ;
        RECT 614.260 2593.930 614.400 2594.210 ;
        RECT 612.880 2593.790 614.400 2593.930 ;
        RECT 648.760 2592.830 648.900 2594.210 ;
        RECT 651.980 2592.830 652.120 2891.710 ;
        RECT 689.700 2891.690 690.760 2891.710 ;
        RECT 689.700 2891.630 690.820 2891.690 ;
        RECT 690.560 2891.370 690.820 2891.630 ;
        RECT 724.600 2891.370 724.860 2891.690 ;
        RECT 724.660 2891.010 724.800 2891.370 ;
        RECT 772.500 2891.010 772.640 2892.050 ;
        RECT 821.260 2891.690 821.400 2892.050 ;
        RECT 869.100 2891.690 869.240 2892.050 ;
        RECT 917.860 2891.690 918.000 2892.050 ;
        RECT 965.700 2891.690 965.840 2892.050 ;
        RECT 1014.460 2891.690 1014.600 2892.050 ;
        RECT 1062.300 2891.690 1062.440 2892.050 ;
        RECT 1111.060 2891.690 1111.200 2892.050 ;
        RECT 1158.900 2891.690 1159.040 2892.050 ;
        RECT 1207.660 2891.690 1207.800 2892.050 ;
        RECT 1255.500 2891.690 1255.640 2892.050 ;
        RECT 1400.860 2891.690 1401.000 2892.050 ;
        RECT 1448.700 2891.690 1448.840 2892.050 ;
        RECT 821.200 2891.370 821.460 2891.690 ;
        RECT 869.040 2891.370 869.300 2891.690 ;
        RECT 917.800 2891.370 918.060 2891.690 ;
        RECT 965.640 2891.370 965.900 2891.690 ;
        RECT 1014.400 2891.370 1014.660 2891.690 ;
        RECT 1062.240 2891.370 1062.500 2891.690 ;
        RECT 1111.000 2891.370 1111.260 2891.690 ;
        RECT 1158.840 2891.370 1159.100 2891.690 ;
        RECT 1207.600 2891.370 1207.860 2891.690 ;
        RECT 1255.440 2891.370 1255.700 2891.690 ;
        RECT 1400.800 2891.370 1401.060 2891.690 ;
        RECT 1448.640 2891.370 1448.900 2891.690 ;
        RECT 724.600 2890.690 724.860 2891.010 ;
        RECT 772.440 2890.690 772.700 2891.010 ;
        RECT 648.700 2592.510 648.960 2592.830 ;
        RECT 651.920 2592.510 652.180 2592.830 ;
        RECT 648.760 1758.810 648.900 2592.510 ;
        RECT 1907.710 1836.835 1907.990 1837.205 ;
        RECT 644.100 1758.490 644.360 1758.810 ;
        RECT 648.700 1758.490 648.960 1758.810 ;
        RECT 651.920 1758.490 652.180 1758.810 ;
        RECT 644.160 1754.925 644.300 1758.490 ;
        RECT 644.090 1754.555 644.370 1754.925 ;
        RECT 651.980 1703.390 652.120 1758.490 ;
        RECT 1401.320 1703.670 1403.300 1703.810 ;
        RECT 1401.320 1703.390 1401.460 1703.670 ;
        RECT 1403.160 1703.390 1403.300 1703.670 ;
        RECT 1642.820 1703.670 1644.800 1703.810 ;
        RECT 1642.820 1703.390 1642.960 1703.670 ;
        RECT 1644.660 1703.390 1644.800 1703.670 ;
        RECT 1907.780 1703.390 1907.920 1836.835 ;
        RECT 651.920 1703.070 652.180 1703.390 ;
        RECT 1401.260 1703.070 1401.520 1703.390 ;
        RECT 1403.100 1703.070 1403.360 1703.390 ;
        RECT 1642.760 1703.070 1643.020 1703.390 ;
        RECT 1644.600 1703.070 1644.860 1703.390 ;
        RECT 1907.720 1703.070 1907.980 1703.390 ;
        RECT 651.980 588.530 652.120 1703.070 ;
        RECT 796.590 600.170 796.870 604.000 ;
        RECT 795.040 600.030 796.870 600.170 ;
        RECT 651.920 588.210 652.180 588.530 ;
        RECT 651.980 22.770 652.120 588.210 ;
        RECT 795.040 588.190 795.180 600.030 ;
        RECT 796.590 600.000 796.870 600.030 ;
        RECT 794.980 587.870 795.240 588.190 ;
        RECT 246.660 22.450 246.920 22.770 ;
        RECT 651.920 22.450 652.180 22.770 ;
        RECT 246.720 2.400 246.860 22.450 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 1907.710 1836.880 1907.990 1837.160 ;
        RECT 644.090 1754.600 644.370 1754.880 ;
      LAYER met3 ;
        RECT 1920.000 1838.440 1924.000 1839.040 ;
        RECT 1907.685 1837.170 1908.015 1837.185 ;
        RECT 1920.350 1837.170 1920.650 1838.440 ;
        RECT 1907.685 1836.870 1920.650 1837.170 ;
        RECT 1907.685 1836.855 1908.015 1836.870 ;
        RECT 627.030 1754.890 631.030 1755.040 ;
        RECT 644.065 1754.890 644.395 1754.905 ;
        RECT 627.030 1754.590 644.395 1754.890 ;
        RECT 627.030 1754.440 631.030 1754.590 ;
        RECT 644.065 1754.575 644.395 1754.590 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 613.710 2900.780 614.030 2900.840 ;
        RECT 1577.410 2900.780 1577.730 2900.840 ;
        RECT 613.710 2900.640 1577.730 2900.780 ;
        RECT 613.710 2900.580 614.030 2900.640 ;
        RECT 1577.410 2900.580 1577.730 2900.640 ;
        RECT 638.550 2594.100 638.870 2594.160 ;
        RECT 614.260 2593.960 638.870 2594.100 ;
        RECT 496.410 2593.760 496.730 2593.820 ;
        RECT 458.780 2593.620 496.730 2593.760 ;
        RECT 432.930 2593.420 433.250 2593.480 ;
        RECT 432.930 2593.280 447.880 2593.420 ;
        RECT 432.930 2593.220 433.250 2593.280 ;
        RECT 447.740 2593.080 447.880 2593.280 ;
        RECT 458.780 2593.080 458.920 2593.620 ;
        RECT 496.410 2593.560 496.730 2593.620 ;
        RECT 496.870 2593.760 497.190 2593.820 ;
        RECT 612.330 2593.760 612.650 2593.820 ;
        RECT 614.260 2593.760 614.400 2593.960 ;
        RECT 638.550 2593.900 638.870 2593.960 ;
        RECT 496.870 2593.620 524.700 2593.760 ;
        RECT 611.895 2593.620 614.400 2593.760 ;
        RECT 496.870 2593.560 497.190 2593.620 ;
        RECT 524.560 2593.420 524.700 2593.620 ;
        RECT 612.330 2593.560 612.650 2593.620 ;
        RECT 545.170 2593.420 545.490 2593.480 ;
        RECT 524.560 2593.280 545.490 2593.420 ;
        RECT 545.170 2593.220 545.490 2593.280 ;
        RECT 545.630 2593.420 545.950 2593.480 ;
        RECT 545.630 2593.280 579.900 2593.420 ;
        RECT 545.630 2593.220 545.950 2593.280 ;
        RECT 447.740 2592.940 458.920 2593.080 ;
        RECT 579.760 2593.080 579.900 2593.280 ;
        RECT 612.420 2593.080 612.560 2593.560 ;
        RECT 579.760 2592.940 612.560 2593.080 ;
        RECT 638.550 1703.640 638.870 1703.700 ;
        RECT 1908.150 1703.640 1908.470 1703.700 ;
        RECT 638.550 1703.500 1908.470 1703.640 ;
        RECT 638.550 1703.440 638.870 1703.500 ;
        RECT 1908.150 1703.440 1908.470 1703.500 ;
        RECT 613.250 1689.360 613.570 1689.420 ;
        RECT 638.550 1689.360 638.870 1689.420 ;
        RECT 613.250 1689.220 638.870 1689.360 ;
        RECT 613.250 1689.160 613.570 1689.220 ;
        RECT 638.550 1689.160 638.870 1689.220 ;
        RECT 612.790 1607.760 613.110 1607.820 ;
        RECT 613.710 1607.760 614.030 1607.820 ;
        RECT 612.790 1607.620 614.030 1607.760 ;
        RECT 612.790 1607.560 613.110 1607.620 ;
        RECT 613.710 1607.560 614.030 1607.620 ;
        RECT 612.330 1593.820 612.650 1593.880 ;
        RECT 613.710 1593.820 614.030 1593.880 ;
        RECT 612.330 1593.680 614.030 1593.820 ;
        RECT 612.330 1593.620 612.650 1593.680 ;
        RECT 613.710 1593.620 614.030 1593.680 ;
        RECT 612.330 1545.880 612.650 1545.940 ;
        RECT 613.250 1545.880 613.570 1545.940 ;
        RECT 612.330 1545.740 613.570 1545.880 ;
        RECT 612.330 1545.680 612.650 1545.740 ;
        RECT 613.250 1545.680 613.570 1545.740 ;
        RECT 612.790 1124.620 613.110 1124.680 ;
        RECT 613.710 1124.620 614.030 1124.680 ;
        RECT 612.790 1124.480 614.030 1124.620 ;
        RECT 612.790 1124.420 613.110 1124.480 ;
        RECT 613.710 1124.420 614.030 1124.480 ;
        RECT 613.710 1077.020 614.030 1077.080 ;
        RECT 613.340 1076.880 614.030 1077.020 ;
        RECT 613.340 1076.400 613.480 1076.880 ;
        RECT 613.710 1076.820 614.030 1076.880 ;
        RECT 613.250 1076.140 613.570 1076.400 ;
        RECT 613.250 1028.740 613.570 1028.800 ;
        RECT 612.880 1028.600 613.570 1028.740 ;
        RECT 612.880 1028.120 613.020 1028.600 ;
        RECT 613.250 1028.540 613.570 1028.600 ;
        RECT 612.790 1027.860 613.110 1028.120 ;
        RECT 611.870 1007.320 612.190 1007.380 ;
        RECT 612.790 1007.320 613.110 1007.380 ;
        RECT 611.870 1007.180 613.110 1007.320 ;
        RECT 611.870 1007.120 612.190 1007.180 ;
        RECT 612.790 1007.120 613.110 1007.180 ;
        RECT 611.870 979.100 612.190 979.160 ;
        RECT 613.250 979.100 613.570 979.160 ;
        RECT 611.870 978.960 613.570 979.100 ;
        RECT 611.870 978.900 612.190 978.960 ;
        RECT 613.250 978.900 613.570 978.960 ;
        RECT 613.710 883.560 614.030 883.620 ;
        RECT 613.340 883.420 614.030 883.560 ;
        RECT 613.340 882.940 613.480 883.420 ;
        RECT 613.710 883.360 614.030 883.420 ;
        RECT 613.250 882.680 613.570 882.940 ;
        RECT 612.790 821.000 613.110 821.060 ;
        RECT 613.710 821.000 614.030 821.060 ;
        RECT 612.790 820.860 614.030 821.000 ;
        RECT 612.790 820.800 613.110 820.860 ;
        RECT 613.710 820.800 614.030 820.860 ;
        RECT 611.410 772.380 611.730 772.440 ;
        RECT 613.250 772.380 613.570 772.440 ;
        RECT 611.410 772.240 613.570 772.380 ;
        RECT 611.410 772.180 611.730 772.240 ;
        RECT 613.250 772.180 613.570 772.240 ;
        RECT 614.170 589.120 614.490 589.180 ;
        RECT 793.570 589.120 793.890 589.180 ;
        RECT 614.170 588.980 793.890 589.120 ;
        RECT 614.170 588.920 614.490 588.980 ;
        RECT 793.570 588.920 793.890 588.980 ;
        RECT 610.490 586.740 610.810 586.800 ;
        RECT 613.250 586.740 613.570 586.800 ;
        RECT 610.490 586.600 613.570 586.740 ;
        RECT 610.490 586.540 610.810 586.600 ;
        RECT 613.250 586.540 613.570 586.600 ;
        RECT 264.110 22.340 264.430 22.400 ;
        RECT 610.490 22.340 610.810 22.400 ;
        RECT 264.110 22.200 610.810 22.340 ;
        RECT 264.110 22.140 264.430 22.200 ;
        RECT 610.490 22.140 610.810 22.200 ;
      LAYER via ;
        RECT 613.740 2900.580 614.000 2900.840 ;
        RECT 1577.440 2900.580 1577.700 2900.840 ;
        RECT 432.960 2593.220 433.220 2593.480 ;
        RECT 496.440 2593.560 496.700 2593.820 ;
        RECT 496.900 2593.560 497.160 2593.820 ;
        RECT 612.360 2593.560 612.620 2593.820 ;
        RECT 638.580 2593.900 638.840 2594.160 ;
        RECT 545.200 2593.220 545.460 2593.480 ;
        RECT 545.660 2593.220 545.920 2593.480 ;
        RECT 638.580 1703.440 638.840 1703.700 ;
        RECT 1908.180 1703.440 1908.440 1703.700 ;
        RECT 613.280 1689.160 613.540 1689.420 ;
        RECT 638.580 1689.160 638.840 1689.420 ;
        RECT 612.820 1607.560 613.080 1607.820 ;
        RECT 613.740 1607.560 614.000 1607.820 ;
        RECT 612.360 1593.620 612.620 1593.880 ;
        RECT 613.740 1593.620 614.000 1593.880 ;
        RECT 612.360 1545.680 612.620 1545.940 ;
        RECT 613.280 1545.680 613.540 1545.940 ;
        RECT 612.820 1124.420 613.080 1124.680 ;
        RECT 613.740 1124.420 614.000 1124.680 ;
        RECT 613.740 1076.820 614.000 1077.080 ;
        RECT 613.280 1076.140 613.540 1076.400 ;
        RECT 613.280 1028.540 613.540 1028.800 ;
        RECT 612.820 1027.860 613.080 1028.120 ;
        RECT 611.900 1007.120 612.160 1007.380 ;
        RECT 612.820 1007.120 613.080 1007.380 ;
        RECT 611.900 978.900 612.160 979.160 ;
        RECT 613.280 978.900 613.540 979.160 ;
        RECT 613.740 883.360 614.000 883.620 ;
        RECT 613.280 882.680 613.540 882.940 ;
        RECT 612.820 820.800 613.080 821.060 ;
        RECT 613.740 820.800 614.000 821.060 ;
        RECT 611.440 772.180 611.700 772.440 ;
        RECT 613.280 772.180 613.540 772.440 ;
        RECT 614.200 588.920 614.460 589.180 ;
        RECT 793.600 588.920 793.860 589.180 ;
        RECT 610.520 586.540 610.780 586.800 ;
        RECT 613.280 586.540 613.540 586.800 ;
        RECT 264.140 22.140 264.400 22.400 ;
        RECT 610.520 22.140 610.780 22.400 ;
      LAYER met2 ;
        RECT 613.740 2900.550 614.000 2900.870 ;
        RECT 1577.440 2900.550 1577.700 2900.870 ;
        RECT 432.850 2600.660 433.130 2604.000 ;
        RECT 432.850 2600.000 433.160 2600.660 ;
        RECT 433.020 2593.510 433.160 2600.000 ;
        RECT 613.800 2598.690 613.940 2900.550 ;
        RECT 1577.500 2900.055 1577.640 2900.550 ;
        RECT 1577.370 2896.055 1577.650 2900.055 ;
        RECT 612.420 2598.550 613.940 2598.690 ;
        RECT 496.500 2593.850 497.100 2593.930 ;
        RECT 612.420 2593.850 612.560 2598.550 ;
        RECT 638.580 2593.870 638.840 2594.190 ;
        RECT 496.440 2593.790 497.160 2593.850 ;
        RECT 496.440 2593.530 496.700 2593.790 ;
        RECT 496.900 2593.530 497.160 2593.790 ;
        RECT 612.360 2593.530 612.620 2593.850 ;
        RECT 432.960 2593.190 433.220 2593.510 ;
        RECT 545.200 2593.250 545.460 2593.510 ;
        RECT 545.660 2593.250 545.920 2593.510 ;
        RECT 545.200 2593.190 545.920 2593.250 ;
        RECT 545.260 2593.110 545.860 2593.190 ;
        RECT 613.090 1700.410 613.370 1704.000 ;
        RECT 638.640 1703.730 638.780 2593.870 ;
        RECT 1908.170 1801.475 1908.450 1801.845 ;
        RECT 1908.240 1703.730 1908.380 1801.475 ;
        RECT 638.580 1703.410 638.840 1703.730 ;
        RECT 1908.180 1703.410 1908.440 1703.730 ;
        RECT 613.090 1700.000 613.480 1700.410 ;
        RECT 613.340 1689.450 613.480 1700.000 ;
        RECT 638.640 1689.450 638.780 1703.410 ;
        RECT 613.280 1689.130 613.540 1689.450 ;
        RECT 638.580 1689.130 638.840 1689.450 ;
        RECT 613.340 1607.930 613.480 1689.130 ;
        RECT 612.880 1607.850 613.480 1607.930 ;
        RECT 612.820 1607.790 613.480 1607.850 ;
        RECT 612.820 1607.530 613.080 1607.790 ;
        RECT 613.740 1607.530 614.000 1607.850 ;
        RECT 612.880 1607.375 613.020 1607.530 ;
        RECT 613.800 1593.910 613.940 1607.530 ;
        RECT 612.360 1593.590 612.620 1593.910 ;
        RECT 613.740 1593.590 614.000 1593.910 ;
        RECT 612.420 1545.970 612.560 1593.590 ;
        RECT 612.360 1545.650 612.620 1545.970 ;
        RECT 613.280 1545.650 613.540 1545.970 ;
        RECT 613.340 1511.370 613.480 1545.650 ;
        RECT 612.880 1511.230 613.480 1511.370 ;
        RECT 612.880 1510.690 613.020 1511.230 ;
        RECT 612.880 1510.550 613.480 1510.690 ;
        RECT 613.340 1463.090 613.480 1510.550 ;
        RECT 613.340 1462.950 613.940 1463.090 ;
        RECT 613.800 1462.410 613.940 1462.950 ;
        RECT 613.340 1462.270 613.940 1462.410 ;
        RECT 613.340 1414.810 613.480 1462.270 ;
        RECT 612.880 1414.670 613.480 1414.810 ;
        RECT 612.880 1414.130 613.020 1414.670 ;
        RECT 612.880 1413.990 613.480 1414.130 ;
        RECT 613.340 1366.530 613.480 1413.990 ;
        RECT 613.340 1366.390 613.940 1366.530 ;
        RECT 613.800 1365.850 613.940 1366.390 ;
        RECT 613.340 1365.710 613.940 1365.850 ;
        RECT 613.340 1318.250 613.480 1365.710 ;
        RECT 612.880 1318.110 613.480 1318.250 ;
        RECT 612.880 1317.570 613.020 1318.110 ;
        RECT 612.880 1317.430 613.480 1317.570 ;
        RECT 613.340 1269.970 613.480 1317.430 ;
        RECT 613.340 1269.830 613.940 1269.970 ;
        RECT 613.800 1269.290 613.940 1269.830 ;
        RECT 613.340 1269.150 613.940 1269.290 ;
        RECT 613.340 1221.690 613.480 1269.150 ;
        RECT 612.880 1221.550 613.480 1221.690 ;
        RECT 612.880 1221.010 613.020 1221.550 ;
        RECT 612.880 1220.870 613.480 1221.010 ;
        RECT 613.340 1173.410 613.480 1220.870 ;
        RECT 613.340 1173.270 613.940 1173.410 ;
        RECT 613.800 1172.730 613.940 1173.270 ;
        RECT 613.340 1172.590 613.940 1172.730 ;
        RECT 613.340 1125.130 613.480 1172.590 ;
        RECT 612.880 1124.990 613.480 1125.130 ;
        RECT 612.880 1124.710 613.020 1124.990 ;
        RECT 612.820 1124.390 613.080 1124.710 ;
        RECT 613.740 1124.390 614.000 1124.710 ;
        RECT 613.800 1077.110 613.940 1124.390 ;
        RECT 613.740 1076.790 614.000 1077.110 ;
        RECT 613.280 1076.110 613.540 1076.430 ;
        RECT 613.340 1028.830 613.480 1076.110 ;
        RECT 613.280 1028.510 613.540 1028.830 ;
        RECT 612.820 1027.830 613.080 1028.150 ;
        RECT 612.880 1007.410 613.020 1027.830 ;
        RECT 611.900 1007.090 612.160 1007.410 ;
        RECT 612.820 1007.090 613.080 1007.410 ;
        RECT 611.960 979.190 612.100 1007.090 ;
        RECT 611.900 978.870 612.160 979.190 ;
        RECT 613.280 978.870 613.540 979.190 ;
        RECT 613.340 932.010 613.480 978.870 ;
        RECT 612.880 931.870 613.480 932.010 ;
        RECT 612.880 931.330 613.020 931.870 ;
        RECT 612.880 931.190 613.480 931.330 ;
        RECT 613.340 917.730 613.480 931.190 ;
        RECT 613.340 917.590 613.940 917.730 ;
        RECT 613.800 883.650 613.940 917.590 ;
        RECT 613.740 883.330 614.000 883.650 ;
        RECT 613.280 882.650 613.540 882.970 ;
        RECT 613.340 835.450 613.480 882.650 ;
        RECT 612.880 835.310 613.480 835.450 ;
        RECT 612.880 821.090 613.020 835.310 ;
        RECT 612.820 820.770 613.080 821.090 ;
        RECT 613.740 820.770 614.000 821.090 ;
        RECT 613.800 785.810 613.940 820.770 ;
        RECT 613.340 785.670 613.940 785.810 ;
        RECT 613.340 772.470 613.480 785.670 ;
        RECT 611.440 772.150 611.700 772.470 ;
        RECT 613.280 772.150 613.540 772.470 ;
        RECT 611.500 724.725 611.640 772.150 ;
        RECT 611.430 724.355 611.710 724.725 ;
        RECT 612.350 724.355 612.630 724.725 ;
        RECT 612.420 689.250 612.560 724.355 ;
        RECT 612.420 689.110 613.480 689.250 ;
        RECT 613.340 589.290 613.480 689.110 ;
        RECT 805.790 600.170 806.070 604.000 ;
        RECT 804.240 600.030 806.070 600.170 ;
        RECT 804.240 589.405 804.380 600.030 ;
        RECT 805.790 600.000 806.070 600.030 ;
        RECT 613.340 589.210 614.400 589.290 ;
        RECT 613.340 589.150 614.460 589.210 ;
        RECT 613.340 586.830 613.480 589.150 ;
        RECT 614.200 588.890 614.460 589.150 ;
        RECT 793.590 589.035 793.870 589.405 ;
        RECT 804.170 589.035 804.450 589.405 ;
        RECT 793.600 588.890 793.860 589.035 ;
        RECT 610.520 586.510 610.780 586.830 ;
        RECT 613.280 586.510 613.540 586.830 ;
        RECT 610.580 22.430 610.720 586.510 ;
        RECT 264.140 22.110 264.400 22.430 ;
        RECT 610.520 22.110 610.780 22.430 ;
        RECT 264.200 2.400 264.340 22.110 ;
        RECT 263.990 -4.800 264.550 2.400 ;
      LAYER via2 ;
        RECT 1908.170 1801.520 1908.450 1801.800 ;
        RECT 611.430 724.400 611.710 724.680 ;
        RECT 612.350 724.400 612.630 724.680 ;
        RECT 793.590 589.080 793.870 589.360 ;
        RECT 804.170 589.080 804.450 589.360 ;
      LAYER met3 ;
        RECT 1920.000 1804.440 1924.000 1805.040 ;
        RECT 1908.145 1801.810 1908.475 1801.825 ;
        RECT 1920.350 1801.810 1920.650 1804.440 ;
        RECT 1908.145 1801.510 1920.650 1801.810 ;
        RECT 1908.145 1801.495 1908.475 1801.510 ;
        RECT 611.405 724.690 611.735 724.705 ;
        RECT 612.325 724.690 612.655 724.705 ;
        RECT 611.405 724.390 612.655 724.690 ;
        RECT 611.405 724.375 611.735 724.390 ;
        RECT 612.325 724.375 612.655 724.390 ;
        RECT 793.565 589.370 793.895 589.385 ;
        RECT 804.145 589.370 804.475 589.385 ;
        RECT 793.565 589.070 804.475 589.370 ;
        RECT 793.565 589.055 793.895 589.070 ;
        RECT 804.145 589.055 804.475 589.070 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 2767.160 562.050 2767.220 ;
        RECT 580.130 2767.160 580.450 2767.220 ;
        RECT 561.730 2767.020 580.450 2767.160 ;
        RECT 561.730 2766.960 562.050 2767.020 ;
        RECT 580.130 2766.960 580.450 2767.020 ;
        RECT 580.130 2490.400 580.450 2490.460 ;
        RECT 1736.570 2490.400 1736.890 2490.460 ;
        RECT 580.130 2490.260 1736.890 2490.400 ;
        RECT 580.130 2490.200 580.450 2490.260 ;
        RECT 1736.570 2490.200 1736.890 2490.260 ;
        RECT 544.710 2488.020 545.030 2488.080 ;
        RECT 580.130 2488.020 580.450 2488.080 ;
        RECT 544.710 2487.880 580.450 2488.020 ;
        RECT 544.710 2487.820 545.030 2487.880 ;
        RECT 580.130 2487.820 580.450 2487.880 ;
        RECT 483.070 1979.380 483.390 1979.440 ;
        RECT 418.760 1979.240 483.390 1979.380 ;
        RECT 357.950 1978.700 358.270 1978.760 ;
        RECT 418.760 1978.700 418.900 1979.240 ;
        RECT 483.070 1979.180 483.390 1979.240 ;
        RECT 357.950 1978.560 418.900 1978.700 ;
        RECT 496.410 1978.700 496.730 1978.760 ;
        RECT 544.710 1978.700 545.030 1978.760 ;
        RECT 629.350 1978.700 629.670 1978.760 ;
        RECT 496.410 1978.560 629.670 1978.700 ;
        RECT 357.950 1978.500 358.270 1978.560 ;
        RECT 496.410 1978.500 496.730 1978.560 ;
        RECT 544.710 1978.500 545.030 1978.560 ;
        RECT 629.350 1978.500 629.670 1978.560 ;
        RECT 282.510 591.500 282.830 591.560 ;
        RECT 629.350 591.500 629.670 591.560 ;
        RECT 282.510 591.360 629.670 591.500 ;
        RECT 282.510 591.300 282.830 591.360 ;
        RECT 629.350 591.300 629.670 591.360 ;
        RECT 629.350 590.480 629.670 590.540 ;
        RECT 664.310 590.480 664.630 590.540 ;
        RECT 629.350 590.340 664.630 590.480 ;
        RECT 629.350 590.280 629.670 590.340 ;
        RECT 664.310 590.280 664.630 590.340 ;
        RECT 665.230 588.780 665.550 588.840 ;
        RECT 794.030 588.780 794.350 588.840 ;
        RECT 665.230 588.640 794.350 588.780 ;
        RECT 665.230 588.580 665.550 588.640 ;
        RECT 794.030 588.580 794.350 588.640 ;
        RECT 794.490 588.780 794.810 588.840 ;
        RECT 813.350 588.780 813.670 588.840 ;
        RECT 794.490 588.640 813.670 588.780 ;
        RECT 794.490 588.580 794.810 588.640 ;
        RECT 813.350 588.580 813.670 588.640 ;
      LAYER via ;
        RECT 561.760 2766.960 562.020 2767.220 ;
        RECT 580.160 2766.960 580.420 2767.220 ;
        RECT 580.160 2490.200 580.420 2490.460 ;
        RECT 1736.600 2490.200 1736.860 2490.460 ;
        RECT 544.740 2487.820 545.000 2488.080 ;
        RECT 580.160 2487.820 580.420 2488.080 ;
        RECT 357.980 1978.500 358.240 1978.760 ;
        RECT 483.100 1979.180 483.360 1979.440 ;
        RECT 496.440 1978.500 496.700 1978.760 ;
        RECT 544.740 1978.500 545.000 1978.760 ;
        RECT 629.380 1978.500 629.640 1978.760 ;
        RECT 282.540 591.300 282.800 591.560 ;
        RECT 629.380 591.300 629.640 591.560 ;
        RECT 629.380 590.280 629.640 590.540 ;
        RECT 664.340 590.280 664.600 590.540 ;
        RECT 665.260 588.580 665.520 588.840 ;
        RECT 794.060 588.580 794.320 588.840 ;
        RECT 794.520 588.580 794.780 588.840 ;
        RECT 813.380 588.580 813.640 588.840 ;
      LAYER met2 ;
        RECT 561.760 2766.930 562.020 2767.250 ;
        RECT 580.160 2766.930 580.420 2767.250 ;
        RECT 561.820 2759.520 561.960 2766.930 ;
        RECT 561.650 2759.100 561.960 2759.520 ;
        RECT 561.650 2755.520 561.930 2759.100 ;
        RECT 580.220 2490.490 580.360 2766.930 ;
        RECT 1736.530 2500.000 1736.810 2504.000 ;
        RECT 1736.660 2490.490 1736.800 2500.000 ;
        RECT 580.160 2490.170 580.420 2490.490 ;
        RECT 1736.600 2490.170 1736.860 2490.490 ;
        RECT 580.220 2488.110 580.360 2490.170 ;
        RECT 544.740 2487.790 545.000 2488.110 ;
        RECT 580.160 2487.790 580.420 2488.110 ;
        RECT 483.100 1979.325 483.360 1979.470 ;
        RECT 483.090 1978.955 483.370 1979.325 ;
        RECT 496.430 1978.955 496.710 1979.325 ;
        RECT 496.500 1978.790 496.640 1978.955 ;
        RECT 544.800 1978.790 544.940 2487.790 ;
        RECT 357.980 1978.470 358.240 1978.790 ;
        RECT 496.440 1978.470 496.700 1978.790 ;
        RECT 544.740 1978.470 545.000 1978.790 ;
        RECT 629.380 1978.470 629.640 1978.790 ;
        RECT 358.040 1814.765 358.180 1978.470 ;
        RECT 357.970 1814.395 358.250 1814.765 ;
        RECT 629.440 591.590 629.580 1978.470 ;
        RECT 814.990 600.170 815.270 604.000 ;
        RECT 813.440 600.030 815.270 600.170 ;
        RECT 282.540 591.270 282.800 591.590 ;
        RECT 629.380 591.270 629.640 591.590 ;
        RECT 282.600 3.130 282.740 591.270 ;
        RECT 629.440 590.570 629.580 591.270 ;
        RECT 629.380 590.250 629.640 590.570 ;
        RECT 664.340 590.250 664.600 590.570 ;
        RECT 664.400 589.970 664.540 590.250 ;
        RECT 664.400 589.830 665.460 589.970 ;
        RECT 665.320 588.870 665.460 589.830 ;
        RECT 813.440 588.870 813.580 600.030 ;
        RECT 814.990 600.000 815.270 600.030 ;
        RECT 665.260 588.550 665.520 588.870 ;
        RECT 794.060 588.780 794.320 588.870 ;
        RECT 794.520 588.780 794.780 588.870 ;
        RECT 794.060 588.640 794.780 588.780 ;
        RECT 794.060 588.550 794.320 588.640 ;
        RECT 794.520 588.550 794.780 588.640 ;
        RECT 813.380 588.550 813.640 588.870 ;
        RECT 282.140 2.990 282.740 3.130 ;
        RECT 282.140 2.400 282.280 2.990 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 483.090 1979.000 483.370 1979.280 ;
        RECT 496.430 1979.000 496.710 1979.280 ;
        RECT 357.970 1814.440 358.250 1814.720 ;
      LAYER met3 ;
        RECT 483.065 1979.290 483.395 1979.305 ;
        RECT 496.405 1979.290 496.735 1979.305 ;
        RECT 483.065 1978.990 496.735 1979.290 ;
        RECT 483.065 1978.975 483.395 1978.990 ;
        RECT 496.405 1978.975 496.735 1978.990 ;
        RECT 357.945 1814.730 358.275 1814.745 ;
        RECT 360.000 1814.730 364.000 1814.880 ;
        RECT 357.945 1814.430 364.000 1814.730 ;
        RECT 357.945 1814.415 358.275 1814.430 ;
        RECT 360.000 1814.280 364.000 1814.430 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.970 2487.340 559.290 2487.400 ;
        RECT 629.810 2487.340 630.130 2487.400 ;
        RECT 1863.530 2487.340 1863.850 2487.400 ;
        RECT 558.970 2487.200 1863.850 2487.340 ;
        RECT 558.970 2487.140 559.290 2487.200 ;
        RECT 629.810 2487.140 630.130 2487.200 ;
        RECT 1863.530 2487.140 1863.850 2487.200 ;
        RECT 413.610 1683.580 413.930 1683.640 ;
        RECT 629.810 1683.580 630.130 1683.640 ;
        RECT 413.610 1683.440 630.130 1683.580 ;
        RECT 413.610 1683.380 413.930 1683.440 ;
        RECT 629.810 1683.380 630.130 1683.440 ;
        RECT 413.610 592.520 413.930 592.580 ;
        RECT 822.550 592.520 822.870 592.580 ;
        RECT 413.610 592.380 822.870 592.520 ;
        RECT 413.610 592.320 413.930 592.380 ;
        RECT 822.550 592.320 822.870 592.380 ;
        RECT 303.210 590.140 303.530 590.200 ;
        RECT 413.610 590.140 413.930 590.200 ;
        RECT 303.210 590.000 413.930 590.140 ;
        RECT 303.210 589.940 303.530 590.000 ;
        RECT 413.610 589.940 413.930 590.000 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 559.000 2487.140 559.260 2487.400 ;
        RECT 629.840 2487.140 630.100 2487.400 ;
        RECT 1863.560 2487.140 1863.820 2487.400 ;
        RECT 413.640 1683.380 413.900 1683.640 ;
        RECT 629.840 1683.380 630.100 1683.640 ;
        RECT 413.640 592.320 413.900 592.580 ;
        RECT 822.580 592.320 822.840 592.580 ;
        RECT 303.240 589.940 303.500 590.200 ;
        RECT 413.640 589.940 413.900 590.200 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 562.570 2600.730 562.850 2604.000 ;
        RECT 559.060 2600.590 562.850 2600.730 ;
        RECT 559.060 2487.430 559.200 2600.590 ;
        RECT 562.570 2600.000 562.850 2600.590 ;
        RECT 1863.490 2500.000 1863.770 2504.000 ;
        RECT 1863.620 2487.430 1863.760 2500.000 ;
        RECT 559.000 2487.110 559.260 2487.430 ;
        RECT 629.840 2487.110 630.100 2487.430 ;
        RECT 1863.560 2487.110 1863.820 2487.430 ;
        RECT 412.530 1700.410 412.810 1704.000 ;
        RECT 412.530 1700.270 413.840 1700.410 ;
        RECT 412.530 1700.000 412.810 1700.270 ;
        RECT 413.700 1683.670 413.840 1700.270 ;
        RECT 629.900 1683.670 630.040 2487.110 ;
        RECT 413.640 1683.350 413.900 1683.670 ;
        RECT 629.840 1683.350 630.100 1683.670 ;
        RECT 413.700 592.610 413.840 1683.350 ;
        RECT 824.190 600.170 824.470 604.000 ;
        RECT 822.640 600.030 824.470 600.170 ;
        RECT 822.640 592.610 822.780 600.030 ;
        RECT 824.190 600.000 824.470 600.030 ;
        RECT 413.640 592.290 413.900 592.610 ;
        RECT 822.580 592.290 822.840 592.610 ;
        RECT 413.700 590.230 413.840 592.290 ;
        RECT 303.240 589.910 303.500 590.230 ;
        RECT 413.640 589.910 413.900 590.230 ;
        RECT 303.300 16.990 303.440 589.910 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 646.370 2899.080 646.690 2899.140 ;
        RECT 1821.210 2899.080 1821.530 2899.140 ;
        RECT 646.370 2898.940 1821.530 2899.080 ;
        RECT 646.370 2898.880 646.690 2898.940 ;
        RECT 1821.210 2898.880 1821.530 2898.940 ;
        RECT 642.690 2626.060 643.010 2626.120 ;
        RECT 646.370 2626.060 646.690 2626.120 ;
        RECT 642.690 2625.920 646.690 2626.060 ;
        RECT 642.690 2625.860 643.010 2625.920 ;
        RECT 646.370 2625.860 646.690 2625.920 ;
        RECT 593.010 2625.380 593.330 2625.440 ;
        RECT 642.690 2625.380 643.010 2625.440 ;
        RECT 593.010 2625.240 643.010 2625.380 ;
        RECT 593.010 2625.180 593.330 2625.240 ;
        RECT 642.690 2625.180 643.010 2625.240 ;
        RECT 666.610 588.440 666.930 588.500 ;
        RECT 793.340 588.440 793.660 588.500 ;
        RECT 666.610 588.300 793.660 588.440 ;
        RECT 666.610 588.240 666.930 588.300 ;
        RECT 793.340 588.240 793.660 588.300 ;
        RECT 645.450 587.080 645.770 587.140 ;
        RECT 666.610 587.080 666.930 587.140 ;
        RECT 645.450 586.940 666.930 587.080 ;
        RECT 645.450 586.880 645.770 586.940 ;
        RECT 666.610 586.880 666.930 586.940 ;
        RECT 317.930 36.280 318.250 36.340 ;
        RECT 645.450 36.280 645.770 36.340 ;
        RECT 317.930 36.140 645.770 36.280 ;
        RECT 317.930 36.080 318.250 36.140 ;
        RECT 645.450 36.080 645.770 36.140 ;
      LAYER via ;
        RECT 646.400 2898.880 646.660 2899.140 ;
        RECT 1821.240 2898.880 1821.500 2899.140 ;
        RECT 642.720 2625.860 642.980 2626.120 ;
        RECT 646.400 2625.860 646.660 2626.120 ;
        RECT 593.040 2625.180 593.300 2625.440 ;
        RECT 642.720 2625.180 642.980 2625.440 ;
        RECT 666.640 588.240 666.900 588.500 ;
        RECT 793.370 588.240 793.630 588.500 ;
        RECT 645.480 586.880 645.740 587.140 ;
        RECT 666.640 586.880 666.900 587.140 ;
        RECT 317.960 36.080 318.220 36.340 ;
        RECT 645.480 36.080 645.740 36.340 ;
      LAYER met2 ;
        RECT 1822.090 2899.250 1822.370 2900.055 ;
        RECT 1821.300 2899.170 1822.370 2899.250 ;
        RECT 646.400 2898.850 646.660 2899.170 ;
        RECT 1821.240 2899.110 1822.370 2899.170 ;
        RECT 1821.240 2898.850 1821.500 2899.110 ;
        RECT 646.460 2626.150 646.600 2898.850 ;
        RECT 1822.090 2896.055 1822.370 2899.110 ;
        RECT 593.030 2625.635 593.310 2626.005 ;
        RECT 642.720 2625.830 642.980 2626.150 ;
        RECT 646.400 2625.830 646.660 2626.150 ;
        RECT 593.100 2625.470 593.240 2625.635 ;
        RECT 642.780 2625.470 642.920 2625.830 ;
        RECT 593.040 2625.150 593.300 2625.470 ;
        RECT 642.720 2625.150 642.980 2625.470 ;
        RECT 642.780 1939.885 642.920 2625.150 ;
        RECT 642.710 1939.515 642.990 1939.885 ;
        RECT 645.470 1939.515 645.750 1939.885 ;
        RECT 645.540 587.170 645.680 1939.515 ;
        RECT 833.390 600.170 833.670 604.000 ;
        RECT 831.840 600.030 833.670 600.170 ;
        RECT 666.640 588.210 666.900 588.530 ;
        RECT 793.370 588.210 793.630 588.530 ;
        RECT 666.700 587.170 666.840 588.210 ;
        RECT 793.430 588.045 793.570 588.210 ;
        RECT 831.840 588.045 831.980 600.030 ;
        RECT 833.390 600.000 833.670 600.030 ;
        RECT 793.360 587.675 793.640 588.045 ;
        RECT 831.770 587.675 832.050 588.045 ;
        RECT 645.480 586.850 645.740 587.170 ;
        RECT 666.640 586.850 666.900 587.170 ;
        RECT 645.540 36.370 645.680 586.850 ;
        RECT 317.960 36.050 318.220 36.370 ;
        RECT 645.480 36.050 645.740 36.370 ;
        RECT 318.020 2.400 318.160 36.050 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 593.030 2625.680 593.310 2625.960 ;
        RECT 642.710 1939.560 642.990 1939.840 ;
        RECT 645.470 1939.560 645.750 1939.840 ;
        RECT 793.360 587.720 793.640 588.000 ;
        RECT 831.770 587.720 832.050 588.000 ;
      LAYER met3 ;
        RECT 574.800 2625.970 578.800 2626.480 ;
        RECT 593.005 2625.970 593.335 2625.985 ;
        RECT 574.800 2625.880 593.335 2625.970 ;
        RECT 578.070 2625.670 593.335 2625.880 ;
        RECT 593.005 2625.655 593.335 2625.670 ;
        RECT 627.030 1939.850 631.030 1940.000 ;
        RECT 642.685 1939.850 643.015 1939.865 ;
        RECT 645.445 1939.850 645.775 1939.865 ;
        RECT 627.030 1939.550 645.775 1939.850 ;
        RECT 627.030 1939.400 631.030 1939.550 ;
        RECT 642.685 1939.535 643.015 1939.550 ;
        RECT 645.445 1939.535 645.775 1939.550 ;
        RECT 793.335 588.010 793.665 588.025 ;
        RECT 831.745 588.010 832.075 588.025 ;
        RECT 793.335 587.710 832.075 588.010 ;
        RECT 793.335 587.695 793.665 587.710 ;
        RECT 831.745 587.695 832.075 587.710 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 2504.000 482.930 2504.060 ;
        RECT 1901.710 2504.000 1902.030 2504.060 ;
        RECT 482.610 2503.860 1902.030 2504.000 ;
        RECT 482.610 2503.800 482.930 2503.860 ;
        RECT 1901.710 2503.800 1902.030 2503.860 ;
        RECT 351.510 2501.280 351.830 2501.340 ;
        RECT 476.170 2501.280 476.490 2501.340 ;
        RECT 482.610 2501.280 482.930 2501.340 ;
        RECT 351.510 2501.140 482.930 2501.280 ;
        RECT 351.510 2501.080 351.830 2501.140 ;
        RECT 476.170 2501.080 476.490 2501.140 ;
        RECT 482.610 2501.080 482.930 2501.140 ;
        RECT 337.710 587.420 338.030 587.480 ;
        RECT 355.190 587.420 355.510 587.480 ;
        RECT 841.870 587.420 842.190 587.480 ;
        RECT 337.710 587.280 842.190 587.420 ;
        RECT 337.710 587.220 338.030 587.280 ;
        RECT 355.190 587.220 355.510 587.280 ;
        RECT 841.870 587.220 842.190 587.280 ;
      LAYER via ;
        RECT 482.640 2503.800 482.900 2504.060 ;
        RECT 1901.740 2503.800 1902.000 2504.060 ;
        RECT 351.540 2501.080 351.800 2501.340 ;
        RECT 476.200 2501.080 476.460 2501.340 ;
        RECT 482.640 2501.080 482.900 2501.340 ;
        RECT 337.740 587.220 338.000 587.480 ;
        RECT 355.220 587.220 355.480 587.480 ;
        RECT 841.900 587.220 842.160 587.480 ;
      LAYER met2 ;
        RECT 476.090 2600.660 476.370 2604.000 ;
        RECT 476.090 2600.000 476.400 2600.660 ;
        RECT 476.260 2501.370 476.400 2600.000 ;
        RECT 1901.730 2532.475 1902.010 2532.845 ;
        RECT 1901.800 2504.090 1901.940 2532.475 ;
        RECT 482.640 2503.770 482.900 2504.090 ;
        RECT 1901.740 2503.770 1902.000 2504.090 ;
        RECT 482.700 2501.370 482.840 2503.770 ;
        RECT 351.540 2501.050 351.800 2501.370 ;
        RECT 476.200 2501.050 476.460 2501.370 ;
        RECT 482.640 2501.050 482.900 2501.370 ;
        RECT 351.600 1889.565 351.740 2501.050 ;
        RECT 351.530 1889.195 351.810 1889.565 ;
        RECT 355.210 1889.195 355.490 1889.565 ;
        RECT 355.280 587.510 355.420 1889.195 ;
        RECT 842.130 600.000 842.410 604.000 ;
        RECT 842.190 598.810 842.330 600.000 ;
        RECT 841.960 598.670 842.330 598.810 ;
        RECT 841.960 587.510 842.100 598.670 ;
        RECT 337.740 587.190 338.000 587.510 ;
        RECT 355.220 587.190 355.480 587.510 ;
        RECT 841.900 587.190 842.160 587.510 ;
        RECT 337.800 17.410 337.940 587.190 ;
        RECT 335.960 17.270 337.940 17.410 ;
        RECT 335.960 2.400 336.100 17.270 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 1901.730 2532.520 1902.010 2532.800 ;
        RECT 351.530 1889.240 351.810 1889.520 ;
        RECT 355.210 1889.240 355.490 1889.520 ;
      LAYER met3 ;
        RECT 1885.335 2534.360 1889.335 2534.640 ;
        RECT 1885.335 2534.040 1889.370 2534.360 ;
        RECT 1889.070 2532.810 1889.370 2534.040 ;
        RECT 1901.705 2532.810 1902.035 2532.825 ;
        RECT 1889.070 2532.510 1902.035 2532.810 ;
        RECT 1901.705 2532.495 1902.035 2532.510 ;
        RECT 351.505 1889.530 351.835 1889.545 ;
        RECT 355.185 1889.530 355.515 1889.545 ;
        RECT 360.000 1889.530 364.000 1889.680 ;
        RECT 351.505 1889.230 364.000 1889.530 ;
        RECT 351.505 1889.215 351.835 1889.230 ;
        RECT 355.185 1889.215 355.515 1889.230 ;
        RECT 360.000 1889.080 364.000 1889.230 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 475.250 2768.860 475.570 2768.920 ;
        RECT 603.590 2768.860 603.910 2768.920 ;
        RECT 475.250 2768.720 603.910 2768.860 ;
        RECT 475.250 2768.660 475.570 2768.720 ;
        RECT 603.590 2768.660 603.910 2768.720 ;
        RECT 603.590 2490.060 603.910 2490.120 ;
        RECT 606.810 2490.060 607.130 2490.120 ;
        RECT 1694.250 2490.060 1694.570 2490.120 ;
        RECT 603.590 2489.920 1694.570 2490.060 ;
        RECT 603.590 2489.860 603.910 2489.920 ;
        RECT 606.810 2489.860 607.130 2489.920 ;
        RECT 1694.250 2489.860 1694.570 2489.920 ;
        RECT 604.510 1994.680 604.830 1994.740 ;
        RECT 606.810 1994.680 607.130 1994.740 ;
        RECT 628.430 1994.680 628.750 1994.740 ;
        RECT 604.510 1994.540 628.750 1994.680 ;
        RECT 604.510 1994.480 604.830 1994.540 ;
        RECT 606.810 1994.480 607.130 1994.540 ;
        RECT 628.430 1994.480 628.750 1994.540 ;
        RECT 628.430 592.180 628.750 592.240 ;
        RECT 850.150 592.180 850.470 592.240 ;
        RECT 628.430 592.040 850.470 592.180 ;
        RECT 628.430 591.980 628.750 592.040 ;
        RECT 850.150 591.980 850.470 592.040 ;
        RECT 603.590 587.080 603.910 587.140 ;
        RECT 628.430 587.080 628.750 587.140 ;
        RECT 603.590 586.940 628.750 587.080 ;
        RECT 603.590 586.880 603.910 586.940 ;
        RECT 628.430 586.880 628.750 586.940 ;
        RECT 353.350 22.000 353.670 22.060 ;
        RECT 603.590 22.000 603.910 22.060 ;
        RECT 353.350 21.860 603.910 22.000 ;
        RECT 353.350 21.800 353.670 21.860 ;
        RECT 603.590 21.800 603.910 21.860 ;
      LAYER via ;
        RECT 475.280 2768.660 475.540 2768.920 ;
        RECT 603.620 2768.660 603.880 2768.920 ;
        RECT 603.620 2489.860 603.880 2490.120 ;
        RECT 606.840 2489.860 607.100 2490.120 ;
        RECT 1694.280 2489.860 1694.540 2490.120 ;
        RECT 604.540 1994.480 604.800 1994.740 ;
        RECT 606.840 1994.480 607.100 1994.740 ;
        RECT 628.460 1994.480 628.720 1994.740 ;
        RECT 628.460 591.980 628.720 592.240 ;
        RECT 850.180 591.980 850.440 592.240 ;
        RECT 603.620 586.880 603.880 587.140 ;
        RECT 628.460 586.880 628.720 587.140 ;
        RECT 353.380 21.800 353.640 22.060 ;
        RECT 603.620 21.800 603.880 22.060 ;
      LAYER met2 ;
        RECT 475.280 2768.630 475.540 2768.950 ;
        RECT 603.620 2768.630 603.880 2768.950 ;
        RECT 475.340 2759.520 475.480 2768.630 ;
        RECT 475.170 2759.100 475.480 2759.520 ;
        RECT 475.170 2755.520 475.450 2759.100 ;
        RECT 603.680 2490.150 603.820 2768.630 ;
        RECT 1694.210 2500.000 1694.490 2504.000 ;
        RECT 1694.340 2490.150 1694.480 2500.000 ;
        RECT 603.620 2489.830 603.880 2490.150 ;
        RECT 606.840 2489.830 607.100 2490.150 ;
        RECT 1694.280 2489.830 1694.540 2490.150 ;
        RECT 606.900 1994.770 607.040 2489.830 ;
        RECT 604.540 1994.450 604.800 1994.770 ;
        RECT 606.840 1994.450 607.100 1994.770 ;
        RECT 628.460 1994.450 628.720 1994.770 ;
        RECT 602.970 1981.250 603.250 1981.750 ;
        RECT 604.600 1981.250 604.740 1994.450 ;
        RECT 602.970 1981.110 604.740 1981.250 ;
        RECT 602.970 1977.750 603.250 1981.110 ;
        RECT 628.520 592.270 628.660 1994.450 ;
        RECT 851.330 600.170 851.610 604.000 ;
        RECT 850.240 600.030 851.610 600.170 ;
        RECT 850.240 592.270 850.380 600.030 ;
        RECT 851.330 600.000 851.610 600.030 ;
        RECT 628.460 591.950 628.720 592.270 ;
        RECT 850.180 591.950 850.440 592.270 ;
        RECT 628.520 587.170 628.660 591.950 ;
        RECT 603.620 586.850 603.880 587.170 ;
        RECT 628.460 586.850 628.720 587.170 ;
        RECT 603.680 22.090 603.820 586.850 ;
        RECT 353.380 21.770 353.640 22.090 ;
        RECT 603.620 21.770 603.880 22.090 ;
        RECT 353.440 2.400 353.580 21.770 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 420.510 2916.080 420.830 2916.140 ;
        RECT 1588.450 2916.080 1588.770 2916.140 ;
        RECT 420.510 2915.940 1588.770 2916.080 ;
        RECT 420.510 2915.880 420.830 2915.940 ;
        RECT 1588.450 2915.880 1588.770 2915.940 ;
        RECT 420.970 1994.480 421.290 1994.740 ;
        RECT 358.410 1994.340 358.730 1994.400 ;
        RECT 421.060 1994.340 421.200 1994.480 ;
        RECT 427.410 1994.340 427.730 1994.400 ;
        RECT 358.410 1994.200 427.730 1994.340 ;
        RECT 358.410 1994.140 358.730 1994.200 ;
        RECT 427.410 1994.140 427.730 1994.200 ;
        RECT 427.410 1993.660 427.730 1993.720 ;
        RECT 451.330 1993.660 451.650 1993.720 ;
        RECT 427.410 1993.520 451.650 1993.660 ;
        RECT 427.410 1993.460 427.730 1993.520 ;
        RECT 451.330 1993.460 451.650 1993.520 ;
        RECT 665.690 589.800 666.010 589.860 ;
        RECT 713.990 589.800 714.310 589.860 ;
        RECT 665.690 589.660 714.310 589.800 ;
        RECT 665.690 589.600 666.010 589.660 ;
        RECT 713.990 589.600 714.310 589.660 ;
        RECT 793.110 589.460 793.430 589.520 ;
        RECT 793.110 589.320 817.260 589.460 ;
        RECT 793.110 589.260 793.430 589.320 ;
        RECT 482.610 589.120 482.930 589.180 ;
        RECT 496.410 589.120 496.730 589.180 ;
        RECT 482.610 588.980 496.730 589.120 ;
        RECT 482.610 588.920 482.930 588.980 ;
        RECT 496.410 588.920 496.730 588.980 ;
        RECT 496.870 589.120 497.190 589.180 ;
        RECT 496.870 588.980 503.080 589.120 ;
        RECT 496.870 588.920 497.190 588.980 ;
        RECT 358.410 588.780 358.730 588.840 ;
        RECT 368.990 588.780 369.310 588.840 ;
        RECT 399.810 588.780 400.130 588.840 ;
        RECT 358.410 588.640 400.130 588.780 ;
        RECT 502.940 588.780 503.080 588.980 ;
        RECT 592.550 588.780 592.870 588.840 ;
        RECT 502.940 588.640 544.940 588.780 ;
        RECT 358.410 588.580 358.730 588.640 ;
        RECT 368.990 588.580 369.310 588.640 ;
        RECT 399.810 588.580 400.130 588.640 ;
        RECT 400.730 588.440 401.050 588.500 ;
        RECT 434.770 588.440 435.090 588.500 ;
        RECT 400.730 588.300 435.090 588.440 ;
        RECT 544.800 588.440 544.940 588.640 ;
        RECT 545.260 588.640 592.870 588.780 ;
        RECT 817.120 588.780 817.260 589.320 ;
        RECT 858.890 588.780 859.210 588.840 ;
        RECT 817.120 588.640 859.210 588.780 ;
        RECT 545.260 588.440 545.400 588.640 ;
        RECT 592.550 588.580 592.870 588.640 ;
        RECT 858.890 588.580 859.210 588.640 ;
        RECT 544.800 588.300 545.400 588.440 ;
        RECT 400.730 588.240 401.050 588.300 ;
        RECT 434.770 588.240 435.090 588.300 ;
        RECT 665.690 588.100 666.010 588.160 ;
        RECT 594.020 587.960 666.010 588.100 ;
        RECT 434.770 587.760 435.090 587.820 ;
        RECT 482.610 587.760 482.930 587.820 ;
        RECT 434.770 587.620 482.930 587.760 ;
        RECT 434.770 587.560 435.090 587.620 ;
        RECT 482.610 587.560 482.930 587.620 ;
        RECT 592.550 587.760 592.870 587.820 ;
        RECT 594.020 587.760 594.160 587.960 ;
        RECT 665.690 587.900 666.010 587.960 ;
        RECT 592.550 587.620 594.160 587.760 ;
        RECT 713.990 587.760 714.310 587.820 ;
        RECT 791.730 587.760 792.050 587.820 ;
        RECT 713.990 587.620 792.050 587.760 ;
        RECT 592.550 587.560 592.870 587.620 ;
        RECT 713.990 587.560 714.310 587.620 ;
        RECT 791.730 587.560 792.050 587.620 ;
        RECT 368.990 20.640 369.310 20.700 ;
        RECT 371.290 20.640 371.610 20.700 ;
        RECT 368.990 20.500 371.610 20.640 ;
        RECT 368.990 20.440 369.310 20.500 ;
        RECT 371.290 20.440 371.610 20.500 ;
      LAYER via ;
        RECT 420.540 2915.880 420.800 2916.140 ;
        RECT 1588.480 2915.880 1588.740 2916.140 ;
        RECT 421.000 1994.480 421.260 1994.740 ;
        RECT 358.440 1994.140 358.700 1994.400 ;
        RECT 427.440 1994.140 427.700 1994.400 ;
        RECT 427.440 1993.460 427.700 1993.720 ;
        RECT 451.360 1993.460 451.620 1993.720 ;
        RECT 665.720 589.600 665.980 589.860 ;
        RECT 714.020 589.600 714.280 589.860 ;
        RECT 793.140 589.260 793.400 589.520 ;
        RECT 482.640 588.920 482.900 589.180 ;
        RECT 496.440 588.920 496.700 589.180 ;
        RECT 496.900 588.920 497.160 589.180 ;
        RECT 358.440 588.580 358.700 588.840 ;
        RECT 369.020 588.580 369.280 588.840 ;
        RECT 399.840 588.580 400.100 588.840 ;
        RECT 400.760 588.240 401.020 588.500 ;
        RECT 434.800 588.240 435.060 588.500 ;
        RECT 592.580 588.580 592.840 588.840 ;
        RECT 858.920 588.580 859.180 588.840 ;
        RECT 434.800 587.560 435.060 587.820 ;
        RECT 482.640 587.560 482.900 587.820 ;
        RECT 592.580 587.560 592.840 587.820 ;
        RECT 665.720 587.900 665.980 588.160 ;
        RECT 714.020 587.560 714.280 587.820 ;
        RECT 791.760 587.560 792.020 587.820 ;
        RECT 369.020 20.440 369.280 20.700 ;
        RECT 371.320 20.440 371.580 20.700 ;
      LAYER met2 ;
        RECT 420.540 2915.850 420.800 2916.170 ;
        RECT 1588.480 2915.850 1588.740 2916.170 ;
        RECT 420.600 2752.485 420.740 2915.850 ;
        RECT 1588.540 2900.055 1588.680 2915.850 ;
        RECT 1588.410 2896.055 1588.690 2900.055 ;
        RECT 420.530 2752.115 420.810 2752.485 ;
        RECT 420.600 2746.930 420.740 2752.115 ;
        RECT 420.600 2746.790 421.200 2746.930 ;
        RECT 421.060 1994.770 421.200 2746.790 ;
        RECT 421.000 1994.450 421.260 1994.770 ;
        RECT 358.440 1994.110 358.700 1994.430 ;
        RECT 427.440 1994.110 427.700 1994.430 ;
        RECT 358.500 588.870 358.640 1994.110 ;
        RECT 427.500 1993.750 427.640 1994.110 ;
        RECT 427.440 1993.430 427.700 1993.750 ;
        RECT 451.360 1993.430 451.620 1993.750 ;
        RECT 451.420 1981.250 451.560 1993.430 ;
        RECT 453.010 1981.250 453.290 1981.750 ;
        RECT 451.420 1981.110 453.290 1981.250 ;
        RECT 453.010 1977.750 453.290 1981.110 ;
        RECT 860.530 600.170 860.810 604.000 ;
        RECT 858.980 600.030 860.810 600.170 ;
        RECT 665.720 589.570 665.980 589.890 ;
        RECT 714.020 589.570 714.280 589.890 ;
        RECT 791.820 589.830 793.340 589.970 ;
        RECT 496.500 589.210 497.100 589.290 ;
        RECT 482.640 588.890 482.900 589.210 ;
        RECT 496.440 589.150 497.160 589.210 ;
        RECT 496.440 588.890 496.700 589.150 ;
        RECT 496.900 588.890 497.160 589.150 ;
        RECT 358.440 588.550 358.700 588.870 ;
        RECT 369.020 588.550 369.280 588.870 ;
        RECT 399.840 588.610 400.100 588.870 ;
        RECT 399.840 588.550 400.960 588.610 ;
        RECT 369.080 20.730 369.220 588.550 ;
        RECT 399.900 588.530 400.960 588.550 ;
        RECT 399.900 588.470 401.020 588.530 ;
        RECT 400.760 588.210 401.020 588.470 ;
        RECT 434.800 588.210 435.060 588.530 ;
        RECT 434.860 587.850 435.000 588.210 ;
        RECT 482.700 587.850 482.840 588.890 ;
        RECT 592.580 588.550 592.840 588.870 ;
        RECT 592.640 587.850 592.780 588.550 ;
        RECT 665.780 588.190 665.920 589.570 ;
        RECT 665.720 587.870 665.980 588.190 ;
        RECT 714.080 587.850 714.220 589.570 ;
        RECT 791.820 587.850 791.960 589.830 ;
        RECT 793.200 589.550 793.340 589.830 ;
        RECT 793.140 589.230 793.400 589.550 ;
        RECT 858.980 588.870 859.120 600.030 ;
        RECT 860.530 600.000 860.810 600.030 ;
        RECT 858.920 588.550 859.180 588.870 ;
        RECT 434.800 587.530 435.060 587.850 ;
        RECT 482.640 587.530 482.900 587.850 ;
        RECT 592.580 587.530 592.840 587.850 ;
        RECT 714.020 587.530 714.280 587.850 ;
        RECT 791.760 587.530 792.020 587.850 ;
        RECT 369.020 20.410 369.280 20.730 ;
        RECT 371.320 20.410 371.580 20.730 ;
        RECT 371.380 2.400 371.520 20.410 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 420.530 2752.160 420.810 2752.440 ;
      LAYER met3 ;
        RECT 430.000 2752.640 434.000 2752.960 ;
        RECT 420.505 2752.450 420.835 2752.465 ;
        RECT 429.950 2752.450 434.000 2752.640 ;
        RECT 420.505 2752.360 434.000 2752.450 ;
        RECT 420.505 2752.150 430.250 2752.360 ;
        RECT 420.505 2752.135 420.835 2752.150 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 503.770 2768.520 504.090 2768.580 ;
        RECT 645.910 2768.520 646.230 2768.580 ;
        RECT 503.770 2768.380 646.230 2768.520 ;
        RECT 503.770 2768.320 504.090 2768.380 ;
        RECT 645.910 2768.320 646.230 2768.380 ;
        RECT 645.910 2490.740 646.230 2490.800 ;
        RECT 1821.210 2490.740 1821.530 2490.800 ;
        RECT 645.910 2490.600 1821.530 2490.740 ;
        RECT 645.910 2490.540 646.230 2490.600 ;
        RECT 1821.210 2490.540 1821.530 2490.600 ;
        RECT 645.910 591.500 646.230 591.560 ;
        RECT 664.310 591.500 664.630 591.560 ;
        RECT 645.910 591.360 664.630 591.500 ;
        RECT 645.910 591.300 646.230 591.360 ;
        RECT 664.310 591.300 664.630 591.360 ;
        RECT 665.230 590.480 665.550 590.540 ;
        RECT 869.930 590.480 870.250 590.540 ;
        RECT 665.230 590.340 870.250 590.480 ;
        RECT 665.230 590.280 665.550 590.340 ;
        RECT 869.930 590.280 870.250 590.340 ;
        RECT 389.230 43.760 389.550 43.820 ;
        RECT 645.910 43.760 646.230 43.820 ;
        RECT 389.230 43.620 646.230 43.760 ;
        RECT 389.230 43.560 389.550 43.620 ;
        RECT 645.910 43.560 646.230 43.620 ;
      LAYER via ;
        RECT 503.800 2768.320 504.060 2768.580 ;
        RECT 645.940 2768.320 646.200 2768.580 ;
        RECT 645.940 2490.540 646.200 2490.800 ;
        RECT 1821.240 2490.540 1821.500 2490.800 ;
        RECT 645.940 591.300 646.200 591.560 ;
        RECT 664.340 591.300 664.600 591.560 ;
        RECT 665.260 590.280 665.520 590.540 ;
        RECT 869.960 590.280 870.220 590.540 ;
        RECT 389.260 43.560 389.520 43.820 ;
        RECT 645.940 43.560 646.200 43.820 ;
      LAYER met2 ;
        RECT 503.800 2768.290 504.060 2768.610 ;
        RECT 645.940 2768.290 646.200 2768.610 ;
        RECT 503.860 2759.520 504.000 2768.290 ;
        RECT 503.690 2759.100 504.000 2759.520 ;
        RECT 503.690 2755.520 503.970 2759.100 ;
        RECT 646.000 2490.830 646.140 2768.290 ;
        RECT 1821.170 2500.000 1821.450 2504.000 ;
        RECT 1821.300 2490.830 1821.440 2500.000 ;
        RECT 645.940 2490.510 646.200 2490.830 ;
        RECT 1821.240 2490.510 1821.500 2490.830 ;
        RECT 646.000 1903.165 646.140 2490.510 ;
        RECT 645.930 1902.795 646.210 1903.165 ;
        RECT 646.000 591.590 646.140 1902.795 ;
        RECT 869.730 600.000 870.010 604.000 ;
        RECT 869.790 598.810 869.930 600.000 ;
        RECT 869.790 598.670 870.160 598.810 ;
        RECT 645.940 591.270 646.200 591.590 ;
        RECT 664.340 591.330 664.600 591.590 ;
        RECT 664.340 591.270 665.460 591.330 ;
        RECT 646.000 43.850 646.140 591.270 ;
        RECT 664.400 591.190 665.460 591.270 ;
        RECT 665.320 590.570 665.460 591.190 ;
        RECT 870.020 590.570 870.160 598.670 ;
        RECT 665.260 590.250 665.520 590.570 ;
        RECT 869.960 590.250 870.220 590.570 ;
        RECT 389.260 43.530 389.520 43.850 ;
        RECT 645.940 43.530 646.200 43.850 ;
        RECT 389.320 2.400 389.460 43.530 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 645.930 1902.840 646.210 1903.120 ;
      LAYER met3 ;
        RECT 627.030 1903.130 631.030 1903.280 ;
        RECT 645.905 1903.130 646.235 1903.145 ;
        RECT 627.030 1902.830 646.235 1903.130 ;
        RECT 627.030 1902.680 631.030 1902.830 ;
        RECT 645.905 1902.815 646.235 1902.830 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 2487.680 419.450 2487.740 ;
        RECT 635.790 2487.680 636.110 2487.740 ;
        RECT 1800.050 2487.680 1800.370 2487.740 ;
        RECT 419.130 2487.540 1800.370 2487.680 ;
        RECT 419.130 2487.480 419.450 2487.540 ;
        RECT 635.790 2487.480 636.110 2487.540 ;
        RECT 1800.050 2487.480 1800.370 2487.540 ;
        RECT 564.030 1689.700 564.350 1689.760 ;
        RECT 565.410 1689.700 565.730 1689.760 ;
        RECT 635.790 1689.700 636.110 1689.760 ;
        RECT 564.030 1689.560 636.110 1689.700 ;
        RECT 564.030 1689.500 564.350 1689.560 ;
        RECT 565.410 1689.500 565.730 1689.560 ;
        RECT 635.790 1689.500 636.110 1689.560 ;
        RECT 565.410 591.160 565.730 591.220 ;
        RECT 877.290 591.160 877.610 591.220 ;
        RECT 565.410 591.020 877.610 591.160 ;
        RECT 565.410 590.960 565.730 591.020 ;
        RECT 877.290 590.960 877.610 591.020 ;
        RECT 548.390 586.740 548.710 586.800 ;
        RECT 565.410 586.740 565.730 586.800 ;
        RECT 548.390 586.600 565.730 586.740 ;
        RECT 548.390 586.540 548.710 586.600 ;
        RECT 565.410 586.540 565.730 586.600 ;
        RECT 407.170 29.140 407.490 29.200 ;
        RECT 548.390 29.140 548.710 29.200 ;
        RECT 407.170 29.000 548.710 29.140 ;
        RECT 407.170 28.940 407.490 29.000 ;
        RECT 548.390 28.940 548.710 29.000 ;
      LAYER via ;
        RECT 419.160 2487.480 419.420 2487.740 ;
        RECT 635.820 2487.480 636.080 2487.740 ;
        RECT 1800.080 2487.480 1800.340 2487.740 ;
        RECT 564.060 1689.500 564.320 1689.760 ;
        RECT 565.440 1689.500 565.700 1689.760 ;
        RECT 635.820 1689.500 636.080 1689.760 ;
        RECT 565.440 590.960 565.700 591.220 ;
        RECT 877.320 590.960 877.580 591.220 ;
        RECT 548.420 586.540 548.680 586.800 ;
        RECT 565.440 586.540 565.700 586.800 ;
        RECT 407.200 28.940 407.460 29.200 ;
        RECT 548.420 28.940 548.680 29.200 ;
      LAYER met2 ;
        RECT 419.150 2643.315 419.430 2643.685 ;
        RECT 419.220 2487.770 419.360 2643.315 ;
        RECT 1800.010 2500.000 1800.290 2504.000 ;
        RECT 1800.140 2487.770 1800.280 2500.000 ;
        RECT 419.160 2487.450 419.420 2487.770 ;
        RECT 635.820 2487.450 636.080 2487.770 ;
        RECT 1800.080 2487.450 1800.340 2487.770 ;
        RECT 562.490 1700.410 562.770 1704.000 ;
        RECT 562.490 1700.270 564.260 1700.410 ;
        RECT 562.490 1700.000 562.770 1700.270 ;
        RECT 564.120 1689.790 564.260 1700.270 ;
        RECT 635.880 1689.790 636.020 2487.450 ;
        RECT 564.060 1689.470 564.320 1689.790 ;
        RECT 565.440 1689.470 565.700 1689.790 ;
        RECT 635.820 1689.470 636.080 1689.790 ;
        RECT 565.500 591.250 565.640 1689.470 ;
        RECT 878.930 600.170 879.210 604.000 ;
        RECT 877.380 600.030 879.210 600.170 ;
        RECT 877.380 591.250 877.520 600.030 ;
        RECT 878.930 600.000 879.210 600.030 ;
        RECT 565.440 590.930 565.700 591.250 ;
        RECT 877.320 590.930 877.580 591.250 ;
        RECT 565.500 586.830 565.640 590.930 ;
        RECT 548.420 586.510 548.680 586.830 ;
        RECT 565.440 586.510 565.700 586.830 ;
        RECT 548.480 29.230 548.620 586.510 ;
        RECT 407.200 28.910 407.460 29.230 ;
        RECT 548.420 28.910 548.680 29.230 ;
        RECT 407.260 2.400 407.400 28.910 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 419.150 2643.360 419.430 2643.640 ;
      LAYER met3 ;
        RECT 430.000 2646.560 434.000 2646.880 ;
        RECT 429.950 2646.280 434.000 2646.560 ;
        RECT 419.125 2643.650 419.455 2643.665 ;
        RECT 429.950 2643.650 430.250 2646.280 ;
        RECT 419.125 2643.350 430.250 2643.650 ;
        RECT 419.125 2643.335 419.455 2643.350 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 596.690 2899.760 597.010 2899.820 ;
        RECT 1683.210 2899.760 1683.530 2899.820 ;
        RECT 596.690 2899.620 1683.530 2899.760 ;
        RECT 596.690 2899.560 597.010 2899.620 ;
        RECT 1683.210 2899.560 1683.530 2899.620 ;
        RECT 589.790 2649.520 590.110 2649.580 ;
        RECT 596.690 2649.520 597.010 2649.580 ;
        RECT 589.790 2649.380 597.010 2649.520 ;
        RECT 589.790 2649.320 590.110 2649.380 ;
        RECT 596.690 2649.320 597.010 2649.380 ;
        RECT 357.490 1983.800 357.810 1983.860 ;
        RECT 589.790 1983.800 590.110 1983.860 ;
        RECT 631.650 1983.800 631.970 1983.860 ;
        RECT 357.490 1983.660 631.970 1983.800 ;
        RECT 357.490 1983.600 357.810 1983.660 ;
        RECT 589.790 1983.600 590.110 1983.660 ;
        RECT 631.650 1983.600 631.970 1983.660 ;
        RECT 631.650 1883.840 631.970 1883.900 ;
        RECT 664.310 1883.840 664.630 1883.900 ;
        RECT 631.650 1883.700 664.630 1883.840 ;
        RECT 631.650 1883.640 631.970 1883.700 ;
        RECT 664.310 1883.640 664.630 1883.700 ;
        RECT 664.310 1849.500 664.630 1849.560 ;
        RECT 663.940 1849.360 664.630 1849.500 ;
        RECT 663.940 1849.220 664.080 1849.360 ;
        RECT 664.310 1849.300 664.630 1849.360 ;
        RECT 663.850 1848.960 664.170 1849.220 ;
        RECT 663.850 1800.880 664.170 1800.940 ;
        RECT 664.770 1800.880 665.090 1800.940 ;
        RECT 663.850 1800.740 665.090 1800.880 ;
        RECT 663.850 1800.680 664.170 1800.740 ;
        RECT 664.770 1800.680 665.090 1800.740 ;
        RECT 664.770 1752.940 665.090 1753.000 ;
        RECT 664.400 1752.800 665.090 1752.940 ;
        RECT 664.400 1752.660 664.540 1752.800 ;
        RECT 664.770 1752.740 665.090 1752.800 ;
        RECT 664.310 1752.400 664.630 1752.660 ;
        RECT 662.470 1738.660 662.790 1738.720 ;
        RECT 664.310 1738.660 664.630 1738.720 ;
        RECT 662.470 1738.520 664.630 1738.660 ;
        RECT 662.470 1738.460 662.790 1738.520 ;
        RECT 664.310 1738.460 664.630 1738.520 ;
        RECT 662.470 1702.960 662.790 1703.020 ;
        RECT 1400.770 1702.960 1401.090 1703.020 ;
        RECT 662.470 1702.820 1401.090 1702.960 ;
        RECT 662.470 1702.760 662.790 1702.820 ;
        RECT 1400.770 1702.760 1401.090 1702.820 ;
        RECT 1402.610 1702.960 1402.930 1703.020 ;
        RECT 1642.270 1702.960 1642.590 1703.020 ;
        RECT 1402.610 1702.820 1642.590 1702.960 ;
        RECT 1402.610 1702.760 1402.930 1702.820 ;
        RECT 1642.270 1702.760 1642.590 1702.820 ;
        RECT 1644.110 1702.960 1644.430 1703.020 ;
        RECT 1918.270 1702.960 1918.590 1703.020 ;
        RECT 1644.110 1702.820 1918.590 1702.960 ;
        RECT 1644.110 1702.760 1644.430 1702.820 ;
        RECT 1918.270 1702.760 1918.590 1702.820 ;
        RECT 662.470 1690.720 662.790 1690.780 ;
        RECT 663.850 1690.720 664.170 1690.780 ;
        RECT 662.470 1690.580 664.170 1690.720 ;
        RECT 662.470 1690.520 662.790 1690.580 ;
        RECT 663.850 1690.520 664.170 1690.580 ;
        RECT 663.390 1642.440 663.710 1642.500 ;
        RECT 664.770 1642.440 665.090 1642.500 ;
        RECT 663.390 1642.300 665.090 1642.440 ;
        RECT 663.390 1642.240 663.710 1642.300 ;
        RECT 664.770 1642.240 665.090 1642.300 ;
        RECT 662.470 1641.760 662.790 1641.820 ;
        RECT 663.390 1641.760 663.710 1641.820 ;
        RECT 662.470 1641.620 663.710 1641.760 ;
        RECT 662.470 1641.560 662.790 1641.620 ;
        RECT 663.390 1641.560 663.710 1641.620 ;
        RECT 662.470 1594.160 662.790 1594.220 ;
        RECT 663.850 1594.160 664.170 1594.220 ;
        RECT 662.470 1594.020 664.170 1594.160 ;
        RECT 662.470 1593.960 662.790 1594.020 ;
        RECT 663.850 1593.960 664.170 1594.020 ;
        RECT 662.470 1497.260 662.790 1497.320 ;
        RECT 663.850 1497.260 664.170 1497.320 ;
        RECT 662.470 1497.120 664.170 1497.260 ;
        RECT 662.470 1497.060 662.790 1497.120 ;
        RECT 663.850 1497.060 664.170 1497.120 ;
        RECT 662.470 1449.320 662.790 1449.380 ;
        RECT 663.390 1449.320 663.710 1449.380 ;
        RECT 662.470 1449.180 663.710 1449.320 ;
        RECT 662.470 1449.120 662.790 1449.180 ;
        RECT 663.390 1449.120 663.710 1449.180 ;
        RECT 662.470 1400.700 662.790 1400.760 ;
        RECT 663.850 1400.700 664.170 1400.760 ;
        RECT 662.470 1400.560 664.170 1400.700 ;
        RECT 662.470 1400.500 662.790 1400.560 ;
        RECT 663.850 1400.500 664.170 1400.560 ;
        RECT 662.470 1352.760 662.790 1352.820 ;
        RECT 663.390 1352.760 663.710 1352.820 ;
        RECT 662.470 1352.620 663.710 1352.760 ;
        RECT 662.470 1352.560 662.790 1352.620 ;
        RECT 663.390 1352.560 663.710 1352.620 ;
        RECT 663.850 1304.140 664.170 1304.200 ;
        RECT 664.770 1304.140 665.090 1304.200 ;
        RECT 663.850 1304.000 665.090 1304.140 ;
        RECT 663.850 1303.940 664.170 1304.000 ;
        RECT 664.770 1303.940 665.090 1304.000 ;
        RECT 664.770 1269.940 665.090 1270.200 ;
        RECT 664.860 1269.180 665.000 1269.940 ;
        RECT 664.770 1268.920 665.090 1269.180 ;
        RECT 663.390 1256.540 663.710 1256.600 ;
        RECT 664.770 1256.540 665.090 1256.600 ;
        RECT 663.390 1256.400 665.090 1256.540 ;
        RECT 663.390 1256.340 663.710 1256.400 ;
        RECT 664.770 1256.340 665.090 1256.400 ;
        RECT 662.470 1160.320 662.790 1160.380 ;
        RECT 663.850 1160.320 664.170 1160.380 ;
        RECT 662.470 1160.180 664.170 1160.320 ;
        RECT 662.470 1160.120 662.790 1160.180 ;
        RECT 663.850 1160.120 664.170 1160.180 ;
        RECT 662.470 1124.960 662.790 1125.020 ;
        RECT 663.850 1124.960 664.170 1125.020 ;
        RECT 662.470 1124.820 664.170 1124.960 ;
        RECT 662.470 1124.760 662.790 1124.820 ;
        RECT 663.850 1124.760 664.170 1124.820 ;
        RECT 663.850 1097.420 664.170 1097.480 ;
        RECT 664.770 1097.420 665.090 1097.480 ;
        RECT 663.850 1097.280 665.090 1097.420 ;
        RECT 663.850 1097.220 664.170 1097.280 ;
        RECT 664.770 1097.220 665.090 1097.280 ;
        RECT 664.770 1052.200 665.090 1052.260 ;
        RECT 668.450 1052.200 668.770 1052.260 ;
        RECT 664.770 1052.060 668.770 1052.200 ;
        RECT 664.770 1052.000 665.090 1052.060 ;
        RECT 668.450 1052.000 668.770 1052.060 ;
        RECT 664.770 1000.860 665.090 1000.920 ;
        RECT 668.450 1000.860 668.770 1000.920 ;
        RECT 664.770 1000.720 668.770 1000.860 ;
        RECT 664.770 1000.660 665.090 1000.720 ;
        RECT 668.450 1000.660 668.770 1000.720 ;
        RECT 665.230 820.660 665.550 820.720 ;
        RECT 665.690 820.660 666.010 820.720 ;
        RECT 665.230 820.520 666.010 820.660 ;
        RECT 665.230 820.460 665.550 820.520 ;
        RECT 665.690 820.460 666.010 820.520 ;
        RECT 664.770 773.060 665.090 773.120 ;
        RECT 665.230 773.060 665.550 773.120 ;
        RECT 664.770 772.920 665.550 773.060 ;
        RECT 664.770 772.860 665.090 772.920 ;
        RECT 665.230 772.860 665.550 772.920 ;
        RECT 664.310 772.720 664.630 772.780 ;
        RECT 664.310 772.580 665.460 772.720 ;
        RECT 664.310 772.520 664.630 772.580 ;
        RECT 665.320 772.440 665.460 772.580 ;
        RECT 665.230 772.180 665.550 772.440 ;
        RECT 663.390 724.440 663.710 724.500 ;
        RECT 664.310 724.440 664.630 724.500 ;
        RECT 663.390 724.300 664.630 724.440 ;
        RECT 663.390 724.240 663.710 724.300 ;
        RECT 664.310 724.240 664.630 724.300 ;
        RECT 663.390 689.080 663.710 689.140 ;
        RECT 665.690 689.080 666.010 689.140 ;
        RECT 663.390 688.940 666.010 689.080 ;
        RECT 663.390 688.880 663.710 688.940 ;
        RECT 665.690 688.880 666.010 688.940 ;
        RECT 666.150 496.780 666.470 497.040 ;
        RECT 666.240 496.360 666.380 496.780 ;
        RECT 666.150 496.100 666.470 496.360 ;
        RECT 665.230 448.700 665.550 448.760 ;
        RECT 666.150 448.700 666.470 448.760 ;
        RECT 665.230 448.560 666.470 448.700 ;
        RECT 665.230 448.500 665.550 448.560 ;
        RECT 666.150 448.500 666.470 448.560 ;
        RECT 664.770 289.580 665.090 289.640 ;
        RECT 666.150 289.580 666.470 289.640 ;
        RECT 664.770 289.440 666.470 289.580 ;
        RECT 664.770 289.380 665.090 289.440 ;
        RECT 666.150 289.380 666.470 289.440 ;
        RECT 68.150 45.460 68.470 45.520 ;
        RECT 665.230 45.460 665.550 45.520 ;
        RECT 68.150 45.320 665.550 45.460 ;
        RECT 68.150 45.260 68.470 45.320 ;
        RECT 665.230 45.260 665.550 45.320 ;
      LAYER via ;
        RECT 596.720 2899.560 596.980 2899.820 ;
        RECT 1683.240 2899.560 1683.500 2899.820 ;
        RECT 589.820 2649.320 590.080 2649.580 ;
        RECT 596.720 2649.320 596.980 2649.580 ;
        RECT 357.520 1983.600 357.780 1983.860 ;
        RECT 589.820 1983.600 590.080 1983.860 ;
        RECT 631.680 1983.600 631.940 1983.860 ;
        RECT 631.680 1883.640 631.940 1883.900 ;
        RECT 664.340 1883.640 664.600 1883.900 ;
        RECT 664.340 1849.300 664.600 1849.560 ;
        RECT 663.880 1848.960 664.140 1849.220 ;
        RECT 663.880 1800.680 664.140 1800.940 ;
        RECT 664.800 1800.680 665.060 1800.940 ;
        RECT 664.800 1752.740 665.060 1753.000 ;
        RECT 664.340 1752.400 664.600 1752.660 ;
        RECT 662.500 1738.460 662.760 1738.720 ;
        RECT 664.340 1738.460 664.600 1738.720 ;
        RECT 662.500 1702.760 662.760 1703.020 ;
        RECT 1400.800 1702.760 1401.060 1703.020 ;
        RECT 1402.640 1702.760 1402.900 1703.020 ;
        RECT 1642.300 1702.760 1642.560 1703.020 ;
        RECT 1644.140 1702.760 1644.400 1703.020 ;
        RECT 1918.300 1702.760 1918.560 1703.020 ;
        RECT 662.500 1690.520 662.760 1690.780 ;
        RECT 663.880 1690.520 664.140 1690.780 ;
        RECT 663.420 1642.240 663.680 1642.500 ;
        RECT 664.800 1642.240 665.060 1642.500 ;
        RECT 662.500 1641.560 662.760 1641.820 ;
        RECT 663.420 1641.560 663.680 1641.820 ;
        RECT 662.500 1593.960 662.760 1594.220 ;
        RECT 663.880 1593.960 664.140 1594.220 ;
        RECT 662.500 1497.060 662.760 1497.320 ;
        RECT 663.880 1497.060 664.140 1497.320 ;
        RECT 662.500 1449.120 662.760 1449.380 ;
        RECT 663.420 1449.120 663.680 1449.380 ;
        RECT 662.500 1400.500 662.760 1400.760 ;
        RECT 663.880 1400.500 664.140 1400.760 ;
        RECT 662.500 1352.560 662.760 1352.820 ;
        RECT 663.420 1352.560 663.680 1352.820 ;
        RECT 663.880 1303.940 664.140 1304.200 ;
        RECT 664.800 1303.940 665.060 1304.200 ;
        RECT 664.800 1269.940 665.060 1270.200 ;
        RECT 664.800 1268.920 665.060 1269.180 ;
        RECT 663.420 1256.340 663.680 1256.600 ;
        RECT 664.800 1256.340 665.060 1256.600 ;
        RECT 662.500 1160.120 662.760 1160.380 ;
        RECT 663.880 1160.120 664.140 1160.380 ;
        RECT 662.500 1124.760 662.760 1125.020 ;
        RECT 663.880 1124.760 664.140 1125.020 ;
        RECT 663.880 1097.220 664.140 1097.480 ;
        RECT 664.800 1097.220 665.060 1097.480 ;
        RECT 664.800 1052.000 665.060 1052.260 ;
        RECT 668.480 1052.000 668.740 1052.260 ;
        RECT 664.800 1000.660 665.060 1000.920 ;
        RECT 668.480 1000.660 668.740 1000.920 ;
        RECT 665.260 820.460 665.520 820.720 ;
        RECT 665.720 820.460 665.980 820.720 ;
        RECT 664.800 772.860 665.060 773.120 ;
        RECT 665.260 772.860 665.520 773.120 ;
        RECT 664.340 772.520 664.600 772.780 ;
        RECT 665.260 772.180 665.520 772.440 ;
        RECT 663.420 724.240 663.680 724.500 ;
        RECT 664.340 724.240 664.600 724.500 ;
        RECT 663.420 688.880 663.680 689.140 ;
        RECT 665.720 688.880 665.980 689.140 ;
        RECT 666.180 496.780 666.440 497.040 ;
        RECT 666.180 496.100 666.440 496.360 ;
        RECT 665.260 448.500 665.520 448.760 ;
        RECT 666.180 448.500 666.440 448.760 ;
        RECT 664.800 289.380 665.060 289.640 ;
        RECT 666.180 289.380 666.440 289.640 ;
        RECT 68.180 45.260 68.440 45.520 ;
        RECT 665.260 45.260 665.520 45.520 ;
      LAYER met2 ;
        RECT 1684.090 2899.930 1684.370 2900.055 ;
        RECT 1683.300 2899.850 1684.370 2899.930 ;
        RECT 596.720 2899.530 596.980 2899.850 ;
        RECT 1683.240 2899.790 1684.370 2899.850 ;
        RECT 1683.240 2899.530 1683.500 2899.790 ;
        RECT 596.780 2649.610 596.920 2899.530 ;
        RECT 1684.090 2896.055 1684.370 2899.790 ;
        RECT 589.820 2649.290 590.080 2649.610 ;
        RECT 596.720 2649.290 596.980 2649.610 ;
        RECT 589.880 2648.445 590.020 2649.290 ;
        RECT 589.810 2648.075 590.090 2648.445 ;
        RECT 589.880 1983.890 590.020 2648.075 ;
        RECT 357.520 1983.570 357.780 1983.890 ;
        RECT 589.820 1983.570 590.080 1983.890 ;
        RECT 631.680 1983.570 631.940 1983.890 ;
        RECT 357.580 1926.285 357.720 1983.570 ;
        RECT 357.510 1925.915 357.790 1926.285 ;
        RECT 631.740 1883.930 631.880 1983.570 ;
        RECT 631.680 1883.610 631.940 1883.930 ;
        RECT 664.340 1883.610 664.600 1883.930 ;
        RECT 664.400 1849.590 664.540 1883.610 ;
        RECT 664.340 1849.270 664.600 1849.590 ;
        RECT 663.880 1848.930 664.140 1849.250 ;
        RECT 663.940 1800.970 664.080 1848.930 ;
        RECT 663.880 1800.650 664.140 1800.970 ;
        RECT 664.800 1800.650 665.060 1800.970 ;
        RECT 664.860 1753.030 665.000 1800.650 ;
        RECT 664.800 1752.710 665.060 1753.030 ;
        RECT 664.340 1752.370 664.600 1752.690 ;
        RECT 664.400 1738.750 664.540 1752.370 ;
        RECT 1922.850 1750.730 1923.130 1754.000 ;
        RECT 1918.360 1750.590 1923.130 1750.730 ;
        RECT 662.500 1738.430 662.760 1738.750 ;
        RECT 664.340 1738.430 664.600 1738.750 ;
        RECT 662.560 1703.050 662.700 1738.430 ;
        RECT 1918.360 1703.050 1918.500 1750.590 ;
        RECT 1922.850 1750.000 1923.130 1750.590 ;
        RECT 662.500 1702.730 662.760 1703.050 ;
        RECT 1400.800 1702.730 1401.060 1703.050 ;
        RECT 1402.640 1702.730 1402.900 1703.050 ;
        RECT 1642.300 1702.730 1642.560 1703.050 ;
        RECT 1644.140 1702.730 1644.400 1703.050 ;
        RECT 1918.300 1702.730 1918.560 1703.050 ;
        RECT 662.560 1690.810 662.700 1702.730 ;
        RECT 1400.860 1702.565 1401.000 1702.730 ;
        RECT 1402.700 1702.565 1402.840 1702.730 ;
        RECT 1642.360 1702.565 1642.500 1702.730 ;
        RECT 1644.200 1702.565 1644.340 1702.730 ;
        RECT 1400.790 1702.195 1401.070 1702.565 ;
        RECT 1402.630 1702.195 1402.910 1702.565 ;
        RECT 1642.290 1702.195 1642.570 1702.565 ;
        RECT 1644.130 1702.195 1644.410 1702.565 ;
        RECT 662.500 1690.490 662.760 1690.810 ;
        RECT 663.880 1690.490 664.140 1690.810 ;
        RECT 663.940 1690.040 664.080 1690.490 ;
        RECT 663.940 1689.900 665.000 1690.040 ;
        RECT 664.860 1642.530 665.000 1689.900 ;
        RECT 663.420 1642.210 663.680 1642.530 ;
        RECT 664.800 1642.210 665.060 1642.530 ;
        RECT 663.480 1641.850 663.620 1642.210 ;
        RECT 662.500 1641.530 662.760 1641.850 ;
        RECT 663.420 1641.530 663.680 1641.850 ;
        RECT 662.560 1594.250 662.700 1641.530 ;
        RECT 662.500 1593.930 662.760 1594.250 ;
        RECT 663.880 1593.930 664.140 1594.250 ;
        RECT 663.940 1593.650 664.080 1593.930 ;
        RECT 663.480 1593.510 664.080 1593.650 ;
        RECT 663.480 1510.690 663.620 1593.510 ;
        RECT 663.480 1510.550 664.080 1510.690 ;
        RECT 663.940 1497.350 664.080 1510.550 ;
        RECT 662.500 1497.030 662.760 1497.350 ;
        RECT 663.880 1497.030 664.140 1497.350 ;
        RECT 662.560 1449.410 662.700 1497.030 ;
        RECT 662.500 1449.090 662.760 1449.410 ;
        RECT 663.420 1449.090 663.680 1449.410 ;
        RECT 663.480 1414.130 663.620 1449.090 ;
        RECT 663.480 1413.990 664.080 1414.130 ;
        RECT 663.940 1400.790 664.080 1413.990 ;
        RECT 662.500 1400.470 662.760 1400.790 ;
        RECT 663.880 1400.470 664.140 1400.790 ;
        RECT 662.560 1352.850 662.700 1400.470 ;
        RECT 662.500 1352.530 662.760 1352.850 ;
        RECT 663.420 1352.530 663.680 1352.850 ;
        RECT 663.480 1317.570 663.620 1352.530 ;
        RECT 663.480 1317.430 664.080 1317.570 ;
        RECT 663.940 1304.230 664.080 1317.430 ;
        RECT 663.880 1303.910 664.140 1304.230 ;
        RECT 664.800 1303.910 665.060 1304.230 ;
        RECT 664.860 1270.230 665.000 1303.910 ;
        RECT 664.800 1269.910 665.060 1270.230 ;
        RECT 664.800 1268.890 665.060 1269.210 ;
        RECT 664.860 1256.630 665.000 1268.890 ;
        RECT 663.420 1256.310 663.680 1256.630 ;
        RECT 664.800 1256.310 665.060 1256.630 ;
        RECT 663.480 1221.010 663.620 1256.310 ;
        RECT 663.480 1220.870 664.080 1221.010 ;
        RECT 663.940 1160.410 664.080 1220.870 ;
        RECT 662.500 1160.090 662.760 1160.410 ;
        RECT 663.880 1160.090 664.140 1160.410 ;
        RECT 662.560 1125.050 662.700 1160.090 ;
        RECT 662.500 1124.730 662.760 1125.050 ;
        RECT 663.880 1124.730 664.140 1125.050 ;
        RECT 663.940 1097.510 664.080 1124.730 ;
        RECT 663.880 1097.190 664.140 1097.510 ;
        RECT 664.800 1097.190 665.060 1097.510 ;
        RECT 664.860 1052.290 665.000 1097.190 ;
        RECT 664.800 1051.970 665.060 1052.290 ;
        RECT 668.480 1051.970 668.740 1052.290 ;
        RECT 668.540 1000.950 668.680 1051.970 ;
        RECT 664.800 1000.630 665.060 1000.950 ;
        RECT 668.480 1000.630 668.740 1000.950 ;
        RECT 664.860 932.125 665.000 1000.630 ;
        RECT 664.790 931.755 665.070 932.125 ;
        RECT 664.790 903.875 665.070 904.245 ;
        RECT 664.860 869.565 665.000 903.875 ;
        RECT 664.790 869.195 665.070 869.565 ;
        RECT 665.710 820.915 665.990 821.285 ;
        RECT 665.780 820.750 665.920 820.915 ;
        RECT 665.260 820.430 665.520 820.750 ;
        RECT 665.720 820.430 665.980 820.750 ;
        RECT 665.320 773.150 665.460 820.430 ;
        RECT 664.800 772.890 665.060 773.150 ;
        RECT 664.400 772.830 665.060 772.890 ;
        RECT 665.260 772.830 665.520 773.150 ;
        RECT 664.400 772.810 665.000 772.830 ;
        RECT 664.340 772.750 665.000 772.810 ;
        RECT 664.340 772.490 664.600 772.750 ;
        RECT 664.400 772.335 664.540 772.490 ;
        RECT 665.260 772.150 665.520 772.470 ;
        RECT 665.320 724.725 665.460 772.150 ;
        RECT 663.420 724.210 663.680 724.530 ;
        RECT 664.330 724.355 664.610 724.725 ;
        RECT 665.250 724.355 665.530 724.725 ;
        RECT 664.340 724.210 664.600 724.355 ;
        RECT 663.480 689.170 663.620 724.210 ;
        RECT 663.420 688.850 663.680 689.170 ;
        RECT 665.720 688.850 665.980 689.170 ;
        RECT 665.780 593.485 665.920 688.850 ;
        RECT 705.050 600.170 705.330 604.000 ;
        RECT 703.960 600.030 705.330 600.170 ;
        RECT 703.960 593.485 704.100 600.030 ;
        RECT 705.050 600.000 705.330 600.030 ;
        RECT 665.710 593.115 665.990 593.485 ;
        RECT 666.630 593.115 666.910 593.485 ;
        RECT 703.890 593.115 704.170 593.485 ;
        RECT 666.700 591.500 666.840 593.115 ;
        RECT 666.240 591.360 666.840 591.500 ;
        RECT 666.240 497.070 666.380 591.360 ;
        RECT 666.180 496.750 666.440 497.070 ;
        RECT 666.180 496.070 666.440 496.390 ;
        RECT 666.240 448.790 666.380 496.070 ;
        RECT 665.260 448.530 665.520 448.790 ;
        RECT 665.260 448.470 665.920 448.530 ;
        RECT 666.180 448.470 666.440 448.790 ;
        RECT 665.320 448.390 665.920 448.470 ;
        RECT 665.780 447.850 665.920 448.390 ;
        RECT 665.780 447.710 666.380 447.850 ;
        RECT 666.240 289.670 666.380 447.710 ;
        RECT 664.800 289.350 665.060 289.670 ;
        RECT 666.180 289.350 666.440 289.670 ;
        RECT 664.860 254.730 665.000 289.350 ;
        RECT 664.860 254.590 665.920 254.730 ;
        RECT 665.780 207.130 665.920 254.590 ;
        RECT 665.780 206.990 666.380 207.130 ;
        RECT 666.240 62.290 666.380 206.990 ;
        RECT 665.320 62.150 666.380 62.290 ;
        RECT 665.320 45.550 665.460 62.150 ;
        RECT 68.180 45.230 68.440 45.550 ;
        RECT 665.260 45.230 665.520 45.550 ;
        RECT 68.240 2.400 68.380 45.230 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 589.810 2648.120 590.090 2648.400 ;
        RECT 357.510 1925.960 357.790 1926.240 ;
        RECT 1400.790 1702.240 1401.070 1702.520 ;
        RECT 1402.630 1702.240 1402.910 1702.520 ;
        RECT 1642.290 1702.240 1642.570 1702.520 ;
        RECT 1644.130 1702.240 1644.410 1702.520 ;
        RECT 664.790 931.800 665.070 932.080 ;
        RECT 664.790 903.920 665.070 904.200 ;
        RECT 664.790 869.240 665.070 869.520 ;
        RECT 665.710 820.960 665.990 821.240 ;
        RECT 664.330 724.400 664.610 724.680 ;
        RECT 665.250 724.400 665.530 724.680 ;
        RECT 665.710 593.160 665.990 593.440 ;
        RECT 666.630 593.160 666.910 593.440 ;
        RECT 703.890 593.160 704.170 593.440 ;
      LAYER met3 ;
        RECT 589.785 2648.410 590.115 2648.425 ;
        RECT 578.070 2648.240 590.115 2648.410 ;
        RECT 574.800 2648.110 590.115 2648.240 ;
        RECT 574.800 2647.640 578.800 2648.110 ;
        RECT 589.785 2648.095 590.115 2648.110 ;
        RECT 357.485 1926.250 357.815 1926.265 ;
        RECT 360.000 1926.250 364.000 1926.400 ;
        RECT 357.485 1925.950 364.000 1926.250 ;
        RECT 357.485 1925.935 357.815 1925.950 ;
        RECT 360.000 1925.800 364.000 1925.950 ;
        RECT 1400.765 1702.530 1401.095 1702.545 ;
        RECT 1402.605 1702.530 1402.935 1702.545 ;
        RECT 1400.765 1702.230 1402.935 1702.530 ;
        RECT 1400.765 1702.215 1401.095 1702.230 ;
        RECT 1402.605 1702.215 1402.935 1702.230 ;
        RECT 1642.265 1702.530 1642.595 1702.545 ;
        RECT 1644.105 1702.530 1644.435 1702.545 ;
        RECT 1642.265 1702.230 1644.435 1702.530 ;
        RECT 1642.265 1702.215 1642.595 1702.230 ;
        RECT 1644.105 1702.215 1644.435 1702.230 ;
        RECT 664.765 932.100 665.095 932.105 ;
        RECT 664.510 932.090 665.095 932.100 ;
        RECT 664.310 931.790 665.095 932.090 ;
        RECT 664.510 931.780 665.095 931.790 ;
        RECT 664.765 931.775 665.095 931.780 ;
        RECT 664.765 904.220 665.095 904.225 ;
        RECT 664.510 904.210 665.095 904.220 ;
        RECT 664.510 903.910 665.320 904.210 ;
        RECT 664.510 903.900 665.095 903.910 ;
        RECT 664.765 903.895 665.095 903.900 ;
        RECT 664.765 869.530 665.095 869.545 ;
        RECT 665.430 869.530 665.810 869.540 ;
        RECT 664.765 869.230 665.810 869.530 ;
        RECT 664.765 869.215 665.095 869.230 ;
        RECT 665.430 869.220 665.810 869.230 ;
        RECT 665.685 821.260 666.015 821.265 ;
        RECT 665.430 821.250 666.015 821.260 ;
        RECT 665.230 820.950 666.015 821.250 ;
        RECT 665.430 820.940 666.015 820.950 ;
        RECT 665.685 820.935 666.015 820.940 ;
        RECT 664.305 724.690 664.635 724.705 ;
        RECT 665.225 724.690 665.555 724.705 ;
        RECT 664.305 724.390 665.555 724.690 ;
        RECT 664.305 724.375 664.635 724.390 ;
        RECT 665.225 724.375 665.555 724.390 ;
        RECT 665.685 593.450 666.015 593.465 ;
        RECT 666.605 593.450 666.935 593.465 ;
        RECT 703.865 593.450 704.195 593.465 ;
        RECT 665.685 593.150 704.195 593.450 ;
        RECT 665.685 593.135 666.015 593.150 ;
        RECT 666.605 593.135 666.935 593.150 ;
        RECT 703.865 593.135 704.195 593.150 ;
      LAYER via3 ;
        RECT 664.540 931.780 664.860 932.100 ;
        RECT 664.540 903.900 664.860 904.220 ;
        RECT 665.460 869.220 665.780 869.540 ;
        RECT 665.460 820.940 665.780 821.260 ;
      LAYER met4 ;
        RECT 664.535 931.775 664.865 932.105 ;
        RECT 664.550 904.225 664.850 931.775 ;
        RECT 664.535 903.895 664.865 904.225 ;
        RECT 665.455 869.215 665.785 869.545 ;
        RECT 665.470 821.265 665.770 869.215 ;
        RECT 665.455 820.935 665.785 821.265 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 645.450 2900.440 645.770 2900.500 ;
        RECT 1651.930 2900.440 1652.250 2900.500 ;
        RECT 645.450 2900.300 1652.250 2900.440 ;
        RECT 645.450 2900.240 645.770 2900.300 ;
        RECT 1651.930 2900.240 1652.250 2900.300 ;
        RECT 642.230 2608.040 642.550 2608.100 ;
        RECT 645.450 2608.040 645.770 2608.100 ;
        RECT 642.230 2607.900 645.770 2608.040 ;
        RECT 642.230 2607.840 642.550 2607.900 ;
        RECT 645.450 2607.840 645.770 2607.900 ;
        RECT 586.570 2604.640 586.890 2604.700 ;
        RECT 642.230 2604.640 642.550 2604.700 ;
        RECT 586.570 2604.500 642.550 2604.640 ;
        RECT 586.570 2604.440 586.890 2604.500 ;
        RECT 642.230 2604.440 642.550 2604.500 ;
        RECT 646.370 588.780 646.690 588.840 ;
        RECT 664.770 588.780 665.090 588.840 ;
        RECT 646.370 588.640 665.090 588.780 ;
        RECT 646.370 588.580 646.690 588.640 ;
        RECT 664.770 588.580 665.090 588.640 ;
        RECT 644.990 587.760 645.310 587.820 ;
        RECT 646.370 587.760 646.690 587.820 ;
        RECT 644.990 587.620 646.690 587.760 ;
        RECT 644.990 587.560 645.310 587.620 ;
        RECT 646.370 587.560 646.690 587.620 ;
        RECT 886.490 587.080 886.810 587.140 ;
        RECT 667.160 586.940 886.810 587.080 ;
        RECT 664.770 586.740 665.090 586.800 ;
        RECT 667.160 586.740 667.300 586.940 ;
        RECT 886.490 586.880 886.810 586.940 ;
        RECT 664.770 586.600 667.300 586.740 ;
        RECT 664.770 586.540 665.090 586.600 ;
        RECT 424.650 21.660 424.970 21.720 ;
        RECT 644.990 21.660 645.310 21.720 ;
        RECT 424.650 21.520 645.310 21.660 ;
        RECT 424.650 21.460 424.970 21.520 ;
        RECT 644.990 21.460 645.310 21.520 ;
      LAYER via ;
        RECT 645.480 2900.240 645.740 2900.500 ;
        RECT 1651.960 2900.240 1652.220 2900.500 ;
        RECT 642.260 2607.840 642.520 2608.100 ;
        RECT 645.480 2607.840 645.740 2608.100 ;
        RECT 586.600 2604.440 586.860 2604.700 ;
        RECT 642.260 2604.440 642.520 2604.700 ;
        RECT 646.400 588.580 646.660 588.840 ;
        RECT 664.800 588.580 665.060 588.840 ;
        RECT 645.020 587.560 645.280 587.820 ;
        RECT 646.400 587.560 646.660 587.820 ;
        RECT 664.800 586.540 665.060 586.800 ;
        RECT 886.520 586.880 886.780 587.140 ;
        RECT 424.680 21.460 424.940 21.720 ;
        RECT 645.020 21.460 645.280 21.720 ;
      LAYER met2 ;
        RECT 645.480 2900.210 645.740 2900.530 ;
        RECT 1651.960 2900.210 1652.220 2900.530 ;
        RECT 645.540 2608.130 645.680 2900.210 ;
        RECT 1652.020 2900.055 1652.160 2900.210 ;
        RECT 1651.890 2896.055 1652.170 2900.055 ;
        RECT 642.260 2607.810 642.520 2608.130 ;
        RECT 645.480 2607.810 645.740 2608.130 ;
        RECT 586.590 2605.235 586.870 2605.605 ;
        RECT 586.660 2604.730 586.800 2605.235 ;
        RECT 642.320 2604.730 642.460 2607.810 ;
        RECT 586.600 2604.410 586.860 2604.730 ;
        RECT 642.260 2604.410 642.520 2604.730 ;
        RECT 642.320 1866.445 642.460 2604.410 ;
        RECT 642.250 1866.075 642.530 1866.445 ;
        RECT 646.390 1866.075 646.670 1866.445 ;
        RECT 646.460 588.870 646.600 1866.075 ;
        RECT 888.130 600.170 888.410 604.000 ;
        RECT 886.580 600.030 888.410 600.170 ;
        RECT 646.400 588.550 646.660 588.870 ;
        RECT 664.800 588.550 665.060 588.870 ;
        RECT 646.460 587.850 646.600 588.550 ;
        RECT 645.020 587.530 645.280 587.850 ;
        RECT 646.400 587.530 646.660 587.850 ;
        RECT 645.080 21.750 645.220 587.530 ;
        RECT 664.860 586.830 665.000 588.550 ;
        RECT 886.580 587.170 886.720 600.030 ;
        RECT 888.130 600.000 888.410 600.030 ;
        RECT 886.520 586.850 886.780 587.170 ;
        RECT 664.800 586.510 665.060 586.830 ;
        RECT 424.680 21.430 424.940 21.750 ;
        RECT 645.020 21.430 645.280 21.750 ;
        RECT 424.740 2.400 424.880 21.430 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 586.590 2605.280 586.870 2605.560 ;
        RECT 642.250 1866.120 642.530 1866.400 ;
        RECT 646.390 1866.120 646.670 1866.400 ;
      LAYER met3 ;
        RECT 574.800 2605.570 578.800 2606.080 ;
        RECT 586.565 2605.570 586.895 2605.585 ;
        RECT 574.800 2605.480 586.895 2605.570 ;
        RECT 578.070 2605.270 586.895 2605.480 ;
        RECT 586.565 2605.255 586.895 2605.270 ;
        RECT 627.030 1866.410 631.030 1866.560 ;
        RECT 642.225 1866.410 642.555 1866.425 ;
        RECT 646.365 1866.410 646.695 1866.425 ;
        RECT 627.030 1866.110 646.695 1866.410 ;
        RECT 627.030 1865.960 631.030 1866.110 ;
        RECT 642.225 1866.095 642.555 1866.110 ;
        RECT 646.365 1866.095 646.695 1866.110 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 2898.740 427.730 2898.800 ;
        RECT 1671.710 2898.740 1672.030 2898.800 ;
        RECT 427.410 2898.600 1672.030 2898.740 ;
        RECT 427.410 2898.540 427.730 2898.600 ;
        RECT 1671.710 2898.540 1672.030 2898.600 ;
        RECT 351.050 2622.320 351.370 2622.380 ;
        RECT 427.410 2622.320 427.730 2622.380 ;
        RECT 351.050 2622.180 427.730 2622.320 ;
        RECT 351.050 2622.120 351.370 2622.180 ;
        RECT 427.410 2622.120 427.730 2622.180 ;
        RECT 357.950 591.840 358.270 591.900 ;
        RECT 441.670 591.840 441.990 591.900 ;
        RECT 357.950 591.700 441.990 591.840 ;
        RECT 357.950 591.640 358.270 591.700 ;
        RECT 441.670 591.640 441.990 591.700 ;
        RECT 441.670 590.140 441.990 590.200 ;
        RECT 897.530 590.140 897.850 590.200 ;
        RECT 441.670 590.000 593.700 590.140 ;
        RECT 441.670 589.940 441.990 590.000 ;
        RECT 593.560 589.800 593.700 590.000 ;
        RECT 629.440 590.000 664.540 590.140 ;
        RECT 629.440 589.800 629.580 590.000 ;
        RECT 593.560 589.660 629.580 589.800 ;
        RECT 664.400 589.800 664.540 590.000 ;
        RECT 665.320 590.000 897.850 590.140 ;
        RECT 665.320 589.800 665.460 590.000 ;
        RECT 897.530 589.940 897.850 590.000 ;
        RECT 664.400 589.660 665.460 589.800 ;
        RECT 441.670 2.960 441.990 3.020 ;
        RECT 442.590 2.960 442.910 3.020 ;
        RECT 441.670 2.820 442.910 2.960 ;
        RECT 441.670 2.760 441.990 2.820 ;
        RECT 442.590 2.760 442.910 2.820 ;
      LAYER via ;
        RECT 427.440 2898.540 427.700 2898.800 ;
        RECT 1671.740 2898.540 1672.000 2898.800 ;
        RECT 351.080 2622.120 351.340 2622.380 ;
        RECT 427.440 2622.120 427.700 2622.380 ;
        RECT 357.980 591.640 358.240 591.900 ;
        RECT 441.700 591.640 441.960 591.900 ;
        RECT 441.700 589.940 441.960 590.200 ;
        RECT 897.560 589.940 897.820 590.200 ;
        RECT 441.700 2.760 441.960 3.020 ;
        RECT 442.620 2.760 442.880 3.020 ;
      LAYER met2 ;
        RECT 427.440 2898.510 427.700 2898.830 ;
        RECT 1671.740 2898.570 1672.000 2898.830 ;
        RECT 1673.050 2898.570 1673.330 2900.055 ;
        RECT 1671.740 2898.510 1673.330 2898.570 ;
        RECT 427.500 2624.985 427.640 2898.510 ;
        RECT 1671.800 2898.430 1673.330 2898.510 ;
        RECT 1673.050 2896.055 1673.330 2898.430 ;
        RECT 427.430 2624.615 427.710 2624.985 ;
        RECT 427.500 2622.410 427.640 2624.615 ;
        RECT 351.080 2622.090 351.340 2622.410 ;
        RECT 427.440 2622.090 427.700 2622.410 ;
        RECT 351.140 1741.325 351.280 2622.090 ;
        RECT 351.070 1740.955 351.350 1741.325 ;
        RECT 357.970 1740.955 358.250 1741.325 ;
        RECT 358.040 591.930 358.180 1740.955 ;
        RECT 897.330 600.000 897.610 604.000 ;
        RECT 897.390 598.810 897.530 600.000 ;
        RECT 897.390 598.670 897.760 598.810 ;
        RECT 357.980 591.610 358.240 591.930 ;
        RECT 441.700 591.610 441.960 591.930 ;
        RECT 441.760 590.230 441.900 591.610 ;
        RECT 897.620 590.230 897.760 598.670 ;
        RECT 441.700 589.910 441.960 590.230 ;
        RECT 897.560 589.910 897.820 590.230 ;
        RECT 441.760 3.050 441.900 589.910 ;
        RECT 441.700 2.730 441.960 3.050 ;
        RECT 442.620 2.730 442.880 3.050 ;
        RECT 442.680 2.400 442.820 2.730 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 427.430 2624.660 427.710 2624.940 ;
        RECT 351.070 1741.000 351.350 1741.280 ;
        RECT 357.970 1741.000 358.250 1741.280 ;
      LAYER met3 ;
        RECT 427.405 2624.950 427.735 2624.965 ;
        RECT 430.000 2624.950 434.000 2625.120 ;
        RECT 427.405 2624.650 434.000 2624.950 ;
        RECT 427.405 2624.635 427.735 2624.650 ;
        RECT 430.000 2624.520 434.000 2624.650 ;
        RECT 351.045 1741.290 351.375 1741.305 ;
        RECT 357.945 1741.290 358.275 1741.305 ;
        RECT 360.000 1741.290 364.000 1741.440 ;
        RECT 351.045 1740.990 364.000 1741.290 ;
        RECT 351.045 1740.975 351.375 1740.990 ;
        RECT 357.945 1740.975 358.275 1740.990 ;
        RECT 360.000 1740.840 364.000 1740.990 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.450 2591.040 461.770 2591.100 ;
        RECT 635.330 2591.040 635.650 2591.100 ;
        RECT 1487.710 2591.040 1488.030 2591.100 ;
        RECT 461.450 2590.900 1488.030 2591.040 ;
        RECT 461.450 2590.840 461.770 2590.900 ;
        RECT 635.330 2590.840 635.650 2590.900 ;
        RECT 1487.710 2590.840 1488.030 2590.900 ;
        RECT 489.510 1690.040 489.830 1690.100 ;
        RECT 635.330 1690.040 635.650 1690.100 ;
        RECT 489.510 1689.900 635.650 1690.040 ;
        RECT 489.510 1689.840 489.830 1689.900 ;
        RECT 635.330 1689.840 635.650 1689.900 ;
        RECT 489.510 592.860 489.830 592.920 ;
        RECT 904.890 592.860 905.210 592.920 ;
        RECT 489.510 592.720 905.210 592.860 ;
        RECT 489.510 592.660 489.830 592.720 ;
        RECT 904.890 592.660 905.210 592.720 ;
        RECT 461.910 586.740 462.230 586.800 ;
        RECT 489.510 586.740 489.830 586.800 ;
        RECT 461.910 586.600 489.830 586.740 ;
        RECT 461.910 586.540 462.230 586.600 ;
        RECT 489.510 586.540 489.830 586.600 ;
        RECT 460.530 2.960 460.850 3.020 ;
        RECT 461.910 2.960 462.230 3.020 ;
        RECT 460.530 2.820 462.230 2.960 ;
        RECT 460.530 2.760 460.850 2.820 ;
        RECT 461.910 2.760 462.230 2.820 ;
      LAYER via ;
        RECT 461.480 2590.840 461.740 2591.100 ;
        RECT 635.360 2590.840 635.620 2591.100 ;
        RECT 1487.740 2590.840 1488.000 2591.100 ;
        RECT 489.540 1689.840 489.800 1690.100 ;
        RECT 635.360 1689.840 635.620 1690.100 ;
        RECT 489.540 592.660 489.800 592.920 ;
        RECT 904.920 592.660 905.180 592.920 ;
        RECT 461.940 586.540 462.200 586.800 ;
        RECT 489.540 586.540 489.800 586.800 ;
        RECT 460.560 2.760 460.820 3.020 ;
        RECT 461.940 2.760 462.200 3.020 ;
      LAYER met2 ;
        RECT 1487.730 2643.995 1488.010 2644.365 ;
        RECT 461.370 2600.660 461.650 2604.000 ;
        RECT 461.370 2600.000 461.680 2600.660 ;
        RECT 461.540 2591.130 461.680 2600.000 ;
        RECT 1487.800 2591.130 1487.940 2643.995 ;
        RECT 461.480 2590.810 461.740 2591.130 ;
        RECT 635.360 2590.810 635.620 2591.130 ;
        RECT 1487.740 2590.810 1488.000 2591.130 ;
        RECT 487.970 1700.410 488.250 1704.000 ;
        RECT 487.970 1700.270 489.740 1700.410 ;
        RECT 487.970 1700.000 488.250 1700.270 ;
        RECT 489.600 1690.130 489.740 1700.270 ;
        RECT 635.420 1690.130 635.560 2590.810 ;
        RECT 489.540 1689.810 489.800 1690.130 ;
        RECT 635.360 1689.810 635.620 1690.130 ;
        RECT 489.600 592.950 489.740 1689.810 ;
        RECT 906.530 600.170 906.810 604.000 ;
        RECT 904.980 600.030 906.810 600.170 ;
        RECT 904.980 592.950 905.120 600.030 ;
        RECT 906.530 600.000 906.810 600.030 ;
        RECT 489.540 592.630 489.800 592.950 ;
        RECT 904.920 592.630 905.180 592.950 ;
        RECT 489.600 586.830 489.740 592.630 ;
        RECT 461.940 586.510 462.200 586.830 ;
        RECT 489.540 586.510 489.800 586.830 ;
        RECT 462.000 3.050 462.140 586.510 ;
        RECT 460.560 2.730 460.820 3.050 ;
        RECT 461.940 2.730 462.200 3.050 ;
        RECT 460.620 2.400 460.760 2.730 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 1487.730 2644.040 1488.010 2644.320 ;
      LAYER met3 ;
        RECT 1500.000 2645.880 1504.000 2646.160 ;
        RECT 1499.910 2645.560 1504.000 2645.880 ;
        RECT 1487.705 2644.330 1488.035 2644.345 ;
        RECT 1499.910 2644.330 1500.210 2645.560 ;
        RECT 1487.705 2644.030 1500.210 2644.330 ;
        RECT 1487.705 2644.015 1488.035 2644.030 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 2900.100 645.310 2900.160 ;
        RECT 1736.110 2900.100 1736.430 2900.160 ;
        RECT 644.990 2899.960 1736.430 2900.100 ;
        RECT 644.990 2899.900 645.310 2899.960 ;
        RECT 1736.110 2899.900 1736.430 2899.960 ;
        RECT 575.530 2769.200 575.850 2769.260 ;
        RECT 641.770 2769.200 642.090 2769.260 ;
        RECT 575.530 2769.060 642.090 2769.200 ;
        RECT 575.530 2769.000 575.850 2769.060 ;
        RECT 641.770 2769.000 642.090 2769.060 ;
        RECT 641.770 2767.160 642.090 2767.220 ;
        RECT 644.990 2767.160 645.310 2767.220 ;
        RECT 641.770 2767.020 645.310 2767.160 ;
        RECT 641.770 2766.960 642.090 2767.020 ;
        RECT 644.990 2766.960 645.310 2767.020 ;
        RECT 667.530 591.500 667.850 591.560 ;
        RECT 914.090 591.500 914.410 591.560 ;
        RECT 667.530 591.360 914.410 591.500 ;
        RECT 667.530 591.300 667.850 591.360 ;
        RECT 914.090 591.300 914.410 591.360 ;
        RECT 644.530 589.800 644.850 589.860 ;
        RECT 646.830 589.800 647.150 589.860 ;
        RECT 661.550 589.800 661.870 589.860 ;
        RECT 644.530 589.660 661.870 589.800 ;
        RECT 644.530 589.600 644.850 589.660 ;
        RECT 646.830 589.600 647.150 589.660 ;
        RECT 661.550 589.600 661.870 589.660 ;
        RECT 478.470 43.420 478.790 43.480 ;
        RECT 646.830 43.420 647.150 43.480 ;
        RECT 478.470 43.280 647.150 43.420 ;
        RECT 478.470 43.220 478.790 43.280 ;
        RECT 646.830 43.220 647.150 43.280 ;
      LAYER via ;
        RECT 645.020 2899.900 645.280 2900.160 ;
        RECT 1736.140 2899.900 1736.400 2900.160 ;
        RECT 575.560 2769.000 575.820 2769.260 ;
        RECT 641.800 2769.000 642.060 2769.260 ;
        RECT 641.800 2766.960 642.060 2767.220 ;
        RECT 645.020 2766.960 645.280 2767.220 ;
        RECT 667.560 591.300 667.820 591.560 ;
        RECT 914.120 591.300 914.380 591.560 ;
        RECT 644.560 589.600 644.820 589.860 ;
        RECT 646.860 589.600 647.120 589.860 ;
        RECT 661.580 589.600 661.840 589.860 ;
        RECT 478.500 43.220 478.760 43.480 ;
        RECT 646.860 43.220 647.120 43.480 ;
      LAYER met2 ;
        RECT 645.020 2899.870 645.280 2900.190 ;
        RECT 1736.140 2899.930 1736.400 2900.190 ;
        RECT 1737.450 2899.930 1737.730 2900.055 ;
        RECT 1736.140 2899.870 1737.730 2899.930 ;
        RECT 575.560 2768.970 575.820 2769.290 ;
        RECT 641.800 2768.970 642.060 2769.290 ;
        RECT 575.620 2759.520 575.760 2768.970 ;
        RECT 641.860 2767.250 642.000 2768.970 ;
        RECT 645.080 2767.250 645.220 2899.870 ;
        RECT 1736.200 2899.790 1737.730 2899.870 ;
        RECT 1737.450 2896.055 1737.730 2899.790 ;
        RECT 641.800 2766.930 642.060 2767.250 ;
        RECT 645.020 2766.930 645.280 2767.250 ;
        RECT 575.450 2759.100 575.760 2759.520 ;
        RECT 575.450 2755.520 575.730 2759.100 ;
        RECT 641.860 1791.645 642.000 2766.930 ;
        RECT 641.790 1791.275 642.070 1791.645 ;
        RECT 644.550 1791.275 644.830 1791.645 ;
        RECT 644.620 589.890 644.760 1791.275 ;
        RECT 915.730 600.170 916.010 604.000 ;
        RECT 914.180 600.030 916.010 600.170 ;
        RECT 914.180 591.590 914.320 600.030 ;
        RECT 915.730 600.000 916.010 600.030 ;
        RECT 667.560 591.270 667.820 591.590 ;
        RECT 914.120 591.270 914.380 591.590 ;
        RECT 644.560 589.570 644.820 589.890 ;
        RECT 646.860 589.570 647.120 589.890 ;
        RECT 661.580 589.570 661.840 589.890 ;
        RECT 646.920 43.510 647.060 589.570 ;
        RECT 661.640 589.405 661.780 589.570 ;
        RECT 667.620 589.405 667.760 591.270 ;
        RECT 661.570 589.035 661.850 589.405 ;
        RECT 667.550 589.035 667.830 589.405 ;
        RECT 478.500 43.190 478.760 43.510 ;
        RECT 646.860 43.190 647.120 43.510 ;
        RECT 478.560 2.400 478.700 43.190 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 641.790 1791.320 642.070 1791.600 ;
        RECT 644.550 1791.320 644.830 1791.600 ;
        RECT 661.570 589.080 661.850 589.360 ;
        RECT 667.550 589.080 667.830 589.360 ;
      LAYER met3 ;
        RECT 627.030 1791.610 631.030 1791.760 ;
        RECT 641.765 1791.610 642.095 1791.625 ;
        RECT 644.525 1791.610 644.855 1791.625 ;
        RECT 627.030 1791.310 644.855 1791.610 ;
        RECT 627.030 1791.160 631.030 1791.310 ;
        RECT 641.765 1791.295 642.095 1791.310 ;
        RECT 644.525 1791.295 644.855 1791.310 ;
        RECT 661.545 589.370 661.875 589.385 ;
        RECT 667.525 589.370 667.855 589.385 ;
        RECT 661.545 589.070 667.855 589.370 ;
        RECT 661.545 589.055 661.875 589.070 ;
        RECT 667.525 589.055 667.855 589.070 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 1687.320 389.550 1687.380 ;
        RECT 496.410 1687.320 496.730 1687.380 ;
        RECT 1649.170 1687.320 1649.490 1687.380 ;
        RECT 389.230 1687.180 1649.490 1687.320 ;
        RECT 389.230 1687.120 389.550 1687.180 ;
        RECT 496.410 1687.120 496.730 1687.180 ;
        RECT 1649.170 1687.120 1649.490 1687.180 ;
        RECT 489.970 16.900 490.290 16.960 ;
        RECT 496.410 16.900 496.730 16.960 ;
        RECT 489.970 16.760 496.730 16.900 ;
        RECT 489.970 16.700 490.290 16.760 ;
        RECT 496.410 16.700 496.730 16.760 ;
      LAYER via ;
        RECT 389.260 1687.120 389.520 1687.380 ;
        RECT 496.440 1687.120 496.700 1687.380 ;
        RECT 1649.200 1687.120 1649.460 1687.380 ;
        RECT 490.000 16.700 490.260 16.960 ;
        RECT 496.440 16.700 496.700 16.960 ;
      LAYER met2 ;
        RECT 1650.970 2500.090 1651.250 2504.000 ;
        RECT 1649.260 2500.000 1651.250 2500.090 ;
        RECT 1649.260 2499.950 1651.170 2500.000 ;
        RECT 387.690 1700.410 387.970 1704.000 ;
        RECT 387.690 1700.270 389.460 1700.410 ;
        RECT 387.690 1700.000 387.970 1700.270 ;
        RECT 389.320 1687.410 389.460 1700.270 ;
        RECT 1649.260 1687.410 1649.400 2499.950 ;
        RECT 389.260 1687.090 389.520 1687.410 ;
        RECT 496.440 1687.090 496.700 1687.410 ;
        RECT 1649.200 1687.090 1649.460 1687.410 ;
        RECT 496.500 590.085 496.640 1687.090 ;
        RECT 924.930 600.000 925.210 604.000 ;
        RECT 924.990 598.810 925.130 600.000 ;
        RECT 924.990 598.670 925.360 598.810 ;
        RECT 489.990 589.715 490.270 590.085 ;
        RECT 496.430 589.715 496.710 590.085 ;
        RECT 490.060 16.990 490.200 589.715 ;
        RECT 925.220 589.405 925.360 598.670 ;
        RECT 744.830 589.035 745.110 589.405 ;
        RECT 925.150 589.035 925.430 589.405 ;
        RECT 565.890 588.355 566.170 588.725 ;
        RECT 695.610 588.355 695.890 588.725 ;
        RECT 565.960 588.045 566.100 588.355 ;
        RECT 695.680 588.045 695.820 588.355 ;
        RECT 565.890 587.675 566.170 588.045 ;
        RECT 649.150 587.675 649.430 588.045 ;
        RECT 695.610 587.675 695.890 588.045 ;
        RECT 648.690 587.250 648.970 587.365 ;
        RECT 649.220 587.250 649.360 587.675 ;
        RECT 744.900 587.365 745.040 589.035 ;
        RECT 648.690 587.110 649.360 587.250 ;
        RECT 648.690 586.995 648.970 587.110 ;
        RECT 744.830 586.995 745.110 587.365 ;
        RECT 490.000 16.670 490.260 16.990 ;
        RECT 496.440 16.670 496.700 16.990 ;
        RECT 496.500 2.400 496.640 16.670 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 489.990 589.760 490.270 590.040 ;
        RECT 496.430 589.760 496.710 590.040 ;
        RECT 744.830 589.080 745.110 589.360 ;
        RECT 925.150 589.080 925.430 589.360 ;
        RECT 565.890 588.400 566.170 588.680 ;
        RECT 695.610 588.400 695.890 588.680 ;
        RECT 565.890 587.720 566.170 588.000 ;
        RECT 649.150 587.720 649.430 588.000 ;
        RECT 695.610 587.720 695.890 588.000 ;
        RECT 648.690 587.040 648.970 587.320 ;
        RECT 744.830 587.040 745.110 587.320 ;
      LAYER met3 ;
        RECT 489.965 590.050 490.295 590.065 ;
        RECT 496.405 590.050 496.735 590.065 ;
        RECT 489.965 589.750 546.170 590.050 ;
        RECT 489.965 589.735 490.295 589.750 ;
        RECT 496.405 589.735 496.735 589.750 ;
        RECT 545.870 588.690 546.170 589.750 ;
        RECT 744.805 589.370 745.135 589.385 ;
        RECT 925.125 589.370 925.455 589.385 ;
        RECT 744.805 589.070 745.810 589.370 ;
        RECT 744.805 589.055 745.135 589.070 ;
        RECT 565.865 588.690 566.195 588.705 ;
        RECT 545.870 588.390 566.195 588.690 ;
        RECT 565.865 588.375 566.195 588.390 ;
        RECT 695.585 588.690 695.915 588.705 ;
        RECT 696.710 588.690 697.090 588.700 ;
        RECT 695.585 588.390 697.090 588.690 ;
        RECT 745.510 588.690 745.810 589.070 ;
        RECT 808.070 589.070 925.455 589.370 ;
        RECT 808.070 588.860 808.370 589.070 ;
        RECT 925.125 589.055 925.455 589.070 ;
        RECT 807.150 588.690 808.370 588.860 ;
        RECT 745.510 588.560 808.370 588.690 ;
        RECT 745.510 588.390 807.450 588.560 ;
        RECT 695.585 588.375 695.915 588.390 ;
        RECT 696.710 588.380 697.090 588.390 ;
        RECT 565.865 588.010 566.195 588.025 ;
        RECT 649.125 588.010 649.455 588.025 ;
        RECT 695.585 588.010 695.915 588.025 ;
        RECT 565.865 587.710 588.490 588.010 ;
        RECT 565.865 587.695 566.195 587.710 ;
        RECT 588.190 587.330 588.490 587.710 ;
        RECT 649.125 587.710 695.915 588.010 ;
        RECT 649.125 587.695 649.455 587.710 ;
        RECT 695.585 587.695 695.915 587.710 ;
        RECT 648.665 587.330 648.995 587.345 ;
        RECT 588.190 587.030 648.995 587.330 ;
        RECT 648.665 587.015 648.995 587.030 ;
        RECT 696.710 587.330 697.090 587.340 ;
        RECT 744.805 587.330 745.135 587.345 ;
        RECT 696.710 587.030 745.135 587.330 ;
        RECT 696.710 587.020 697.090 587.030 ;
        RECT 744.805 587.015 745.135 587.030 ;
      LAYER via3 ;
        RECT 696.740 588.380 697.060 588.700 ;
        RECT 696.740 587.020 697.060 587.340 ;
      LAYER met4 ;
        RECT 696.735 588.375 697.065 588.705 ;
        RECT 696.750 587.345 697.050 588.375 ;
        RECT 696.735 587.015 697.065 587.345 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1497.830 2452.320 1498.150 2452.380 ;
        RECT 1502.890 2452.320 1503.210 2452.380 ;
        RECT 1497.830 2452.180 1503.210 2452.320 ;
        RECT 1497.830 2452.120 1498.150 2452.180 ;
        RECT 1502.890 2452.120 1503.210 2452.180 ;
        RECT 364.390 1687.660 364.710 1687.720 ;
        RECT 650.970 1687.660 651.290 1687.720 ;
        RECT 1497.830 1687.660 1498.150 1687.720 ;
        RECT 364.390 1687.520 1498.150 1687.660 ;
        RECT 364.390 1687.460 364.710 1687.520 ;
        RECT 650.970 1687.460 651.290 1687.520 ;
        RECT 1497.830 1687.460 1498.150 1687.520 ;
        RECT 650.970 670.380 651.290 670.440 ;
        RECT 660.170 670.380 660.490 670.440 ;
        RECT 650.970 670.240 660.490 670.380 ;
        RECT 650.970 670.180 651.290 670.240 ;
        RECT 660.170 670.180 660.490 670.240 ;
        RECT 851.990 601.700 852.310 601.760 ;
        RECT 932.030 601.700 932.350 601.760 ;
        RECT 933.410 601.700 933.730 601.760 ;
        RECT 738.000 601.560 756.080 601.700 ;
        RECT 738.000 601.360 738.140 601.560 ;
        RECT 714.540 601.220 738.140 601.360 ;
        RECT 755.940 601.360 756.080 601.560 ;
        RECT 851.990 601.560 933.730 601.700 ;
        RECT 851.990 601.500 852.310 601.560 ;
        RECT 932.030 601.500 932.350 601.560 ;
        RECT 933.410 601.500 933.730 601.560 ;
        RECT 834.970 601.360 835.290 601.420 ;
        RECT 755.940 601.220 835.290 601.360 ;
        RECT 660.630 600.000 660.950 600.060 ;
        RECT 714.540 600.000 714.680 601.220 ;
        RECT 834.970 601.160 835.290 601.220 ;
        RECT 660.630 599.860 714.680 600.000 ;
        RECT 834.970 600.000 835.290 600.060 ;
        RECT 851.990 600.000 852.310 600.060 ;
        RECT 834.970 599.860 852.310 600.000 ;
        RECT 660.630 599.800 660.950 599.860 ;
        RECT 834.970 599.800 835.290 599.860 ;
        RECT 851.990 599.800 852.310 599.860 ;
        RECT 931.110 572.460 931.430 572.520 ;
        RECT 932.030 572.460 932.350 572.520 ;
        RECT 931.110 572.320 932.350 572.460 ;
        RECT 931.110 572.260 931.430 572.320 ;
        RECT 932.030 572.260 932.350 572.320 ;
        RECT 931.110 524.520 931.430 524.580 ;
        RECT 932.490 524.520 932.810 524.580 ;
        RECT 931.110 524.380 932.810 524.520 ;
        RECT 931.110 524.320 931.430 524.380 ;
        RECT 932.490 524.320 932.810 524.380 ;
        RECT 931.110 186.220 931.430 186.280 ;
        RECT 932.490 186.220 932.810 186.280 ;
        RECT 931.110 186.080 932.810 186.220 ;
        RECT 931.110 186.020 931.430 186.080 ;
        RECT 932.490 186.020 932.810 186.080 ;
        RECT 931.110 138.280 931.430 138.340 ;
        RECT 932.030 138.280 932.350 138.340 ;
        RECT 931.110 138.140 932.350 138.280 ;
        RECT 931.110 138.080 931.430 138.140 ;
        RECT 932.030 138.080 932.350 138.140 ;
        RECT 932.030 110.540 932.350 110.800 ;
        RECT 932.120 110.400 932.260 110.540 ;
        RECT 932.490 110.400 932.810 110.460 ;
        RECT 932.120 110.260 932.810 110.400 ;
        RECT 932.490 110.200 932.810 110.260 ;
        RECT 513.890 34.240 514.210 34.300 ;
        RECT 932.490 34.240 932.810 34.300 ;
        RECT 513.890 34.100 932.810 34.240 ;
        RECT 513.890 34.040 514.210 34.100 ;
        RECT 932.490 34.040 932.810 34.100 ;
      LAYER via ;
        RECT 1497.860 2452.120 1498.120 2452.380 ;
        RECT 1502.920 2452.120 1503.180 2452.380 ;
        RECT 364.420 1687.460 364.680 1687.720 ;
        RECT 651.000 1687.460 651.260 1687.720 ;
        RECT 1497.860 1687.460 1498.120 1687.720 ;
        RECT 651.000 670.180 651.260 670.440 ;
        RECT 660.200 670.180 660.460 670.440 ;
        RECT 852.020 601.500 852.280 601.760 ;
        RECT 932.060 601.500 932.320 601.760 ;
        RECT 933.440 601.500 933.700 601.760 ;
        RECT 660.660 599.800 660.920 600.060 ;
        RECT 835.000 601.160 835.260 601.420 ;
        RECT 835.000 599.800 835.260 600.060 ;
        RECT 852.020 599.800 852.280 600.060 ;
        RECT 931.140 572.260 931.400 572.520 ;
        RECT 932.060 572.260 932.320 572.520 ;
        RECT 931.140 524.320 931.400 524.580 ;
        RECT 932.520 524.320 932.780 524.580 ;
        RECT 931.140 186.020 931.400 186.280 ;
        RECT 932.520 186.020 932.780 186.280 ;
        RECT 931.140 138.080 931.400 138.340 ;
        RECT 932.060 138.080 932.320 138.340 ;
        RECT 932.060 110.540 932.320 110.800 ;
        RECT 932.520 110.200 932.780 110.460 ;
        RECT 513.920 34.040 514.180 34.300 ;
        RECT 932.520 34.040 932.780 34.300 ;
      LAYER met2 ;
        RECT 1502.850 2500.000 1503.130 2504.000 ;
        RECT 1502.980 2452.410 1503.120 2500.000 ;
        RECT 1497.860 2452.090 1498.120 2452.410 ;
        RECT 1502.920 2452.090 1503.180 2452.410 ;
        RECT 362.850 1700.410 363.130 1704.000 ;
        RECT 362.850 1700.270 364.620 1700.410 ;
        RECT 362.850 1700.000 363.130 1700.270 ;
        RECT 364.480 1687.750 364.620 1700.270 ;
        RECT 1497.920 1687.750 1498.060 2452.090 ;
        RECT 364.420 1687.430 364.680 1687.750 ;
        RECT 651.000 1687.430 651.260 1687.750 ;
        RECT 1497.860 1687.430 1498.120 1687.750 ;
        RECT 651.060 670.470 651.200 1687.430 ;
        RECT 651.000 670.150 651.260 670.470 ;
        RECT 660.200 670.150 660.460 670.470 ;
        RECT 660.260 665.450 660.400 670.150 ;
        RECT 660.260 665.310 660.860 665.450 ;
        RECT 660.720 600.090 660.860 665.310 ;
        RECT 852.020 601.470 852.280 601.790 ;
        RECT 932.060 601.470 932.320 601.790 ;
        RECT 933.440 601.530 933.700 601.790 ;
        RECT 934.130 601.530 934.410 604.000 ;
        RECT 933.440 601.470 934.410 601.530 ;
        RECT 835.000 601.130 835.260 601.450 ;
        RECT 835.060 600.090 835.200 601.130 ;
        RECT 852.080 600.090 852.220 601.470 ;
        RECT 660.660 599.770 660.920 600.090 ;
        RECT 835.000 599.770 835.260 600.090 ;
        RECT 852.020 599.770 852.280 600.090 ;
        RECT 932.120 572.550 932.260 601.470 ;
        RECT 933.500 601.390 934.410 601.470 ;
        RECT 934.130 600.000 934.410 601.390 ;
        RECT 931.140 572.230 931.400 572.550 ;
        RECT 932.060 572.230 932.320 572.550 ;
        RECT 931.200 524.610 931.340 572.230 ;
        RECT 931.140 524.290 931.400 524.610 ;
        RECT 932.520 524.290 932.780 524.610 ;
        RECT 932.580 314.570 932.720 524.290 ;
        RECT 932.120 314.430 932.720 314.570 ;
        RECT 932.120 313.210 932.260 314.430 ;
        RECT 932.120 313.070 932.720 313.210 ;
        RECT 932.580 207.130 932.720 313.070 ;
        RECT 932.120 206.990 932.720 207.130 ;
        RECT 932.120 206.450 932.260 206.990 ;
        RECT 932.120 206.310 932.720 206.450 ;
        RECT 932.580 186.310 932.720 206.310 ;
        RECT 931.140 185.990 931.400 186.310 ;
        RECT 932.520 185.990 932.780 186.310 ;
        RECT 931.200 138.370 931.340 185.990 ;
        RECT 931.140 138.050 931.400 138.370 ;
        RECT 932.060 138.050 932.320 138.370 ;
        RECT 932.120 110.830 932.260 138.050 ;
        RECT 932.060 110.510 932.320 110.830 ;
        RECT 932.520 110.170 932.780 110.490 ;
        RECT 932.580 34.330 932.720 110.170 ;
        RECT 513.920 34.010 514.180 34.330 ;
        RECT 932.520 34.010 932.780 34.330 ;
        RECT 513.980 2.400 514.120 34.010 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 941.690 2039.220 942.010 2039.280 ;
        RECT 1902.630 2039.220 1902.950 2039.280 ;
        RECT 941.690 2039.080 1902.950 2039.220 ;
        RECT 941.690 2039.020 942.010 2039.080 ;
        RECT 1902.630 2039.020 1902.950 2039.080 ;
        RECT 927.890 1780.140 928.210 1780.200 ;
        RECT 941.690 1780.140 942.010 1780.200 ;
        RECT 927.890 1780.000 942.010 1780.140 ;
        RECT 927.890 1779.940 928.210 1780.000 ;
        RECT 941.690 1779.940 942.010 1780.000 ;
        RECT 350.590 1707.720 350.910 1707.780 ;
        RECT 651.430 1707.720 651.750 1707.780 ;
        RECT 927.890 1707.720 928.210 1707.780 ;
        RECT 350.590 1707.580 928.210 1707.720 ;
        RECT 350.590 1707.520 350.910 1707.580 ;
        RECT 651.430 1707.520 651.750 1707.580 ;
        RECT 927.890 1707.520 928.210 1707.580 ;
        RECT 651.430 624.820 651.750 624.880 ;
        RECT 659.710 624.820 660.030 624.880 ;
        RECT 651.430 624.680 660.030 624.820 ;
        RECT 651.430 624.620 651.750 624.680 ;
        RECT 659.710 624.620 660.030 624.680 ;
        RECT 695.680 602.240 834.740 602.380 ;
        RECT 659.710 600.680 660.030 600.740 ;
        RECT 695.680 600.680 695.820 602.240 ;
        RECT 834.600 601.760 834.740 602.240 ;
        RECT 851.390 602.240 893.620 602.380 ;
        RECT 834.510 601.500 834.830 601.760 ;
        RECT 834.510 601.020 834.830 601.080 ;
        RECT 851.390 601.020 851.530 602.240 ;
        RECT 893.480 602.040 893.620 602.240 ;
        RECT 893.480 601.900 938.700 602.040 ;
        RECT 938.560 601.760 938.700 601.900 ;
        RECT 938.470 601.500 938.790 601.760 ;
        RECT 834.510 600.880 851.530 601.020 ;
        RECT 834.510 600.820 834.830 600.880 ;
        RECT 659.710 600.540 695.820 600.680 ;
        RECT 938.470 600.680 938.790 600.740 ;
        RECT 941.690 600.680 942.010 600.740 ;
        RECT 938.470 600.540 942.010 600.680 ;
        RECT 659.710 600.480 660.030 600.540 ;
        RECT 938.470 600.480 938.790 600.540 ;
        RECT 941.690 600.480 942.010 600.540 ;
        RECT 531.830 29.480 532.150 29.540 ;
        RECT 938.470 29.480 938.790 29.540 ;
        RECT 531.830 29.340 938.790 29.480 ;
        RECT 531.830 29.280 532.150 29.340 ;
        RECT 938.470 29.280 938.790 29.340 ;
      LAYER via ;
        RECT 941.720 2039.020 941.980 2039.280 ;
        RECT 1902.660 2039.020 1902.920 2039.280 ;
        RECT 927.920 1779.940 928.180 1780.200 ;
        RECT 941.720 1779.940 941.980 1780.200 ;
        RECT 350.620 1707.520 350.880 1707.780 ;
        RECT 651.460 1707.520 651.720 1707.780 ;
        RECT 927.920 1707.520 928.180 1707.780 ;
        RECT 651.460 624.620 651.720 624.880 ;
        RECT 659.740 624.620 660.000 624.880 ;
        RECT 659.740 600.480 660.000 600.740 ;
        RECT 834.540 601.500 834.800 601.760 ;
        RECT 834.540 600.820 834.800 601.080 ;
        RECT 938.500 601.500 938.760 601.760 ;
        RECT 938.500 600.480 938.760 600.740 ;
        RECT 941.720 600.480 941.980 600.740 ;
        RECT 531.860 29.280 532.120 29.540 ;
        RECT 938.500 29.280 938.760 29.540 ;
      LAYER met2 ;
        RECT 1902.650 2877.235 1902.930 2877.605 ;
        RECT 1902.720 2039.310 1902.860 2877.235 ;
        RECT 941.720 2038.990 941.980 2039.310 ;
        RECT 1902.660 2038.990 1902.920 2039.310 ;
        RECT 941.780 1780.230 941.920 2038.990 ;
        RECT 927.920 1779.910 928.180 1780.230 ;
        RECT 941.720 1779.910 941.980 1780.230 ;
        RECT 350.610 1777.675 350.890 1778.045 ;
        RECT 350.680 1707.810 350.820 1777.675 ;
        RECT 927.980 1707.810 928.120 1779.910 ;
        RECT 350.620 1707.490 350.880 1707.810 ;
        RECT 651.460 1707.490 651.720 1707.810 ;
        RECT 927.920 1707.490 928.180 1707.810 ;
        RECT 651.520 624.910 651.660 1707.490 ;
        RECT 651.460 624.590 651.720 624.910 ;
        RECT 659.740 624.590 660.000 624.910 ;
        RECT 659.800 600.770 659.940 624.590 ;
        RECT 834.540 601.470 834.800 601.790 ;
        RECT 938.500 601.470 938.760 601.790 ;
        RECT 834.600 601.110 834.740 601.470 ;
        RECT 834.540 600.790 834.800 601.110 ;
        RECT 938.560 600.770 938.700 601.470 ;
        RECT 943.330 600.850 943.610 604.000 ;
        RECT 941.780 600.770 943.610 600.850 ;
        RECT 659.740 600.450 660.000 600.770 ;
        RECT 938.500 600.450 938.760 600.770 ;
        RECT 941.720 600.710 943.610 600.770 ;
        RECT 941.720 600.450 941.980 600.710 ;
        RECT 938.560 29.570 938.700 600.450 ;
        RECT 943.330 600.000 943.610 600.710 ;
        RECT 531.860 29.250 532.120 29.570 ;
        RECT 938.500 29.250 938.760 29.570 ;
        RECT 531.920 2.400 532.060 29.250 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 1902.650 2877.280 1902.930 2877.560 ;
        RECT 350.610 1777.720 350.890 1778.000 ;
      LAYER met3 ;
        RECT 1885.335 2879.800 1889.335 2880.080 ;
        RECT 1885.335 2879.480 1889.370 2879.800 ;
        RECT 1889.070 2877.570 1889.370 2879.480 ;
        RECT 1902.625 2877.570 1902.955 2877.585 ;
        RECT 1889.070 2877.270 1902.955 2877.570 ;
        RECT 1902.625 2877.255 1902.955 2877.270 ;
        RECT 350.585 1778.010 350.915 1778.025 ;
        RECT 360.000 1778.010 364.000 1778.160 ;
        RECT 350.585 1777.710 364.000 1778.010 ;
        RECT 350.585 1777.695 350.915 1777.710 ;
        RECT 360.000 1777.560 364.000 1777.710 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 589.790 1688.000 590.110 1688.060 ;
        RECT 640.850 1688.000 641.170 1688.060 ;
        RECT 1486.330 1688.000 1486.650 1688.060 ;
        RECT 589.790 1687.860 1486.650 1688.000 ;
        RECT 589.790 1687.800 590.110 1687.860 ;
        RECT 640.850 1687.800 641.170 1687.860 ;
        RECT 1486.330 1687.800 1486.650 1687.860 ;
        RECT 638.090 586.740 638.410 586.800 ;
        RECT 640.850 586.740 641.170 586.800 ;
        RECT 952.730 586.740 953.050 586.800 ;
        RECT 638.090 586.600 664.540 586.740 ;
        RECT 638.090 586.540 638.410 586.600 ;
        RECT 640.850 586.540 641.170 586.600 ;
        RECT 664.400 586.060 664.540 586.600 ;
        RECT 668.080 586.600 953.050 586.740 ;
        RECT 668.080 586.060 668.220 586.600 ;
        RECT 952.730 586.540 953.050 586.600 ;
        RECT 664.400 585.920 668.220 586.060 ;
        RECT 549.770 36.620 550.090 36.680 ;
        RECT 638.090 36.620 638.410 36.680 ;
        RECT 549.770 36.480 638.410 36.620 ;
        RECT 549.770 36.420 550.090 36.480 ;
        RECT 638.090 36.420 638.410 36.480 ;
      LAYER via ;
        RECT 589.820 1687.800 590.080 1688.060 ;
        RECT 640.880 1687.800 641.140 1688.060 ;
        RECT 1486.360 1687.800 1486.620 1688.060 ;
        RECT 638.120 586.540 638.380 586.800 ;
        RECT 640.880 586.540 641.140 586.800 ;
        RECT 952.760 586.540 953.020 586.800 ;
        RECT 549.800 36.420 550.060 36.680 ;
        RECT 638.120 36.420 638.380 36.680 ;
      LAYER met2 ;
        RECT 1486.350 2705.195 1486.630 2705.565 ;
        RECT 588.250 1700.410 588.530 1704.000 ;
        RECT 588.250 1700.270 590.020 1700.410 ;
        RECT 588.250 1700.000 588.530 1700.270 ;
        RECT 589.880 1688.090 590.020 1700.270 ;
        RECT 1486.420 1688.090 1486.560 2705.195 ;
        RECT 589.820 1687.770 590.080 1688.090 ;
        RECT 640.880 1687.770 641.140 1688.090 ;
        RECT 1486.360 1687.770 1486.620 1688.090 ;
        RECT 640.940 586.830 641.080 1687.770 ;
        RECT 952.530 600.000 952.810 604.000 ;
        RECT 952.590 598.810 952.730 600.000 ;
        RECT 952.590 598.670 952.960 598.810 ;
        RECT 952.820 586.830 952.960 598.670 ;
        RECT 638.120 586.510 638.380 586.830 ;
        RECT 640.880 586.510 641.140 586.830 ;
        RECT 952.760 586.510 953.020 586.830 ;
        RECT 638.180 36.710 638.320 586.510 ;
        RECT 549.800 36.390 550.060 36.710 ;
        RECT 638.120 36.390 638.380 36.710 ;
        RECT 549.860 2.400 550.000 36.390 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 1486.350 2705.240 1486.630 2705.520 ;
      LAYER met3 ;
        RECT 1500.000 2708.440 1504.000 2708.720 ;
        RECT 1499.910 2708.120 1504.000 2708.440 ;
        RECT 1486.325 2705.530 1486.655 2705.545 ;
        RECT 1499.910 2705.530 1500.210 2708.120 ;
        RECT 1486.325 2705.230 1500.210 2705.530 ;
        RECT 1486.325 2705.215 1486.655 2705.230 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 962.390 2532.560 962.710 2532.620 ;
        RECT 1487.710 2532.560 1488.030 2532.620 ;
        RECT 962.390 2532.420 1488.030 2532.560 ;
        RECT 962.390 2532.360 962.710 2532.420 ;
        RECT 1487.710 2532.360 1488.030 2532.420 ;
        RECT 675.810 1714.520 676.130 1714.580 ;
        RECT 962.390 1714.520 962.710 1714.580 ;
        RECT 675.810 1714.380 962.710 1714.520 ;
        RECT 675.810 1714.320 676.130 1714.380 ;
        RECT 962.390 1714.320 962.710 1714.380 ;
        RECT 644.070 1712.480 644.390 1712.540 ;
        RECT 675.810 1712.480 676.130 1712.540 ;
        RECT 644.070 1712.340 676.130 1712.480 ;
        RECT 644.070 1712.280 644.390 1712.340 ;
        RECT 675.810 1712.280 676.130 1712.340 ;
        RECT 668.450 737.360 668.770 737.420 ;
        RECT 669.370 737.360 669.690 737.420 ;
        RECT 668.450 737.220 669.690 737.360 ;
        RECT 668.450 737.160 668.770 737.220 ;
        RECT 669.370 737.160 669.690 737.220 ;
        RECT 665.690 690.440 666.010 690.500 ;
        RECT 669.370 690.440 669.690 690.500 ;
        RECT 665.690 690.300 669.690 690.440 ;
        RECT 665.690 690.240 666.010 690.300 ;
        RECT 669.370 690.240 669.690 690.300 ;
        RECT 665.690 689.760 666.010 689.820 ;
        RECT 669.370 689.760 669.690 689.820 ;
        RECT 665.690 689.620 669.690 689.760 ;
        RECT 665.690 689.560 666.010 689.620 ;
        RECT 669.370 689.560 669.690 689.620 ;
        RECT 668.450 609.520 668.770 609.580 ;
        RECT 669.370 609.520 669.690 609.580 ;
        RECT 668.450 609.380 669.690 609.520 ;
        RECT 668.450 609.320 668.770 609.380 ;
        RECT 669.370 609.320 669.690 609.380 ;
        RECT 850.700 602.580 894.080 602.720 ;
        RECT 786.300 601.900 807.600 602.040 ;
        RECT 786.300 601.760 786.440 601.900 ;
        RECT 807.460 601.760 807.600 601.900 ;
        RECT 850.700 601.760 850.840 602.580 ;
        RECT 893.940 602.380 894.080 602.580 ;
        RECT 893.940 602.240 952.960 602.380 ;
        RECT 731.470 601.700 731.790 601.760 ;
        RECT 714.080 601.560 731.790 601.700 ;
        RECT 668.450 600.340 668.770 600.400 ;
        RECT 714.080 600.340 714.220 601.560 ;
        RECT 731.470 601.500 731.790 601.560 ;
        RECT 786.210 601.500 786.530 601.760 ;
        RECT 807.370 601.500 807.690 601.760 ;
        RECT 850.610 601.500 850.930 601.760 ;
        RECT 952.820 601.700 952.960 602.240 ;
        RECT 961.930 601.700 962.250 601.760 ;
        RECT 952.820 601.560 962.250 601.700 ;
        RECT 961.930 601.500 962.250 601.560 ;
        RECT 731.470 601.020 731.790 601.080 ;
        RECT 786.210 601.020 786.530 601.080 ;
        RECT 731.470 600.880 786.530 601.020 ;
        RECT 731.470 600.820 731.790 600.880 ;
        RECT 786.210 600.820 786.530 600.880 ;
        RECT 668.450 600.200 714.220 600.340 ;
        RECT 668.450 600.140 668.770 600.200 ;
        RECT 959.170 591.840 959.490 591.900 ;
        RECT 961.930 591.840 962.250 591.900 ;
        RECT 959.170 591.700 962.250 591.840 ;
        RECT 959.170 591.640 959.490 591.700 ;
        RECT 961.930 591.640 962.250 591.700 ;
        RECT 959.170 572.460 959.490 572.520 ;
        RECT 960.090 572.460 960.410 572.520 ;
        RECT 959.170 572.320 960.410 572.460 ;
        RECT 959.170 572.260 959.490 572.320 ;
        RECT 960.090 572.260 960.410 572.320 ;
        RECT 959.170 410.620 959.490 410.680 ;
        RECT 960.090 410.620 960.410 410.680 ;
        RECT 959.170 410.480 960.410 410.620 ;
        RECT 959.170 410.420 959.490 410.480 ;
        RECT 960.090 410.420 960.410 410.480 ;
        RECT 959.170 386.480 959.490 386.540 ;
        RECT 959.630 386.480 959.950 386.540 ;
        RECT 959.170 386.340 959.950 386.480 ;
        RECT 959.170 386.280 959.490 386.340 ;
        RECT 959.630 386.280 959.950 386.340 ;
        RECT 959.630 337.860 959.950 337.920 ;
        RECT 960.550 337.860 960.870 337.920 ;
        RECT 959.630 337.720 960.870 337.860 ;
        RECT 959.630 337.660 959.950 337.720 ;
        RECT 960.550 337.660 960.870 337.720 ;
        RECT 959.630 289.920 959.950 289.980 ;
        RECT 960.550 289.920 960.870 289.980 ;
        RECT 959.630 289.780 960.870 289.920 ;
        RECT 959.630 289.720 959.950 289.780 ;
        RECT 960.550 289.720 960.870 289.780 ;
        RECT 959.170 186.220 959.490 186.280 ;
        RECT 960.090 186.220 960.410 186.280 ;
        RECT 959.170 186.080 960.410 186.220 ;
        RECT 959.170 186.020 959.490 186.080 ;
        RECT 960.090 186.020 960.410 186.080 ;
        RECT 959.170 138.280 959.490 138.340 ;
        RECT 959.630 138.280 959.950 138.340 ;
        RECT 959.170 138.140 959.950 138.280 ;
        RECT 959.170 138.080 959.490 138.140 ;
        RECT 959.630 138.080 959.950 138.140 ;
        RECT 567.710 44.100 568.030 44.160 ;
        RECT 959.630 44.100 959.950 44.160 ;
        RECT 567.710 43.960 959.950 44.100 ;
        RECT 567.710 43.900 568.030 43.960 ;
        RECT 959.630 43.900 959.950 43.960 ;
      LAYER via ;
        RECT 962.420 2532.360 962.680 2532.620 ;
        RECT 1487.740 2532.360 1488.000 2532.620 ;
        RECT 675.840 1714.320 676.100 1714.580 ;
        RECT 962.420 1714.320 962.680 1714.580 ;
        RECT 644.100 1712.280 644.360 1712.540 ;
        RECT 675.840 1712.280 676.100 1712.540 ;
        RECT 668.480 737.160 668.740 737.420 ;
        RECT 669.400 737.160 669.660 737.420 ;
        RECT 665.720 690.240 665.980 690.500 ;
        RECT 669.400 690.240 669.660 690.500 ;
        RECT 665.720 689.560 665.980 689.820 ;
        RECT 669.400 689.560 669.660 689.820 ;
        RECT 668.480 609.320 668.740 609.580 ;
        RECT 669.400 609.320 669.660 609.580 ;
        RECT 668.480 600.140 668.740 600.400 ;
        RECT 731.500 601.500 731.760 601.760 ;
        RECT 786.240 601.500 786.500 601.760 ;
        RECT 807.400 601.500 807.660 601.760 ;
        RECT 850.640 601.500 850.900 601.760 ;
        RECT 961.960 601.500 962.220 601.760 ;
        RECT 731.500 600.820 731.760 601.080 ;
        RECT 786.240 600.820 786.500 601.080 ;
        RECT 959.200 591.640 959.460 591.900 ;
        RECT 961.960 591.640 962.220 591.900 ;
        RECT 959.200 572.260 959.460 572.520 ;
        RECT 960.120 572.260 960.380 572.520 ;
        RECT 959.200 410.420 959.460 410.680 ;
        RECT 960.120 410.420 960.380 410.680 ;
        RECT 959.200 386.280 959.460 386.540 ;
        RECT 959.660 386.280 959.920 386.540 ;
        RECT 959.660 337.660 959.920 337.920 ;
        RECT 960.580 337.660 960.840 337.920 ;
        RECT 959.660 289.720 959.920 289.980 ;
        RECT 960.580 289.720 960.840 289.980 ;
        RECT 959.200 186.020 959.460 186.280 ;
        RECT 960.120 186.020 960.380 186.280 ;
        RECT 959.200 138.080 959.460 138.340 ;
        RECT 959.660 138.080 959.920 138.340 ;
        RECT 567.740 43.900 568.000 44.160 ;
        RECT 959.660 43.900 959.920 44.160 ;
      LAYER met2 ;
        RECT 962.420 2532.330 962.680 2532.650 ;
        RECT 1487.730 2532.475 1488.010 2532.845 ;
        RECT 1487.740 2532.330 1488.000 2532.475 ;
        RECT 644.090 1717.835 644.370 1718.205 ;
        RECT 644.160 1712.570 644.300 1717.835 ;
        RECT 962.480 1714.610 962.620 2532.330 ;
        RECT 675.840 1714.290 676.100 1714.610 ;
        RECT 962.420 1714.290 962.680 1714.610 ;
        RECT 675.900 1712.570 676.040 1714.290 ;
        RECT 644.100 1712.250 644.360 1712.570 ;
        RECT 675.840 1712.250 676.100 1712.570 ;
        RECT 675.900 999.445 676.040 1712.250 ;
        RECT 675.830 999.075 676.110 999.445 ;
        RECT 668.470 787.595 668.750 787.965 ;
        RECT 668.540 737.450 668.680 787.595 ;
        RECT 668.480 737.130 668.740 737.450 ;
        RECT 669.400 737.130 669.660 737.450 ;
        RECT 669.460 690.530 669.600 737.130 ;
        RECT 665.720 690.210 665.980 690.530 ;
        RECT 669.400 690.210 669.660 690.530 ;
        RECT 665.780 689.850 665.920 690.210 ;
        RECT 665.720 689.530 665.980 689.850 ;
        RECT 669.400 689.530 669.660 689.850 ;
        RECT 669.460 609.610 669.600 689.530 ;
        RECT 668.480 609.290 668.740 609.610 ;
        RECT 669.400 609.290 669.660 609.610 ;
        RECT 668.540 600.430 668.680 609.290 ;
        RECT 731.500 601.470 731.760 601.790 ;
        RECT 786.240 601.470 786.500 601.790 ;
        RECT 807.400 601.645 807.660 601.790 ;
        RECT 850.640 601.645 850.900 601.790 ;
        RECT 731.560 601.110 731.700 601.470 ;
        RECT 786.300 601.110 786.440 601.470 ;
        RECT 807.390 601.275 807.670 601.645 ;
        RECT 850.630 601.275 850.910 601.645 ;
        RECT 961.270 601.530 961.550 604.000 ;
        RECT 962.020 601.790 962.160 601.945 ;
        RECT 961.960 601.530 962.220 601.790 ;
        RECT 961.270 601.470 962.220 601.530 ;
        RECT 961.270 601.390 962.160 601.470 ;
        RECT 731.500 600.790 731.760 601.110 ;
        RECT 786.240 600.790 786.500 601.110 ;
        RECT 668.480 600.110 668.740 600.430 ;
        RECT 961.270 600.000 961.550 601.390 ;
        RECT 962.020 591.930 962.160 601.390 ;
        RECT 959.200 591.610 959.460 591.930 ;
        RECT 961.960 591.610 962.220 591.930 ;
        RECT 959.260 572.550 959.400 591.610 ;
        RECT 959.200 572.230 959.460 572.550 ;
        RECT 960.120 572.230 960.380 572.550 ;
        RECT 960.180 410.710 960.320 572.230 ;
        RECT 959.200 410.390 959.460 410.710 ;
        RECT 960.120 410.390 960.380 410.710 ;
        RECT 959.260 386.570 959.400 410.390 ;
        RECT 959.200 386.250 959.460 386.570 ;
        RECT 959.660 386.250 959.920 386.570 ;
        RECT 959.720 337.950 959.860 386.250 ;
        RECT 959.660 337.630 959.920 337.950 ;
        RECT 960.580 337.630 960.840 337.950 ;
        RECT 960.640 290.010 960.780 337.630 ;
        RECT 959.660 289.690 959.920 290.010 ;
        RECT 960.580 289.690 960.840 290.010 ;
        RECT 959.720 265.610 959.860 289.690 ;
        RECT 959.720 265.470 960.780 265.610 ;
        RECT 960.640 241.810 960.780 265.470 ;
        RECT 960.180 241.670 960.780 241.810 ;
        RECT 960.180 186.310 960.320 241.670 ;
        RECT 959.200 185.990 959.460 186.310 ;
        RECT 960.120 185.990 960.380 186.310 ;
        RECT 959.260 138.370 959.400 185.990 ;
        RECT 959.200 138.050 959.460 138.370 ;
        RECT 959.660 138.050 959.920 138.370 ;
        RECT 959.720 44.190 959.860 138.050 ;
        RECT 567.740 43.870 568.000 44.190 ;
        RECT 959.660 43.870 959.920 44.190 ;
        RECT 567.800 2.400 567.940 43.870 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1487.730 2532.520 1488.010 2532.800 ;
        RECT 644.090 1717.880 644.370 1718.160 ;
        RECT 675.830 999.120 676.110 999.400 ;
        RECT 668.470 787.640 668.750 787.920 ;
        RECT 807.390 601.320 807.670 601.600 ;
        RECT 850.630 601.320 850.910 601.600 ;
      LAYER met3 ;
        RECT 1500.000 2535.720 1504.000 2536.000 ;
        RECT 1499.910 2535.400 1504.000 2535.720 ;
        RECT 1487.705 2532.810 1488.035 2532.825 ;
        RECT 1499.910 2532.810 1500.210 2535.400 ;
        RECT 1487.705 2532.510 1500.210 2532.810 ;
        RECT 1487.705 2532.495 1488.035 2532.510 ;
        RECT 627.030 1718.170 631.030 1718.320 ;
        RECT 644.065 1718.170 644.395 1718.185 ;
        RECT 627.030 1717.870 644.395 1718.170 ;
        RECT 627.030 1717.720 631.030 1717.870 ;
        RECT 644.065 1717.855 644.395 1717.870 ;
        RECT 669.110 999.410 669.490 999.420 ;
        RECT 675.805 999.410 676.135 999.425 ;
        RECT 669.110 999.110 676.135 999.410 ;
        RECT 669.110 999.100 669.490 999.110 ;
        RECT 675.805 999.095 676.135 999.110 ;
        RECT 668.445 787.930 668.775 787.945 ;
        RECT 669.110 787.930 669.490 787.940 ;
        RECT 668.445 787.630 669.490 787.930 ;
        RECT 668.445 787.615 668.775 787.630 ;
        RECT 669.110 787.620 669.490 787.630 ;
        RECT 807.365 601.610 807.695 601.625 ;
        RECT 850.605 601.610 850.935 601.625 ;
        RECT 807.365 601.310 850.935 601.610 ;
        RECT 807.365 601.295 807.695 601.310 ;
        RECT 850.605 601.295 850.935 601.310 ;
      LAYER via3 ;
        RECT 669.140 999.100 669.460 999.420 ;
        RECT 669.140 787.620 669.460 787.940 ;
      LAYER met4 ;
        RECT 669.135 999.095 669.465 999.425 ;
        RECT 669.150 787.945 669.450 999.095 ;
        RECT 669.135 787.615 669.465 787.945 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 438.910 1686.980 439.230 1687.040 ;
        RECT 586.110 1686.980 586.430 1687.040 ;
        RECT 1902.170 1686.980 1902.490 1687.040 ;
        RECT 438.910 1686.840 1902.490 1686.980 ;
        RECT 438.910 1686.780 439.230 1686.840 ;
        RECT 586.110 1686.780 586.430 1686.840 ;
        RECT 1902.170 1686.780 1902.490 1686.840 ;
        RECT 579.670 15.880 579.990 15.940 ;
        RECT 585.650 15.880 585.970 15.940 ;
        RECT 579.670 15.740 585.970 15.880 ;
        RECT 579.670 15.680 579.990 15.740 ;
        RECT 585.650 15.680 585.970 15.740 ;
      LAYER via ;
        RECT 438.940 1686.780 439.200 1687.040 ;
        RECT 586.140 1686.780 586.400 1687.040 ;
        RECT 1902.200 1686.780 1902.460 1687.040 ;
        RECT 579.700 15.680 579.960 15.940 ;
        RECT 585.680 15.680 585.940 15.940 ;
      LAYER met2 ;
        RECT 1902.190 2643.315 1902.470 2643.685 ;
        RECT 437.370 1700.410 437.650 1704.000 ;
        RECT 437.370 1700.270 439.140 1700.410 ;
        RECT 437.370 1700.000 437.650 1700.270 ;
        RECT 439.000 1687.070 439.140 1700.270 ;
        RECT 1902.260 1687.070 1902.400 2643.315 ;
        RECT 438.940 1686.750 439.200 1687.070 ;
        RECT 586.140 1686.750 586.400 1687.070 ;
        RECT 1902.200 1686.750 1902.460 1687.070 ;
        RECT 586.200 592.805 586.340 1686.750 ;
        RECT 970.470 600.170 970.750 604.000 ;
        RECT 968.920 600.030 970.750 600.170 ;
        RECT 968.920 592.805 969.060 600.030 ;
        RECT 970.470 600.000 970.750 600.030 ;
        RECT 586.130 592.435 586.410 592.805 ;
        RECT 968.850 592.435 969.130 592.805 ;
        RECT 586.200 586.685 586.340 592.435 ;
        RECT 579.690 586.315 579.970 586.685 ;
        RECT 586.130 586.315 586.410 586.685 ;
        RECT 579.760 15.970 579.900 586.315 ;
        RECT 579.700 15.650 579.960 15.970 ;
        RECT 585.680 15.650 585.940 15.970 ;
        RECT 585.740 2.400 585.880 15.650 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 1902.190 2643.360 1902.470 2643.640 ;
        RECT 586.130 592.480 586.410 592.760 ;
        RECT 968.850 592.480 969.130 592.760 ;
        RECT 579.690 586.360 579.970 586.640 ;
        RECT 586.130 586.360 586.410 586.640 ;
      LAYER met3 ;
        RECT 1885.335 2644.520 1889.335 2644.800 ;
        RECT 1885.335 2644.200 1889.370 2644.520 ;
        RECT 1889.070 2643.650 1889.370 2644.200 ;
        RECT 1902.165 2643.650 1902.495 2643.665 ;
        RECT 1889.070 2643.350 1902.495 2643.650 ;
        RECT 1902.165 2643.335 1902.495 2643.350 ;
        RECT 586.105 592.770 586.435 592.785 ;
        RECT 968.825 592.770 969.155 592.785 ;
        RECT 586.105 592.470 969.155 592.770 ;
        RECT 586.105 592.455 586.435 592.470 ;
        RECT 968.825 592.455 969.155 592.470 ;
        RECT 579.665 586.650 579.995 586.665 ;
        RECT 586.105 586.650 586.435 586.665 ;
        RECT 579.665 586.350 586.435 586.650 ;
        RECT 579.665 586.335 579.995 586.350 ;
        RECT 586.105 586.335 586.435 586.350 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1438.490 2666.860 1438.810 2666.920 ;
        RECT 1487.710 2666.860 1488.030 2666.920 ;
        RECT 1438.490 2666.720 1488.030 2666.860 ;
        RECT 1438.490 2666.660 1438.810 2666.720 ;
        RECT 1487.710 2666.660 1488.030 2666.720 ;
        RECT 426.950 2606.340 427.270 2606.400 ;
        RECT 1435.270 2606.340 1435.590 2606.400 ;
        RECT 1438.490 2606.340 1438.810 2606.400 ;
        RECT 426.950 2606.200 1438.810 2606.340 ;
        RECT 426.950 2606.140 427.270 2606.200 ;
        RECT 1435.270 2606.140 1435.590 2606.200 ;
        RECT 1438.490 2606.140 1438.810 2606.200 ;
        RECT 989.070 2032.760 989.390 2032.820 ;
        RECT 1435.270 2032.760 1435.590 2032.820 ;
        RECT 1438.490 2032.760 1438.810 2032.820 ;
        RECT 989.070 2032.620 1438.810 2032.760 ;
        RECT 989.070 2032.560 989.390 2032.620 ;
        RECT 1435.270 2032.560 1435.590 2032.620 ;
        RECT 1438.490 2032.560 1438.810 2032.620 ;
        RECT 1438.490 1928.380 1438.810 1928.440 ;
        RECT 1941.270 1928.380 1941.590 1928.440 ;
        RECT 1438.490 1928.240 1941.590 1928.380 ;
        RECT 1438.490 1928.180 1438.810 1928.240 ;
        RECT 1941.270 1928.180 1941.590 1928.240 ;
        RECT 644.530 1828.760 644.850 1828.820 ;
        RECT 644.530 1828.620 648.900 1828.760 ;
        RECT 644.530 1828.560 644.850 1828.620 ;
        RECT 648.760 1828.420 648.900 1828.620 ;
        RECT 652.350 1828.420 652.670 1828.480 ;
        RECT 989.070 1828.420 989.390 1828.480 ;
        RECT 648.760 1828.280 989.390 1828.420 ;
        RECT 652.350 1828.220 652.670 1828.280 ;
        RECT 989.070 1828.220 989.390 1828.280 ;
        RECT 652.350 587.760 652.670 587.820 ;
        RECT 677.190 587.760 677.510 587.820 ;
        RECT 713.530 587.760 713.850 587.820 ;
        RECT 652.350 587.620 713.850 587.760 ;
        RECT 652.350 587.560 652.670 587.620 ;
        RECT 677.190 587.560 677.510 587.620 ;
        RECT 713.530 587.560 713.850 587.620 ;
        RECT 91.610 31.180 91.930 31.240 ;
        RECT 677.190 31.180 677.510 31.240 ;
        RECT 91.610 31.040 677.510 31.180 ;
        RECT 91.610 30.980 91.930 31.040 ;
        RECT 677.190 30.980 677.510 31.040 ;
      LAYER via ;
        RECT 1438.520 2666.660 1438.780 2666.920 ;
        RECT 1487.740 2666.660 1488.000 2666.920 ;
        RECT 426.980 2606.140 427.240 2606.400 ;
        RECT 1435.300 2606.140 1435.560 2606.400 ;
        RECT 1438.520 2606.140 1438.780 2606.400 ;
        RECT 989.100 2032.560 989.360 2032.820 ;
        RECT 1435.300 2032.560 1435.560 2032.820 ;
        RECT 1438.520 2032.560 1438.780 2032.820 ;
        RECT 1438.520 1928.180 1438.780 1928.440 ;
        RECT 1941.300 1928.180 1941.560 1928.440 ;
        RECT 644.560 1828.560 644.820 1828.820 ;
        RECT 652.380 1828.220 652.640 1828.480 ;
        RECT 989.100 1828.220 989.360 1828.480 ;
        RECT 652.380 587.560 652.640 587.820 ;
        RECT 677.220 587.560 677.480 587.820 ;
        RECT 713.560 587.560 713.820 587.820 ;
        RECT 91.640 30.980 91.900 31.240 ;
        RECT 677.220 30.980 677.480 31.240 ;
      LAYER met2 ;
        RECT 1487.730 2864.315 1488.010 2864.685 ;
        RECT 1487.800 2666.950 1487.940 2864.315 ;
        RECT 1438.520 2666.630 1438.780 2666.950 ;
        RECT 1487.740 2666.630 1488.000 2666.950 ;
        RECT 426.970 2665.075 427.250 2665.445 ;
        RECT 427.040 2606.430 427.180 2665.075 ;
        RECT 1438.580 2606.430 1438.720 2666.630 ;
        RECT 426.980 2606.110 427.240 2606.430 ;
        RECT 1435.300 2606.110 1435.560 2606.430 ;
        RECT 1438.520 2606.110 1438.780 2606.430 ;
        RECT 1435.360 2032.850 1435.500 2606.110 ;
        RECT 989.100 2032.530 989.360 2032.850 ;
        RECT 1435.300 2032.530 1435.560 2032.850 ;
        RECT 1438.520 2032.530 1438.780 2032.850 ;
        RECT 644.550 1829.355 644.830 1829.725 ;
        RECT 644.620 1828.850 644.760 1829.355 ;
        RECT 644.560 1828.530 644.820 1828.850 ;
        RECT 989.160 1828.510 989.300 2032.530 ;
        RECT 1438.580 1928.470 1438.720 2032.530 ;
        RECT 1438.520 1928.150 1438.780 1928.470 ;
        RECT 1941.300 1928.150 1941.560 1928.470 ;
        RECT 1941.360 1917.095 1941.500 1928.150 ;
        RECT 1941.250 1913.095 1941.530 1917.095 ;
        RECT 652.380 1828.190 652.640 1828.510 ;
        RECT 989.100 1828.190 989.360 1828.510 ;
        RECT 652.440 587.850 652.580 1828.190 ;
        RECT 717.010 600.170 717.290 604.000 ;
        RECT 715.460 600.030 717.290 600.170 ;
        RECT 715.460 590.650 715.600 600.030 ;
        RECT 717.010 600.000 717.290 600.030 ;
        RECT 713.620 590.510 715.600 590.650 ;
        RECT 713.620 587.850 713.760 590.510 ;
        RECT 652.380 587.530 652.640 587.850 ;
        RECT 677.220 587.530 677.480 587.850 ;
        RECT 713.560 587.530 713.820 587.850 ;
        RECT 677.280 31.270 677.420 587.530 ;
        RECT 91.640 30.950 91.900 31.270 ;
        RECT 677.220 30.950 677.480 31.270 ;
        RECT 91.700 2.400 91.840 30.950 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 1487.730 2864.360 1488.010 2864.640 ;
        RECT 426.970 2665.120 427.250 2665.400 ;
        RECT 644.550 1829.400 644.830 1829.680 ;
      LAYER met3 ;
        RECT 1500.000 2864.840 1504.000 2865.120 ;
        RECT 1487.705 2864.650 1488.035 2864.665 ;
        RECT 1499.910 2864.650 1504.000 2864.840 ;
        RECT 1487.705 2864.520 1504.000 2864.650 ;
        RECT 1487.705 2864.350 1500.210 2864.520 ;
        RECT 1487.705 2864.335 1488.035 2864.350 ;
        RECT 430.000 2668.320 434.000 2668.640 ;
        RECT 429.950 2668.040 434.000 2668.320 ;
        RECT 426.945 2665.410 427.275 2665.425 ;
        RECT 429.950 2665.410 430.250 2668.040 ;
        RECT 426.945 2665.110 430.250 2665.410 ;
        RECT 426.945 2665.095 427.275 2665.110 ;
        RECT 627.030 1829.690 631.030 1829.840 ;
        RECT 644.525 1829.690 644.855 1829.705 ;
        RECT 627.030 1829.390 644.855 1829.690 ;
        RECT 627.030 1829.240 631.030 1829.390 ;
        RECT 644.525 1829.375 644.855 1829.390 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 631.190 2918.120 631.510 2918.180 ;
        RECT 1513.930 2918.120 1514.250 2918.180 ;
        RECT 631.190 2917.980 1514.250 2918.120 ;
        RECT 631.190 2917.920 631.510 2917.980 ;
        RECT 1513.930 2917.920 1514.250 2917.980 ;
        RECT 479.390 1988.220 479.710 1988.280 ;
        RECT 631.190 1988.220 631.510 1988.280 ;
        RECT 479.390 1988.080 631.510 1988.220 ;
        RECT 479.390 1988.020 479.710 1988.080 ;
        RECT 631.190 1988.020 631.510 1988.080 ;
        RECT 603.130 43.080 603.450 43.140 ;
        RECT 631.190 43.080 631.510 43.140 ;
        RECT 603.130 42.940 631.510 43.080 ;
        RECT 603.130 42.880 603.450 42.940 ;
        RECT 631.190 42.880 631.510 42.940 ;
      LAYER via ;
        RECT 631.220 2917.920 631.480 2918.180 ;
        RECT 1513.960 2917.920 1514.220 2918.180 ;
        RECT 479.420 1988.020 479.680 1988.280 ;
        RECT 631.220 1988.020 631.480 1988.280 ;
        RECT 603.160 42.880 603.420 43.140 ;
        RECT 631.220 42.880 631.480 43.140 ;
      LAYER met2 ;
        RECT 631.220 2917.890 631.480 2918.210 ;
        RECT 1513.960 2917.890 1514.220 2918.210 ;
        RECT 631.280 1988.310 631.420 2917.890 ;
        RECT 1514.020 2900.055 1514.160 2917.890 ;
        RECT 1513.890 2896.055 1514.170 2900.055 ;
        RECT 479.420 1987.990 479.680 1988.310 ;
        RECT 631.220 1987.990 631.480 1988.310 ;
        RECT 477.850 1981.250 478.130 1981.750 ;
        RECT 479.480 1981.250 479.620 1987.990 ;
        RECT 477.850 1981.110 479.620 1981.250 ;
        RECT 477.850 1977.750 478.130 1981.110 ;
        RECT 631.280 591.445 631.420 1987.990 ;
        RECT 979.670 600.000 979.950 604.000 ;
        RECT 979.730 598.810 979.870 600.000 ;
        RECT 979.730 598.670 980.100 598.810 ;
        RECT 979.960 591.445 980.100 598.670 ;
        RECT 631.210 591.075 631.490 591.445 ;
        RECT 979.890 591.075 980.170 591.445 ;
        RECT 631.280 43.170 631.420 591.075 ;
        RECT 603.160 42.850 603.420 43.170 ;
        RECT 631.220 42.850 631.480 43.170 ;
        RECT 603.220 2.400 603.360 42.850 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 631.210 591.120 631.490 591.400 ;
        RECT 979.890 591.120 980.170 591.400 ;
      LAYER met3 ;
        RECT 631.185 591.410 631.515 591.425 ;
        RECT 979.865 591.410 980.195 591.425 ;
        RECT 631.185 591.110 980.195 591.410 ;
        RECT 631.185 591.095 631.515 591.110 ;
        RECT 979.865 591.095 980.195 591.110 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 624.290 2916.420 624.610 2916.480 ;
        RECT 1620.650 2916.420 1620.970 2916.480 ;
        RECT 624.290 2916.280 1620.970 2916.420 ;
        RECT 624.290 2916.220 624.610 2916.280 ;
        RECT 1620.650 2916.220 1620.970 2916.280 ;
        RECT 403.950 1988.900 404.270 1988.960 ;
        RECT 620.610 1988.900 620.930 1988.960 ;
        RECT 403.950 1988.760 620.930 1988.900 ;
        RECT 403.950 1988.700 404.270 1988.760 ;
        RECT 620.610 1988.700 620.930 1988.760 ;
        RECT 620.610 1987.200 620.930 1987.260 ;
        RECT 624.290 1987.200 624.610 1987.260 ;
        RECT 628.890 1987.200 629.210 1987.260 ;
        RECT 620.610 1987.060 629.210 1987.200 ;
        RECT 620.610 1987.000 620.930 1987.060 ;
        RECT 624.290 1987.000 624.610 1987.060 ;
        RECT 628.890 1987.000 629.210 1987.060 ;
        RECT 621.070 15.540 621.390 15.600 ;
        RECT 627.510 15.540 627.830 15.600 ;
        RECT 621.070 15.400 627.830 15.540 ;
        RECT 621.070 15.340 621.390 15.400 ;
        RECT 627.510 15.340 627.830 15.400 ;
      LAYER via ;
        RECT 624.320 2916.220 624.580 2916.480 ;
        RECT 1620.680 2916.220 1620.940 2916.480 ;
        RECT 403.980 1988.700 404.240 1988.960 ;
        RECT 620.640 1988.700 620.900 1988.960 ;
        RECT 620.640 1987.000 620.900 1987.260 ;
        RECT 624.320 1987.000 624.580 1987.260 ;
        RECT 628.920 1987.000 629.180 1987.260 ;
        RECT 621.100 15.340 621.360 15.600 ;
        RECT 627.540 15.340 627.800 15.600 ;
      LAYER met2 ;
        RECT 624.320 2916.190 624.580 2916.510 ;
        RECT 1620.680 2916.190 1620.940 2916.510 ;
        RECT 403.980 1988.670 404.240 1988.990 ;
        RECT 620.640 1988.670 620.900 1988.990 ;
        RECT 402.410 1981.250 402.690 1981.750 ;
        RECT 404.040 1981.250 404.180 1988.670 ;
        RECT 620.700 1987.290 620.840 1988.670 ;
        RECT 624.380 1987.290 624.520 2916.190 ;
        RECT 1620.740 2900.055 1620.880 2916.190 ;
        RECT 1620.610 2896.055 1620.890 2900.055 ;
        RECT 620.640 1986.970 620.900 1987.290 ;
        RECT 624.320 1986.970 624.580 1987.290 ;
        RECT 628.920 1986.970 629.180 1987.290 ;
        RECT 402.410 1981.110 404.180 1981.250 ;
        RECT 402.410 1977.750 402.690 1981.110 ;
        RECT 628.980 592.125 629.120 1986.970 ;
        RECT 988.870 600.170 989.150 604.000 ;
        RECT 987.320 600.030 989.150 600.170 ;
        RECT 987.320 592.125 987.460 600.030 ;
        RECT 988.870 600.000 989.150 600.030 ;
        RECT 628.910 591.755 629.190 592.125 ;
        RECT 987.250 591.755 987.530 592.125 ;
        RECT 628.980 586.570 629.120 591.755 ;
        RECT 627.600 586.430 629.120 586.570 ;
        RECT 627.600 15.630 627.740 586.430 ;
        RECT 621.100 15.310 621.360 15.630 ;
        RECT 627.540 15.310 627.800 15.630 ;
        RECT 621.160 2.400 621.300 15.310 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 628.910 591.800 629.190 592.080 ;
        RECT 987.250 591.800 987.530 592.080 ;
      LAYER met3 ;
        RECT 628.885 592.090 629.215 592.105 ;
        RECT 987.225 592.090 987.555 592.105 ;
        RECT 628.885 591.790 987.555 592.090 ;
        RECT 628.885 591.775 629.215 591.790 ;
        RECT 987.225 591.775 987.555 591.790 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 2877.660 551.930 2877.720 ;
        RECT 1483.570 2877.660 1483.890 2877.720 ;
        RECT 551.610 2877.520 1483.890 2877.660 ;
        RECT 551.610 2877.460 551.930 2877.520 ;
        RECT 1483.570 2877.460 1483.890 2877.520 ;
        RECT 547.010 2773.960 547.330 2774.020 ;
        RECT 551.610 2773.960 551.930 2774.020 ;
        RECT 579.670 2773.960 579.990 2774.020 ;
        RECT 547.010 2773.820 579.990 2773.960 ;
        RECT 547.010 2773.760 547.330 2773.820 ;
        RECT 551.610 2773.760 551.930 2773.820 ;
        RECT 579.670 2773.760 579.990 2773.820 ;
        RECT 379.110 1990.600 379.430 1990.660 ;
        RECT 579.670 1990.600 579.990 1990.660 ;
        RECT 636.250 1990.600 636.570 1990.660 ;
        RECT 379.110 1990.460 636.570 1990.600 ;
        RECT 379.110 1990.400 379.430 1990.460 ;
        RECT 579.670 1990.400 579.990 1990.460 ;
        RECT 636.250 1990.400 636.570 1990.460 ;
        RECT 636.250 1703.980 636.570 1704.040 ;
        RECT 2021.770 1703.980 2022.090 1704.040 ;
        RECT 636.250 1703.840 2022.090 1703.980 ;
        RECT 636.250 1703.780 636.570 1703.840 ;
        RECT 2021.770 1703.780 2022.090 1703.840 ;
        RECT 551.610 1700.920 551.930 1700.980 ;
        RECT 636.250 1700.920 636.570 1700.980 ;
        RECT 551.610 1700.780 636.570 1700.920 ;
        RECT 551.610 1700.720 551.930 1700.780 ;
        RECT 636.250 1700.720 636.570 1700.780 ;
        RECT 551.610 591.840 551.930 591.900 ;
        RECT 727.790 591.840 728.110 591.900 ;
        RECT 551.610 591.700 728.110 591.840 ;
        RECT 551.610 591.640 551.930 591.700 ;
        RECT 727.790 591.640 728.110 591.700 ;
        RECT 116.910 590.480 117.230 590.540 ;
        RECT 551.610 590.480 551.930 590.540 ;
        RECT 116.910 590.340 551.930 590.480 ;
        RECT 116.910 590.280 117.230 590.340 ;
        RECT 551.610 590.280 551.930 590.340 ;
      LAYER via ;
        RECT 551.640 2877.460 551.900 2877.720 ;
        RECT 1483.600 2877.460 1483.860 2877.720 ;
        RECT 547.040 2773.760 547.300 2774.020 ;
        RECT 551.640 2773.760 551.900 2774.020 ;
        RECT 579.700 2773.760 579.960 2774.020 ;
        RECT 379.140 1990.400 379.400 1990.660 ;
        RECT 579.700 1990.400 579.960 1990.660 ;
        RECT 636.280 1990.400 636.540 1990.660 ;
        RECT 636.280 1703.780 636.540 1704.040 ;
        RECT 2021.800 1703.780 2022.060 1704.040 ;
        RECT 551.640 1700.720 551.900 1700.980 ;
        RECT 636.280 1700.720 636.540 1700.980 ;
        RECT 551.640 591.640 551.900 591.900 ;
        RECT 727.820 591.640 728.080 591.900 ;
        RECT 116.940 590.280 117.200 590.540 ;
        RECT 551.640 590.280 551.900 590.540 ;
      LAYER met2 ;
        RECT 1483.590 2878.595 1483.870 2878.965 ;
        RECT 1483.660 2877.750 1483.800 2878.595 ;
        RECT 551.640 2877.430 551.900 2877.750 ;
        RECT 1483.600 2877.430 1483.860 2877.750 ;
        RECT 551.700 2774.050 551.840 2877.430 ;
        RECT 547.040 2773.730 547.300 2774.050 ;
        RECT 551.640 2773.730 551.900 2774.050 ;
        RECT 579.700 2773.730 579.960 2774.050 ;
        RECT 547.100 2759.520 547.240 2773.730 ;
        RECT 546.930 2759.100 547.240 2759.520 ;
        RECT 546.930 2755.520 547.210 2759.100 ;
        RECT 579.760 1990.690 579.900 2773.730 ;
        RECT 379.140 1990.370 379.400 1990.690 ;
        RECT 579.700 1990.370 579.960 1990.690 ;
        RECT 636.280 1990.370 636.540 1990.690 ;
        RECT 377.570 1981.250 377.850 1981.750 ;
        RECT 379.200 1981.250 379.340 1990.370 ;
        RECT 377.570 1981.110 379.340 1981.250 ;
        RECT 377.570 1977.750 377.850 1981.110 ;
        RECT 636.340 1704.070 636.480 1990.370 ;
        RECT 2025.890 1750.730 2026.170 1754.000 ;
        RECT 2021.860 1750.590 2026.170 1750.730 ;
        RECT 2021.860 1704.070 2022.000 1750.590 ;
        RECT 2025.890 1750.000 2026.170 1750.590 ;
        RECT 636.280 1703.750 636.540 1704.070 ;
        RECT 2021.800 1703.750 2022.060 1704.070 ;
        RECT 636.340 1701.010 636.480 1703.750 ;
        RECT 551.640 1700.690 551.900 1701.010 ;
        RECT 636.280 1700.690 636.540 1701.010 ;
        RECT 551.700 591.930 551.840 1700.690 ;
        RECT 729.430 600.170 729.710 604.000 ;
        RECT 727.880 600.030 729.710 600.170 ;
        RECT 727.880 591.930 728.020 600.030 ;
        RECT 729.430 600.000 729.710 600.030 ;
        RECT 551.640 591.610 551.900 591.930 ;
        RECT 727.820 591.610 728.080 591.930 ;
        RECT 551.700 590.570 551.840 591.610 ;
        RECT 116.940 590.250 117.200 590.570 ;
        RECT 551.640 590.250 551.900 590.570 ;
        RECT 117.000 17.410 117.140 590.250 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 1483.590 2878.640 1483.870 2878.920 ;
      LAYER met3 ;
        RECT 1500.000 2881.160 1504.000 2881.440 ;
        RECT 1499.910 2880.840 1504.000 2881.160 ;
        RECT 1483.565 2878.930 1483.895 2878.945 ;
        RECT 1499.910 2878.930 1500.210 2880.840 ;
        RECT 1483.565 2878.630 1500.210 2878.930 ;
        RECT 1483.565 2878.615 1483.895 2878.630 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 460.530 2769.880 460.850 2769.940 ;
        RECT 576.450 2769.880 576.770 2769.940 ;
        RECT 460.530 2769.740 576.770 2769.880 ;
        RECT 460.530 2769.680 460.850 2769.740 ;
        RECT 576.450 2769.680 576.770 2769.740 ;
        RECT 558.510 2489.380 558.830 2489.440 ;
        RECT 576.450 2489.380 576.770 2489.440 ;
        RECT 1566.370 2489.380 1566.690 2489.440 ;
        RECT 558.510 2489.240 1566.690 2489.380 ;
        RECT 558.510 2489.180 558.830 2489.240 ;
        RECT 576.450 2489.180 576.770 2489.240 ;
        RECT 1566.370 2489.180 1566.690 2489.240 ;
        RECT 554.830 1994.340 555.150 1994.400 ;
        RECT 558.510 1994.340 558.830 1994.400 ;
        RECT 630.270 1994.340 630.590 1994.400 ;
        RECT 554.830 1994.200 630.590 1994.340 ;
        RECT 554.830 1994.140 555.150 1994.200 ;
        RECT 558.510 1994.140 558.830 1994.200 ;
        RECT 630.270 1994.140 630.590 1994.200 ;
        RECT 630.270 1704.320 630.590 1704.380 ;
        RECT 2042.470 1704.320 2042.790 1704.380 ;
        RECT 630.270 1704.180 2042.790 1704.320 ;
        RECT 630.270 1704.120 630.590 1704.180 ;
        RECT 2042.470 1704.120 2042.790 1704.180 ;
        RECT 572.310 1701.260 572.630 1701.320 ;
        RECT 630.270 1701.260 630.590 1701.320 ;
        RECT 572.310 1701.120 630.590 1701.260 ;
        RECT 572.310 1701.060 572.630 1701.120 ;
        RECT 630.270 1701.060 630.590 1701.120 ;
        RECT 144.510 590.820 144.830 590.880 ;
        RECT 572.310 590.820 572.630 590.880 ;
        RECT 739.750 590.820 740.070 590.880 ;
        RECT 144.510 590.680 740.070 590.820 ;
        RECT 144.510 590.620 144.830 590.680 ;
        RECT 572.310 590.620 572.630 590.680 ;
        RECT 739.750 590.620 740.070 590.680 ;
        RECT 139.450 16.900 139.770 16.960 ;
        RECT 144.510 16.900 144.830 16.960 ;
        RECT 139.450 16.760 144.830 16.900 ;
        RECT 139.450 16.700 139.770 16.760 ;
        RECT 144.510 16.700 144.830 16.760 ;
      LAYER via ;
        RECT 460.560 2769.680 460.820 2769.940 ;
        RECT 576.480 2769.680 576.740 2769.940 ;
        RECT 558.540 2489.180 558.800 2489.440 ;
        RECT 576.480 2489.180 576.740 2489.440 ;
        RECT 1566.400 2489.180 1566.660 2489.440 ;
        RECT 554.860 1994.140 555.120 1994.400 ;
        RECT 558.540 1994.140 558.800 1994.400 ;
        RECT 630.300 1994.140 630.560 1994.400 ;
        RECT 630.300 1704.120 630.560 1704.380 ;
        RECT 2042.500 1704.120 2042.760 1704.380 ;
        RECT 572.340 1701.060 572.600 1701.320 ;
        RECT 630.300 1701.060 630.560 1701.320 ;
        RECT 144.540 590.620 144.800 590.880 ;
        RECT 572.340 590.620 572.600 590.880 ;
        RECT 739.780 590.620 740.040 590.880 ;
        RECT 139.480 16.700 139.740 16.960 ;
        RECT 144.540 16.700 144.800 16.960 ;
      LAYER met2 ;
        RECT 460.560 2769.650 460.820 2769.970 ;
        RECT 576.480 2769.650 576.740 2769.970 ;
        RECT 460.620 2759.520 460.760 2769.650 ;
        RECT 460.450 2759.100 460.760 2759.520 ;
        RECT 460.450 2755.520 460.730 2759.100 ;
        RECT 576.540 2489.470 576.680 2769.650 ;
        RECT 1566.330 2500.000 1566.610 2504.000 ;
        RECT 1566.460 2489.470 1566.600 2500.000 ;
        RECT 558.540 2489.150 558.800 2489.470 ;
        RECT 576.480 2489.150 576.740 2489.470 ;
        RECT 1566.400 2489.150 1566.660 2489.470 ;
        RECT 558.600 1994.430 558.740 2489.150 ;
        RECT 554.860 1994.110 555.120 1994.430 ;
        RECT 558.540 1994.110 558.800 1994.430 ;
        RECT 630.300 1994.110 630.560 1994.430 ;
        RECT 553.290 1981.250 553.570 1981.750 ;
        RECT 554.920 1981.250 555.060 1994.110 ;
        RECT 553.290 1981.110 555.060 1981.250 ;
        RECT 553.290 1977.750 553.570 1981.110 ;
        RECT 630.360 1704.410 630.500 1994.110 ;
        RECT 2048.890 1750.730 2049.170 1754.000 ;
        RECT 2042.560 1750.590 2049.170 1750.730 ;
        RECT 2042.560 1704.410 2042.700 1750.590 ;
        RECT 2048.890 1750.000 2049.170 1750.590 ;
        RECT 630.300 1704.090 630.560 1704.410 ;
        RECT 2042.500 1704.090 2042.760 1704.410 ;
        RECT 630.360 1701.350 630.500 1704.090 ;
        RECT 572.340 1701.030 572.600 1701.350 ;
        RECT 630.300 1701.030 630.560 1701.350 ;
        RECT 572.400 590.910 572.540 1701.030 ;
        RECT 741.390 600.170 741.670 604.000 ;
        RECT 739.840 600.030 741.670 600.170 ;
        RECT 739.840 590.910 739.980 600.030 ;
        RECT 741.390 600.000 741.670 600.030 ;
        RECT 144.540 590.590 144.800 590.910 ;
        RECT 572.340 590.590 572.600 590.910 ;
        RECT 739.780 590.590 740.040 590.910 ;
        RECT 144.600 16.990 144.740 590.590 ;
        RECT 139.480 16.670 139.740 16.990 ;
        RECT 144.540 16.670 144.800 16.990 ;
        RECT 139.540 2.400 139.680 16.670 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 590.250 2497.540 590.570 2497.600 ;
        RECT 1514.390 2497.540 1514.710 2497.600 ;
        RECT 590.250 2497.400 1514.710 2497.540 ;
        RECT 590.250 2497.340 590.570 2497.400 ;
        RECT 1514.390 2497.340 1514.710 2497.400 ;
        RECT 1514.390 1907.640 1514.710 1907.700 ;
        RECT 1904.470 1907.640 1904.790 1907.700 ;
        RECT 1514.390 1907.500 1904.790 1907.640 ;
        RECT 1514.390 1907.440 1514.710 1907.500 ;
        RECT 1904.470 1907.440 1904.790 1907.500 ;
        RECT 537.810 1690.380 538.130 1690.440 ;
        RECT 1351.550 1690.380 1351.870 1690.440 ;
        RECT 537.810 1690.240 1351.870 1690.380 ;
        RECT 537.810 1690.180 538.130 1690.240 ;
        RECT 1351.550 1690.180 1351.870 1690.240 ;
        RECT 1355.690 1690.380 1356.010 1690.440 ;
        RECT 1514.390 1690.380 1514.710 1690.440 ;
        RECT 1355.690 1690.240 1514.710 1690.380 ;
        RECT 1355.690 1690.180 1356.010 1690.240 ;
        RECT 1514.390 1690.180 1514.710 1690.240 ;
        RECT 1351.550 1689.700 1351.870 1689.760 ;
        RECT 1355.690 1689.700 1356.010 1689.760 ;
        RECT 1351.550 1689.560 1356.010 1689.700 ;
        RECT 1351.550 1689.500 1351.870 1689.560 ;
        RECT 1355.690 1689.500 1356.010 1689.560 ;
        RECT 158.310 591.160 158.630 591.220 ;
        RECT 537.810 591.160 538.130 591.220 ;
        RECT 158.310 591.020 538.130 591.160 ;
        RECT 158.310 590.960 158.630 591.020 ;
        RECT 537.810 590.960 538.130 591.020 ;
        RECT 537.810 589.460 538.130 589.520 ;
        RECT 748.950 589.460 749.270 589.520 ;
        RECT 537.810 589.320 749.270 589.460 ;
        RECT 537.810 589.260 538.130 589.320 ;
        RECT 748.950 589.260 749.270 589.320 ;
      LAYER via ;
        RECT 590.280 2497.340 590.540 2497.600 ;
        RECT 1514.420 2497.340 1514.680 2497.600 ;
        RECT 1514.420 1907.440 1514.680 1907.700 ;
        RECT 1904.500 1907.440 1904.760 1907.700 ;
        RECT 537.840 1690.180 538.100 1690.440 ;
        RECT 1351.580 1690.180 1351.840 1690.440 ;
        RECT 1355.720 1690.180 1355.980 1690.440 ;
        RECT 1514.420 1690.180 1514.680 1690.440 ;
        RECT 1351.580 1689.500 1351.840 1689.760 ;
        RECT 1355.720 1689.500 1355.980 1689.760 ;
        RECT 158.340 590.960 158.600 591.220 ;
        RECT 537.840 590.960 538.100 591.220 ;
        RECT 537.840 589.260 538.100 589.520 ;
        RECT 748.980 589.260 749.240 589.520 ;
      LAYER met2 ;
        RECT 590.270 2732.395 590.550 2732.765 ;
        RECT 590.340 2497.630 590.480 2732.395 ;
        RECT 1512.970 2500.770 1513.250 2504.000 ;
        RECT 1512.970 2500.630 1514.620 2500.770 ;
        RECT 1512.970 2500.000 1513.250 2500.630 ;
        RECT 1514.480 2497.630 1514.620 2500.630 ;
        RECT 590.280 2497.310 590.540 2497.630 ;
        RECT 1514.420 2497.310 1514.680 2497.630 ;
        RECT 1514.480 1907.730 1514.620 2497.310 ;
        RECT 1514.420 1907.410 1514.680 1907.730 ;
        RECT 1904.500 1907.410 1904.760 1907.730 ;
        RECT 537.650 1700.410 537.930 1704.000 ;
        RECT 537.650 1700.000 538.040 1700.410 ;
        RECT 537.900 1690.470 538.040 1700.000 ;
        RECT 1514.480 1690.470 1514.620 1907.410 ;
        RECT 1904.560 1907.245 1904.700 1907.410 ;
        RECT 1904.490 1906.875 1904.770 1907.245 ;
        RECT 537.840 1690.150 538.100 1690.470 ;
        RECT 1351.580 1690.150 1351.840 1690.470 ;
        RECT 1355.720 1690.150 1355.980 1690.470 ;
        RECT 1514.420 1690.150 1514.680 1690.470 ;
        RECT 537.900 591.250 538.040 1690.150 ;
        RECT 1351.640 1689.790 1351.780 1690.150 ;
        RECT 1355.780 1689.790 1355.920 1690.150 ;
        RECT 1351.580 1689.470 1351.840 1689.790 ;
        RECT 1355.720 1689.470 1355.980 1689.790 ;
        RECT 750.590 600.170 750.870 604.000 ;
        RECT 749.040 600.030 750.870 600.170 ;
        RECT 158.340 590.930 158.600 591.250 ;
        RECT 537.840 590.930 538.100 591.250 ;
        RECT 158.400 17.410 158.540 590.930 ;
        RECT 537.900 589.550 538.040 590.930 ;
        RECT 749.040 589.550 749.180 600.030 ;
        RECT 750.590 600.000 750.870 600.030 ;
        RECT 537.840 589.230 538.100 589.550 ;
        RECT 748.980 589.230 749.240 589.550 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 590.270 2732.440 590.550 2732.720 ;
        RECT 1904.490 1906.920 1904.770 1907.200 ;
      LAYER met3 ;
        RECT 574.800 2733.320 578.800 2733.920 ;
        RECT 578.070 2732.730 578.370 2733.320 ;
        RECT 590.245 2732.730 590.575 2732.745 ;
        RECT 578.070 2732.430 590.575 2732.730 ;
        RECT 590.245 2732.415 590.575 2732.430 ;
        RECT 1904.465 1907.210 1904.795 1907.225 ;
        RECT 1904.465 1907.040 1920.650 1907.210 ;
        RECT 1904.465 1906.910 1924.000 1907.040 ;
        RECT 1904.465 1906.895 1904.795 1906.910 ;
        RECT 1920.000 1906.440 1924.000 1906.910 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 575.990 2899.420 576.310 2899.480 ;
        RECT 1714.950 2899.420 1715.270 2899.480 ;
        RECT 575.990 2899.280 1715.270 2899.420 ;
        RECT 575.990 2899.220 576.310 2899.280 ;
        RECT 1714.950 2899.220 1715.270 2899.280 ;
        RECT 547.930 2594.100 548.250 2594.160 ;
        RECT 569.090 2594.100 569.410 2594.160 ;
        RECT 575.990 2594.100 576.310 2594.160 ;
        RECT 547.930 2593.960 576.310 2594.100 ;
        RECT 547.930 2593.900 548.250 2593.960 ;
        RECT 569.090 2593.900 569.410 2593.960 ;
        RECT 575.990 2593.900 576.310 2593.960 ;
        RECT 639.010 2035.820 639.330 2035.880 ;
        RECT 2056.270 2035.820 2056.590 2035.880 ;
        RECT 639.010 2035.680 2056.590 2035.820 ;
        RECT 639.010 2035.620 639.330 2035.680 ;
        RECT 2056.270 2035.620 2056.590 2035.680 ;
        RECT 567.710 1994.000 568.030 1994.060 ;
        RECT 569.090 1994.000 569.410 1994.060 ;
        RECT 634.870 1994.000 635.190 1994.060 ;
        RECT 639.010 1994.000 639.330 1994.060 ;
        RECT 567.710 1993.860 639.330 1994.000 ;
        RECT 567.710 1993.800 568.030 1993.860 ;
        RECT 569.090 1993.800 569.410 1993.860 ;
        RECT 634.870 1993.800 635.190 1993.860 ;
        RECT 639.010 1993.800 639.330 1993.860 ;
        RECT 503.310 1990.940 503.630 1991.000 ;
        RECT 567.710 1990.940 568.030 1991.000 ;
        RECT 503.310 1990.800 568.030 1990.940 ;
        RECT 503.310 1990.740 503.630 1990.800 ;
        RECT 567.710 1990.740 568.030 1990.800 ;
        RECT 575.990 590.480 576.310 590.540 ;
        RECT 627.970 590.480 628.290 590.540 ;
        RECT 575.990 590.340 628.290 590.480 ;
        RECT 575.990 590.280 576.310 590.340 ;
        RECT 627.970 590.280 628.290 590.340 ;
        RECT 627.970 588.780 628.290 588.840 ;
        RECT 634.870 588.780 635.190 588.840 ;
        RECT 627.970 588.640 635.190 588.780 ;
        RECT 627.970 588.580 628.290 588.640 ;
        RECT 634.870 588.580 635.190 588.640 ;
        RECT 174.870 41.380 175.190 41.440 ;
        RECT 575.990 41.380 576.310 41.440 ;
        RECT 174.870 41.240 576.310 41.380 ;
        RECT 174.870 41.180 175.190 41.240 ;
        RECT 575.990 41.180 576.310 41.240 ;
      LAYER via ;
        RECT 576.020 2899.220 576.280 2899.480 ;
        RECT 1714.980 2899.220 1715.240 2899.480 ;
        RECT 547.960 2593.900 548.220 2594.160 ;
        RECT 569.120 2593.900 569.380 2594.160 ;
        RECT 576.020 2593.900 576.280 2594.160 ;
        RECT 639.040 2035.620 639.300 2035.880 ;
        RECT 2056.300 2035.620 2056.560 2035.880 ;
        RECT 567.740 1993.800 568.000 1994.060 ;
        RECT 569.120 1993.800 569.380 1994.060 ;
        RECT 634.900 1993.800 635.160 1994.060 ;
        RECT 639.040 1993.800 639.300 1994.060 ;
        RECT 503.340 1990.740 503.600 1991.000 ;
        RECT 567.740 1990.740 568.000 1991.000 ;
        RECT 576.020 590.280 576.280 590.540 ;
        RECT 628.000 590.280 628.260 590.540 ;
        RECT 628.000 588.580 628.260 588.840 ;
        RECT 634.900 588.580 635.160 588.840 ;
        RECT 174.900 41.180 175.160 41.440 ;
        RECT 576.020 41.180 576.280 41.440 ;
      LAYER met2 ;
        RECT 576.020 2899.190 576.280 2899.510 ;
        RECT 1714.980 2899.250 1715.240 2899.510 ;
        RECT 1716.290 2899.250 1716.570 2900.055 ;
        RECT 1714.980 2899.190 1716.570 2899.250 ;
        RECT 547.850 2600.660 548.130 2604.000 ;
        RECT 547.850 2600.000 548.160 2600.660 ;
        RECT 548.020 2594.190 548.160 2600.000 ;
        RECT 576.080 2594.190 576.220 2899.190 ;
        RECT 1715.040 2899.110 1716.570 2899.190 ;
        RECT 1716.290 2896.055 1716.570 2899.110 ;
        RECT 547.960 2593.870 548.220 2594.190 ;
        RECT 569.120 2593.870 569.380 2594.190 ;
        RECT 576.020 2593.870 576.280 2594.190 ;
        RECT 569.180 1994.090 569.320 2593.870 ;
        RECT 639.040 2035.590 639.300 2035.910 ;
        RECT 2056.300 2035.590 2056.560 2035.910 ;
        RECT 639.100 1994.090 639.240 2035.590 ;
        RECT 567.740 1993.770 568.000 1994.090 ;
        RECT 569.120 1993.770 569.380 1994.090 ;
        RECT 634.900 1993.770 635.160 1994.090 ;
        RECT 639.040 1993.770 639.300 1994.090 ;
        RECT 567.800 1991.030 567.940 1993.770 ;
        RECT 503.340 1990.710 503.600 1991.030 ;
        RECT 567.740 1990.710 568.000 1991.030 ;
        RECT 502.690 1981.250 502.970 1981.750 ;
        RECT 503.400 1981.250 503.540 1990.710 ;
        RECT 502.690 1981.110 503.540 1981.250 ;
        RECT 502.690 1977.750 502.970 1981.110 ;
        RECT 634.960 590.765 635.100 1993.770 ;
        RECT 2056.360 1917.095 2056.500 2035.590 ;
        RECT 2056.250 1913.095 2056.530 1917.095 ;
        RECT 759.790 600.170 760.070 604.000 ;
        RECT 759.160 600.030 760.070 600.170 ;
        RECT 759.160 590.765 759.300 600.030 ;
        RECT 759.790 600.000 760.070 600.030 ;
        RECT 576.020 590.250 576.280 590.570 ;
        RECT 628.000 590.250 628.260 590.570 ;
        RECT 634.890 590.395 635.170 590.765 ;
        RECT 759.090 590.395 759.370 590.765 ;
        RECT 576.080 41.470 576.220 590.250 ;
        RECT 628.060 588.870 628.200 590.250 ;
        RECT 634.960 588.870 635.100 590.395 ;
        RECT 628.000 588.550 628.260 588.870 ;
        RECT 634.900 588.550 635.160 588.870 ;
        RECT 174.900 41.150 175.160 41.470 ;
        RECT 576.020 41.150 576.280 41.470 ;
        RECT 174.960 2.400 175.100 41.150 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 634.890 590.440 635.170 590.720 ;
        RECT 759.090 590.440 759.370 590.720 ;
      LAYER met3 ;
        RECT 634.865 590.730 635.195 590.745 ;
        RECT 759.065 590.730 759.395 590.745 ;
        RECT 634.865 590.430 759.395 590.730 ;
        RECT 634.865 590.415 635.195 590.430 ;
        RECT 759.065 590.415 759.395 590.430 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.870 2901.460 428.190 2901.520 ;
        RECT 1726.450 2901.460 1726.770 2901.520 ;
        RECT 427.870 2901.320 1726.770 2901.460 ;
        RECT 427.870 2901.260 428.190 2901.320 ;
        RECT 1726.450 2901.260 1726.770 2901.320 ;
        RECT 996.890 2032.420 997.210 2032.480 ;
        RECT 2014.870 2032.420 2015.190 2032.480 ;
        RECT 996.890 2032.280 2015.190 2032.420 ;
        RECT 996.890 2032.220 997.210 2032.280 ;
        RECT 2014.870 2032.220 2015.190 2032.280 ;
        RECT 419.590 1980.060 419.910 1980.120 ;
        RECT 422.810 1980.060 423.130 1980.120 ;
        RECT 419.590 1979.920 423.130 1980.060 ;
        RECT 419.590 1979.860 419.910 1979.920 ;
        RECT 422.810 1979.860 423.130 1979.920 ;
        RECT 422.810 1978.700 423.130 1978.760 ;
        RECT 422.810 1978.560 496.180 1978.700 ;
        RECT 422.810 1978.500 423.130 1978.560 ;
        RECT 418.670 1978.160 418.990 1978.420 ;
        RECT 496.040 1978.360 496.180 1978.560 ;
        RECT 634.410 1978.360 634.730 1978.420 ;
        RECT 496.040 1978.220 634.730 1978.360 ;
        RECT 634.410 1978.160 634.730 1978.220 ;
        RECT 361.630 1977.680 361.950 1977.740 ;
        RECT 418.760 1977.680 418.900 1978.160 ;
        RECT 361.630 1977.540 418.900 1977.680 ;
        RECT 361.630 1977.480 361.950 1977.540 ;
        RECT 2014.870 1966.460 2015.190 1966.520 ;
        RECT 2019.470 1966.460 2019.790 1966.520 ;
        RECT 2014.870 1966.320 2019.790 1966.460 ;
        RECT 2014.870 1966.260 2015.190 1966.320 ;
        RECT 2019.470 1966.260 2019.790 1966.320 ;
        RECT 634.410 1959.660 634.730 1959.720 ;
        RECT 996.890 1959.660 997.210 1959.720 ;
        RECT 634.410 1959.520 997.210 1959.660 ;
        RECT 634.410 1959.460 634.730 1959.520 ;
        RECT 996.890 1959.460 997.210 1959.520 ;
        RECT 733.310 591.840 733.630 591.900 ;
        RECT 767.350 591.840 767.670 591.900 ;
        RECT 733.310 591.700 767.670 591.840 ;
        RECT 733.310 591.640 733.630 591.700 ;
        RECT 767.350 591.640 767.670 591.700 ;
        RECT 192.810 46.140 193.130 46.200 ;
        RECT 732.390 46.140 732.710 46.200 ;
        RECT 192.810 46.000 732.710 46.140 ;
        RECT 192.810 45.940 193.130 46.000 ;
        RECT 732.390 45.940 732.710 46.000 ;
      LAYER via ;
        RECT 427.900 2901.260 428.160 2901.520 ;
        RECT 1726.480 2901.260 1726.740 2901.520 ;
        RECT 996.920 2032.220 997.180 2032.480 ;
        RECT 2014.900 2032.220 2015.160 2032.480 ;
        RECT 419.620 1979.860 419.880 1980.120 ;
        RECT 422.840 1979.860 423.100 1980.120 ;
        RECT 422.840 1978.500 423.100 1978.760 ;
        RECT 418.700 1978.160 418.960 1978.420 ;
        RECT 634.440 1978.160 634.700 1978.420 ;
        RECT 361.660 1977.480 361.920 1977.740 ;
        RECT 2014.900 1966.260 2015.160 1966.520 ;
        RECT 2019.500 1966.260 2019.760 1966.520 ;
        RECT 634.440 1959.460 634.700 1959.720 ;
        RECT 996.920 1959.460 997.180 1959.720 ;
        RECT 733.340 591.640 733.600 591.900 ;
        RECT 767.380 591.640 767.640 591.900 ;
        RECT 192.840 45.940 193.100 46.200 ;
        RECT 732.420 45.940 732.680 46.200 ;
      LAYER met2 ;
        RECT 427.900 2901.230 428.160 2901.550 ;
        RECT 1726.480 2901.230 1726.740 2901.550 ;
        RECT 427.960 2688.905 428.100 2901.230 ;
        RECT 1726.540 2900.055 1726.680 2901.230 ;
        RECT 1726.410 2896.055 1726.690 2900.055 ;
        RECT 427.890 2688.535 428.170 2688.905 ;
        RECT 419.610 2685.475 419.890 2685.845 ;
        RECT 419.680 1980.150 419.820 2685.475 ;
        RECT 996.920 2032.190 997.180 2032.510 ;
        RECT 2014.900 2032.190 2015.160 2032.510 ;
        RECT 419.620 1979.830 419.880 1980.150 ;
        RECT 422.840 1979.830 423.100 1980.150 ;
        RECT 419.680 1978.530 419.820 1979.830 ;
        RECT 422.900 1978.790 423.040 1979.830 ;
        RECT 418.760 1978.450 419.820 1978.530 ;
        RECT 422.840 1978.470 423.100 1978.790 ;
        RECT 418.700 1978.390 419.820 1978.450 ;
        RECT 418.700 1978.130 418.960 1978.390 ;
        RECT 634.440 1978.130 634.700 1978.450 ;
        RECT 361.660 1977.450 361.920 1977.770 ;
        RECT 361.720 1965.045 361.860 1977.450 ;
        RECT 361.650 1964.675 361.930 1965.045 ;
        RECT 634.500 1959.750 634.640 1978.130 ;
        RECT 996.980 1959.750 997.120 2032.190 ;
        RECT 2014.960 1966.550 2015.100 2032.190 ;
        RECT 2014.900 1966.230 2015.160 1966.550 ;
        RECT 2019.500 1966.230 2019.760 1966.550 ;
        RECT 634.440 1959.430 634.700 1959.750 ;
        RECT 996.920 1959.430 997.180 1959.750 ;
        RECT 634.500 590.085 634.640 1959.430 ;
        RECT 2019.560 1916.650 2019.700 1966.230 ;
        RECT 2021.290 1916.650 2021.570 1917.095 ;
        RECT 2019.560 1916.510 2021.570 1916.650 ;
        RECT 2021.290 1913.095 2021.570 1916.510 ;
        RECT 768.990 600.170 769.270 604.000 ;
        RECT 767.440 600.030 769.270 600.170 ;
        RECT 767.440 591.930 767.580 600.030 ;
        RECT 768.990 600.000 769.270 600.030 ;
        RECT 733.340 591.610 733.600 591.930 ;
        RECT 767.380 591.610 767.640 591.930 ;
        RECT 733.400 590.085 733.540 591.610 ;
        RECT 634.430 589.715 634.710 590.085 ;
        RECT 732.410 589.715 732.690 590.085 ;
        RECT 733.330 589.715 733.610 590.085 ;
        RECT 732.480 46.230 732.620 589.715 ;
        RECT 192.840 45.910 193.100 46.230 ;
        RECT 732.420 45.910 732.680 46.230 ;
        RECT 192.900 2.400 193.040 45.910 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 427.890 2688.580 428.170 2688.860 ;
        RECT 419.610 2685.520 419.890 2685.800 ;
        RECT 361.650 1964.720 361.930 1965.000 ;
        RECT 634.430 589.760 634.710 590.040 ;
        RECT 732.410 589.760 732.690 590.040 ;
        RECT 733.330 589.760 733.610 590.040 ;
      LAYER met3 ;
        RECT 427.865 2688.870 428.195 2688.885 ;
        RECT 430.000 2688.870 434.000 2689.040 ;
        RECT 427.865 2688.570 434.000 2688.870 ;
        RECT 427.865 2688.555 428.195 2688.570 ;
        RECT 429.950 2688.440 434.000 2688.570 ;
        RECT 419.585 2685.810 419.915 2685.825 ;
        RECT 429.950 2685.810 430.250 2688.440 ;
        RECT 419.585 2685.510 430.250 2685.810 ;
        RECT 419.585 2685.495 419.915 2685.510 ;
        RECT 361.625 1965.010 361.955 1965.025 ;
        RECT 361.625 1964.695 362.170 1965.010 ;
        RECT 361.870 1963.120 362.170 1964.695 ;
        RECT 360.000 1962.520 364.000 1963.120 ;
        RECT 634.405 590.050 634.735 590.065 ;
        RECT 732.385 590.050 732.715 590.065 ;
        RECT 733.305 590.050 733.635 590.065 ;
        RECT 634.405 589.750 733.635 590.050 ;
        RECT 634.405 589.735 634.735 589.750 ;
        RECT 732.385 589.735 732.715 589.750 ;
        RECT 733.305 589.735 733.635 589.750 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 593.010 2712.080 593.330 2712.140 ;
        RECT 776.090 2712.080 776.410 2712.140 ;
        RECT 593.010 2711.940 776.410 2712.080 ;
        RECT 593.010 2711.880 593.330 2711.940 ;
        RECT 776.090 2711.880 776.410 2711.940 ;
        RECT 776.090 2489.040 776.410 2489.100 ;
        RECT 1598.570 2489.040 1598.890 2489.100 ;
        RECT 776.090 2488.900 1598.890 2489.040 ;
        RECT 776.090 2488.840 776.410 2488.900 ;
        RECT 1598.570 2488.840 1598.890 2488.900 ;
        RECT 776.090 2484.620 776.410 2484.680 ;
        RECT 779.310 2484.620 779.630 2484.680 ;
        RECT 776.090 2484.480 779.630 2484.620 ;
        RECT 776.090 2484.420 776.410 2484.480 ;
        RECT 779.310 2484.420 779.630 2484.480 ;
        RECT 776.090 2038.200 776.410 2038.260 ;
        RECT 779.310 2038.200 779.630 2038.260 ;
        RECT 776.090 2038.060 779.630 2038.200 ;
        RECT 776.090 2038.000 776.410 2038.060 ;
        RECT 779.310 2038.000 779.630 2038.060 ;
        RECT 779.310 2036.160 779.630 2036.220 ;
        RECT 2084.330 2036.160 2084.650 2036.220 ;
        RECT 779.310 2036.020 2084.650 2036.160 ;
        RECT 779.310 2035.960 779.630 2036.020 ;
        RECT 2084.330 2035.960 2084.650 2036.020 ;
        RECT 641.310 1990.600 641.630 1990.660 ;
        RECT 776.090 1990.600 776.410 1990.660 ;
        RECT 641.310 1990.460 776.410 1990.600 ;
        RECT 641.310 1990.400 641.630 1990.460 ;
        RECT 776.090 1990.400 776.410 1990.460 ;
        RECT 429.710 1987.880 430.030 1987.940 ;
        RECT 641.310 1987.880 641.630 1987.940 ;
        RECT 429.710 1987.740 641.630 1987.880 ;
        RECT 429.710 1987.680 430.030 1987.740 ;
        RECT 641.310 1987.680 641.630 1987.740 ;
        RECT 641.310 593.540 641.630 593.600 ;
        RECT 773.330 593.540 773.650 593.600 ;
        RECT 776.550 593.540 776.870 593.600 ;
        RECT 641.310 593.400 776.870 593.540 ;
        RECT 641.310 593.340 641.630 593.400 ;
        RECT 773.330 593.340 773.650 593.400 ;
        RECT 776.550 593.340 776.870 593.400 ;
        RECT 213.510 52.260 213.830 52.320 ;
        RECT 773.330 52.260 773.650 52.320 ;
        RECT 213.510 52.120 773.650 52.260 ;
        RECT 213.510 52.060 213.830 52.120 ;
        RECT 773.330 52.060 773.650 52.120 ;
        RECT 210.750 16.900 211.070 16.960 ;
        RECT 213.510 16.900 213.830 16.960 ;
        RECT 210.750 16.760 213.830 16.900 ;
        RECT 210.750 16.700 211.070 16.760 ;
        RECT 213.510 16.700 213.830 16.760 ;
      LAYER via ;
        RECT 593.040 2711.880 593.300 2712.140 ;
        RECT 776.120 2711.880 776.380 2712.140 ;
        RECT 776.120 2488.840 776.380 2489.100 ;
        RECT 1598.600 2488.840 1598.860 2489.100 ;
        RECT 776.120 2484.420 776.380 2484.680 ;
        RECT 779.340 2484.420 779.600 2484.680 ;
        RECT 776.120 2038.000 776.380 2038.260 ;
        RECT 779.340 2038.000 779.600 2038.260 ;
        RECT 779.340 2035.960 779.600 2036.220 ;
        RECT 2084.360 2035.960 2084.620 2036.220 ;
        RECT 641.340 1990.400 641.600 1990.660 ;
        RECT 776.120 1990.400 776.380 1990.660 ;
        RECT 429.740 1987.680 430.000 1987.940 ;
        RECT 641.340 1987.680 641.600 1987.940 ;
        RECT 641.340 593.340 641.600 593.600 ;
        RECT 773.360 593.340 773.620 593.600 ;
        RECT 776.580 593.340 776.840 593.600 ;
        RECT 213.540 52.060 213.800 52.320 ;
        RECT 773.360 52.060 773.620 52.320 ;
        RECT 210.780 16.700 211.040 16.960 ;
        RECT 213.540 16.700 213.800 16.960 ;
      LAYER met2 ;
        RECT 593.030 2711.995 593.310 2712.365 ;
        RECT 593.040 2711.850 593.300 2711.995 ;
        RECT 776.120 2711.850 776.380 2712.170 ;
        RECT 776.180 2489.130 776.320 2711.850 ;
        RECT 1598.530 2500.000 1598.810 2504.000 ;
        RECT 1598.660 2489.130 1598.800 2500.000 ;
        RECT 776.120 2488.810 776.380 2489.130 ;
        RECT 1598.600 2488.810 1598.860 2489.130 ;
        RECT 776.180 2484.710 776.320 2488.810 ;
        RECT 776.120 2484.390 776.380 2484.710 ;
        RECT 779.340 2484.390 779.600 2484.710 ;
        RECT 779.400 2038.290 779.540 2484.390 ;
        RECT 776.120 2037.970 776.380 2038.290 ;
        RECT 779.340 2037.970 779.600 2038.290 ;
        RECT 776.180 1990.690 776.320 2037.970 ;
        RECT 779.400 2036.250 779.540 2037.970 ;
        RECT 779.340 2035.930 779.600 2036.250 ;
        RECT 2084.360 2035.930 2084.620 2036.250 ;
        RECT 641.340 1990.370 641.600 1990.690 ;
        RECT 776.120 1990.370 776.380 1990.690 ;
        RECT 641.400 1987.970 641.540 1990.370 ;
        RECT 429.740 1987.650 430.000 1987.970 ;
        RECT 641.340 1987.650 641.600 1987.970 ;
        RECT 428.170 1981.250 428.450 1981.750 ;
        RECT 429.800 1981.250 429.940 1987.650 ;
        RECT 428.170 1981.110 429.940 1981.250 ;
        RECT 428.170 1977.750 428.450 1981.110 ;
        RECT 641.400 593.630 641.540 1987.650 ;
        RECT 2084.420 1904.525 2084.560 2035.930 ;
        RECT 2084.350 1904.155 2084.630 1904.525 ;
        RECT 778.190 600.170 778.470 604.000 ;
        RECT 776.640 600.030 778.470 600.170 ;
        RECT 776.640 593.630 776.780 600.030 ;
        RECT 778.190 600.000 778.470 600.030 ;
        RECT 641.340 593.310 641.600 593.630 ;
        RECT 773.360 593.310 773.620 593.630 ;
        RECT 776.580 593.310 776.840 593.630 ;
        RECT 773.420 52.350 773.560 593.310 ;
        RECT 213.540 52.030 213.800 52.350 ;
        RECT 773.360 52.030 773.620 52.350 ;
        RECT 213.600 16.990 213.740 52.030 ;
        RECT 210.780 16.670 211.040 16.990 ;
        RECT 213.540 16.670 213.800 16.990 ;
        RECT 210.840 2.400 210.980 16.670 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 593.030 2712.040 593.310 2712.320 ;
        RECT 2084.350 1904.200 2084.630 1904.480 ;
      LAYER met3 ;
        RECT 593.005 2712.330 593.335 2712.345 ;
        RECT 578.070 2712.160 593.335 2712.330 ;
        RECT 574.800 2712.030 593.335 2712.160 ;
        RECT 574.800 2711.560 578.800 2712.030 ;
        RECT 593.005 2712.015 593.335 2712.030 ;
        RECT 2084.325 1904.490 2084.655 1904.505 ;
        RECT 2075.830 1904.320 2084.655 1904.490 ;
        RECT 2072.375 1904.190 2084.655 1904.320 ;
        RECT 2072.375 1903.720 2076.375 1904.190 ;
        RECT 2084.325 1904.175 2084.655 1904.190 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 489.970 2592.060 490.290 2592.120 ;
        RECT 638.090 2592.060 638.410 2592.120 ;
        RECT 489.970 2591.920 638.410 2592.060 ;
        RECT 489.970 2591.860 490.290 2591.920 ;
        RECT 638.090 2591.860 638.410 2591.920 ;
        RECT 641.310 2489.720 641.630 2489.780 ;
        RECT 1672.170 2489.720 1672.490 2489.780 ;
        RECT 641.310 2489.580 1672.490 2489.720 ;
        RECT 641.310 2489.520 641.630 2489.580 ;
        RECT 1672.170 2489.520 1672.490 2489.580 ;
        RECT 638.090 2488.020 638.410 2488.080 ;
        RECT 641.310 2488.020 641.630 2488.080 ;
        RECT 638.090 2487.880 641.630 2488.020 ;
        RECT 638.090 2487.820 638.410 2487.880 ;
        RECT 641.310 2487.820 641.630 2487.880 ;
        RECT 627.970 1991.280 628.290 1991.340 ;
        RECT 641.310 1991.280 641.630 1991.340 ;
        RECT 690.070 1991.280 690.390 1991.340 ;
        RECT 627.970 1991.140 690.390 1991.280 ;
        RECT 627.970 1991.080 628.290 1991.140 ;
        RECT 641.310 1991.080 641.630 1991.140 ;
        RECT 690.070 1991.080 690.390 1991.140 ;
        RECT 644.070 1702.620 644.390 1702.680 ;
        RECT 689.610 1702.620 689.930 1702.680 ;
        RECT 869.470 1702.620 869.790 1702.680 ;
        RECT 644.070 1702.480 689.930 1702.620 ;
        RECT 644.070 1702.420 644.390 1702.480 ;
        RECT 689.610 1702.420 689.930 1702.480 ;
        RECT 834.600 1702.480 869.790 1702.620 ;
        RECT 785.750 1702.280 786.070 1702.340 ;
        RECT 772.500 1702.140 786.070 1702.280 ;
        RECT 691.450 1701.940 691.770 1702.000 ;
        RECT 724.570 1701.940 724.890 1702.000 ;
        RECT 691.450 1701.800 724.890 1701.940 ;
        RECT 691.450 1701.740 691.770 1701.800 ;
        RECT 724.570 1701.740 724.890 1701.800 ;
        RECT 738.830 1701.940 739.150 1702.000 ;
        RECT 772.500 1701.940 772.640 1702.140 ;
        RECT 785.750 1702.080 786.070 1702.140 ;
        RECT 787.130 1702.280 787.450 1702.340 ;
        RECT 834.600 1702.280 834.740 1702.480 ;
        RECT 869.470 1702.420 869.790 1702.480 ;
        RECT 966.070 1702.620 966.390 1702.680 ;
        RECT 1279.790 1702.620 1280.110 1702.680 ;
        RECT 1303.710 1702.620 1304.030 1702.680 ;
        RECT 1400.310 1702.620 1400.630 1702.680 ;
        RECT 1641.810 1702.620 1642.130 1702.680 ;
        RECT 1642.730 1702.620 1643.050 1702.680 ;
        RECT 1751.290 1702.620 1751.610 1702.680 ;
        RECT 966.070 1702.480 1028.400 1702.620 ;
        RECT 966.070 1702.420 966.390 1702.480 ;
        RECT 787.130 1702.140 834.740 1702.280 ;
        RECT 917.310 1702.280 917.630 1702.340 ;
        RECT 1028.260 1702.280 1028.400 1702.480 ;
        RECT 1279.790 1702.480 1304.030 1702.620 ;
        RECT 1279.790 1702.420 1280.110 1702.480 ;
        RECT 1303.710 1702.420 1304.030 1702.480 ;
        RECT 1366.820 1702.480 1400.630 1702.620 ;
        RECT 1076.010 1702.280 1076.330 1702.340 ;
        RECT 917.310 1702.140 931.340 1702.280 ;
        RECT 1028.260 1702.140 1076.330 1702.280 ;
        RECT 787.130 1702.080 787.450 1702.140 ;
        RECT 917.310 1702.080 917.630 1702.140 ;
        RECT 738.830 1701.800 772.640 1701.940 ;
        RECT 931.200 1701.940 931.340 1702.140 ;
        RECT 1076.010 1702.080 1076.330 1702.140 ;
        RECT 1200.210 1702.280 1200.530 1702.340 ;
        RECT 1200.210 1702.140 1268.980 1702.280 ;
        RECT 1200.210 1702.080 1200.530 1702.140 ;
        RECT 966.070 1701.940 966.390 1702.000 ;
        RECT 931.200 1701.800 966.390 1701.940 ;
        RECT 738.830 1701.740 739.150 1701.800 ;
        RECT 966.070 1701.740 966.390 1701.800 ;
        RECT 1124.770 1701.940 1125.090 1702.000 ;
        RECT 1152.370 1701.940 1152.690 1702.000 ;
        RECT 1124.770 1701.800 1152.690 1701.940 ;
        RECT 1268.840 1701.940 1268.980 1702.140 ;
        RECT 1279.790 1701.940 1280.110 1702.000 ;
        RECT 1268.840 1701.800 1280.110 1701.940 ;
        RECT 1124.770 1701.740 1125.090 1701.800 ;
        RECT 1152.370 1701.740 1152.690 1701.800 ;
        RECT 1279.790 1701.740 1280.110 1701.800 ;
        RECT 1304.170 1701.940 1304.490 1702.000 ;
        RECT 1304.170 1701.800 1351.780 1701.940 ;
        RECT 1304.170 1701.740 1304.490 1701.800 ;
        RECT 869.930 1701.600 870.250 1701.660 ;
        RECT 917.310 1701.600 917.630 1701.660 ;
        RECT 869.930 1701.460 917.630 1701.600 ;
        RECT 869.930 1701.400 870.250 1701.460 ;
        RECT 917.310 1701.400 917.630 1701.460 ;
        RECT 1076.930 1701.600 1077.250 1701.660 ;
        RECT 1124.310 1701.600 1124.630 1701.660 ;
        RECT 1076.930 1701.460 1124.630 1701.600 ;
        RECT 1351.640 1701.600 1351.780 1701.800 ;
        RECT 1366.820 1701.600 1366.960 1702.480 ;
        RECT 1400.310 1702.420 1400.630 1702.480 ;
        RECT 1510.800 1702.480 1511.400 1702.620 ;
        RECT 1401.230 1702.280 1401.550 1702.340 ;
        RECT 1510.800 1702.280 1510.940 1702.480 ;
        RECT 1401.230 1702.140 1441.940 1702.280 ;
        RECT 1401.230 1702.080 1401.550 1702.140 ;
        RECT 1351.640 1701.460 1366.960 1701.600 ;
        RECT 1441.800 1701.600 1441.940 1702.140 ;
        RECT 1468.940 1702.140 1510.940 1702.280 ;
        RECT 1511.260 1702.280 1511.400 1702.480 ;
        RECT 1641.810 1702.480 1643.050 1702.620 ;
        RECT 1641.810 1702.420 1642.130 1702.480 ;
        RECT 1642.730 1702.420 1643.050 1702.480 ;
        RECT 1738.500 1702.480 1751.610 1702.620 ;
        RECT 1565.450 1702.280 1565.770 1702.340 ;
        RECT 1690.570 1702.280 1690.890 1702.340 ;
        RECT 1511.260 1702.140 1565.770 1702.280 ;
        RECT 1462.410 1701.940 1462.730 1702.000 ;
        RECT 1448.700 1701.800 1462.730 1701.940 ;
        RECT 1448.700 1701.600 1448.840 1701.800 ;
        RECT 1462.410 1701.740 1462.730 1701.800 ;
        RECT 1462.870 1701.940 1463.190 1702.000 ;
        RECT 1468.940 1701.940 1469.080 1702.140 ;
        RECT 1565.450 1702.080 1565.770 1702.140 ;
        RECT 1658.000 1702.140 1690.890 1702.280 ;
        RECT 1462.870 1701.800 1469.080 1701.940 ;
        RECT 1565.910 1701.940 1566.230 1702.000 ;
        RECT 1593.970 1701.940 1594.290 1702.000 ;
        RECT 1565.910 1701.800 1594.290 1701.940 ;
        RECT 1462.870 1701.740 1463.190 1701.800 ;
        RECT 1565.910 1701.740 1566.230 1701.800 ;
        RECT 1593.970 1701.740 1594.290 1701.800 ;
        RECT 1642.730 1701.940 1643.050 1702.000 ;
        RECT 1658.000 1701.940 1658.140 1702.140 ;
        RECT 1690.570 1702.080 1690.890 1702.140 ;
        RECT 1709.430 1702.280 1709.750 1702.340 ;
        RECT 1738.500 1702.280 1738.640 1702.480 ;
        RECT 1751.290 1702.420 1751.610 1702.480 ;
        RECT 1709.430 1702.140 1738.640 1702.280 ;
        RECT 1835.010 1702.280 1835.330 1702.340 ;
        RECT 1848.350 1702.280 1848.670 1702.340 ;
        RECT 1835.010 1702.140 1848.670 1702.280 ;
        RECT 1709.430 1702.080 1709.750 1702.140 ;
        RECT 1835.010 1702.080 1835.330 1702.140 ;
        RECT 1848.350 1702.080 1848.670 1702.140 ;
        RECT 1642.730 1701.800 1658.140 1701.940 ;
        RECT 1786.710 1701.940 1787.030 1702.000 ;
        RECT 1849.730 1701.940 1850.050 1702.000 ;
        RECT 1883.770 1701.940 1884.090 1702.000 ;
        RECT 1786.710 1701.800 1787.400 1701.940 ;
        RECT 1642.730 1701.740 1643.050 1701.800 ;
        RECT 1786.710 1701.740 1787.030 1701.800 ;
        RECT 1787.260 1701.660 1787.400 1701.800 ;
        RECT 1849.730 1701.800 1884.090 1701.940 ;
        RECT 1849.730 1701.740 1850.050 1701.800 ;
        RECT 1883.770 1701.740 1884.090 1701.800 ;
        RECT 1441.800 1701.460 1448.840 1701.600 ;
        RECT 1076.930 1701.400 1077.250 1701.460 ;
        RECT 1124.310 1701.400 1124.630 1701.460 ;
        RECT 1787.170 1701.400 1787.490 1701.660 ;
        RECT 1593.970 1701.260 1594.290 1701.320 ;
        RECT 1641.810 1701.260 1642.130 1701.320 ;
        RECT 1593.970 1701.120 1642.130 1701.260 ;
        RECT 1593.970 1701.060 1594.290 1701.120 ;
        RECT 1641.810 1701.060 1642.130 1701.120 ;
        RECT 644.070 596.940 644.390 597.000 ;
        RECT 696.970 596.940 697.290 597.000 ;
        RECT 644.070 596.800 697.290 596.940 ;
        RECT 644.070 596.740 644.390 596.800 ;
        RECT 696.970 596.740 697.290 596.800 ;
        RECT 693.750 593.200 694.070 593.260 ;
        RECT 696.970 593.200 697.290 593.260 ;
        RECT 786.670 593.200 786.990 593.260 ;
        RECT 693.750 593.060 786.990 593.200 ;
        RECT 693.750 593.000 694.070 593.060 ;
        RECT 696.970 593.000 697.290 593.060 ;
        RECT 786.670 593.000 786.990 593.060 ;
        RECT 228.690 47.840 229.010 47.900 ;
        RECT 693.290 47.840 693.610 47.900 ;
        RECT 228.690 47.700 693.610 47.840 ;
        RECT 228.690 47.640 229.010 47.700 ;
        RECT 693.290 47.640 693.610 47.700 ;
      LAYER via ;
        RECT 490.000 2591.860 490.260 2592.120 ;
        RECT 638.120 2591.860 638.380 2592.120 ;
        RECT 641.340 2489.520 641.600 2489.780 ;
        RECT 1672.200 2489.520 1672.460 2489.780 ;
        RECT 638.120 2487.820 638.380 2488.080 ;
        RECT 641.340 2487.820 641.600 2488.080 ;
        RECT 628.000 1991.080 628.260 1991.340 ;
        RECT 641.340 1991.080 641.600 1991.340 ;
        RECT 690.100 1991.080 690.360 1991.340 ;
        RECT 644.100 1702.420 644.360 1702.680 ;
        RECT 689.640 1702.420 689.900 1702.680 ;
        RECT 691.480 1701.740 691.740 1702.000 ;
        RECT 724.600 1701.740 724.860 1702.000 ;
        RECT 738.860 1701.740 739.120 1702.000 ;
        RECT 785.780 1702.080 786.040 1702.340 ;
        RECT 787.160 1702.080 787.420 1702.340 ;
        RECT 869.500 1702.420 869.760 1702.680 ;
        RECT 966.100 1702.420 966.360 1702.680 ;
        RECT 917.340 1702.080 917.600 1702.340 ;
        RECT 1279.820 1702.420 1280.080 1702.680 ;
        RECT 1303.740 1702.420 1304.000 1702.680 ;
        RECT 1076.040 1702.080 1076.300 1702.340 ;
        RECT 1200.240 1702.080 1200.500 1702.340 ;
        RECT 966.100 1701.740 966.360 1702.000 ;
        RECT 1124.800 1701.740 1125.060 1702.000 ;
        RECT 1152.400 1701.740 1152.660 1702.000 ;
        RECT 1279.820 1701.740 1280.080 1702.000 ;
        RECT 1304.200 1701.740 1304.460 1702.000 ;
        RECT 869.960 1701.400 870.220 1701.660 ;
        RECT 917.340 1701.400 917.600 1701.660 ;
        RECT 1076.960 1701.400 1077.220 1701.660 ;
        RECT 1124.340 1701.400 1124.600 1701.660 ;
        RECT 1400.340 1702.420 1400.600 1702.680 ;
        RECT 1401.260 1702.080 1401.520 1702.340 ;
        RECT 1641.840 1702.420 1642.100 1702.680 ;
        RECT 1642.760 1702.420 1643.020 1702.680 ;
        RECT 1462.440 1701.740 1462.700 1702.000 ;
        RECT 1462.900 1701.740 1463.160 1702.000 ;
        RECT 1565.480 1702.080 1565.740 1702.340 ;
        RECT 1565.940 1701.740 1566.200 1702.000 ;
        RECT 1594.000 1701.740 1594.260 1702.000 ;
        RECT 1642.760 1701.740 1643.020 1702.000 ;
        RECT 1690.600 1702.080 1690.860 1702.340 ;
        RECT 1709.460 1702.080 1709.720 1702.340 ;
        RECT 1751.320 1702.420 1751.580 1702.680 ;
        RECT 1835.040 1702.080 1835.300 1702.340 ;
        RECT 1848.380 1702.080 1848.640 1702.340 ;
        RECT 1786.740 1701.740 1787.000 1702.000 ;
        RECT 1849.760 1701.740 1850.020 1702.000 ;
        RECT 1883.800 1701.740 1884.060 1702.000 ;
        RECT 1787.200 1701.400 1787.460 1701.660 ;
        RECT 1594.000 1701.060 1594.260 1701.320 ;
        RECT 1641.840 1701.060 1642.100 1701.320 ;
        RECT 644.100 596.740 644.360 597.000 ;
        RECT 697.000 596.740 697.260 597.000 ;
        RECT 693.780 593.000 694.040 593.260 ;
        RECT 697.000 593.000 697.260 593.260 ;
        RECT 786.700 593.000 786.960 593.260 ;
        RECT 228.720 47.640 228.980 47.900 ;
        RECT 693.320 47.640 693.580 47.900 ;
      LAYER met2 ;
        RECT 489.890 2600.660 490.170 2604.000 ;
        RECT 489.890 2600.000 490.200 2600.660 ;
        RECT 490.060 2592.150 490.200 2600.000 ;
        RECT 490.000 2591.830 490.260 2592.150 ;
        RECT 638.120 2591.830 638.380 2592.150 ;
        RECT 638.180 2488.110 638.320 2591.830 ;
        RECT 1672.130 2500.000 1672.410 2504.000 ;
        RECT 1672.260 2489.810 1672.400 2500.000 ;
        RECT 641.340 2489.490 641.600 2489.810 ;
        RECT 1672.200 2489.490 1672.460 2489.810 ;
        RECT 641.400 2488.110 641.540 2489.490 ;
        RECT 638.120 2487.790 638.380 2488.110 ;
        RECT 641.340 2487.790 641.600 2488.110 ;
        RECT 641.400 1991.370 641.540 2487.790 ;
        RECT 628.000 1991.050 628.260 1991.370 ;
        RECT 641.340 1991.050 641.600 1991.370 ;
        RECT 690.100 1991.050 690.360 1991.370 ;
        RECT 628.060 1981.750 628.200 1991.050 ;
        RECT 627.810 1981.110 628.200 1981.750 ;
        RECT 627.810 1977.750 628.090 1981.110 ;
        RECT 644.100 1702.390 644.360 1702.710 ;
        RECT 689.640 1702.390 689.900 1702.710 ;
        RECT 644.160 597.030 644.300 1702.390 ;
        RECT 689.700 1701.940 689.840 1702.390 ;
        RECT 690.160 1701.940 690.300 1991.050 ;
        RECT 1908.630 1783.795 1908.910 1784.165 ;
        RECT 869.560 1702.990 870.160 1703.130 ;
        RECT 869.560 1702.710 869.700 1702.990 ;
        RECT 785.840 1702.370 787.360 1702.450 ;
        RECT 869.500 1702.390 869.760 1702.710 ;
        RECT 785.780 1702.310 787.420 1702.370 ;
        RECT 785.780 1702.050 786.040 1702.310 ;
        RECT 787.160 1702.050 787.420 1702.310 ;
        RECT 691.480 1701.940 691.740 1702.030 ;
        RECT 689.700 1701.800 691.740 1701.940 ;
        RECT 724.600 1701.885 724.860 1702.030 ;
        RECT 738.860 1701.885 739.120 1702.030 ;
        RECT 691.480 1701.710 691.740 1701.800 ;
        RECT 724.590 1701.515 724.870 1701.885 ;
        RECT 738.850 1701.515 739.130 1701.885 ;
        RECT 870.020 1701.690 870.160 1702.990 ;
        RECT 966.100 1702.390 966.360 1702.710 ;
        RECT 1279.820 1702.390 1280.080 1702.710 ;
        RECT 1303.740 1702.450 1304.000 1702.710 ;
        RECT 1303.740 1702.390 1304.400 1702.450 ;
        RECT 1400.340 1702.390 1400.600 1702.710 ;
        RECT 917.340 1702.050 917.600 1702.370 ;
        RECT 917.400 1701.690 917.540 1702.050 ;
        RECT 966.160 1702.030 966.300 1702.390 ;
        RECT 1076.040 1702.050 1076.300 1702.370 ;
        RECT 1200.240 1702.050 1200.500 1702.370 ;
        RECT 966.100 1701.710 966.360 1702.030 ;
        RECT 1076.100 1701.770 1076.240 1702.050 ;
        RECT 1124.800 1701.770 1125.060 1702.030 ;
        RECT 1152.400 1701.885 1152.660 1702.030 ;
        RECT 1200.300 1701.885 1200.440 1702.050 ;
        RECT 1279.880 1702.030 1280.020 1702.390 ;
        RECT 1303.800 1702.310 1304.400 1702.390 ;
        RECT 1304.260 1702.030 1304.400 1702.310 ;
        RECT 1076.100 1701.690 1077.160 1701.770 ;
        RECT 1124.400 1701.710 1125.060 1701.770 ;
        RECT 1124.400 1701.690 1125.000 1701.710 ;
        RECT 869.960 1701.370 870.220 1701.690 ;
        RECT 917.340 1701.370 917.600 1701.690 ;
        RECT 1076.100 1701.630 1077.220 1701.690 ;
        RECT 1076.960 1701.370 1077.220 1701.630 ;
        RECT 1124.340 1701.630 1125.000 1701.690 ;
        RECT 1124.340 1701.370 1124.600 1701.630 ;
        RECT 1152.390 1701.515 1152.670 1701.885 ;
        RECT 1200.230 1701.515 1200.510 1701.885 ;
        RECT 1279.820 1701.710 1280.080 1702.030 ;
        RECT 1304.200 1701.710 1304.460 1702.030 ;
        RECT 1400.400 1701.770 1400.540 1702.390 ;
        RECT 1565.540 1702.370 1566.140 1702.450 ;
        RECT 1641.840 1702.390 1642.100 1702.710 ;
        RECT 1642.760 1702.390 1643.020 1702.710 ;
        RECT 1751.320 1702.565 1751.580 1702.710 ;
        RECT 1401.260 1702.050 1401.520 1702.370 ;
        RECT 1565.480 1702.310 1566.140 1702.370 ;
        RECT 1565.480 1702.050 1565.740 1702.310 ;
        RECT 1401.320 1701.770 1401.460 1702.050 ;
        RECT 1566.000 1702.030 1566.140 1702.310 ;
        RECT 1400.400 1701.630 1401.460 1701.770 ;
        RECT 1462.440 1701.770 1462.700 1702.030 ;
        RECT 1462.900 1701.770 1463.160 1702.030 ;
        RECT 1462.440 1701.710 1463.160 1701.770 ;
        RECT 1565.940 1701.710 1566.200 1702.030 ;
        RECT 1594.000 1701.710 1594.260 1702.030 ;
        RECT 1462.500 1701.630 1463.100 1701.710 ;
        RECT 1594.060 1701.350 1594.200 1701.710 ;
        RECT 1641.900 1701.350 1642.040 1702.390 ;
        RECT 1642.820 1702.030 1642.960 1702.390 ;
        RECT 1690.590 1702.195 1690.870 1702.565 ;
        RECT 1709.450 1702.195 1709.730 1702.565 ;
        RECT 1751.310 1702.195 1751.590 1702.565 ;
        RECT 1786.730 1702.195 1787.010 1702.565 ;
        RECT 1690.600 1702.050 1690.860 1702.195 ;
        RECT 1709.460 1702.050 1709.720 1702.195 ;
        RECT 1786.800 1702.030 1786.940 1702.195 ;
        RECT 1835.040 1702.050 1835.300 1702.370 ;
        RECT 1848.370 1702.195 1848.650 1702.565 ;
        RECT 1849.750 1702.195 1850.030 1702.565 ;
        RECT 1848.380 1702.050 1848.640 1702.195 ;
        RECT 1642.760 1701.710 1643.020 1702.030 ;
        RECT 1786.740 1701.710 1787.000 1702.030 ;
        RECT 1835.100 1701.885 1835.240 1702.050 ;
        RECT 1849.820 1702.030 1849.960 1702.195 ;
        RECT 1787.190 1701.515 1787.470 1701.885 ;
        RECT 1835.030 1701.515 1835.310 1701.885 ;
        RECT 1849.760 1701.710 1850.020 1702.030 ;
        RECT 1883.800 1701.885 1884.060 1702.030 ;
        RECT 1908.700 1701.885 1908.840 1783.795 ;
        RECT 1883.790 1701.515 1884.070 1701.885 ;
        RECT 1908.630 1701.515 1908.910 1701.885 ;
        RECT 1787.200 1701.370 1787.460 1701.515 ;
        RECT 1594.000 1701.030 1594.260 1701.350 ;
        RECT 1641.840 1701.030 1642.100 1701.350 ;
        RECT 787.390 600.170 787.670 604.000 ;
        RECT 786.760 600.030 787.670 600.170 ;
        RECT 644.100 596.710 644.360 597.030 ;
        RECT 697.000 596.710 697.260 597.030 ;
        RECT 697.060 593.290 697.200 596.710 ;
        RECT 786.760 593.290 786.900 600.030 ;
        RECT 787.390 600.000 787.670 600.030 ;
        RECT 693.780 592.970 694.040 593.290 ;
        RECT 697.000 592.970 697.260 593.290 ;
        RECT 786.700 592.970 786.960 593.290 ;
        RECT 693.840 592.690 693.980 592.970 ;
        RECT 693.380 592.550 693.980 592.690 ;
        RECT 693.380 47.930 693.520 592.550 ;
        RECT 228.720 47.610 228.980 47.930 ;
        RECT 693.320 47.610 693.580 47.930 ;
        RECT 228.780 2.400 228.920 47.610 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 1908.630 1783.840 1908.910 1784.120 ;
        RECT 724.590 1701.560 724.870 1701.840 ;
        RECT 738.850 1701.560 739.130 1701.840 ;
        RECT 1152.390 1701.560 1152.670 1701.840 ;
        RECT 1200.230 1701.560 1200.510 1701.840 ;
        RECT 1690.590 1702.240 1690.870 1702.520 ;
        RECT 1709.450 1702.240 1709.730 1702.520 ;
        RECT 1751.310 1702.240 1751.590 1702.520 ;
        RECT 1786.730 1702.240 1787.010 1702.520 ;
        RECT 1848.370 1702.240 1848.650 1702.520 ;
        RECT 1849.750 1702.240 1850.030 1702.520 ;
        RECT 1787.190 1701.560 1787.470 1701.840 ;
        RECT 1835.030 1701.560 1835.310 1701.840 ;
        RECT 1883.790 1701.560 1884.070 1701.840 ;
        RECT 1908.630 1701.560 1908.910 1701.840 ;
      LAYER met3 ;
        RECT 1920.000 1786.760 1924.000 1787.360 ;
        RECT 1908.605 1784.130 1908.935 1784.145 ;
        RECT 1920.350 1784.130 1920.650 1786.760 ;
        RECT 1908.605 1783.830 1920.650 1784.130 ;
        RECT 1908.605 1783.815 1908.935 1783.830 ;
        RECT 1690.565 1702.530 1690.895 1702.545 ;
        RECT 1709.425 1702.530 1709.755 1702.545 ;
        RECT 1690.565 1702.230 1709.755 1702.530 ;
        RECT 1690.565 1702.215 1690.895 1702.230 ;
        RECT 1709.425 1702.215 1709.755 1702.230 ;
        RECT 1751.285 1702.530 1751.615 1702.545 ;
        RECT 1786.705 1702.530 1787.035 1702.545 ;
        RECT 1751.285 1702.230 1787.035 1702.530 ;
        RECT 1751.285 1702.215 1751.615 1702.230 ;
        RECT 1786.705 1702.215 1787.035 1702.230 ;
        RECT 1848.345 1702.530 1848.675 1702.545 ;
        RECT 1849.725 1702.530 1850.055 1702.545 ;
        RECT 1848.345 1702.230 1850.055 1702.530 ;
        RECT 1848.345 1702.215 1848.675 1702.230 ;
        RECT 1849.725 1702.215 1850.055 1702.230 ;
        RECT 724.565 1701.850 724.895 1701.865 ;
        RECT 738.825 1701.850 739.155 1701.865 ;
        RECT 724.565 1701.550 739.155 1701.850 ;
        RECT 724.565 1701.535 724.895 1701.550 ;
        RECT 738.825 1701.535 739.155 1701.550 ;
        RECT 1152.365 1701.850 1152.695 1701.865 ;
        RECT 1200.205 1701.850 1200.535 1701.865 ;
        RECT 1152.365 1701.550 1200.535 1701.850 ;
        RECT 1152.365 1701.535 1152.695 1701.550 ;
        RECT 1200.205 1701.535 1200.535 1701.550 ;
        RECT 1787.165 1701.850 1787.495 1701.865 ;
        RECT 1835.005 1701.850 1835.335 1701.865 ;
        RECT 1787.165 1701.550 1835.335 1701.850 ;
        RECT 1787.165 1701.535 1787.495 1701.550 ;
        RECT 1835.005 1701.535 1835.335 1701.550 ;
        RECT 1883.765 1701.850 1884.095 1701.865 ;
        RECT 1908.605 1701.850 1908.935 1701.865 ;
        RECT 1883.765 1701.550 1908.935 1701.850 ;
        RECT 1883.765 1701.535 1884.095 1701.550 ;
        RECT 1908.605 1701.535 1908.935 1701.550 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 690.530 497.120 690.850 497.380 ;
        RECT 690.620 496.700 690.760 497.120 ;
        RECT 690.530 496.440 690.850 496.700 ;
        RECT 689.150 355.540 689.470 355.600 ;
        RECT 690.530 355.540 690.850 355.600 ;
        RECT 689.150 355.400 690.850 355.540 ;
        RECT 689.150 355.340 689.470 355.400 ;
        RECT 690.530 355.340 690.850 355.400 ;
        RECT 690.530 276.320 690.850 276.380 ;
        RECT 691.450 276.320 691.770 276.380 ;
        RECT 690.530 276.180 691.770 276.320 ;
        RECT 690.530 276.120 690.850 276.180 ;
        RECT 691.450 276.120 691.770 276.180 ;
        RECT 690.530 159.360 690.850 159.420 ;
        RECT 691.450 159.360 691.770 159.420 ;
        RECT 690.530 159.220 691.770 159.360 ;
        RECT 690.530 159.160 690.850 159.220 ;
        RECT 691.450 159.160 691.770 159.220 ;
        RECT 690.530 131.480 690.850 131.540 ;
        RECT 691.450 131.480 691.770 131.540 ;
        RECT 690.530 131.340 691.770 131.480 ;
        RECT 690.530 131.280 690.850 131.340 ;
        RECT 691.450 131.280 691.770 131.340 ;
        RECT 689.610 107.000 689.930 107.060 ;
        RECT 690.530 107.000 690.850 107.060 ;
        RECT 689.610 106.860 690.850 107.000 ;
        RECT 689.610 106.800 689.930 106.860 ;
        RECT 690.530 106.800 690.850 106.860 ;
        RECT 689.610 83.200 689.930 83.260 ;
        RECT 690.070 83.200 690.390 83.260 ;
        RECT 689.610 83.060 690.390 83.200 ;
        RECT 689.610 83.000 689.930 83.060 ;
        RECT 690.070 83.000 690.390 83.060 ;
        RECT 50.210 45.120 50.530 45.180 ;
        RECT 690.070 45.120 690.390 45.180 ;
        RECT 50.210 44.980 690.390 45.120 ;
        RECT 50.210 44.920 50.530 44.980 ;
        RECT 690.070 44.920 690.390 44.980 ;
      LAYER via ;
        RECT 690.560 497.120 690.820 497.380 ;
        RECT 690.560 496.440 690.820 496.700 ;
        RECT 689.180 355.340 689.440 355.600 ;
        RECT 690.560 355.340 690.820 355.600 ;
        RECT 690.560 276.120 690.820 276.380 ;
        RECT 691.480 276.120 691.740 276.380 ;
        RECT 690.560 159.160 690.820 159.420 ;
        RECT 691.480 159.160 691.740 159.420 ;
        RECT 690.560 131.280 690.820 131.540 ;
        RECT 691.480 131.280 691.740 131.540 ;
        RECT 689.640 106.800 689.900 107.060 ;
        RECT 690.560 106.800 690.820 107.060 ;
        RECT 689.640 83.000 689.900 83.260 ;
        RECT 690.100 83.000 690.360 83.260 ;
        RECT 50.240 44.920 50.500 45.180 ;
        RECT 690.100 44.920 690.360 45.180 ;
      LAYER met2 ;
        RECT 695.850 600.170 696.130 604.000 ;
        RECT 693.380 600.030 696.130 600.170 ;
        RECT 693.380 593.370 693.520 600.030 ;
        RECT 695.850 600.000 696.130 600.030 ;
        RECT 691.540 593.230 693.520 593.370 ;
        RECT 691.540 569.400 691.680 593.230 ;
        RECT 690.620 569.260 691.680 569.400 ;
        RECT 690.620 497.410 690.760 569.260 ;
        RECT 690.560 497.090 690.820 497.410 ;
        RECT 690.560 496.410 690.820 496.730 ;
        RECT 690.620 355.630 690.760 496.410 ;
        RECT 689.180 355.310 689.440 355.630 ;
        RECT 690.560 355.310 690.820 355.630 ;
        RECT 689.240 340.410 689.380 355.310 ;
        RECT 689.240 340.270 690.300 340.410 ;
        RECT 690.160 300.970 690.300 340.270 ;
        RECT 690.160 300.830 691.680 300.970 ;
        RECT 691.540 276.410 691.680 300.830 ;
        RECT 690.560 276.090 690.820 276.410 ;
        RECT 691.480 276.090 691.740 276.410 ;
        RECT 690.620 159.450 690.760 276.090 ;
        RECT 690.560 159.130 690.820 159.450 ;
        RECT 691.480 159.130 691.740 159.450 ;
        RECT 691.540 131.570 691.680 159.130 ;
        RECT 690.560 131.250 690.820 131.570 ;
        RECT 691.480 131.250 691.740 131.570 ;
        RECT 690.620 107.090 690.760 131.250 ;
        RECT 689.640 106.770 689.900 107.090 ;
        RECT 690.560 106.770 690.820 107.090 ;
        RECT 689.700 83.290 689.840 106.770 ;
        RECT 689.640 82.970 689.900 83.290 ;
        RECT 690.100 82.970 690.360 83.290 ;
        RECT 690.160 45.210 690.300 82.970 ;
        RECT 50.240 44.890 50.500 45.210 ;
        RECT 690.100 44.890 690.360 45.210 ;
        RECT 50.300 2.400 50.440 44.890 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 795.410 593.540 795.730 593.600 ;
        RECT 798.170 593.540 798.490 593.600 ;
        RECT 795.410 593.400 798.490 593.540 ;
        RECT 795.410 593.340 795.730 593.400 ;
        RECT 798.170 593.340 798.490 593.400 ;
        RECT 794.950 558.860 795.270 558.920 ;
        RECT 796.790 558.860 797.110 558.920 ;
        RECT 794.950 558.720 797.110 558.860 ;
        RECT 794.950 558.660 795.270 558.720 ;
        RECT 796.790 558.660 797.110 558.720 ;
        RECT 795.410 510.580 795.730 510.640 ;
        RECT 795.870 510.580 796.190 510.640 ;
        RECT 795.410 510.440 796.190 510.580 ;
        RECT 795.410 510.380 795.730 510.440 ;
        RECT 795.870 510.380 796.190 510.440 ;
        RECT 794.490 455.500 794.810 455.560 ;
        RECT 795.410 455.500 795.730 455.560 ;
        RECT 794.490 455.360 795.730 455.500 ;
        RECT 794.490 455.300 794.810 455.360 ;
        RECT 795.410 455.300 795.730 455.360 ;
        RECT 794.490 414.360 794.810 414.420 ;
        RECT 794.950 414.360 795.270 414.420 ;
        RECT 794.490 414.220 795.270 414.360 ;
        RECT 794.490 414.160 794.810 414.220 ;
        RECT 794.950 414.160 795.270 414.220 ;
        RECT 794.950 234.840 795.270 234.900 ;
        RECT 795.870 234.840 796.190 234.900 ;
        RECT 794.950 234.700 796.190 234.840 ;
        RECT 794.950 234.640 795.270 234.700 ;
        RECT 795.870 234.640 796.190 234.700 ;
        RECT 795.870 227.700 796.190 227.760 ;
        RECT 796.790 227.700 797.110 227.760 ;
        RECT 795.870 227.560 797.110 227.700 ;
        RECT 795.870 227.500 796.190 227.560 ;
        RECT 796.790 227.500 797.110 227.560 ;
        RECT 795.870 179.760 796.190 179.820 ;
        RECT 796.790 179.760 797.110 179.820 ;
        RECT 795.870 179.620 797.110 179.760 ;
        RECT 795.870 179.560 796.190 179.620 ;
        RECT 796.790 179.560 797.110 179.620 ;
        RECT 793.570 162.080 793.890 162.140 ;
        RECT 795.870 162.080 796.190 162.140 ;
        RECT 793.570 161.940 796.190 162.080 ;
        RECT 793.570 161.880 793.890 161.940 ;
        RECT 795.870 161.880 796.190 161.940 ;
        RECT 794.950 137.940 795.270 138.000 ;
        RECT 795.870 137.940 796.190 138.000 ;
        RECT 794.950 137.800 796.190 137.940 ;
        RECT 794.950 137.740 795.270 137.800 ;
        RECT 795.870 137.740 796.190 137.800 ;
        RECT 794.950 90.000 795.270 90.060 ;
        RECT 795.870 90.000 796.190 90.060 ;
        RECT 794.950 89.860 796.190 90.000 ;
        RECT 794.950 89.800 795.270 89.860 ;
        RECT 795.870 89.800 796.190 89.860 ;
        RECT 794.950 62.460 795.270 62.520 ;
        RECT 794.580 62.320 795.270 62.460 ;
        RECT 794.580 62.180 794.720 62.320 ;
        RECT 794.950 62.260 795.270 62.320 ;
        RECT 794.490 61.920 794.810 62.180 ;
        RECT 252.610 32.200 252.930 32.260 ;
        RECT 794.490 32.200 794.810 32.260 ;
        RECT 252.610 32.060 794.810 32.200 ;
        RECT 252.610 32.000 252.930 32.060 ;
        RECT 794.490 32.000 794.810 32.060 ;
      LAYER via ;
        RECT 795.440 593.340 795.700 593.600 ;
        RECT 798.200 593.340 798.460 593.600 ;
        RECT 794.980 558.660 795.240 558.920 ;
        RECT 796.820 558.660 797.080 558.920 ;
        RECT 795.440 510.380 795.700 510.640 ;
        RECT 795.900 510.380 796.160 510.640 ;
        RECT 794.520 455.300 794.780 455.560 ;
        RECT 795.440 455.300 795.700 455.560 ;
        RECT 794.520 414.160 794.780 414.420 ;
        RECT 794.980 414.160 795.240 414.420 ;
        RECT 794.980 234.640 795.240 234.900 ;
        RECT 795.900 234.640 796.160 234.900 ;
        RECT 795.900 227.500 796.160 227.760 ;
        RECT 796.820 227.500 797.080 227.760 ;
        RECT 795.900 179.560 796.160 179.820 ;
        RECT 796.820 179.560 797.080 179.820 ;
        RECT 793.600 161.880 793.860 162.140 ;
        RECT 795.900 161.880 796.160 162.140 ;
        RECT 794.980 137.740 795.240 138.000 ;
        RECT 795.900 137.740 796.160 138.000 ;
        RECT 794.980 89.800 795.240 90.060 ;
        RECT 795.900 89.800 796.160 90.060 ;
        RECT 794.980 62.260 795.240 62.520 ;
        RECT 794.520 61.920 794.780 62.180 ;
        RECT 252.640 32.000 252.900 32.260 ;
        RECT 794.520 32.000 794.780 32.260 ;
      LAYER met2 ;
        RECT 799.350 600.170 799.630 604.000 ;
        RECT 798.260 600.030 799.630 600.170 ;
        RECT 798.260 593.630 798.400 600.030 ;
        RECT 799.350 600.000 799.630 600.030 ;
        RECT 795.440 593.310 795.700 593.630 ;
        RECT 798.200 593.310 798.460 593.630 ;
        RECT 795.500 569.570 795.640 593.310 ;
        RECT 795.040 569.430 795.640 569.570 ;
        RECT 795.040 558.950 795.180 569.430 ;
        RECT 794.980 558.630 795.240 558.950 ;
        RECT 796.820 558.630 797.080 558.950 ;
        RECT 796.880 511.205 797.020 558.630 ;
        RECT 795.430 510.835 795.710 511.205 ;
        RECT 796.810 510.835 797.090 511.205 ;
        RECT 795.500 510.670 795.640 510.835 ;
        RECT 795.440 510.350 795.700 510.670 ;
        RECT 795.900 510.350 796.160 510.670 ;
        RECT 795.960 503.610 796.100 510.350 ;
        RECT 795.500 503.470 796.100 503.610 ;
        RECT 795.500 455.590 795.640 503.470 ;
        RECT 794.520 455.270 794.780 455.590 ;
        RECT 795.440 455.270 795.700 455.590 ;
        RECT 794.580 414.450 794.720 455.270 ;
        RECT 794.520 414.130 794.780 414.450 ;
        RECT 794.980 414.130 795.240 414.450 ;
        RECT 795.040 362.170 795.180 414.130 ;
        RECT 795.040 362.030 795.640 362.170 ;
        RECT 795.500 305.050 795.640 362.030 ;
        RECT 795.040 304.910 795.640 305.050 ;
        RECT 795.040 303.690 795.180 304.910 ;
        RECT 795.040 303.550 795.640 303.690 ;
        RECT 795.500 264.250 795.640 303.550 ;
        RECT 795.040 264.110 795.640 264.250 ;
        RECT 795.040 234.930 795.180 264.110 ;
        RECT 794.980 234.610 795.240 234.930 ;
        RECT 795.900 234.610 796.160 234.930 ;
        RECT 795.960 227.790 796.100 234.610 ;
        RECT 795.900 227.470 796.160 227.790 ;
        RECT 796.820 227.470 797.080 227.790 ;
        RECT 796.880 179.850 797.020 227.470 ;
        RECT 795.900 179.530 796.160 179.850 ;
        RECT 796.820 179.530 797.080 179.850 ;
        RECT 795.960 162.170 796.100 179.530 ;
        RECT 793.600 161.850 793.860 162.170 ;
        RECT 795.900 161.850 796.160 162.170 ;
        RECT 793.660 138.565 793.800 161.850 ;
        RECT 793.590 138.195 793.870 138.565 ;
        RECT 794.970 138.195 795.250 138.565 ;
        RECT 795.040 138.030 795.180 138.195 ;
        RECT 794.980 137.710 795.240 138.030 ;
        RECT 795.900 137.710 796.160 138.030 ;
        RECT 795.960 90.090 796.100 137.710 ;
        RECT 794.980 89.770 795.240 90.090 ;
        RECT 795.900 89.770 796.160 90.090 ;
        RECT 795.040 62.550 795.180 89.770 ;
        RECT 794.980 62.230 795.240 62.550 ;
        RECT 794.520 61.890 794.780 62.210 ;
        RECT 794.580 32.290 794.720 61.890 ;
        RECT 252.640 31.970 252.900 32.290 ;
        RECT 794.520 31.970 794.780 32.290 ;
        RECT 252.700 2.400 252.840 31.970 ;
        RECT 252.490 -4.800 253.050 2.400 ;
      LAYER via2 ;
        RECT 795.430 510.880 795.710 511.160 ;
        RECT 796.810 510.880 797.090 511.160 ;
        RECT 793.590 138.240 793.870 138.520 ;
        RECT 794.970 138.240 795.250 138.520 ;
      LAYER met3 ;
        RECT 795.405 511.170 795.735 511.185 ;
        RECT 796.785 511.170 797.115 511.185 ;
        RECT 795.405 510.870 797.115 511.170 ;
        RECT 795.405 510.855 795.735 510.870 ;
        RECT 796.785 510.855 797.115 510.870 ;
        RECT 793.565 138.530 793.895 138.545 ;
        RECT 794.945 138.530 795.275 138.545 ;
        RECT 793.565 138.230 795.275 138.530 ;
        RECT 793.565 138.215 793.895 138.230 ;
        RECT 794.945 138.215 795.275 138.230 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 32.540 270.410 32.600 ;
        RECT 807.370 32.540 807.690 32.600 ;
        RECT 270.090 32.400 807.690 32.540 ;
        RECT 270.090 32.340 270.410 32.400 ;
        RECT 807.370 32.340 807.690 32.400 ;
      LAYER via ;
        RECT 270.120 32.340 270.380 32.600 ;
        RECT 807.400 32.340 807.660 32.600 ;
      LAYER met2 ;
        RECT 808.550 600.170 808.830 604.000 ;
        RECT 807.460 600.030 808.830 600.170 ;
        RECT 807.460 32.630 807.600 600.030 ;
        RECT 808.550 600.000 808.830 600.030 ;
        RECT 270.120 32.310 270.380 32.630 ;
        RECT 807.400 32.310 807.660 32.630 ;
        RECT 270.180 2.400 270.320 32.310 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 814.730 497.120 815.050 497.380 ;
        RECT 814.820 496.700 814.960 497.120 ;
        RECT 814.730 496.440 815.050 496.700 ;
        RECT 814.730 351.940 815.050 352.200 ;
        RECT 814.820 351.520 814.960 351.940 ;
        RECT 814.730 351.260 815.050 351.520 ;
        RECT 815.190 282.780 815.510 282.840 ;
        RECT 816.110 282.780 816.430 282.840 ;
        RECT 815.190 282.640 816.430 282.780 ;
        RECT 815.190 282.580 815.510 282.640 ;
        RECT 816.110 282.580 816.430 282.640 ;
        RECT 814.730 234.840 815.050 234.900 ;
        RECT 816.110 234.840 816.430 234.900 ;
        RECT 814.730 234.700 816.430 234.840 ;
        RECT 814.730 234.640 815.050 234.700 ;
        RECT 816.110 234.640 816.430 234.700 ;
        RECT 814.270 96.460 814.590 96.520 ;
        RECT 814.730 96.460 815.050 96.520 ;
        RECT 814.270 96.320 815.050 96.460 ;
        RECT 814.270 96.260 814.590 96.320 ;
        RECT 814.730 96.260 815.050 96.320 ;
        RECT 288.030 32.880 288.350 32.940 ;
        RECT 814.270 32.880 814.590 32.940 ;
        RECT 288.030 32.740 814.590 32.880 ;
        RECT 288.030 32.680 288.350 32.740 ;
        RECT 814.270 32.680 814.590 32.740 ;
      LAYER via ;
        RECT 814.760 497.120 815.020 497.380 ;
        RECT 814.760 496.440 815.020 496.700 ;
        RECT 814.760 351.940 815.020 352.200 ;
        RECT 814.760 351.260 815.020 351.520 ;
        RECT 815.220 282.580 815.480 282.840 ;
        RECT 816.140 282.580 816.400 282.840 ;
        RECT 814.760 234.640 815.020 234.900 ;
        RECT 816.140 234.640 816.400 234.900 ;
        RECT 814.300 96.260 814.560 96.520 ;
        RECT 814.760 96.260 815.020 96.520 ;
        RECT 288.060 32.680 288.320 32.940 ;
        RECT 814.300 32.680 814.560 32.940 ;
      LAYER met2 ;
        RECT 817.750 600.170 818.030 604.000 ;
        RECT 816.660 600.030 818.030 600.170 ;
        RECT 816.660 596.770 816.800 600.030 ;
        RECT 817.750 600.000 818.030 600.030 ;
        RECT 814.820 596.630 816.800 596.770 ;
        RECT 814.820 497.410 814.960 596.630 ;
        RECT 814.760 497.090 815.020 497.410 ;
        RECT 814.760 496.410 815.020 496.730 ;
        RECT 814.820 352.230 814.960 496.410 ;
        RECT 814.760 351.910 815.020 352.230 ;
        RECT 814.760 351.230 815.020 351.550 ;
        RECT 814.820 312.530 814.960 351.230 ;
        RECT 814.360 312.390 814.960 312.530 ;
        RECT 814.360 283.405 814.500 312.390 ;
        RECT 814.290 283.035 814.570 283.405 ;
        RECT 815.210 283.035 815.490 283.405 ;
        RECT 815.280 282.870 815.420 283.035 ;
        RECT 815.220 282.550 815.480 282.870 ;
        RECT 816.140 282.550 816.400 282.870 ;
        RECT 816.200 234.930 816.340 282.550 ;
        RECT 814.760 234.610 815.020 234.930 ;
        RECT 816.140 234.610 816.400 234.930 ;
        RECT 814.820 96.550 814.960 234.610 ;
        RECT 814.300 96.230 814.560 96.550 ;
        RECT 814.760 96.230 815.020 96.550 ;
        RECT 814.360 32.970 814.500 96.230 ;
        RECT 288.060 32.650 288.320 32.970 ;
        RECT 814.300 32.650 814.560 32.970 ;
        RECT 288.120 2.400 288.260 32.650 ;
        RECT 287.910 -4.800 288.470 2.400 ;
      LAYER via2 ;
        RECT 814.290 283.080 814.570 283.360 ;
        RECT 815.210 283.080 815.490 283.360 ;
      LAYER met3 ;
        RECT 814.265 283.370 814.595 283.385 ;
        RECT 815.185 283.370 815.515 283.385 ;
        RECT 814.265 283.070 815.515 283.370 ;
        RECT 814.265 283.055 814.595 283.070 ;
        RECT 815.185 283.055 815.515 283.070 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 823.010 593.540 823.330 593.600 ;
        RECT 825.770 593.540 826.090 593.600 ;
        RECT 823.010 593.400 826.090 593.540 ;
        RECT 823.010 593.340 823.330 593.400 ;
        RECT 825.770 593.340 826.090 593.400 ;
        RECT 822.550 410.420 822.870 410.680 ;
        RECT 822.640 410.280 822.780 410.420 ;
        RECT 823.010 410.280 823.330 410.340 ;
        RECT 822.640 410.140 823.330 410.280 ;
        RECT 823.010 410.080 823.330 410.140 ;
        RECT 822.550 331.060 822.870 331.120 ;
        RECT 823.010 331.060 823.330 331.120 ;
        RECT 822.550 330.920 823.330 331.060 ;
        RECT 822.550 330.860 822.870 330.920 ;
        RECT 823.010 330.860 823.330 330.920 ;
        RECT 823.010 283.120 823.330 283.180 ;
        RECT 823.930 283.120 824.250 283.180 ;
        RECT 823.010 282.980 824.250 283.120 ;
        RECT 823.010 282.920 823.330 282.980 ;
        RECT 823.930 282.920 824.250 282.980 ;
        RECT 823.010 241.640 823.330 241.700 ;
        RECT 823.930 241.640 824.250 241.700 ;
        RECT 823.010 241.500 824.250 241.640 ;
        RECT 823.010 241.440 823.330 241.500 ;
        RECT 823.930 241.440 824.250 241.500 ;
        RECT 822.550 193.020 822.870 193.080 ;
        RECT 823.010 193.020 823.330 193.080 ;
        RECT 822.550 192.880 823.330 193.020 ;
        RECT 822.550 192.820 822.870 192.880 ;
        RECT 823.010 192.820 823.330 192.880 ;
        RECT 821.170 137.940 821.490 138.000 ;
        RECT 822.550 137.940 822.870 138.000 ;
        RECT 821.170 137.800 822.870 137.940 ;
        RECT 821.170 137.740 821.490 137.800 ;
        RECT 822.550 137.740 822.870 137.800 ;
        RECT 821.170 48.520 821.490 48.580 ;
        RECT 822.090 48.520 822.410 48.580 ;
        RECT 821.170 48.380 822.410 48.520 ;
        RECT 821.170 48.320 821.490 48.380 ;
        RECT 822.090 48.320 822.410 48.380 ;
        RECT 305.970 33.220 306.290 33.280 ;
        RECT 822.090 33.220 822.410 33.280 ;
        RECT 305.970 33.080 822.410 33.220 ;
        RECT 305.970 33.020 306.290 33.080 ;
        RECT 822.090 33.020 822.410 33.080 ;
      LAYER via ;
        RECT 823.040 593.340 823.300 593.600 ;
        RECT 825.800 593.340 826.060 593.600 ;
        RECT 822.580 410.420 822.840 410.680 ;
        RECT 823.040 410.080 823.300 410.340 ;
        RECT 822.580 330.860 822.840 331.120 ;
        RECT 823.040 330.860 823.300 331.120 ;
        RECT 823.040 282.920 823.300 283.180 ;
        RECT 823.960 282.920 824.220 283.180 ;
        RECT 823.040 241.440 823.300 241.700 ;
        RECT 823.960 241.440 824.220 241.700 ;
        RECT 822.580 192.820 822.840 193.080 ;
        RECT 823.040 192.820 823.300 193.080 ;
        RECT 821.200 137.740 821.460 138.000 ;
        RECT 822.580 137.740 822.840 138.000 ;
        RECT 821.200 48.320 821.460 48.580 ;
        RECT 822.120 48.320 822.380 48.580 ;
        RECT 306.000 33.020 306.260 33.280 ;
        RECT 822.120 33.020 822.380 33.280 ;
      LAYER met2 ;
        RECT 826.950 600.170 827.230 604.000 ;
        RECT 825.860 600.030 827.230 600.170 ;
        RECT 825.860 593.630 826.000 600.030 ;
        RECT 826.950 600.000 827.230 600.030 ;
        RECT 823.040 593.310 823.300 593.630 ;
        RECT 825.800 593.310 826.060 593.630 ;
        RECT 823.100 569.570 823.240 593.310 ;
        RECT 822.640 569.430 823.240 569.570 ;
        RECT 822.640 410.710 822.780 569.430 ;
        RECT 822.580 410.390 822.840 410.710 ;
        RECT 823.040 410.050 823.300 410.370 ;
        RECT 823.100 386.650 823.240 410.050 ;
        RECT 822.640 386.510 823.240 386.650 ;
        RECT 822.640 385.970 822.780 386.510 ;
        RECT 822.640 385.830 823.240 385.970 ;
        RECT 823.100 339.165 823.240 385.830 ;
        RECT 823.030 338.795 823.310 339.165 ;
        RECT 822.570 338.115 822.850 338.485 ;
        RECT 822.640 331.150 822.780 338.115 ;
        RECT 822.580 330.830 822.840 331.150 ;
        RECT 823.040 330.830 823.300 331.150 ;
        RECT 823.100 283.210 823.240 330.830 ;
        RECT 823.040 282.890 823.300 283.210 ;
        RECT 823.960 282.890 824.220 283.210 ;
        RECT 824.020 241.730 824.160 282.890 ;
        RECT 823.040 241.410 823.300 241.730 ;
        RECT 823.960 241.410 824.220 241.730 ;
        RECT 823.100 207.925 823.240 241.410 ;
        RECT 823.030 207.555 823.310 207.925 ;
        RECT 822.570 193.275 822.850 193.645 ;
        RECT 822.640 193.110 822.780 193.275 ;
        RECT 822.580 192.790 822.840 193.110 ;
        RECT 823.040 192.790 823.300 193.110 ;
        RECT 823.100 145.250 823.240 192.790 ;
        RECT 822.640 145.110 823.240 145.250 ;
        RECT 822.640 138.030 822.780 145.110 ;
        RECT 821.200 137.710 821.460 138.030 ;
        RECT 822.580 137.710 822.840 138.030 ;
        RECT 821.260 48.610 821.400 137.710 ;
        RECT 821.200 48.290 821.460 48.610 ;
        RECT 822.120 48.290 822.380 48.610 ;
        RECT 822.180 33.310 822.320 48.290 ;
        RECT 306.000 32.990 306.260 33.310 ;
        RECT 822.120 32.990 822.380 33.310 ;
        RECT 306.060 2.400 306.200 32.990 ;
        RECT 305.850 -4.800 306.410 2.400 ;
      LAYER via2 ;
        RECT 823.030 338.840 823.310 339.120 ;
        RECT 822.570 338.160 822.850 338.440 ;
        RECT 823.030 207.600 823.310 207.880 ;
        RECT 822.570 193.320 822.850 193.600 ;
      LAYER met3 ;
        RECT 823.005 339.130 823.335 339.145 ;
        RECT 821.870 338.830 823.335 339.130 ;
        RECT 821.870 338.450 822.170 338.830 ;
        RECT 823.005 338.815 823.335 338.830 ;
        RECT 822.545 338.450 822.875 338.465 ;
        RECT 821.870 338.150 822.875 338.450 ;
        RECT 822.545 338.135 822.875 338.150 ;
        RECT 823.005 207.900 823.335 207.905 ;
        RECT 822.750 207.890 823.335 207.900 ;
        RECT 822.550 207.590 823.335 207.890 ;
        RECT 822.750 207.580 823.335 207.590 ;
        RECT 823.005 207.575 823.335 207.580 ;
        RECT 822.545 193.620 822.875 193.625 ;
        RECT 822.545 193.610 823.130 193.620 ;
        RECT 822.545 193.310 823.330 193.610 ;
        RECT 822.545 193.300 823.130 193.310 ;
        RECT 822.545 193.295 822.875 193.300 ;
      LAYER via3 ;
        RECT 822.780 207.580 823.100 207.900 ;
        RECT 822.780 193.300 823.100 193.620 ;
      LAYER met4 ;
        RECT 822.775 207.575 823.105 207.905 ;
        RECT 822.790 193.625 823.090 207.575 ;
        RECT 822.775 193.295 823.105 193.625 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 52.600 324.230 52.660 ;
        RECT 835.430 52.600 835.750 52.660 ;
        RECT 323.910 52.460 835.750 52.600 ;
        RECT 323.910 52.400 324.230 52.460 ;
        RECT 835.430 52.400 835.750 52.460 ;
      LAYER via ;
        RECT 323.940 52.400 324.200 52.660 ;
        RECT 835.460 52.400 835.720 52.660 ;
      LAYER met2 ;
        RECT 836.150 600.170 836.430 604.000 ;
        RECT 835.520 600.030 836.430 600.170 ;
        RECT 835.520 52.690 835.660 600.030 ;
        RECT 836.150 600.000 836.430 600.030 ;
        RECT 323.940 52.370 324.200 52.690 ;
        RECT 835.460 52.370 835.720 52.690 ;
        RECT 324.000 2.400 324.140 52.370 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 842.790 483.040 843.110 483.100 ;
        RECT 843.710 483.040 844.030 483.100 ;
        RECT 842.790 482.900 844.030 483.040 ;
        RECT 842.790 482.840 843.110 482.900 ;
        RECT 843.710 482.840 844.030 482.900 ;
        RECT 842.330 241.640 842.650 241.700 ;
        RECT 842.790 241.640 843.110 241.700 ;
        RECT 842.330 241.500 843.110 241.640 ;
        RECT 842.330 241.440 842.650 241.500 ;
        RECT 842.790 241.440 843.110 241.500 ;
        RECT 841.410 193.020 841.730 193.080 ;
        RECT 842.790 193.020 843.110 193.080 ;
        RECT 841.410 192.880 843.110 193.020 ;
        RECT 841.410 192.820 841.730 192.880 ;
        RECT 842.790 192.820 843.110 192.880 ;
        RECT 341.390 39.680 341.710 39.740 ;
        RECT 841.870 39.680 842.190 39.740 ;
        RECT 341.390 39.540 842.190 39.680 ;
        RECT 341.390 39.480 341.710 39.540 ;
        RECT 841.870 39.480 842.190 39.540 ;
      LAYER via ;
        RECT 842.820 482.840 843.080 483.100 ;
        RECT 843.740 482.840 844.000 483.100 ;
        RECT 842.360 241.440 842.620 241.700 ;
        RECT 842.820 241.440 843.080 241.700 ;
        RECT 841.440 192.820 841.700 193.080 ;
        RECT 842.820 192.820 843.080 193.080 ;
        RECT 341.420 39.480 341.680 39.740 ;
        RECT 841.900 39.480 842.160 39.740 ;
      LAYER met2 ;
        RECT 845.350 600.170 845.630 604.000 ;
        RECT 843.340 600.030 845.630 600.170 ;
        RECT 843.340 583.170 843.480 600.030 ;
        RECT 845.350 600.000 845.630 600.030 ;
        RECT 842.420 583.030 843.480 583.170 ;
        RECT 842.420 497.490 842.560 583.030 ;
        RECT 841.960 497.350 842.560 497.490 ;
        RECT 841.960 496.810 842.100 497.350 ;
        RECT 841.960 496.670 843.020 496.810 ;
        RECT 842.880 483.130 843.020 496.670 ;
        RECT 842.820 482.810 843.080 483.130 ;
        RECT 843.740 482.810 844.000 483.130 ;
        RECT 843.800 434.930 843.940 482.810 ;
        RECT 842.880 434.790 843.940 434.930 ;
        RECT 842.880 351.290 843.020 434.790 ;
        RECT 842.420 351.150 843.020 351.290 ;
        RECT 842.420 303.690 842.560 351.150 ;
        RECT 842.420 303.550 843.020 303.690 ;
        RECT 842.880 241.730 843.020 303.550 ;
        RECT 842.360 241.410 842.620 241.730 ;
        RECT 842.820 241.410 843.080 241.730 ;
        RECT 842.420 207.130 842.560 241.410 ;
        RECT 842.420 206.990 843.020 207.130 ;
        RECT 842.880 193.110 843.020 206.990 ;
        RECT 841.440 192.790 841.700 193.110 ;
        RECT 842.820 192.790 843.080 193.110 ;
        RECT 841.500 158.170 841.640 192.790 ;
        RECT 841.500 158.030 842.560 158.170 ;
        RECT 842.420 110.570 842.560 158.030 ;
        RECT 842.420 110.430 843.020 110.570 ;
        RECT 842.880 62.290 843.020 110.430 ;
        RECT 841.960 62.150 843.020 62.290 ;
        RECT 841.960 39.770 842.100 62.150 ;
        RECT 341.420 39.450 341.680 39.770 ;
        RECT 841.900 39.450 842.160 39.770 ;
        RECT 341.480 2.400 341.620 39.450 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 849.230 583.000 849.550 583.060 ;
        RECT 852.910 583.000 853.230 583.060 ;
        RECT 849.230 582.860 853.230 583.000 ;
        RECT 849.230 582.800 849.550 582.860 ;
        RECT 852.910 582.800 853.230 582.860 ;
        RECT 359.330 52.940 359.650 53.000 ;
        RECT 849.230 52.940 849.550 53.000 ;
        RECT 359.330 52.800 849.550 52.940 ;
        RECT 359.330 52.740 359.650 52.800 ;
        RECT 849.230 52.740 849.550 52.800 ;
      LAYER via ;
        RECT 849.260 582.800 849.520 583.060 ;
        RECT 852.940 582.800 853.200 583.060 ;
        RECT 359.360 52.740 359.620 53.000 ;
        RECT 849.260 52.740 849.520 53.000 ;
      LAYER met2 ;
        RECT 854.550 600.170 854.830 604.000 ;
        RECT 853.000 600.030 854.830 600.170 ;
        RECT 853.000 583.090 853.140 600.030 ;
        RECT 854.550 600.000 854.830 600.030 ;
        RECT 849.260 582.770 849.520 583.090 ;
        RECT 852.940 582.770 853.200 583.090 ;
        RECT 849.320 53.030 849.460 582.770 ;
        RECT 359.360 52.710 359.620 53.030 ;
        RECT 849.260 52.710 849.520 53.030 ;
        RECT 359.420 2.400 359.560 52.710 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 377.270 40.020 377.590 40.080 ;
        RECT 863.030 40.020 863.350 40.080 ;
        RECT 377.270 39.880 863.350 40.020 ;
        RECT 377.270 39.820 377.590 39.880 ;
        RECT 863.030 39.820 863.350 39.880 ;
      LAYER via ;
        RECT 377.300 39.820 377.560 40.080 ;
        RECT 863.060 39.820 863.320 40.080 ;
      LAYER met2 ;
        RECT 863.750 600.170 864.030 604.000 ;
        RECT 863.120 600.030 864.030 600.170 ;
        RECT 863.120 40.110 863.260 600.030 ;
        RECT 863.750 600.000 864.030 600.030 ;
        RECT 377.300 39.790 377.560 40.110 ;
        RECT 863.060 39.790 863.320 40.110 ;
        RECT 377.360 2.400 377.500 39.790 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 53.280 395.530 53.340 ;
        RECT 869.930 53.280 870.250 53.340 ;
        RECT 395.210 53.140 870.250 53.280 ;
        RECT 395.210 53.080 395.530 53.140 ;
        RECT 869.930 53.080 870.250 53.140 ;
      LAYER via ;
        RECT 395.240 53.080 395.500 53.340 ;
        RECT 869.960 53.080 870.220 53.340 ;
      LAYER met2 ;
        RECT 872.950 600.170 873.230 604.000 ;
        RECT 870.480 600.030 873.230 600.170 ;
        RECT 870.480 583.170 870.620 600.030 ;
        RECT 872.950 600.000 873.230 600.030 ;
        RECT 870.020 583.030 870.620 583.170 ;
        RECT 870.020 53.370 870.160 583.030 ;
        RECT 395.240 53.050 395.500 53.370 ;
        RECT 869.960 53.050 870.220 53.370 ;
        RECT 395.300 2.400 395.440 53.050 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.150 40.360 413.470 40.420 ;
        RECT 876.830 40.360 877.150 40.420 ;
        RECT 413.150 40.220 877.150 40.360 ;
        RECT 413.150 40.160 413.470 40.220 ;
        RECT 876.830 40.160 877.150 40.220 ;
      LAYER via ;
        RECT 413.180 40.160 413.440 40.420 ;
        RECT 876.860 40.160 877.120 40.420 ;
      LAYER met2 ;
        RECT 882.150 600.170 882.430 604.000 ;
        RECT 880.140 600.030 882.430 600.170 ;
        RECT 880.140 583.170 880.280 600.030 ;
        RECT 882.150 600.000 882.430 600.030 ;
        RECT 876.920 583.030 880.280 583.170 ;
        RECT 876.920 40.450 877.060 583.030 ;
        RECT 413.180 40.130 413.440 40.450 ;
        RECT 876.860 40.130 877.120 40.450 ;
        RECT 413.240 2.400 413.380 40.130 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 704.330 545.400 704.650 545.660 ;
        RECT 704.420 544.980 704.560 545.400 ;
        RECT 704.330 544.720 704.650 544.980 ;
        RECT 703.870 524.520 704.190 524.580 ;
        RECT 704.330 524.520 704.650 524.580 ;
        RECT 703.870 524.380 704.650 524.520 ;
        RECT 703.870 524.320 704.190 524.380 ;
        RECT 704.330 524.320 704.650 524.380 ;
        RECT 703.870 523.840 704.190 523.900 ;
        RECT 704.790 523.840 705.110 523.900 ;
        RECT 703.870 523.700 705.110 523.840 ;
        RECT 703.870 523.640 704.190 523.700 ;
        RECT 704.790 523.640 705.110 523.700 ;
        RECT 704.330 331.200 704.650 331.460 ;
        RECT 703.870 331.060 704.190 331.120 ;
        RECT 704.420 331.060 704.560 331.200 ;
        RECT 703.870 330.920 704.560 331.060 ;
        RECT 703.870 330.860 704.190 330.920 ;
        RECT 703.870 324.600 704.190 324.660 ;
        RECT 704.330 324.600 704.650 324.660 ;
        RECT 703.870 324.460 704.650 324.600 ;
        RECT 703.870 324.400 704.190 324.460 ;
        RECT 704.330 324.400 704.650 324.460 ;
        RECT 703.410 280.400 703.730 280.460 ;
        RECT 705.250 280.400 705.570 280.460 ;
        RECT 703.410 280.260 705.570 280.400 ;
        RECT 703.410 280.200 703.730 280.260 ;
        RECT 705.250 280.200 705.570 280.260 ;
        RECT 703.410 234.840 703.730 234.900 ;
        RECT 703.870 234.840 704.190 234.900 ;
        RECT 703.410 234.700 704.190 234.840 ;
        RECT 703.410 234.640 703.730 234.700 ;
        RECT 703.870 234.640 704.190 234.700 ;
        RECT 703.410 159.020 703.730 159.080 ;
        RECT 704.330 159.020 704.650 159.080 ;
        RECT 703.410 158.880 704.650 159.020 ;
        RECT 703.410 158.820 703.730 158.880 ;
        RECT 704.330 158.820 704.650 158.880 ;
        RECT 703.410 131.480 703.730 131.540 ;
        RECT 704.790 131.480 705.110 131.540 ;
        RECT 703.410 131.340 705.110 131.480 ;
        RECT 703.410 131.280 703.730 131.340 ;
        RECT 704.790 131.280 705.110 131.340 ;
        RECT 74.130 17.920 74.450 17.980 ;
        RECT 648.210 17.920 648.530 17.980 ;
        RECT 74.130 17.780 648.530 17.920 ;
        RECT 74.130 17.720 74.450 17.780 ;
        RECT 648.210 17.720 648.530 17.780 ;
        RECT 648.210 15.200 648.530 15.260 ;
        RECT 704.790 15.200 705.110 15.260 ;
        RECT 648.210 15.060 705.110 15.200 ;
        RECT 648.210 15.000 648.530 15.060 ;
        RECT 704.790 15.000 705.110 15.060 ;
      LAYER via ;
        RECT 704.360 545.400 704.620 545.660 ;
        RECT 704.360 544.720 704.620 544.980 ;
        RECT 703.900 524.320 704.160 524.580 ;
        RECT 704.360 524.320 704.620 524.580 ;
        RECT 703.900 523.640 704.160 523.900 ;
        RECT 704.820 523.640 705.080 523.900 ;
        RECT 704.360 331.200 704.620 331.460 ;
        RECT 703.900 330.860 704.160 331.120 ;
        RECT 703.900 324.400 704.160 324.660 ;
        RECT 704.360 324.400 704.620 324.660 ;
        RECT 703.440 280.200 703.700 280.460 ;
        RECT 705.280 280.200 705.540 280.460 ;
        RECT 703.440 234.640 703.700 234.900 ;
        RECT 703.900 234.640 704.160 234.900 ;
        RECT 703.440 158.820 703.700 159.080 ;
        RECT 704.360 158.820 704.620 159.080 ;
        RECT 703.440 131.280 703.700 131.540 ;
        RECT 704.820 131.280 705.080 131.540 ;
        RECT 74.160 17.720 74.420 17.980 ;
        RECT 648.240 17.720 648.500 17.980 ;
        RECT 648.240 15.000 648.500 15.260 ;
        RECT 704.820 15.000 705.080 15.260 ;
      LAYER met2 ;
        RECT 707.810 600.170 708.090 604.000 ;
        RECT 706.260 600.030 708.090 600.170 ;
        RECT 706.260 596.770 706.400 600.030 ;
        RECT 707.810 600.000 708.090 600.030 ;
        RECT 704.420 596.630 706.400 596.770 ;
        RECT 704.420 545.690 704.560 596.630 ;
        RECT 704.360 545.370 704.620 545.690 ;
        RECT 704.360 544.690 704.620 545.010 ;
        RECT 704.420 524.610 704.560 544.690 ;
        RECT 703.900 524.290 704.160 524.610 ;
        RECT 704.360 524.290 704.620 524.610 ;
        RECT 703.960 523.930 704.100 524.290 ;
        RECT 703.900 523.610 704.160 523.930 ;
        RECT 704.820 523.610 705.080 523.930 ;
        RECT 704.880 496.130 705.020 523.610 ;
        RECT 704.420 495.990 705.020 496.130 ;
        RECT 704.420 331.490 704.560 495.990 ;
        RECT 704.360 331.170 704.620 331.490 ;
        RECT 703.900 330.830 704.160 331.150 ;
        RECT 703.960 324.690 704.100 330.830 ;
        RECT 703.900 324.370 704.160 324.690 ;
        RECT 704.360 324.370 704.620 324.690 ;
        RECT 704.420 324.205 704.560 324.370 ;
        RECT 704.350 323.835 704.630 324.205 ;
        RECT 705.270 323.835 705.550 324.205 ;
        RECT 705.340 280.490 705.480 323.835 ;
        RECT 703.440 280.170 703.700 280.490 ;
        RECT 705.280 280.170 705.540 280.490 ;
        RECT 703.500 234.930 703.640 280.170 ;
        RECT 703.440 234.610 703.700 234.930 ;
        RECT 703.900 234.610 704.160 234.930 ;
        RECT 703.960 206.450 704.100 234.610 ;
        RECT 703.960 206.310 704.560 206.450 ;
        RECT 704.420 159.110 704.560 206.310 ;
        RECT 703.440 158.790 703.700 159.110 ;
        RECT 704.360 158.790 704.620 159.110 ;
        RECT 703.500 131.570 703.640 158.790 ;
        RECT 703.440 131.250 703.700 131.570 ;
        RECT 704.820 131.250 705.080 131.570 ;
        RECT 74.160 17.690 74.420 18.010 ;
        RECT 648.240 17.690 648.500 18.010 ;
        RECT 74.220 2.400 74.360 17.690 ;
        RECT 648.300 15.290 648.440 17.690 ;
        RECT 704.880 15.290 705.020 131.250 ;
        RECT 648.240 14.970 648.500 15.290 ;
        RECT 704.820 14.970 705.080 15.290 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 704.350 323.880 704.630 324.160 ;
        RECT 705.270 323.880 705.550 324.160 ;
      LAYER met3 ;
        RECT 704.325 324.170 704.655 324.185 ;
        RECT 705.245 324.170 705.575 324.185 ;
        RECT 704.325 323.870 705.575 324.170 ;
        RECT 704.325 323.855 704.655 323.870 ;
        RECT 705.245 323.855 705.575 323.870 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.310 53.620 434.630 53.680 ;
        RECT 890.630 53.620 890.950 53.680 ;
        RECT 434.310 53.480 890.950 53.620 ;
        RECT 434.310 53.420 434.630 53.480 ;
        RECT 890.630 53.420 890.950 53.480 ;
        RECT 430.630 16.900 430.950 16.960 ;
        RECT 434.310 16.900 434.630 16.960 ;
        RECT 430.630 16.760 434.630 16.900 ;
        RECT 430.630 16.700 430.950 16.760 ;
        RECT 434.310 16.700 434.630 16.760 ;
      LAYER via ;
        RECT 434.340 53.420 434.600 53.680 ;
        RECT 890.660 53.420 890.920 53.680 ;
        RECT 430.660 16.700 430.920 16.960 ;
        RECT 434.340 16.700 434.600 16.960 ;
      LAYER met2 ;
        RECT 891.350 600.170 891.630 604.000 ;
        RECT 890.720 600.030 891.630 600.170 ;
        RECT 890.720 53.710 890.860 600.030 ;
        RECT 891.350 600.000 891.630 600.030 ;
        RECT 434.340 53.390 434.600 53.710 ;
        RECT 890.660 53.390 890.920 53.710 ;
        RECT 434.400 16.990 434.540 53.390 ;
        RECT 430.660 16.670 430.920 16.990 ;
        RECT 434.340 16.670 434.600 16.990 ;
        RECT 430.720 2.400 430.860 16.670 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 40.700 448.890 40.760 ;
        RECT 897.990 40.700 898.310 40.760 ;
        RECT 448.570 40.560 898.310 40.700 ;
        RECT 448.570 40.500 448.890 40.560 ;
        RECT 897.990 40.500 898.310 40.560 ;
      LAYER via ;
        RECT 448.600 40.500 448.860 40.760 ;
        RECT 898.020 40.500 898.280 40.760 ;
      LAYER met2 ;
        RECT 900.550 600.170 900.830 604.000 ;
        RECT 898.080 600.030 900.830 600.170 ;
        RECT 898.080 40.790 898.220 600.030 ;
        RECT 900.550 600.000 900.830 600.030 ;
        RECT 448.600 40.470 448.860 40.790 ;
        RECT 898.020 40.470 898.280 40.790 ;
        RECT 448.660 2.400 448.800 40.470 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 903.970 386.480 904.290 386.540 ;
        RECT 904.890 386.480 905.210 386.540 ;
        RECT 903.970 386.340 905.210 386.480 ;
        RECT 903.970 386.280 904.290 386.340 ;
        RECT 904.890 386.280 905.210 386.340 ;
        RECT 904.430 303.520 904.750 303.580 ;
        RECT 905.350 303.520 905.670 303.580 ;
        RECT 904.430 303.380 905.670 303.520 ;
        RECT 904.430 303.320 904.750 303.380 ;
        RECT 905.350 303.320 905.670 303.380 ;
        RECT 904.430 289.580 904.750 289.640 ;
        RECT 905.350 289.580 905.670 289.640 ;
        RECT 904.430 289.440 905.670 289.580 ;
        RECT 904.430 289.380 904.750 289.440 ;
        RECT 905.350 289.380 905.670 289.440 ;
        RECT 863.030 21.320 863.350 21.380 ;
        RECT 904.430 21.320 904.750 21.380 ;
        RECT 863.030 21.180 904.750 21.320 ;
        RECT 863.030 21.120 863.350 21.180 ;
        RECT 904.430 21.120 904.750 21.180 ;
        RECT 466.510 20.640 466.830 20.700 ;
        RECT 469.270 20.640 469.590 20.700 ;
        RECT 466.510 20.500 469.590 20.640 ;
        RECT 466.510 20.440 466.830 20.500 ;
        RECT 469.270 20.440 469.590 20.500 ;
        RECT 517.110 20.640 517.430 20.700 ;
        RECT 565.870 20.640 566.190 20.700 ;
        RECT 517.110 20.500 566.190 20.640 ;
        RECT 517.110 20.440 517.430 20.500 ;
        RECT 565.870 20.440 566.190 20.500 ;
        RECT 613.710 20.640 614.030 20.700 ;
        RECT 665.690 20.640 666.010 20.700 ;
        RECT 613.710 20.500 666.010 20.640 ;
        RECT 613.710 20.440 614.030 20.500 ;
        RECT 665.690 20.440 666.010 20.500 ;
        RECT 810.590 19.620 810.910 19.680 ;
        RECT 862.570 19.620 862.890 19.680 ;
        RECT 810.590 19.480 862.890 19.620 ;
        RECT 810.590 19.420 810.910 19.480 ;
        RECT 862.570 19.420 862.890 19.480 ;
        RECT 810.590 17.920 810.910 17.980 ;
        RECT 714.080 17.780 810.910 17.920 ;
        RECT 665.690 17.580 666.010 17.640 ;
        RECT 714.080 17.580 714.220 17.780 ;
        RECT 810.590 17.720 810.910 17.780 ;
        RECT 665.690 17.440 714.220 17.580 ;
        RECT 665.690 17.380 666.010 17.440 ;
        RECT 469.270 16.560 469.590 16.620 ;
        RECT 517.110 16.560 517.430 16.620 ;
        RECT 469.270 16.420 517.430 16.560 ;
        RECT 469.270 16.360 469.590 16.420 ;
        RECT 517.110 16.360 517.430 16.420 ;
        RECT 565.870 15.200 566.190 15.260 ;
        RECT 613.710 15.200 614.030 15.260 ;
        RECT 565.870 15.060 614.030 15.200 ;
        RECT 565.870 15.000 566.190 15.060 ;
        RECT 613.710 15.000 614.030 15.060 ;
      LAYER via ;
        RECT 904.000 386.280 904.260 386.540 ;
        RECT 904.920 386.280 905.180 386.540 ;
        RECT 904.460 303.320 904.720 303.580 ;
        RECT 905.380 303.320 905.640 303.580 ;
        RECT 904.460 289.380 904.720 289.640 ;
        RECT 905.380 289.380 905.640 289.640 ;
        RECT 863.060 21.120 863.320 21.380 ;
        RECT 904.460 21.120 904.720 21.380 ;
        RECT 466.540 20.440 466.800 20.700 ;
        RECT 469.300 20.440 469.560 20.700 ;
        RECT 517.140 20.440 517.400 20.700 ;
        RECT 565.900 20.440 566.160 20.700 ;
        RECT 613.740 20.440 614.000 20.700 ;
        RECT 665.720 20.440 665.980 20.700 ;
        RECT 810.620 19.420 810.880 19.680 ;
        RECT 862.600 19.420 862.860 19.680 ;
        RECT 665.720 17.380 665.980 17.640 ;
        RECT 810.620 17.720 810.880 17.980 ;
        RECT 469.300 16.360 469.560 16.620 ;
        RECT 517.140 16.360 517.400 16.620 ;
        RECT 565.900 15.000 566.160 15.260 ;
        RECT 613.740 15.000 614.000 15.260 ;
      LAYER met2 ;
        RECT 909.750 600.850 910.030 604.000 ;
        RECT 907.280 600.710 910.030 600.850 ;
        RECT 907.280 596.770 907.420 600.710 ;
        RECT 909.750 600.000 910.030 600.710 ;
        RECT 905.440 596.630 907.420 596.770 ;
        RECT 905.440 569.400 905.580 596.630 ;
        RECT 904.980 569.260 905.580 569.400 ;
        RECT 904.980 386.570 905.120 569.260 ;
        RECT 904.000 386.250 904.260 386.570 ;
        RECT 904.920 386.250 905.180 386.570 ;
        RECT 904.060 351.290 904.200 386.250 ;
        RECT 904.060 351.150 904.660 351.290 ;
        RECT 904.520 303.610 904.660 351.150 ;
        RECT 904.460 303.290 904.720 303.610 ;
        RECT 905.380 303.290 905.640 303.610 ;
        RECT 905.440 289.670 905.580 303.290 ;
        RECT 904.460 289.350 904.720 289.670 ;
        RECT 905.380 289.350 905.640 289.670 ;
        RECT 904.520 252.010 904.660 289.350 ;
        RECT 904.520 251.870 905.580 252.010 ;
        RECT 905.440 207.810 905.580 251.870 ;
        RECT 904.980 207.670 905.580 207.810 ;
        RECT 904.980 207.130 905.120 207.670 ;
        RECT 904.520 206.990 905.120 207.130 ;
        RECT 904.520 206.450 904.660 206.990 ;
        RECT 904.520 206.310 905.120 206.450 ;
        RECT 904.980 110.570 905.120 206.310 ;
        RECT 904.520 110.430 905.120 110.570 ;
        RECT 904.520 21.410 904.660 110.430 ;
        RECT 863.060 21.090 863.320 21.410 ;
        RECT 904.460 21.090 904.720 21.410 ;
        RECT 466.540 20.410 466.800 20.730 ;
        RECT 469.300 20.410 469.560 20.730 ;
        RECT 517.140 20.410 517.400 20.730 ;
        RECT 565.900 20.410 566.160 20.730 ;
        RECT 613.740 20.410 614.000 20.730 ;
        RECT 665.720 20.410 665.980 20.730 ;
        RECT 466.600 2.400 466.740 20.410 ;
        RECT 469.360 16.650 469.500 20.410 ;
        RECT 517.200 16.650 517.340 20.410 ;
        RECT 469.300 16.330 469.560 16.650 ;
        RECT 517.140 16.330 517.400 16.650 ;
        RECT 565.960 15.290 566.100 20.410 ;
        RECT 613.800 15.290 613.940 20.410 ;
        RECT 665.780 17.670 665.920 20.410 ;
        RECT 810.620 19.390 810.880 19.710 ;
        RECT 862.600 19.450 862.860 19.710 ;
        RECT 863.120 19.450 863.260 21.090 ;
        RECT 862.600 19.390 863.260 19.450 ;
        RECT 810.680 18.010 810.820 19.390 ;
        RECT 862.660 19.310 863.260 19.390 ;
        RECT 810.620 17.690 810.880 18.010 ;
        RECT 665.720 17.350 665.980 17.670 ;
        RECT 565.900 14.970 566.160 15.290 ;
        RECT 613.740 14.970 614.000 15.290 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 41.040 484.770 41.100 ;
        RECT 918.230 41.040 918.550 41.100 ;
        RECT 484.450 40.900 918.550 41.040 ;
        RECT 484.450 40.840 484.770 40.900 ;
        RECT 918.230 40.840 918.550 40.900 ;
      LAYER via ;
        RECT 484.480 40.840 484.740 41.100 ;
        RECT 918.260 40.840 918.520 41.100 ;
      LAYER met2 ;
        RECT 918.490 600.000 918.770 604.000 ;
        RECT 918.550 598.810 918.690 600.000 ;
        RECT 918.320 598.670 918.690 598.810 ;
        RECT 918.320 41.130 918.460 598.670 ;
        RECT 484.480 40.810 484.740 41.130 ;
        RECT 918.260 40.810 918.520 41.130 ;
        RECT 484.540 2.400 484.680 40.810 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 888.790 18.940 889.110 19.000 ;
        RECT 924.670 18.940 924.990 19.000 ;
        RECT 888.790 18.800 924.990 18.940 ;
        RECT 888.790 18.740 889.110 18.800 ;
        RECT 924.670 18.740 924.990 18.800 ;
        RECT 502.390 16.900 502.710 16.960 ;
        RECT 888.790 16.900 889.110 16.960 ;
        RECT 502.390 16.760 889.110 16.900 ;
        RECT 502.390 16.700 502.710 16.760 ;
        RECT 888.790 16.700 889.110 16.760 ;
      LAYER via ;
        RECT 888.820 18.740 889.080 19.000 ;
        RECT 924.700 18.740 924.960 19.000 ;
        RECT 502.420 16.700 502.680 16.960 ;
        RECT 888.820 16.700 889.080 16.960 ;
      LAYER met2 ;
        RECT 927.690 600.170 927.970 604.000 ;
        RECT 925.680 600.030 927.970 600.170 ;
        RECT 925.680 569.400 925.820 600.030 ;
        RECT 927.690 600.000 927.970 600.030 ;
        RECT 924.760 569.260 925.820 569.400 ;
        RECT 924.760 19.030 924.900 569.260 ;
        RECT 888.820 18.710 889.080 19.030 ;
        RECT 924.700 18.710 924.960 19.030 ;
        RECT 888.880 16.990 889.020 18.710 ;
        RECT 502.420 16.670 502.680 16.990 ;
        RECT 888.820 16.670 889.080 16.990 ;
        RECT 502.480 2.400 502.620 16.670 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 931.570 569.400 931.890 569.460 ;
        RECT 935.250 569.400 935.570 569.460 ;
        RECT 931.570 569.260 935.570 569.400 ;
        RECT 931.570 569.200 931.890 569.260 ;
        RECT 935.250 569.200 935.570 569.260 ;
        RECT 519.870 16.560 520.190 16.620 ;
        RECT 519.870 16.420 908.340 16.560 ;
        RECT 519.870 16.360 520.190 16.420 ;
        RECT 908.200 16.220 908.340 16.420 ;
        RECT 931.570 16.220 931.890 16.280 ;
        RECT 908.200 16.080 931.890 16.220 ;
        RECT 931.570 16.020 931.890 16.080 ;
      LAYER via ;
        RECT 931.600 569.200 931.860 569.460 ;
        RECT 935.280 569.200 935.540 569.460 ;
        RECT 519.900 16.360 520.160 16.620 ;
        RECT 931.600 16.020 931.860 16.280 ;
      LAYER met2 ;
        RECT 936.890 600.170 937.170 604.000 ;
        RECT 935.340 600.030 937.170 600.170 ;
        RECT 935.340 569.490 935.480 600.030 ;
        RECT 936.890 600.000 937.170 600.030 ;
        RECT 931.600 569.170 931.860 569.490 ;
        RECT 935.280 569.170 935.540 569.490 ;
        RECT 519.900 16.330 520.160 16.650 ;
        RECT 519.960 2.400 520.100 16.330 ;
        RECT 931.660 16.310 931.800 569.170 ;
        RECT 931.600 15.990 931.860 16.310 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 16.220 538.130 16.280 ;
        RECT 907.650 16.220 907.970 16.280 ;
        RECT 537.810 16.080 907.970 16.220 ;
        RECT 537.810 16.020 538.130 16.080 ;
        RECT 907.650 16.020 907.970 16.080 ;
        RECT 907.650 15.200 907.970 15.260 ;
        RECT 946.290 15.200 946.610 15.260 ;
        RECT 907.650 15.060 946.610 15.200 ;
        RECT 907.650 15.000 907.970 15.060 ;
        RECT 946.290 15.000 946.610 15.060 ;
      LAYER via ;
        RECT 537.840 16.020 538.100 16.280 ;
        RECT 907.680 16.020 907.940 16.280 ;
        RECT 907.680 15.000 907.940 15.260 ;
        RECT 946.320 15.000 946.580 15.260 ;
      LAYER met2 ;
        RECT 946.090 600.000 946.370 604.000 ;
        RECT 946.150 598.810 946.290 600.000 ;
        RECT 946.150 598.670 946.520 598.810 ;
        RECT 537.840 15.990 538.100 16.310 ;
        RECT 907.680 15.990 907.940 16.310 ;
        RECT 537.900 2.400 538.040 15.990 ;
        RECT 907.740 15.290 907.880 15.990 ;
        RECT 946.380 15.290 946.520 598.670 ;
        RECT 907.680 14.970 907.940 15.290 ;
        RECT 946.320 14.970 946.580 15.290 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 952.270 596.940 952.590 597.000 ;
        RECT 953.650 596.940 953.970 597.000 ;
        RECT 952.270 596.800 953.970 596.940 ;
        RECT 952.270 596.740 952.590 596.800 ;
        RECT 953.650 596.740 953.970 596.800 ;
        RECT 555.750 37.640 556.070 37.700 ;
        RECT 952.730 37.640 953.050 37.700 ;
        RECT 555.750 37.500 953.050 37.640 ;
        RECT 555.750 37.440 556.070 37.500 ;
        RECT 952.730 37.440 953.050 37.500 ;
      LAYER via ;
        RECT 952.300 596.740 952.560 597.000 ;
        RECT 953.680 596.740 953.940 597.000 ;
        RECT 555.780 37.440 556.040 37.700 ;
        RECT 952.760 37.440 953.020 37.700 ;
      LAYER met2 ;
        RECT 955.290 600.170 955.570 604.000 ;
        RECT 953.740 600.030 955.570 600.170 ;
        RECT 953.740 597.030 953.880 600.030 ;
        RECT 955.290 600.000 955.570 600.030 ;
        RECT 952.300 596.710 952.560 597.030 ;
        RECT 953.680 596.710 953.940 597.030 ;
        RECT 952.360 569.570 952.500 596.710 ;
        RECT 952.360 569.430 952.960 569.570 ;
        RECT 952.820 37.730 952.960 569.430 ;
        RECT 555.780 37.410 556.040 37.730 ;
        RECT 952.760 37.410 953.020 37.730 ;
        RECT 555.840 2.400 555.980 37.410 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 838.190 589.120 838.510 589.180 ;
        RECT 962.850 589.120 963.170 589.180 ;
        RECT 838.190 588.980 963.170 589.120 ;
        RECT 838.190 588.920 838.510 588.980 ;
        RECT 962.850 588.920 963.170 588.980 ;
        RECT 838.190 15.880 838.510 15.940 ;
        RECT 586.200 15.740 838.510 15.880 ;
        RECT 573.690 15.540 574.010 15.600 ;
        RECT 586.200 15.540 586.340 15.740 ;
        RECT 838.190 15.680 838.510 15.740 ;
        RECT 573.690 15.400 586.340 15.540 ;
        RECT 573.690 15.340 574.010 15.400 ;
      LAYER via ;
        RECT 838.220 588.920 838.480 589.180 ;
        RECT 962.880 588.920 963.140 589.180 ;
        RECT 573.720 15.340 573.980 15.600 ;
        RECT 838.220 15.680 838.480 15.940 ;
      LAYER met2 ;
        RECT 964.490 600.170 964.770 604.000 ;
        RECT 962.940 600.030 964.770 600.170 ;
        RECT 962.940 589.210 963.080 600.030 ;
        RECT 964.490 600.000 964.770 600.030 ;
        RECT 838.220 588.890 838.480 589.210 ;
        RECT 962.880 588.890 963.140 589.210 ;
        RECT 838.280 15.970 838.420 588.890 ;
        RECT 838.220 15.650 838.480 15.970 ;
        RECT 573.720 15.310 573.980 15.630 ;
        RECT 573.780 2.400 573.920 15.310 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 591.170 41.380 591.490 41.440 ;
        RECT 973.430 41.380 973.750 41.440 ;
        RECT 591.170 41.240 925.360 41.380 ;
        RECT 591.170 41.180 591.490 41.240 ;
        RECT 925.220 41.040 925.360 41.240 ;
        RECT 926.140 41.240 973.750 41.380 ;
        RECT 926.140 41.040 926.280 41.240 ;
        RECT 973.430 41.180 973.750 41.240 ;
        RECT 925.220 40.900 926.280 41.040 ;
      LAYER via ;
        RECT 591.200 41.180 591.460 41.440 ;
        RECT 973.460 41.180 973.720 41.440 ;
      LAYER met2 ;
        RECT 973.690 600.000 973.970 604.000 ;
        RECT 973.750 598.810 973.890 600.000 ;
        RECT 973.520 598.670 973.890 598.810 ;
        RECT 973.520 41.470 973.660 598.670 ;
        RECT 591.200 41.150 591.460 41.470 ;
        RECT 973.460 41.150 973.720 41.470 ;
        RECT 591.260 2.400 591.400 41.150 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 18.260 97.910 18.320 ;
        RECT 718.590 18.260 718.910 18.320 ;
        RECT 97.590 18.120 718.910 18.260 ;
        RECT 97.590 18.060 97.910 18.120 ;
        RECT 718.590 18.060 718.910 18.120 ;
      LAYER via ;
        RECT 97.620 18.060 97.880 18.320 ;
        RECT 718.620 18.060 718.880 18.320 ;
      LAYER met2 ;
        RECT 720.230 600.170 720.510 604.000 ;
        RECT 717.760 600.030 720.510 600.170 ;
        RECT 717.760 41.325 717.900 600.030 ;
        RECT 720.230 600.000 720.510 600.030 ;
        RECT 717.690 40.955 717.970 41.325 ;
        RECT 718.610 40.275 718.890 40.645 ;
        RECT 718.680 18.350 718.820 40.275 ;
        RECT 97.620 18.030 97.880 18.350 ;
        RECT 718.620 18.030 718.880 18.350 ;
        RECT 97.680 2.400 97.820 18.030 ;
        RECT 97.470 -4.800 98.030 2.400 ;
      LAYER via2 ;
        RECT 717.690 41.000 717.970 41.280 ;
        RECT 718.610 40.320 718.890 40.600 ;
      LAYER met3 ;
        RECT 717.665 41.290 717.995 41.305 ;
        RECT 717.665 40.975 718.210 41.290 ;
        RECT 717.910 40.610 718.210 40.975 ;
        RECT 718.585 40.610 718.915 40.625 ;
        RECT 717.910 40.310 718.915 40.610 ;
        RECT 718.585 40.295 718.915 40.310 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 37.300 609.430 37.360 ;
        RECT 980.330 37.300 980.650 37.360 ;
        RECT 609.110 37.160 980.650 37.300 ;
        RECT 609.110 37.100 609.430 37.160 ;
        RECT 980.330 37.100 980.650 37.160 ;
      LAYER via ;
        RECT 609.140 37.100 609.400 37.360 ;
        RECT 980.360 37.100 980.620 37.360 ;
      LAYER met2 ;
        RECT 982.890 600.170 983.170 604.000 ;
        RECT 980.420 600.030 983.170 600.170 ;
        RECT 980.420 37.390 980.560 600.030 ;
        RECT 982.890 600.000 983.170 600.030 ;
        RECT 609.140 37.070 609.400 37.390 ;
        RECT 980.360 37.070 980.620 37.390 ;
        RECT 609.200 2.400 609.340 37.070 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 845.090 589.460 845.410 589.520 ;
        RECT 990.450 589.460 990.770 589.520 ;
        RECT 845.090 589.320 990.770 589.460 ;
        RECT 845.090 589.260 845.410 589.320 ;
        RECT 990.450 589.260 990.770 589.320 ;
        RECT 845.090 15.540 845.410 15.600 ;
        RECT 628.060 15.400 845.410 15.540 ;
        RECT 627.050 15.200 627.370 15.260 ;
        RECT 628.060 15.200 628.200 15.400 ;
        RECT 845.090 15.340 845.410 15.400 ;
        RECT 627.050 15.060 628.200 15.200 ;
        RECT 627.050 15.000 627.370 15.060 ;
      LAYER via ;
        RECT 845.120 589.260 845.380 589.520 ;
        RECT 990.480 589.260 990.740 589.520 ;
        RECT 627.080 15.000 627.340 15.260 ;
        RECT 845.120 15.340 845.380 15.600 ;
      LAYER met2 ;
        RECT 992.090 600.170 992.370 604.000 ;
        RECT 990.540 600.030 992.370 600.170 ;
        RECT 990.540 589.550 990.680 600.030 ;
        RECT 992.090 600.000 992.370 600.030 ;
        RECT 845.120 589.230 845.380 589.550 ;
        RECT 990.480 589.230 990.740 589.550 ;
        RECT 845.180 15.630 845.320 589.230 ;
        RECT 845.120 15.310 845.380 15.630 ;
        RECT 627.080 14.970 627.340 15.290 ;
        RECT 627.140 2.400 627.280 14.970 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 18.940 121.830 19.000 ;
        RECT 731.470 18.940 731.790 19.000 ;
        RECT 121.510 18.800 731.790 18.940 ;
        RECT 121.510 18.740 121.830 18.800 ;
        RECT 731.470 18.740 731.790 18.800 ;
      LAYER via ;
        RECT 121.540 18.740 121.800 19.000 ;
        RECT 731.500 18.740 731.760 19.000 ;
      LAYER met2 ;
        RECT 732.190 600.170 732.470 604.000 ;
        RECT 731.560 600.030 732.470 600.170 ;
        RECT 731.560 19.030 731.700 600.030 ;
        RECT 732.190 600.000 732.470 600.030 ;
        RECT 121.540 18.710 121.800 19.030 ;
        RECT 731.500 18.710 731.760 19.030 ;
        RECT 121.600 2.400 121.740 18.710 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 739.290 517.720 739.610 517.780 ;
        RECT 742.050 517.720 742.370 517.780 ;
        RECT 739.290 517.580 742.370 517.720 ;
        RECT 739.290 517.520 739.610 517.580 ;
        RECT 742.050 517.520 742.370 517.580 ;
        RECT 739.290 469.440 739.610 469.500 ;
        RECT 739.750 469.440 740.070 469.500 ;
        RECT 739.290 469.300 740.070 469.440 ;
        RECT 739.290 469.240 739.610 469.300 ;
        RECT 739.750 469.240 740.070 469.300 ;
        RECT 739.290 448.500 739.610 448.760 ;
        RECT 739.380 448.020 739.520 448.500 ;
        RECT 739.750 448.020 740.070 448.080 ;
        RECT 739.380 447.880 740.070 448.020 ;
        RECT 739.750 447.820 740.070 447.880 ;
        RECT 738.370 427.620 738.690 427.680 ;
        RECT 739.750 427.620 740.070 427.680 ;
        RECT 738.370 427.480 740.070 427.620 ;
        RECT 738.370 427.420 738.690 427.480 ;
        RECT 739.750 427.420 740.070 427.480 ;
        RECT 738.370 379.340 738.690 379.400 ;
        RECT 739.290 379.340 739.610 379.400 ;
        RECT 738.370 379.200 739.610 379.340 ;
        RECT 738.370 379.140 738.690 379.200 ;
        RECT 739.290 379.140 739.610 379.200 ;
        RECT 739.290 338.000 739.610 338.260 ;
        RECT 739.380 337.580 739.520 338.000 ;
        RECT 739.290 337.320 739.610 337.580 ;
        RECT 739.290 289.240 739.610 289.300 ;
        RECT 740.210 289.240 740.530 289.300 ;
        RECT 739.290 289.100 740.530 289.240 ;
        RECT 739.290 289.040 739.610 289.100 ;
        RECT 740.210 289.040 740.530 289.100 ;
        RECT 739.290 144.740 739.610 144.800 ;
        RECT 739.750 144.740 740.070 144.800 ;
        RECT 739.290 144.600 740.070 144.740 ;
        RECT 739.290 144.540 739.610 144.600 ;
        RECT 739.750 144.540 740.070 144.600 ;
        RECT 739.290 96.800 739.610 96.860 ;
        RECT 739.750 96.800 740.070 96.860 ;
        RECT 739.290 96.660 740.070 96.800 ;
        RECT 739.290 96.600 739.610 96.660 ;
        RECT 739.750 96.600 740.070 96.660 ;
        RECT 145.430 19.280 145.750 19.340 ;
        RECT 739.290 19.280 739.610 19.340 ;
        RECT 145.430 19.140 739.610 19.280 ;
        RECT 145.430 19.080 145.750 19.140 ;
        RECT 739.290 19.080 739.610 19.140 ;
      LAYER via ;
        RECT 739.320 517.520 739.580 517.780 ;
        RECT 742.080 517.520 742.340 517.780 ;
        RECT 739.320 469.240 739.580 469.500 ;
        RECT 739.780 469.240 740.040 469.500 ;
        RECT 739.320 448.500 739.580 448.760 ;
        RECT 739.780 447.820 740.040 448.080 ;
        RECT 738.400 427.420 738.660 427.680 ;
        RECT 739.780 427.420 740.040 427.680 ;
        RECT 738.400 379.140 738.660 379.400 ;
        RECT 739.320 379.140 739.580 379.400 ;
        RECT 739.320 338.000 739.580 338.260 ;
        RECT 739.320 337.320 739.580 337.580 ;
        RECT 739.320 289.040 739.580 289.300 ;
        RECT 740.240 289.040 740.500 289.300 ;
        RECT 739.320 144.540 739.580 144.800 ;
        RECT 739.780 144.540 740.040 144.800 ;
        RECT 739.320 96.600 739.580 96.860 ;
        RECT 739.780 96.600 740.040 96.860 ;
        RECT 145.460 19.080 145.720 19.340 ;
        RECT 739.320 19.080 739.580 19.340 ;
      LAYER met2 ;
        RECT 744.610 600.170 744.890 604.000 ;
        RECT 742.140 600.030 744.890 600.170 ;
        RECT 742.140 517.810 742.280 600.030 ;
        RECT 744.610 600.000 744.890 600.030 ;
        RECT 739.320 517.490 739.580 517.810 ;
        RECT 742.080 517.490 742.340 517.810 ;
        RECT 739.380 517.210 739.520 517.490 ;
        RECT 739.380 517.070 739.980 517.210 ;
        RECT 739.840 469.530 739.980 517.070 ;
        RECT 739.320 469.210 739.580 469.530 ;
        RECT 739.780 469.210 740.040 469.530 ;
        RECT 739.380 448.790 739.520 469.210 ;
        RECT 739.320 448.470 739.580 448.790 ;
        RECT 739.780 447.790 740.040 448.110 ;
        RECT 739.840 427.710 739.980 447.790 ;
        RECT 738.400 427.390 738.660 427.710 ;
        RECT 739.780 427.390 740.040 427.710 ;
        RECT 738.460 379.430 738.600 427.390 ;
        RECT 738.400 379.110 738.660 379.430 ;
        RECT 739.320 379.110 739.580 379.430 ;
        RECT 739.380 338.290 739.520 379.110 ;
        RECT 739.320 337.970 739.580 338.290 ;
        RECT 739.320 337.290 739.580 337.610 ;
        RECT 739.380 289.330 739.520 337.290 ;
        RECT 739.320 289.010 739.580 289.330 ;
        RECT 740.240 289.010 740.500 289.330 ;
        RECT 740.300 254.730 740.440 289.010 ;
        RECT 739.840 254.590 740.440 254.730 ;
        RECT 739.840 217.330 739.980 254.590 ;
        RECT 739.380 217.190 739.980 217.330 ;
        RECT 739.380 144.830 739.520 217.190 ;
        RECT 739.320 144.510 739.580 144.830 ;
        RECT 739.780 144.510 740.040 144.830 ;
        RECT 739.840 96.890 739.980 144.510 ;
        RECT 739.320 96.570 739.580 96.890 ;
        RECT 739.780 96.570 740.040 96.890 ;
        RECT 739.380 19.370 739.520 96.570 ;
        RECT 145.460 19.050 145.720 19.370 ;
        RECT 739.320 19.050 739.580 19.370 ;
        RECT 145.520 2.400 145.660 19.050 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 30.840 163.690 30.900 ;
        RECT 752.630 30.840 752.950 30.900 ;
        RECT 163.370 30.700 752.950 30.840 ;
        RECT 163.370 30.640 163.690 30.700 ;
        RECT 752.630 30.640 752.950 30.700 ;
      LAYER via ;
        RECT 163.400 30.640 163.660 30.900 ;
        RECT 752.660 30.640 752.920 30.900 ;
      LAYER met2 ;
        RECT 753.810 600.170 754.090 604.000 ;
        RECT 752.720 600.030 754.090 600.170 ;
        RECT 752.720 30.930 752.860 600.030 ;
        RECT 753.810 600.000 754.090 600.030 ;
        RECT 163.400 30.610 163.660 30.930 ;
        RECT 752.660 30.610 752.920 30.930 ;
        RECT 163.460 2.400 163.600 30.610 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 760.450 598.980 760.770 599.040 ;
        RECT 762.980 598.980 763.300 599.040 ;
        RECT 760.450 598.840 763.300 598.980 ;
        RECT 760.450 598.780 760.770 598.840 ;
        RECT 762.980 598.780 763.300 598.840 ;
        RECT 760.450 517.720 760.770 517.780 ;
        RECT 760.910 517.720 761.230 517.780 ;
        RECT 760.450 517.580 761.230 517.720 ;
        RECT 760.450 517.520 760.770 517.580 ;
        RECT 760.910 517.520 761.230 517.580 ;
        RECT 759.070 469.440 759.390 469.500 ;
        RECT 760.910 469.440 761.230 469.500 ;
        RECT 759.070 469.300 761.230 469.440 ;
        RECT 759.070 469.240 759.390 469.300 ;
        RECT 760.910 469.240 761.230 469.300 ;
        RECT 759.070 427.620 759.390 427.680 ;
        RECT 759.530 427.620 759.850 427.680 ;
        RECT 759.070 427.480 759.850 427.620 ;
        RECT 759.070 427.420 759.390 427.480 ;
        RECT 759.530 427.420 759.850 427.480 ;
        RECT 468.810 20.980 469.130 21.040 ;
        RECT 466.140 20.840 469.130 20.980 ;
        RECT 324.370 20.640 324.690 20.700 ;
        RECT 368.530 20.640 368.850 20.700 ;
        RECT 324.370 20.500 368.850 20.640 ;
        RECT 324.370 20.440 324.690 20.500 ;
        RECT 368.530 20.440 368.850 20.500 ;
        RECT 420.970 20.640 421.290 20.700 ;
        RECT 466.140 20.640 466.280 20.840 ;
        RECT 468.810 20.780 469.130 20.840 ;
        RECT 420.970 20.500 466.280 20.640 ;
        RECT 420.970 20.440 421.290 20.500 ;
        RECT 759.070 19.960 759.390 20.020 ;
        RECT 739.840 19.820 759.390 19.960 ;
        RECT 180.850 19.620 181.170 19.680 ;
        RECT 324.370 19.620 324.690 19.680 ;
        RECT 180.850 19.480 324.690 19.620 ;
        RECT 180.850 19.420 181.170 19.480 ;
        RECT 324.370 19.420 324.690 19.480 ;
        RECT 368.530 19.620 368.850 19.680 ;
        RECT 420.970 19.620 421.290 19.680 ;
        RECT 368.530 19.480 421.290 19.620 ;
        RECT 368.530 19.420 368.850 19.480 ;
        RECT 420.970 19.420 421.290 19.480 ;
        RECT 468.810 19.620 469.130 19.680 ;
        RECT 517.570 19.620 517.890 19.680 ;
        RECT 468.810 19.480 517.890 19.620 ;
        RECT 468.810 19.420 469.130 19.480 ;
        RECT 517.570 19.420 517.890 19.480 ;
        RECT 565.410 19.620 565.730 19.680 ;
        RECT 614.170 19.620 614.490 19.680 ;
        RECT 565.410 19.480 614.490 19.620 ;
        RECT 565.410 19.420 565.730 19.480 ;
        RECT 614.170 19.420 614.490 19.480 ;
        RECT 665.230 19.620 665.550 19.680 ;
        RECT 739.840 19.620 739.980 19.820 ;
        RECT 759.070 19.760 759.390 19.820 ;
        RECT 665.230 19.480 739.980 19.620 ;
        RECT 665.230 19.420 665.550 19.480 ;
        RECT 517.570 15.880 517.890 15.940 ;
        RECT 565.410 15.880 565.730 15.940 ;
        RECT 517.570 15.740 565.730 15.880 ;
        RECT 517.570 15.680 517.890 15.740 ;
        RECT 565.410 15.680 565.730 15.740 ;
        RECT 614.170 14.860 614.490 14.920 ;
        RECT 665.230 14.860 665.550 14.920 ;
        RECT 614.170 14.720 665.550 14.860 ;
        RECT 614.170 14.660 614.490 14.720 ;
        RECT 665.230 14.660 665.550 14.720 ;
      LAYER via ;
        RECT 760.480 598.780 760.740 599.040 ;
        RECT 763.010 598.780 763.270 599.040 ;
        RECT 760.480 517.520 760.740 517.780 ;
        RECT 760.940 517.520 761.200 517.780 ;
        RECT 759.100 469.240 759.360 469.500 ;
        RECT 760.940 469.240 761.200 469.500 ;
        RECT 759.100 427.420 759.360 427.680 ;
        RECT 759.560 427.420 759.820 427.680 ;
        RECT 324.400 20.440 324.660 20.700 ;
        RECT 368.560 20.440 368.820 20.700 ;
        RECT 421.000 20.440 421.260 20.700 ;
        RECT 468.840 20.780 469.100 21.040 ;
        RECT 180.880 19.420 181.140 19.680 ;
        RECT 324.400 19.420 324.660 19.680 ;
        RECT 368.560 19.420 368.820 19.680 ;
        RECT 421.000 19.420 421.260 19.680 ;
        RECT 468.840 19.420 469.100 19.680 ;
        RECT 517.600 19.420 517.860 19.680 ;
        RECT 565.440 19.420 565.700 19.680 ;
        RECT 614.200 19.420 614.460 19.680 ;
        RECT 665.260 19.420 665.520 19.680 ;
        RECT 759.100 19.760 759.360 20.020 ;
        RECT 517.600 15.680 517.860 15.940 ;
        RECT 565.440 15.680 565.700 15.940 ;
        RECT 614.200 14.660 614.460 14.920 ;
        RECT 665.260 14.660 665.520 14.920 ;
      LAYER met2 ;
        RECT 763.010 600.000 763.290 604.000 ;
        RECT 763.070 599.070 763.210 600.000 ;
        RECT 760.480 598.750 760.740 599.070 ;
        RECT 763.010 598.750 763.270 599.070 ;
        RECT 760.540 517.810 760.680 598.750 ;
        RECT 760.480 517.490 760.740 517.810 ;
        RECT 760.940 517.490 761.200 517.810 ;
        RECT 761.000 469.530 761.140 517.490 ;
        RECT 759.100 469.210 759.360 469.530 ;
        RECT 760.940 469.210 761.200 469.530 ;
        RECT 759.160 451.930 759.300 469.210 ;
        RECT 759.160 451.790 759.760 451.930 ;
        RECT 759.620 427.710 759.760 451.790 ;
        RECT 759.100 427.390 759.360 427.710 ;
        RECT 759.560 427.390 759.820 427.710 ;
        RECT 468.840 20.750 469.100 21.070 ;
        RECT 324.400 20.410 324.660 20.730 ;
        RECT 368.560 20.410 368.820 20.730 ;
        RECT 421.000 20.410 421.260 20.730 ;
        RECT 324.460 19.710 324.600 20.410 ;
        RECT 368.620 19.710 368.760 20.410 ;
        RECT 421.060 19.710 421.200 20.410 ;
        RECT 468.900 19.710 469.040 20.750 ;
        RECT 759.160 20.050 759.300 427.390 ;
        RECT 759.100 19.730 759.360 20.050 ;
        RECT 180.880 19.390 181.140 19.710 ;
        RECT 324.400 19.390 324.660 19.710 ;
        RECT 368.560 19.390 368.820 19.710 ;
        RECT 421.000 19.390 421.260 19.710 ;
        RECT 468.840 19.390 469.100 19.710 ;
        RECT 517.600 19.390 517.860 19.710 ;
        RECT 565.440 19.390 565.700 19.710 ;
        RECT 614.200 19.390 614.460 19.710 ;
        RECT 665.260 19.390 665.520 19.710 ;
        RECT 180.940 2.400 181.080 19.390 ;
        RECT 517.660 15.970 517.800 19.390 ;
        RECT 565.500 15.970 565.640 19.390 ;
        RECT 517.600 15.650 517.860 15.970 ;
        RECT 565.440 15.650 565.700 15.970 ;
        RECT 614.260 14.950 614.400 19.390 ;
        RECT 665.320 14.950 665.460 19.390 ;
        RECT 614.200 14.630 614.460 14.950 ;
        RECT 665.260 14.630 665.520 14.950 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 766.430 550.700 766.750 550.760 ;
        RECT 770.570 550.700 770.890 550.760 ;
        RECT 766.430 550.560 770.890 550.700 ;
        RECT 766.430 550.500 766.750 550.560 ;
        RECT 770.570 550.500 770.890 550.560 ;
        RECT 198.790 31.520 199.110 31.580 ;
        RECT 766.430 31.520 766.750 31.580 ;
        RECT 198.790 31.380 766.750 31.520 ;
        RECT 198.790 31.320 199.110 31.380 ;
        RECT 766.430 31.320 766.750 31.380 ;
      LAYER via ;
        RECT 766.460 550.500 766.720 550.760 ;
        RECT 770.600 550.500 770.860 550.760 ;
        RECT 198.820 31.320 199.080 31.580 ;
        RECT 766.460 31.320 766.720 31.580 ;
      LAYER met2 ;
        RECT 772.210 600.170 772.490 604.000 ;
        RECT 770.660 600.030 772.490 600.170 ;
        RECT 770.660 550.790 770.800 600.030 ;
        RECT 772.210 600.000 772.490 600.030 ;
        RECT 766.460 550.470 766.720 550.790 ;
        RECT 770.600 550.470 770.860 550.790 ;
        RECT 766.520 31.610 766.660 550.470 ;
        RECT 198.820 31.290 199.080 31.610 ;
        RECT 766.460 31.290 766.720 31.610 ;
        RECT 198.880 2.400 199.020 31.290 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 19.960 217.050 20.020 ;
        RECT 738.830 19.960 739.150 20.020 ;
        RECT 216.730 19.820 739.150 19.960 ;
        RECT 216.730 19.760 217.050 19.820 ;
        RECT 738.830 19.760 739.150 19.820 ;
        RECT 738.830 18.940 739.150 19.000 ;
        RECT 779.770 18.940 780.090 19.000 ;
        RECT 738.830 18.800 780.090 18.940 ;
        RECT 738.830 18.740 739.150 18.800 ;
        RECT 779.770 18.740 780.090 18.800 ;
      LAYER via ;
        RECT 216.760 19.760 217.020 20.020 ;
        RECT 738.860 19.760 739.120 20.020 ;
        RECT 738.860 18.740 739.120 19.000 ;
        RECT 779.800 18.740 780.060 19.000 ;
      LAYER met2 ;
        RECT 781.410 600.170 781.690 604.000 ;
        RECT 779.860 600.030 781.690 600.170 ;
        RECT 216.760 19.730 217.020 20.050 ;
        RECT 738.860 19.730 739.120 20.050 ;
        RECT 216.820 2.400 216.960 19.730 ;
        RECT 738.920 19.030 739.060 19.730 ;
        RECT 779.860 19.030 780.000 600.030 ;
        RECT 781.410 600.000 781.690 600.030 ;
        RECT 738.860 18.710 739.120 19.030 ;
        RECT 779.800 18.710 780.060 19.030 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 787.130 144.740 787.450 144.800 ;
        RECT 787.590 144.740 787.910 144.800 ;
        RECT 787.130 144.600 787.910 144.740 ;
        RECT 787.130 144.540 787.450 144.600 ;
        RECT 787.590 144.540 787.910 144.600 ;
        RECT 787.130 96.800 787.450 96.860 ;
        RECT 787.590 96.800 787.910 96.860 ;
        RECT 787.130 96.660 787.910 96.800 ;
        RECT 787.130 96.600 787.450 96.660 ;
        RECT 787.590 96.600 787.910 96.660 ;
        RECT 234.670 20.300 234.990 20.360 ;
        RECT 786.670 20.300 786.990 20.360 ;
        RECT 234.670 20.160 786.990 20.300 ;
        RECT 234.670 20.100 234.990 20.160 ;
        RECT 786.670 20.100 786.990 20.160 ;
      LAYER via ;
        RECT 787.160 144.540 787.420 144.800 ;
        RECT 787.620 144.540 787.880 144.800 ;
        RECT 787.160 96.600 787.420 96.860 ;
        RECT 787.620 96.600 787.880 96.860 ;
        RECT 234.700 20.100 234.960 20.360 ;
        RECT 786.700 20.100 786.960 20.360 ;
      LAYER met2 ;
        RECT 790.610 600.850 790.890 604.000 ;
        RECT 788.140 600.710 790.890 600.850 ;
        RECT 788.140 596.770 788.280 600.710 ;
        RECT 790.610 600.000 790.890 600.710 ;
        RECT 787.220 596.630 788.280 596.770 ;
        RECT 787.220 144.830 787.360 596.630 ;
        RECT 787.160 144.510 787.420 144.830 ;
        RECT 787.620 144.510 787.880 144.830 ;
        RECT 787.680 96.890 787.820 144.510 ;
        RECT 787.160 96.570 787.420 96.890 ;
        RECT 787.620 96.570 787.880 96.890 ;
        RECT 787.220 72.490 787.360 96.570 ;
        RECT 786.760 72.350 787.360 72.490 ;
        RECT 786.760 20.390 786.900 72.350 ;
        RECT 234.700 20.070 234.960 20.390 ;
        RECT 786.700 20.070 786.960 20.390 ;
        RECT 234.760 2.400 234.900 20.070 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 697.890 17.920 698.210 17.980 ;
        RECT 648.760 17.780 698.210 17.920 ;
        RECT 56.190 17.580 56.510 17.640 ;
        RECT 648.760 17.580 648.900 17.780 ;
        RECT 697.890 17.720 698.210 17.780 ;
        RECT 56.190 17.440 648.900 17.580 ;
        RECT 56.190 17.380 56.510 17.440 ;
      LAYER via ;
        RECT 56.220 17.380 56.480 17.640 ;
        RECT 697.920 17.720 698.180 17.980 ;
      LAYER met2 ;
        RECT 698.610 600.170 698.890 604.000 ;
        RECT 697.980 600.030 698.890 600.170 ;
        RECT 697.980 18.010 698.120 600.030 ;
        RECT 698.610 600.000 698.890 600.030 ;
        RECT 697.920 17.690 698.180 18.010 ;
        RECT 56.220 17.350 56.480 17.670 ;
        RECT 56.280 2.400 56.420 17.350 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 51.580 82.730 51.640 ;
        RECT 711.690 51.580 712.010 51.640 ;
        RECT 82.410 51.440 712.010 51.580 ;
        RECT 82.410 51.380 82.730 51.440 ;
        RECT 711.690 51.380 712.010 51.440 ;
        RECT 80.110 16.900 80.430 16.960 ;
        RECT 82.410 16.900 82.730 16.960 ;
        RECT 80.110 16.760 82.730 16.900 ;
        RECT 80.110 16.700 80.430 16.760 ;
        RECT 82.410 16.700 82.730 16.760 ;
      LAYER via ;
        RECT 82.440 51.380 82.700 51.640 ;
        RECT 711.720 51.380 711.980 51.640 ;
        RECT 80.140 16.700 80.400 16.960 ;
        RECT 82.440 16.700 82.700 16.960 ;
      LAYER met2 ;
        RECT 711.030 600.170 711.310 604.000 ;
        RECT 711.030 600.030 711.920 600.170 ;
        RECT 711.030 600.000 711.310 600.030 ;
        RECT 711.780 51.670 711.920 600.030 ;
        RECT 82.440 51.350 82.700 51.670 ;
        RECT 711.720 51.350 711.980 51.670 ;
        RECT 82.500 16.990 82.640 51.350 ;
        RECT 80.140 16.670 80.400 16.990 ;
        RECT 82.440 16.670 82.700 16.990 ;
        RECT 80.200 2.400 80.340 16.670 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 718.130 596.940 718.450 597.000 ;
        RECT 721.810 596.940 722.130 597.000 ;
        RECT 718.130 596.800 722.130 596.940 ;
        RECT 718.130 596.740 718.450 596.800 ;
        RECT 721.810 596.740 722.130 596.800 ;
        RECT 717.210 469.100 717.530 469.160 ;
        RECT 718.130 469.100 718.450 469.160 ;
        RECT 717.210 468.960 718.450 469.100 ;
        RECT 717.210 468.900 717.530 468.960 ;
        RECT 718.130 468.900 718.450 468.960 ;
        RECT 718.590 420.820 718.910 420.880 ;
        RECT 719.510 420.820 719.830 420.880 ;
        RECT 718.590 420.680 719.830 420.820 ;
        RECT 718.590 420.620 718.910 420.680 ;
        RECT 719.510 420.620 719.830 420.680 ;
        RECT 719.510 414.020 719.830 414.080 ;
        RECT 720.430 414.020 720.750 414.080 ;
        RECT 719.510 413.880 720.750 414.020 ;
        RECT 719.510 413.820 719.830 413.880 ;
        RECT 720.430 413.820 720.750 413.880 ;
        RECT 719.510 366.080 719.830 366.140 ;
        RECT 720.430 366.080 720.750 366.140 ;
        RECT 719.510 365.940 720.750 366.080 ;
        RECT 719.510 365.880 719.830 365.940 ;
        RECT 720.430 365.880 720.750 365.940 ;
        RECT 718.130 324.600 718.450 324.660 ;
        RECT 719.970 324.600 720.290 324.660 ;
        RECT 718.130 324.460 720.290 324.600 ;
        RECT 718.130 324.400 718.450 324.460 ;
        RECT 719.970 324.400 720.290 324.460 ;
        RECT 718.130 317.460 718.450 317.520 ;
        RECT 719.050 317.460 719.370 317.520 ;
        RECT 718.130 317.320 719.370 317.460 ;
        RECT 718.130 317.260 718.450 317.320 ;
        RECT 719.050 317.260 719.370 317.320 ;
        RECT 718.590 210.020 718.910 210.080 ;
        RECT 718.220 209.880 718.910 210.020 ;
        RECT 718.220 209.740 718.360 209.880 ;
        RECT 718.590 209.820 718.910 209.880 ;
        RECT 718.130 209.480 718.450 209.740 ;
        RECT 103.570 18.600 103.890 18.660 ;
        RECT 719.510 18.600 719.830 18.660 ;
        RECT 103.570 18.460 719.830 18.600 ;
        RECT 103.570 18.400 103.890 18.460 ;
        RECT 719.510 18.400 719.830 18.460 ;
      LAYER via ;
        RECT 718.160 596.740 718.420 597.000 ;
        RECT 721.840 596.740 722.100 597.000 ;
        RECT 717.240 468.900 717.500 469.160 ;
        RECT 718.160 468.900 718.420 469.160 ;
        RECT 718.620 420.620 718.880 420.880 ;
        RECT 719.540 420.620 719.800 420.880 ;
        RECT 719.540 413.820 719.800 414.080 ;
        RECT 720.460 413.820 720.720 414.080 ;
        RECT 719.540 365.880 719.800 366.140 ;
        RECT 720.460 365.880 720.720 366.140 ;
        RECT 718.160 324.400 718.420 324.660 ;
        RECT 720.000 324.400 720.260 324.660 ;
        RECT 718.160 317.260 718.420 317.520 ;
        RECT 719.080 317.260 719.340 317.520 ;
        RECT 718.620 209.820 718.880 210.080 ;
        RECT 718.160 209.480 718.420 209.740 ;
        RECT 103.600 18.400 103.860 18.660 ;
        RECT 719.540 18.400 719.800 18.660 ;
      LAYER met2 ;
        RECT 722.990 600.170 723.270 604.000 ;
        RECT 721.900 600.030 723.270 600.170 ;
        RECT 721.900 597.030 722.040 600.030 ;
        RECT 722.990 600.000 723.270 600.030 ;
        RECT 718.160 596.710 718.420 597.030 ;
        RECT 721.840 596.710 722.100 597.030 ;
        RECT 718.220 469.190 718.360 596.710 ;
        RECT 717.240 468.870 717.500 469.190 ;
        RECT 718.160 468.870 718.420 469.190 ;
        RECT 717.300 421.445 717.440 468.870 ;
        RECT 717.230 421.075 717.510 421.445 ;
        RECT 718.610 421.075 718.890 421.445 ;
        RECT 718.680 420.910 718.820 421.075 ;
        RECT 718.620 420.590 718.880 420.910 ;
        RECT 719.540 420.590 719.800 420.910 ;
        RECT 719.600 414.110 719.740 420.590 ;
        RECT 719.540 413.790 719.800 414.110 ;
        RECT 720.460 413.790 720.720 414.110 ;
        RECT 720.520 366.170 720.660 413.790 ;
        RECT 719.540 365.850 719.800 366.170 ;
        RECT 720.460 365.850 720.720 366.170 ;
        RECT 719.600 331.570 719.740 365.850 ;
        RECT 719.600 331.430 720.200 331.570 ;
        RECT 720.060 324.690 720.200 331.430 ;
        RECT 718.160 324.370 718.420 324.690 ;
        RECT 720.000 324.370 720.260 324.690 ;
        RECT 718.220 317.550 718.360 324.370 ;
        RECT 718.160 317.230 718.420 317.550 ;
        RECT 719.080 317.230 719.340 317.550 ;
        RECT 719.140 241.130 719.280 317.230 ;
        RECT 718.680 240.990 719.280 241.130 ;
        RECT 718.680 210.110 718.820 240.990 ;
        RECT 718.620 209.790 718.880 210.110 ;
        RECT 718.160 209.450 718.420 209.770 ;
        RECT 718.220 41.210 718.360 209.450 ;
        RECT 718.220 41.070 719.740 41.210 ;
        RECT 719.600 18.690 719.740 41.070 ;
        RECT 103.600 18.370 103.860 18.690 ;
        RECT 719.540 18.370 719.800 18.690 ;
        RECT 103.660 2.400 103.800 18.370 ;
        RECT 103.450 -4.800 104.010 2.400 ;
      LAYER via2 ;
        RECT 717.230 421.120 717.510 421.400 ;
        RECT 718.610 421.120 718.890 421.400 ;
      LAYER met3 ;
        RECT 717.205 421.410 717.535 421.425 ;
        RECT 718.585 421.410 718.915 421.425 ;
        RECT 717.205 421.110 718.915 421.410 ;
        RECT 717.205 421.095 717.535 421.110 ;
        RECT 718.585 421.095 718.915 421.110 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 130.710 51.920 131.030 51.980 ;
        RECT 731.930 51.920 732.250 51.980 ;
        RECT 130.710 51.780 732.250 51.920 ;
        RECT 130.710 51.720 131.030 51.780 ;
        RECT 731.930 51.720 732.250 51.780 ;
        RECT 127.490 16.900 127.810 16.960 ;
        RECT 130.710 16.900 131.030 16.960 ;
        RECT 127.490 16.760 131.030 16.900 ;
        RECT 127.490 16.700 127.810 16.760 ;
        RECT 130.710 16.700 131.030 16.760 ;
      LAYER via ;
        RECT 130.740 51.720 131.000 51.980 ;
        RECT 731.960 51.720 732.220 51.980 ;
        RECT 127.520 16.700 127.780 16.960 ;
        RECT 130.740 16.700 131.000 16.960 ;
      LAYER met2 ;
        RECT 735.410 600.170 735.690 604.000 ;
        RECT 732.940 600.030 735.690 600.170 ;
        RECT 732.940 590.650 733.080 600.030 ;
        RECT 735.410 600.000 735.690 600.030 ;
        RECT 732.020 590.510 733.080 590.650 ;
        RECT 732.020 52.010 732.160 590.510 ;
        RECT 130.740 51.690 131.000 52.010 ;
        RECT 731.960 51.690 732.220 52.010 ;
        RECT 130.800 16.990 130.940 51.690 ;
        RECT 127.520 16.670 127.780 16.990 ;
        RECT 130.740 16.670 131.000 16.990 ;
        RECT 127.580 2.400 127.720 16.670 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 684.550 255.380 684.870 255.640 ;
        RECT 684.640 254.960 684.780 255.380 ;
        RECT 684.550 254.700 684.870 254.960 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 684.550 17.240 684.870 17.300 ;
        RECT 26.290 17.100 684.870 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 684.550 17.040 684.870 17.100 ;
      LAYER via ;
        RECT 684.580 255.380 684.840 255.640 ;
        RECT 684.580 254.700 684.840 254.960 ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 684.580 17.040 684.840 17.300 ;
      LAYER met2 ;
        RECT 683.430 600.170 683.710 604.000 ;
        RECT 683.430 600.030 684.780 600.170 ;
        RECT 683.430 600.000 683.710 600.030 ;
        RECT 684.640 255.670 684.780 600.030 ;
        RECT 684.580 255.350 684.840 255.670 ;
        RECT 684.580 254.670 684.840 254.990 ;
        RECT 684.640 17.330 684.780 254.670 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 684.580 17.010 684.840 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 685.010 524.520 685.330 524.580 ;
        RECT 685.930 524.520 686.250 524.580 ;
        RECT 685.010 524.380 686.250 524.520 ;
        RECT 685.010 524.320 685.330 524.380 ;
        RECT 685.930 524.320 686.250 524.380 ;
        RECT 684.090 496.980 684.410 497.040 ;
        RECT 685.010 496.980 685.330 497.040 ;
        RECT 684.090 496.840 685.330 496.980 ;
        RECT 684.090 496.780 684.410 496.840 ;
        RECT 685.010 496.780 685.330 496.840 ;
        RECT 684.090 255.920 684.410 255.980 ;
        RECT 684.090 255.780 685.240 255.920 ;
        RECT 684.090 255.720 684.410 255.780 ;
        RECT 685.100 255.300 685.240 255.780 ;
        RECT 685.010 255.040 685.330 255.300 ;
        RECT 684.090 207.300 684.410 207.360 ;
        RECT 685.010 207.300 685.330 207.360 ;
        RECT 684.090 207.160 685.330 207.300 ;
        RECT 684.090 207.100 684.410 207.160 ;
        RECT 685.010 207.100 685.330 207.160 ;
        RECT 673.970 89.660 674.290 89.720 ;
        RECT 684.090 89.660 684.410 89.720 ;
        RECT 673.970 89.520 684.410 89.660 ;
        RECT 673.970 89.460 674.290 89.520 ;
        RECT 684.090 89.460 684.410 89.520 ;
        RECT 32.270 44.780 32.590 44.840 ;
        RECT 673.970 44.780 674.290 44.840 ;
        RECT 32.270 44.640 674.290 44.780 ;
        RECT 32.270 44.580 32.590 44.640 ;
        RECT 673.970 44.580 674.290 44.640 ;
      LAYER via ;
        RECT 685.040 524.320 685.300 524.580 ;
        RECT 685.960 524.320 686.220 524.580 ;
        RECT 684.120 496.780 684.380 497.040 ;
        RECT 685.040 496.780 685.300 497.040 ;
        RECT 684.120 255.720 684.380 255.980 ;
        RECT 685.040 255.040 685.300 255.300 ;
        RECT 684.120 207.100 684.380 207.360 ;
        RECT 685.040 207.100 685.300 207.360 ;
        RECT 674.000 89.460 674.260 89.720 ;
        RECT 684.120 89.460 684.380 89.720 ;
        RECT 32.300 44.580 32.560 44.840 ;
        RECT 674.000 44.580 674.260 44.840 ;
      LAYER met2 ;
        RECT 686.650 600.170 686.930 604.000 ;
        RECT 686.020 600.030 686.930 600.170 ;
        RECT 686.020 524.610 686.160 600.030 ;
        RECT 686.650 600.000 686.930 600.030 ;
        RECT 685.040 524.290 685.300 524.610 ;
        RECT 685.960 524.290 686.220 524.610 ;
        RECT 685.100 497.070 685.240 524.290 ;
        RECT 684.120 496.750 684.380 497.070 ;
        RECT 685.040 496.750 685.300 497.070 ;
        RECT 684.180 256.010 684.320 496.750 ;
        RECT 684.120 255.690 684.380 256.010 ;
        RECT 685.040 255.010 685.300 255.330 ;
        RECT 685.100 207.390 685.240 255.010 ;
        RECT 684.120 207.070 684.380 207.390 ;
        RECT 685.040 207.070 685.300 207.390 ;
        RECT 684.180 89.750 684.320 207.070 ;
        RECT 674.000 89.430 674.260 89.750 ;
        RECT 684.120 89.430 684.380 89.750 ;
        RECT 674.060 44.870 674.200 89.430 ;
        RECT 32.300 44.550 32.560 44.870 ;
        RECT 674.000 44.550 674.260 44.870 ;
        RECT 32.360 2.400 32.500 44.550 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 1982.750 367.020 3529.000 ;
        RECT 544.020 2760.520 547.020 3529.000 ;
        RECT 457.645 2610.640 459.245 2747.120 ;
        RECT 544.020 1982.750 547.020 2599.000 ;
        RECT 381.040 1710.640 382.640 1969.520 ;
        RECT 364.020 -9.320 367.020 1699.000 ;
        RECT 544.020 -9.320 547.020 1699.000 ;
        RECT 724.020 1001.000 727.020 3529.000 ;
        RECT 904.020 1001.000 907.020 3529.000 ;
        RECT 1084.020 2801.000 1087.020 3529.000 ;
        RECT 1019.545 2610.640 1021.145 2787.920 ;
        RECT 1084.020 2045.110 1087.020 2599.000 ;
        RECT 1264.020 2045.110 1267.020 3529.000 ;
        RECT 1021.040 1710.640 1022.640 2032.080 ;
        RECT 1084.020 1001.000 1087.020 1699.000 ;
        RECT 1264.020 1001.000 1267.020 1699.000 ;
        RECT 1444.020 1001.000 1447.020 3529.000 ;
        RECT 1624.020 2901.055 1627.020 3529.000 ;
        RECT 1804.020 2901.055 1807.020 3529.000 ;
        RECT 1521.040 2510.640 1522.640 2889.200 ;
        RECT 1624.020 1001.000 1627.020 2499.000 ;
        RECT 1804.020 1001.000 1807.020 2499.000 ;
        RECT 1984.020 1918.095 1987.020 3529.000 ;
        RECT 1948.870 1760.640 1950.470 1905.280 ;
        RECT 1984.020 1001.000 1987.020 1749.000 ;
        RECT 2164.020 1001.000 2167.020 3529.000 ;
        RECT 2344.020 1940.270 2347.020 3529.000 ;
        RECT 2524.020 2774.820 2527.020 3529.000 ;
        RECT 2427.190 2610.640 2428.790 2760.720 ;
        RECT 2524.020 1940.270 2527.020 2599.000 ;
        RECT 2321.040 1710.640 2322.640 1926.000 ;
        RECT 691.040 610.640 692.640 989.200 ;
        RECT 724.020 -9.320 727.020 599.000 ;
        RECT 904.020 -9.320 907.020 599.000 ;
        RECT 1084.020 -9.320 1087.020 599.000 ;
        RECT 1264.020 -9.320 1267.020 599.000 ;
        RECT 1444.020 -9.320 1447.020 599.000 ;
        RECT 1624.020 -9.320 1627.020 599.000 ;
        RECT 1804.020 -9.320 1807.020 599.000 ;
        RECT 1984.020 -9.320 1987.020 599.000 ;
        RECT 2164.020 -9.320 2167.020 599.000 ;
        RECT 2344.020 -9.320 2347.020 1699.000 ;
        RECT 2524.020 -9.320 2527.020 1699.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 457.855 2711.090 459.035 2712.270 ;
        RECT 457.855 2709.490 459.035 2710.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 381.250 1811.090 382.430 1812.270 ;
        RECT 381.250 1809.490 382.430 1810.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 1019.755 2711.090 1020.935 2712.270 ;
        RECT 1019.755 2709.490 1020.935 2710.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1521.250 2711.090 1522.430 2712.270 ;
        RECT 1521.250 2709.490 1522.430 2710.670 ;
        RECT 1521.250 2531.090 1522.430 2532.270 ;
        RECT 1521.250 2529.490 1522.430 2530.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 1021.250 1991.090 1022.430 1992.270 ;
        RECT 1021.250 1989.490 1022.430 1990.670 ;
        RECT 1021.250 1811.090 1022.430 1812.270 ;
        RECT 1021.250 1809.490 1022.430 1810.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1949.080 1811.090 1950.260 1812.270 ;
        RECT 1949.080 1809.490 1950.260 1810.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2427.400 2711.090 2428.580 2712.270 ;
        RECT 2427.400 2709.490 2428.580 2710.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 2321.250 1811.090 2322.430 1812.270 ;
        RECT 2321.250 1809.490 2322.430 1810.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 691.250 911.090 692.430 912.270 ;
        RECT 691.250 909.490 692.430 910.670 ;
        RECT 691.250 731.090 692.430 732.270 ;
        RECT 691.250 729.490 692.430 730.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 457.645 2712.380 459.245 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1019.545 2712.380 1021.145 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1521.040 2712.380 1522.640 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2427.190 2712.380 2428.790 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 457.645 2709.370 459.245 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1019.545 2709.370 1021.145 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1521.040 2709.370 1522.640 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2427.190 2709.370 2428.790 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1521.040 2532.380 1522.640 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1521.040 2529.370 1522.640 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1021.040 1992.380 1022.640 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1021.040 1989.370 1022.640 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 381.040 1812.380 382.640 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1021.040 1812.380 1022.640 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1948.870 1812.380 1950.470 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2321.040 1812.380 2322.640 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 381.040 1809.370 382.640 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1021.040 1809.370 1022.640 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1948.870 1809.370 1950.470 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2321.040 1809.370 2322.640 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 691.040 912.380 692.640 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 691.040 909.370 692.640 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 691.040 732.380 692.640 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 691.040 729.370 692.640 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 2760.520 457.020 3529.000 ;
        RECT 480.565 2610.640 482.165 2747.120 ;
        RECT 454.020 1982.750 457.020 2599.000 ;
        RECT 457.840 1710.640 459.440 1969.520 ;
        RECT 454.020 -9.320 457.020 1699.000 ;
        RECT 634.020 -9.320 637.020 3529.000 ;
        RECT 814.020 1001.000 817.020 3529.000 ;
        RECT 994.020 1001.000 997.020 3529.000 ;
        RECT 1034.375 2610.640 1035.975 2787.920 ;
        RECT 1174.020 2045.110 1177.020 3529.000 ;
        RECT 1097.840 1710.640 1099.440 2032.080 ;
        RECT 1174.020 1001.000 1177.020 1699.000 ;
        RECT 1354.020 1001.000 1357.020 3529.000 ;
        RECT 1534.020 2901.055 1537.020 3529.000 ;
        RECT 1714.020 2901.055 1717.020 3529.000 ;
        RECT 1597.840 2510.640 1599.440 2889.200 ;
        RECT 1534.020 1001.000 1537.020 2499.000 ;
        RECT 1714.020 1001.000 1717.020 2499.000 ;
        RECT 1894.020 1001.000 1897.020 3529.000 ;
        RECT 2074.020 1918.095 2077.020 3529.000 ;
        RECT 1973.020 1760.640 1974.620 1905.280 ;
        RECT 2074.020 1001.000 2077.020 1749.000 ;
        RECT 767.840 610.640 769.440 989.200 ;
        RECT 814.020 -9.320 817.020 599.000 ;
        RECT 994.020 -9.320 997.020 599.000 ;
        RECT 1174.020 -9.320 1177.020 599.000 ;
        RECT 1354.020 -9.320 1357.020 599.000 ;
        RECT 1534.020 -9.320 1537.020 599.000 ;
        RECT 1714.020 -9.320 1717.020 599.000 ;
        RECT 1894.020 -9.320 1897.020 599.000 ;
        RECT 2074.020 -9.320 2077.020 599.000 ;
        RECT 2254.020 -9.320 2257.020 3529.000 ;
        RECT 2434.020 2774.820 2437.020 3529.000 ;
        RECT 2452.490 2610.640 2454.090 2760.720 ;
        RECT 2434.020 1940.270 2437.020 2599.000 ;
        RECT 2397.840 1710.640 2399.440 1926.000 ;
        RECT 2434.020 -9.320 2437.020 1699.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 480.775 2621.090 481.955 2622.270 ;
        RECT 480.775 2619.490 481.955 2620.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 458.050 1901.090 459.230 1902.270 ;
        RECT 458.050 1899.490 459.230 1900.670 ;
        RECT 458.050 1721.090 459.230 1722.270 ;
        RECT 458.050 1719.490 459.230 1720.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 1034.585 2621.090 1035.765 2622.270 ;
        RECT 1034.585 2619.490 1035.765 2620.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1598.050 2801.090 1599.230 2802.270 ;
        RECT 1598.050 2799.490 1599.230 2800.670 ;
        RECT 1598.050 2621.090 1599.230 2622.270 ;
        RECT 1598.050 2619.490 1599.230 2620.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 1098.050 1901.090 1099.230 1902.270 ;
        RECT 1098.050 1899.490 1099.230 1900.670 ;
        RECT 1098.050 1721.090 1099.230 1722.270 ;
        RECT 1098.050 1719.490 1099.230 1720.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2452.700 2621.090 2453.880 2622.270 ;
        RECT 2452.700 2619.490 2453.880 2620.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1973.230 1901.090 1974.410 1902.270 ;
        RECT 1973.230 1899.490 1974.410 1900.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2398.050 1901.090 2399.230 1902.270 ;
        RECT 2398.050 1899.490 2399.230 1900.670 ;
        RECT 2398.050 1721.090 2399.230 1722.270 ;
        RECT 2398.050 1719.490 2399.230 1720.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 768.050 821.090 769.230 822.270 ;
        RECT 768.050 819.490 769.230 820.670 ;
        RECT 768.050 641.090 769.230 642.270 ;
        RECT 768.050 639.490 769.230 640.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1597.840 2802.380 1599.440 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1597.840 2799.370 1599.440 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 480.565 2622.380 482.165 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1034.375 2622.380 1035.975 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1597.840 2622.380 1599.440 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2452.490 2622.380 2454.090 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 480.565 2619.370 482.165 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1034.375 2619.370 1035.975 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1597.840 2619.370 1599.440 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2452.490 2619.370 2454.090 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 457.840 1902.380 459.440 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1097.840 1902.380 1099.440 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 1973.020 1902.380 1974.620 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2397.840 1902.380 2399.440 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 457.840 1899.370 459.440 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1097.840 1899.370 1099.440 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 1973.020 1899.370 1974.620 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2397.840 1899.370 2399.440 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 457.840 1722.380 459.440 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1097.840 1722.380 1099.440 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2397.840 1722.380 2399.440 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 457.840 1719.370 459.440 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1097.840 1719.370 1099.440 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2397.840 1719.370 2399.440 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 767.840 822.380 769.440 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 767.840 819.370 769.440 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 767.840 642.380 769.440 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 767.840 639.370 769.440 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 382.020 1982.750 385.020 3538.400 ;
        RECT 562.020 2760.520 565.020 3538.400 ;
        RECT 562.020 1982.750 565.020 2599.000 ;
        RECT 382.020 -18.720 385.020 1699.000 ;
        RECT 562.020 -18.720 565.020 1699.000 ;
        RECT 742.020 1001.000 745.020 3538.400 ;
        RECT 922.020 1001.000 925.020 3538.400 ;
        RECT 1102.020 2045.110 1105.020 3538.400 ;
        RECT 1282.020 2045.110 1285.020 3538.400 ;
        RECT 1102.020 1001.000 1105.020 1699.000 ;
        RECT 1282.020 1001.000 1285.020 1699.000 ;
        RECT 1462.020 1001.000 1465.020 3538.400 ;
        RECT 1642.020 2901.055 1645.020 3538.400 ;
        RECT 1822.020 2901.055 1825.020 3538.400 ;
        RECT 1642.020 1001.000 1645.020 2499.000 ;
        RECT 1822.020 1001.000 1825.020 2499.000 ;
        RECT 2002.020 1918.095 2005.020 3538.400 ;
        RECT 2002.020 1001.000 2005.020 1749.000 ;
        RECT 742.020 -18.720 745.020 599.000 ;
        RECT 922.020 -18.720 925.020 599.000 ;
        RECT 1102.020 -18.720 1105.020 599.000 ;
        RECT 1282.020 -18.720 1285.020 599.000 ;
        RECT 1462.020 -18.720 1465.020 599.000 ;
        RECT 1642.020 -18.720 1645.020 599.000 ;
        RECT 1822.020 -18.720 1825.020 599.000 ;
        RECT 2002.020 -18.720 2005.020 599.000 ;
        RECT 2182.020 -18.720 2185.020 3538.400 ;
        RECT 2362.020 1940.270 2365.020 3538.400 ;
        RECT 2542.020 2774.820 2545.020 3538.400 ;
        RECT 2362.020 -18.720 2365.020 1699.000 ;
        RECT 2542.020 -18.720 2545.020 2599.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 292.020 -18.720 295.020 3538.400 ;
        RECT 472.020 2760.520 475.020 3538.400 ;
        RECT 472.020 1982.750 475.020 2599.000 ;
        RECT 472.020 -18.720 475.020 1699.000 ;
        RECT 652.020 -18.720 655.020 3538.400 ;
        RECT 832.020 1001.000 835.020 3538.400 ;
        RECT 1012.020 2801.000 1015.020 3538.400 ;
        RECT 1012.020 2045.110 1015.020 2599.000 ;
        RECT 1192.020 2045.110 1195.020 3538.400 ;
        RECT 1012.020 1001.000 1015.020 1699.000 ;
        RECT 1192.020 1001.000 1195.020 1699.000 ;
        RECT 1372.020 1001.000 1375.020 3538.400 ;
        RECT 1552.020 2901.055 1555.020 3538.400 ;
        RECT 1732.020 2901.055 1735.020 3538.400 ;
        RECT 1552.020 1001.000 1555.020 2499.000 ;
        RECT 1732.020 1001.000 1735.020 2499.000 ;
        RECT 1912.020 1001.000 1915.020 3538.400 ;
        RECT 2092.020 1001.000 2095.020 3538.400 ;
        RECT 832.020 -18.720 835.020 599.000 ;
        RECT 1012.020 -18.720 1015.020 599.000 ;
        RECT 1192.020 -18.720 1195.020 599.000 ;
        RECT 1372.020 -18.720 1375.020 599.000 ;
        RECT 1552.020 -18.720 1555.020 599.000 ;
        RECT 1732.020 -18.720 1735.020 599.000 ;
        RECT 1912.020 -18.720 1915.020 599.000 ;
        RECT 2092.020 -18.720 2095.020 599.000 ;
        RECT 2272.020 -18.720 2275.020 3538.400 ;
        RECT 2452.020 2774.820 2455.020 3538.400 ;
        RECT 2452.020 1940.270 2455.020 2599.000 ;
        RECT 2452.020 -18.720 2455.020 1699.000 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 400.020 1982.750 403.020 3547.800 ;
        RECT 580.020 1982.750 583.020 3547.800 ;
        RECT 400.020 -28.120 403.020 1699.000 ;
        RECT 580.020 -28.120 583.020 1699.000 ;
        RECT 760.020 1001.000 763.020 3547.800 ;
        RECT 940.020 1001.000 943.020 3547.800 ;
        RECT 1120.020 2045.110 1123.020 3547.800 ;
        RECT 1300.020 2045.110 1303.020 3547.800 ;
        RECT 1120.020 1001.000 1123.020 1699.000 ;
        RECT 1300.020 1001.000 1303.020 1699.000 ;
        RECT 1480.020 1001.000 1483.020 3547.800 ;
        RECT 1660.020 2901.055 1663.020 3547.800 ;
        RECT 1840.020 2901.055 1843.020 3547.800 ;
        RECT 1660.020 1001.000 1663.020 2499.000 ;
        RECT 1840.020 1001.000 1843.020 2499.000 ;
        RECT 2020.020 1918.095 2023.020 3547.800 ;
        RECT 2020.020 1001.000 2023.020 1749.000 ;
        RECT 760.020 -28.120 763.020 599.000 ;
        RECT 940.020 -28.120 943.020 599.000 ;
        RECT 1120.020 -28.120 1123.020 599.000 ;
        RECT 1300.020 -28.120 1303.020 599.000 ;
        RECT 1480.020 -28.120 1483.020 599.000 ;
        RECT 1660.020 -28.120 1663.020 599.000 ;
        RECT 1840.020 -28.120 1843.020 599.000 ;
        RECT 2020.020 -28.120 2023.020 599.000 ;
        RECT 2200.020 -28.120 2203.020 3547.800 ;
        RECT 2380.020 1940.270 2383.020 3547.800 ;
        RECT 2380.020 -28.120 2383.020 1699.000 ;
        RECT 2560.020 -28.120 2563.020 3547.800 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 310.020 -28.120 313.020 3547.800 ;
        RECT 490.020 2760.520 493.020 3547.800 ;
        RECT 490.020 1982.750 493.020 2599.000 ;
        RECT 490.020 -28.120 493.020 1699.000 ;
        RECT 670.020 1001.000 673.020 3547.800 ;
        RECT 850.020 1001.000 853.020 3547.800 ;
        RECT 1030.020 2801.000 1033.020 3547.800 ;
        RECT 1030.020 2045.110 1033.020 2599.000 ;
        RECT 1210.020 2045.110 1213.020 3547.800 ;
        RECT 1030.020 1001.000 1033.020 1699.000 ;
        RECT 1210.020 1001.000 1213.020 1699.000 ;
        RECT 1390.020 1001.000 1393.020 3547.800 ;
        RECT 1570.020 2901.055 1573.020 3547.800 ;
        RECT 1750.020 2901.055 1753.020 3547.800 ;
        RECT 1570.020 1001.000 1573.020 2499.000 ;
        RECT 1750.020 1001.000 1753.020 2499.000 ;
        RECT 1930.020 1918.095 1933.020 3547.800 ;
        RECT 1930.020 1001.000 1933.020 1749.000 ;
        RECT 2110.020 1001.000 2113.020 3547.800 ;
        RECT 670.020 -28.120 673.020 599.000 ;
        RECT 850.020 -28.120 853.020 599.000 ;
        RECT 1030.020 -28.120 1033.020 599.000 ;
        RECT 1210.020 -28.120 1213.020 599.000 ;
        RECT 1390.020 -28.120 1393.020 599.000 ;
        RECT 1570.020 -28.120 1573.020 599.000 ;
        RECT 1750.020 -28.120 1753.020 599.000 ;
        RECT 1930.020 -28.120 1933.020 599.000 ;
        RECT 2110.020 -28.120 2113.020 599.000 ;
        RECT 2290.020 -28.120 2293.020 3547.800 ;
        RECT 2470.020 2774.820 2473.020 3547.800 ;
        RECT 2470.020 1940.270 2473.020 2599.000 ;
        RECT 2470.020 -28.120 2473.020 1699.000 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 418.020 1982.750 421.020 3557.200 ;
        RECT 598.020 1982.750 601.020 3557.200 ;
        RECT 418.020 -37.520 421.020 1699.000 ;
        RECT 598.020 -37.520 601.020 1699.000 ;
        RECT 778.020 1001.000 781.020 3557.200 ;
        RECT 958.020 1001.000 961.020 3557.200 ;
        RECT 1138.020 2045.110 1141.020 3557.200 ;
        RECT 1318.020 2045.110 1321.020 3557.200 ;
        RECT 1498.020 2901.055 1501.020 3557.200 ;
        RECT 1678.020 2901.055 1681.020 3557.200 ;
        RECT 1858.020 2901.055 1861.020 3557.200 ;
        RECT 1138.020 1001.000 1141.020 1699.000 ;
        RECT 1318.020 1001.000 1321.020 1699.000 ;
        RECT 1498.020 1001.000 1501.020 2499.000 ;
        RECT 1678.020 1001.000 1681.020 2499.000 ;
        RECT 1858.020 1001.000 1861.020 2499.000 ;
        RECT 2038.020 1918.095 2041.020 3557.200 ;
        RECT 2038.020 1001.000 2041.020 1749.000 ;
        RECT 778.020 -37.520 781.020 599.000 ;
        RECT 958.020 -37.520 961.020 599.000 ;
        RECT 1138.020 -37.520 1141.020 599.000 ;
        RECT 1318.020 -37.520 1321.020 599.000 ;
        RECT 1498.020 -37.520 1501.020 599.000 ;
        RECT 1678.020 -37.520 1681.020 599.000 ;
        RECT 1858.020 -37.520 1861.020 599.000 ;
        RECT 2038.020 -37.520 2041.020 599.000 ;
        RECT 2218.020 -37.520 2221.020 3557.200 ;
        RECT 2398.020 2774.820 2401.020 3557.200 ;
        RECT 2398.020 1940.270 2401.020 2599.000 ;
        RECT 2398.020 -37.520 2401.020 1699.000 ;
        RECT 2578.020 -37.520 2581.020 3557.200 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 328.020 -37.520 331.020 3557.200 ;
        RECT 508.020 2760.520 511.020 3557.200 ;
        RECT 508.020 1982.750 511.020 2599.000 ;
        RECT 508.020 -37.520 511.020 1699.000 ;
        RECT 688.020 1001.000 691.020 3557.200 ;
        RECT 868.020 1001.000 871.020 3557.200 ;
        RECT 1048.020 2801.000 1051.020 3557.200 ;
        RECT 1048.020 2045.110 1051.020 2599.000 ;
        RECT 1228.020 2045.110 1231.020 3557.200 ;
        RECT 1048.020 1001.000 1051.020 1699.000 ;
        RECT 1228.020 1001.000 1231.020 1699.000 ;
        RECT 1408.020 1001.000 1411.020 3557.200 ;
        RECT 1588.020 2901.055 1591.020 3557.200 ;
        RECT 1768.020 2901.055 1771.020 3557.200 ;
        RECT 1588.020 1001.000 1591.020 2499.000 ;
        RECT 1768.020 1001.000 1771.020 2499.000 ;
        RECT 1948.020 1918.095 1951.020 3557.200 ;
        RECT 1948.020 1001.000 1951.020 1749.000 ;
        RECT 2128.020 1001.000 2131.020 3557.200 ;
        RECT 2308.020 1940.270 2311.020 3557.200 ;
        RECT 2488.020 2774.820 2491.020 3557.200 ;
        RECT 2488.020 1940.270 2491.020 2599.000 ;
        RECT 688.020 -37.520 691.020 599.000 ;
        RECT 868.020 -37.520 871.020 599.000 ;
        RECT 1048.020 -37.520 1051.020 599.000 ;
        RECT 1228.020 -37.520 1231.020 599.000 ;
        RECT 1408.020 -37.520 1411.020 599.000 ;
        RECT 1588.020 -37.520 1591.020 599.000 ;
        RECT 1768.020 -37.520 1771.020 599.000 ;
        RECT 1948.020 -37.520 1951.020 599.000 ;
        RECT 2128.020 -37.520 2131.020 599.000 ;
        RECT 2308.020 -37.520 2311.020 1699.000 ;
        RECT 2488.020 -37.520 2491.020 1699.000 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 435.520 2610.795 573.060 2746.965 ;
        RECT 1005.520 2610.795 1094.300 2787.765 ;
        RECT 1505.520 2510.795 1884.415 2889.045 ;
        RECT 2402.690 2610.795 2554.490 2760.565 ;
        RECT 365.520 1710.795 625.420 1969.365 ;
        RECT 1005.520 1710.795 1327.520 2031.925 ;
        RECT 1925.520 1760.795 2070.420 1905.125 ;
        RECT 2305.520 1710.795 2522.640 1925.845 ;
        RECT 675.520 610.795 2164.080 998.055 ;
      LAYER met1 ;
        RECT 1351.090 2917.780 1351.410 2917.840 ;
        RECT 1535.090 2917.780 1535.410 2917.840 ;
        RECT 1351.090 2917.640 1535.410 2917.780 ;
        RECT 1351.090 2917.580 1351.410 2917.640 ;
        RECT 1535.090 2917.580 1535.410 2917.640 ;
        RECT 1501.510 2917.440 1501.830 2917.500 ;
        RECT 1546.130 2917.440 1546.450 2917.500 ;
        RECT 1501.510 2917.300 1546.450 2917.440 ;
        RECT 1501.510 2917.240 1501.830 2917.300 ;
        RECT 1546.130 2917.240 1546.450 2917.300 ;
        RECT 1414.110 2917.100 1414.430 2917.160 ;
        RECT 1567.290 2917.100 1567.610 2917.160 ;
        RECT 1414.110 2916.960 1567.610 2917.100 ;
        RECT 1414.110 2916.900 1414.430 2916.960 ;
        RECT 1567.290 2916.900 1567.610 2916.960 ;
        RECT 1479.890 2915.740 1480.210 2915.800 ;
        RECT 1641.810 2915.740 1642.130 2915.800 ;
        RECT 1479.890 2915.600 1642.130 2915.740 ;
        RECT 1479.890 2915.540 1480.210 2915.600 ;
        RECT 1641.810 2915.540 1642.130 2915.600 ;
        RECT 1495.530 2915.400 1495.850 2915.460 ;
        RECT 1705.290 2915.400 1705.610 2915.460 ;
        RECT 1495.530 2915.260 1705.610 2915.400 ;
        RECT 1495.530 2915.200 1495.850 2915.260 ;
        RECT 1705.290 2915.200 1705.610 2915.260 ;
        RECT 1379.610 2915.060 1379.930 2915.120 ;
        RECT 1598.570 2915.060 1598.890 2915.120 ;
        RECT 1379.610 2914.920 1598.890 2915.060 ;
        RECT 1379.610 2914.860 1379.930 2914.920 ;
        RECT 1598.570 2914.860 1598.890 2914.920 ;
        RECT 1407.210 2914.720 1407.530 2914.780 ;
        RECT 1630.770 2914.720 1631.090 2914.780 ;
        RECT 1407.210 2914.580 1631.090 2914.720 ;
        RECT 1407.210 2914.520 1407.530 2914.580 ;
        RECT 1630.770 2914.520 1631.090 2914.580 ;
        RECT 1461.490 2914.380 1461.810 2914.440 ;
        RECT 1694.250 2914.380 1694.570 2914.440 ;
        RECT 1461.490 2914.240 1694.570 2914.380 ;
        RECT 1461.490 2914.180 1461.810 2914.240 ;
        RECT 1694.250 2914.180 1694.570 2914.240 ;
        RECT 1494.610 2914.040 1494.930 2914.100 ;
        RECT 1768.770 2914.040 1769.090 2914.100 ;
        RECT 1494.610 2913.900 1769.090 2914.040 ;
        RECT 1494.610 2913.840 1494.930 2913.900 ;
        RECT 1768.770 2913.840 1769.090 2913.900 ;
        RECT 1789.930 2914.040 1790.250 2914.100 ;
        RECT 1895.270 2914.040 1895.590 2914.100 ;
        RECT 1789.930 2913.900 1895.590 2914.040 ;
        RECT 1789.930 2913.840 1790.250 2913.900 ;
        RECT 1895.270 2913.840 1895.590 2913.900 ;
        RECT 1501.970 2913.700 1502.290 2913.760 ;
        RECT 1812.010 2913.700 1812.330 2913.760 ;
        RECT 1501.970 2913.560 1812.330 2913.700 ;
        RECT 1501.970 2913.500 1502.290 2913.560 ;
        RECT 1812.010 2913.500 1812.330 2913.560 ;
        RECT 1372.710 2913.360 1373.030 2913.420 ;
        RECT 1843.290 2913.360 1843.610 2913.420 ;
        RECT 1372.710 2913.220 1843.610 2913.360 ;
        RECT 1372.710 2913.160 1373.030 2913.220 ;
        RECT 1843.290 2913.160 1843.610 2913.220 ;
        RECT 1493.690 2913.020 1494.010 2913.080 ;
        RECT 1800.970 2913.020 1801.290 2913.080 ;
        RECT 1493.690 2912.880 1801.290 2913.020 ;
        RECT 1493.690 2912.820 1494.010 2912.880 ;
        RECT 1800.970 2912.820 1801.290 2912.880 ;
        RECT 1833.170 2913.020 1833.490 2913.080 ;
        RECT 1887.450 2913.020 1887.770 2913.080 ;
        RECT 1833.170 2912.880 1887.770 2913.020 ;
        RECT 1833.170 2912.820 1833.490 2912.880 ;
        RECT 1887.450 2912.820 1887.770 2912.880 ;
        RECT 1496.910 2912.680 1497.230 2912.740 ;
        RECT 1662.970 2912.680 1663.290 2912.740 ;
        RECT 1496.910 2912.540 1663.290 2912.680 ;
        RECT 1496.910 2912.480 1497.230 2912.540 ;
        RECT 1662.970 2912.480 1663.290 2912.540 ;
        RECT 1854.330 2912.680 1854.650 2912.740 ;
        RECT 1886.530 2912.680 1886.850 2912.740 ;
        RECT 1854.330 2912.540 1886.850 2912.680 ;
        RECT 1854.330 2912.480 1854.650 2912.540 ;
        RECT 1886.530 2912.480 1886.850 2912.540 ;
        RECT 1495.070 2912.340 1495.390 2912.400 ;
        RECT 1609.610 2912.340 1609.930 2912.400 ;
        RECT 1495.070 2912.200 1609.930 2912.340 ;
        RECT 1495.070 2912.140 1495.390 2912.200 ;
        RECT 1609.610 2912.140 1609.930 2912.200 ;
        RECT 1351.090 2911.800 1351.410 2912.060 ;
        RECT 1502.430 2912.000 1502.750 2912.060 ;
        RECT 1779.810 2912.000 1780.130 2912.060 ;
        RECT 1502.430 2911.860 1780.130 2912.000 ;
        RECT 1502.430 2911.800 1502.750 2911.860 ;
        RECT 1779.810 2911.800 1780.130 2911.860 ;
        RECT 1864.450 2912.000 1864.770 2912.060 ;
        RECT 1894.810 2912.000 1895.130 2912.060 ;
        RECT 1864.450 2911.860 1895.130 2912.000 ;
        RECT 1864.450 2911.800 1864.770 2911.860 ;
        RECT 1894.810 2911.800 1895.130 2911.860 ;
        RECT 1351.180 2911.380 1351.320 2911.800 ;
        RECT 1351.090 2911.120 1351.410 2911.380 ;
        RECT 1455.510 2901.120 1455.830 2901.180 ;
        RECT 1758.650 2901.120 1758.970 2901.180 ;
        RECT 1455.510 2900.980 1758.970 2901.120 ;
        RECT 1455.510 2900.920 1455.830 2900.980 ;
        RECT 1758.650 2900.920 1758.970 2900.980 ;
        RECT 1496.450 2898.400 1496.770 2898.460 ;
        RECT 1524.050 2898.400 1524.370 2898.460 ;
        RECT 1496.450 2898.260 1524.370 2898.400 ;
        RECT 1496.450 2898.200 1496.770 2898.260 ;
        RECT 1524.050 2898.200 1524.370 2898.260 ;
        RECT 1497.370 2896.700 1497.690 2896.760 ;
        RECT 1503.350 2896.700 1503.670 2896.760 ;
        RECT 1497.370 2896.560 1503.670 2896.700 ;
        RECT 1497.370 2896.500 1497.690 2896.560 ;
        RECT 1503.350 2896.500 1503.670 2896.560 ;
        RECT 1876.870 2896.700 1877.190 2896.760 ;
        RECT 1887.910 2896.700 1888.230 2896.760 ;
        RECT 1876.870 2896.560 1888.230 2896.700 ;
        RECT 1876.870 2896.500 1877.190 2896.560 ;
        RECT 1887.910 2896.500 1888.230 2896.560 ;
        RECT 1351.090 2849.920 1351.410 2850.180 ;
        RECT 1351.180 2849.500 1351.320 2849.920 ;
        RECT 1357.990 2849.780 1358.310 2849.840 ;
        RECT 1490.010 2849.780 1490.330 2849.840 ;
        RECT 1357.990 2849.640 1490.330 2849.780 ;
        RECT 1357.990 2849.580 1358.310 2849.640 ;
        RECT 1490.010 2849.580 1490.330 2849.640 ;
        RECT 1351.090 2849.240 1351.410 2849.500 ;
        RECT 1350.630 2842.980 1350.950 2843.040 ;
        RECT 1351.090 2842.980 1351.410 2843.040 ;
        RECT 1350.630 2842.840 1351.410 2842.980 ;
        RECT 1350.630 2842.780 1350.950 2842.840 ;
        RECT 1351.090 2842.780 1351.410 2842.840 ;
        RECT 1476.210 2829.380 1476.530 2829.440 ;
        RECT 1490.010 2829.380 1490.330 2829.440 ;
        RECT 1476.210 2829.240 1490.330 2829.380 ;
        RECT 1476.210 2829.180 1476.530 2829.240 ;
        RECT 1490.010 2829.180 1490.330 2829.240 ;
        RECT 1000.570 2810.680 1000.890 2810.740 ;
        RECT 1048.410 2810.680 1048.730 2810.740 ;
        RECT 1000.570 2810.540 1048.730 2810.680 ;
        RECT 1000.570 2810.480 1000.890 2810.540 ;
        RECT 1048.410 2810.480 1048.730 2810.540 ;
        RECT 985.390 2810.340 985.710 2810.400 ;
        RECT 1073.710 2810.340 1074.030 2810.400 ;
        RECT 985.390 2810.200 1074.030 2810.340 ;
        RECT 985.390 2810.140 985.710 2810.200 ;
        RECT 1073.710 2810.140 1074.030 2810.200 ;
        RECT 978.490 2810.000 978.810 2810.060 ;
        RECT 1027.710 2810.000 1028.030 2810.060 ;
        RECT 978.490 2809.860 1028.030 2810.000 ;
        RECT 978.490 2809.800 978.810 2809.860 ;
        RECT 1027.710 2809.800 1028.030 2809.860 ;
        RECT 978.950 2809.660 979.270 2809.720 ;
        RECT 1043.350 2809.660 1043.670 2809.720 ;
        RECT 978.950 2809.520 1043.670 2809.660 ;
        RECT 978.950 2809.460 979.270 2809.520 ;
        RECT 1043.350 2809.460 1043.670 2809.520 ;
        RECT 985.850 2809.320 986.170 2809.380 ;
        RECT 1058.070 2809.320 1058.390 2809.380 ;
        RECT 985.850 2809.180 1058.390 2809.320 ;
        RECT 985.850 2809.120 986.170 2809.180 ;
        RECT 1058.070 2809.120 1058.390 2809.180 ;
        RECT 979.410 2808.980 979.730 2809.040 ;
        RECT 1000.570 2808.980 1000.890 2809.040 ;
        RECT 979.410 2808.840 1000.890 2808.980 ;
        RECT 979.410 2808.780 979.730 2808.840 ;
        RECT 1000.570 2808.780 1000.890 2808.840 ;
        RECT 1048.410 2808.640 1048.730 2808.700 ;
        RECT 1089.350 2808.640 1089.670 2808.700 ;
        RECT 1048.410 2808.500 1089.670 2808.640 ;
        RECT 1048.410 2808.440 1048.730 2808.500 ;
        RECT 1089.350 2808.440 1089.670 2808.500 ;
        RECT 986.310 2801.160 986.630 2801.220 ;
        RECT 1010.230 2801.160 1010.550 2801.220 ;
        RECT 986.310 2801.020 1010.550 2801.160 ;
        RECT 986.310 2800.960 986.630 2801.020 ;
        RECT 1010.230 2800.960 1010.550 2801.020 ;
        RECT 1351.550 2795.040 1351.870 2795.100 ;
        RECT 1352.930 2795.040 1353.250 2795.100 ;
        RECT 1351.550 2794.900 1353.250 2795.040 ;
        RECT 1351.550 2794.840 1351.870 2794.900 ;
        RECT 1352.930 2794.840 1353.250 2794.900 ;
        RECT 445.810 2769.540 446.130 2769.600 ;
        RECT 796.790 2769.540 797.110 2769.600 ;
        RECT 445.810 2769.400 797.110 2769.540 ;
        RECT 445.810 2769.340 446.130 2769.400 ;
        RECT 796.790 2769.340 797.110 2769.400 ;
        RECT 532.290 2768.180 532.610 2768.240 ;
        RECT 707.090 2768.180 707.410 2768.240 ;
        RECT 532.290 2768.040 707.410 2768.180 ;
        RECT 532.290 2767.980 532.610 2768.040 ;
        RECT 707.090 2767.980 707.410 2768.040 ;
        RECT 518.490 2767.840 518.810 2767.900 ;
        RECT 755.390 2767.840 755.710 2767.900 ;
        RECT 518.490 2767.700 755.710 2767.840 ;
        RECT 518.490 2767.640 518.810 2767.700 ;
        RECT 755.390 2767.640 755.710 2767.700 ;
        RECT 489.050 2767.500 489.370 2767.560 ;
        RECT 769.190 2767.500 769.510 2767.560 ;
        RECT 489.050 2767.360 769.510 2767.500 ;
        RECT 489.050 2767.300 489.370 2767.360 ;
        RECT 769.190 2767.300 769.510 2767.360 ;
      LAYER met1 ;
        RECT 432.830 2606.500 575.750 2752.620 ;
      LAYER met1 ;
        RECT 588.870 2684.200 589.190 2684.260 ;
        RECT 720.890 2684.200 721.210 2684.260 ;
        RECT 588.870 2684.060 721.210 2684.200 ;
        RECT 588.870 2684.000 589.190 2684.060 ;
        RECT 720.890 2684.000 721.210 2684.060 ;
        RECT 588.870 2663.800 589.190 2663.860 ;
        RECT 789.890 2663.800 790.210 2663.860 ;
        RECT 588.870 2663.660 790.210 2663.800 ;
        RECT 588.870 2663.600 589.190 2663.660 ;
        RECT 789.890 2663.600 790.210 2663.660 ;
        RECT 978.030 2644.080 978.350 2644.140 ;
        RECT 987.230 2644.080 987.550 2644.140 ;
        RECT 978.030 2643.940 987.550 2644.080 ;
        RECT 978.030 2643.880 978.350 2643.940 ;
        RECT 987.230 2643.880 987.550 2643.940 ;
      LAYER met1 ;
        RECT 1002.830 2610.640 1095.150 2787.920 ;
      LAYER met1 ;
        RECT 1358.450 2781.100 1358.770 2781.160 ;
        RECT 1485.410 2781.100 1485.730 2781.160 ;
        RECT 1358.450 2780.960 1485.730 2781.100 ;
        RECT 1358.450 2780.900 1358.770 2780.960 ;
        RECT 1485.410 2780.900 1485.730 2780.960 ;
        RECT 1351.550 2767.500 1351.870 2767.560 ;
        RECT 1351.180 2767.360 1351.870 2767.500 ;
        RECT 1351.180 2766.880 1351.320 2767.360 ;
        RECT 1351.550 2767.300 1351.870 2767.360 ;
        RECT 1351.090 2766.620 1351.410 2766.880 ;
        RECT 1350.630 2739.280 1350.950 2739.340 ;
        RECT 1351.090 2739.280 1351.410 2739.340 ;
        RECT 1350.630 2739.140 1351.410 2739.280 ;
        RECT 1350.630 2739.080 1350.950 2739.140 ;
        RECT 1351.090 2739.080 1351.410 2739.140 ;
        RECT 1350.170 2691.340 1350.490 2691.400 ;
        RECT 1350.630 2691.340 1350.950 2691.400 ;
        RECT 1350.170 2691.200 1350.950 2691.340 ;
        RECT 1350.170 2691.140 1350.490 2691.200 ;
        RECT 1350.630 2691.140 1350.950 2691.200 ;
        RECT 1434.350 2691.340 1434.670 2691.400 ;
        RECT 1489.090 2691.340 1489.410 2691.400 ;
        RECT 1434.350 2691.200 1489.410 2691.340 ;
        RECT 1434.350 2691.140 1434.670 2691.200 ;
        RECT 1489.090 2691.140 1489.410 2691.200 ;
        RECT 1350.170 2670.260 1350.490 2670.320 ;
        RECT 1351.090 2670.260 1351.410 2670.320 ;
        RECT 1350.170 2670.120 1351.410 2670.260 ;
        RECT 1350.170 2670.060 1350.490 2670.120 ;
        RECT 1351.090 2670.060 1351.410 2670.120 ;
        RECT 1351.090 2622.460 1351.410 2622.720 ;
        RECT 1351.180 2622.040 1351.320 2622.460 ;
        RECT 1351.090 2621.780 1351.410 2622.040 ;
        RECT 1393.410 2608.380 1393.730 2608.440 ;
        RECT 1488.630 2608.380 1488.950 2608.440 ;
        RECT 1393.410 2608.240 1488.950 2608.380 ;
        RECT 1393.410 2608.180 1393.730 2608.240 ;
        RECT 1488.630 2608.180 1488.950 2608.240 ;
        RECT 999.190 2605.660 999.510 2605.720 ;
        RECT 1111.890 2605.660 1112.210 2605.720 ;
        RECT 999.190 2605.520 1112.210 2605.660 ;
        RECT 999.190 2605.460 999.510 2605.520 ;
        RECT 1111.890 2605.460 1112.210 2605.520 ;
        RECT 999.650 2605.320 999.970 2605.380 ;
        RECT 1112.810 2605.320 1113.130 2605.380 ;
        RECT 999.650 2605.180 1113.130 2605.320 ;
        RECT 999.650 2605.120 999.970 2605.180 ;
        RECT 1112.810 2605.120 1113.130 2605.180 ;
        RECT 982.170 2604.980 982.490 2605.040 ;
        RECT 1113.270 2604.980 1113.590 2605.040 ;
        RECT 982.170 2604.840 1113.590 2604.980 ;
        RECT 982.170 2604.780 982.490 2604.840 ;
        RECT 1113.270 2604.780 1113.590 2604.840 ;
        RECT 975.270 2604.640 975.590 2604.700 ;
        RECT 1112.350 2604.640 1112.670 2604.700 ;
        RECT 975.270 2604.500 1112.670 2604.640 ;
        RECT 975.270 2604.440 975.590 2604.500 ;
        RECT 1112.350 2604.440 1112.670 2604.500 ;
        RECT 1392.950 2594.780 1393.270 2594.840 ;
        RECT 1488.170 2594.780 1488.490 2594.840 ;
        RECT 1392.950 2594.640 1488.490 2594.780 ;
        RECT 1392.950 2594.580 1393.270 2594.640 ;
        RECT 1488.170 2594.580 1488.490 2594.640 ;
        RECT 533.210 2591.720 533.530 2591.780 ;
        RECT 762.290 2591.720 762.610 2591.780 ;
        RECT 533.210 2591.580 762.610 2591.720 ;
        RECT 533.210 2591.520 533.530 2591.580 ;
        RECT 762.290 2591.520 762.610 2591.580 ;
        RECT 984.930 2591.720 985.250 2591.780 ;
        RECT 1048.870 2591.720 1049.190 2591.780 ;
        RECT 984.930 2591.580 1049.190 2591.720 ;
        RECT 984.930 2591.520 985.250 2591.580 ;
        RECT 1048.870 2591.520 1049.190 2591.580 ;
        RECT 504.690 2591.380 505.010 2591.440 ;
        RECT 782.990 2591.380 783.310 2591.440 ;
        RECT 504.690 2591.240 783.310 2591.380 ;
        RECT 504.690 2591.180 505.010 2591.240 ;
        RECT 782.990 2591.180 783.310 2591.240 ;
        RECT 974.810 2591.380 975.130 2591.440 ;
        RECT 1094.870 2591.380 1095.190 2591.440 ;
        RECT 974.810 2591.240 1095.190 2591.380 ;
        RECT 974.810 2591.180 975.130 2591.240 ;
        RECT 1094.870 2591.180 1095.190 2591.240 ;
        RECT 1028.170 2587.640 1028.490 2587.700 ;
        RECT 1033.230 2587.640 1033.550 2587.700 ;
        RECT 1028.170 2587.500 1033.550 2587.640 ;
        RECT 1028.170 2587.440 1028.490 2587.500 ;
        RECT 1033.230 2587.440 1033.550 2587.500 ;
        RECT 1413.650 2580.840 1413.970 2580.900 ;
        RECT 1488.170 2580.840 1488.490 2580.900 ;
        RECT 1413.650 2580.700 1488.490 2580.840 ;
        RECT 1413.650 2580.640 1413.970 2580.700 ;
        RECT 1488.170 2580.640 1488.490 2580.700 ;
        RECT 1468.850 2546.500 1469.170 2546.560 ;
        RECT 1484.490 2546.500 1484.810 2546.560 ;
        RECT 1468.850 2546.360 1484.810 2546.500 ;
        RECT 1468.850 2546.300 1469.170 2546.360 ;
        RECT 1484.490 2546.300 1484.810 2546.360 ;
        RECT 1350.170 2511.820 1350.490 2511.880 ;
        RECT 1352.010 2511.820 1352.330 2511.880 ;
        RECT 1350.170 2511.680 1352.330 2511.820 ;
        RECT 1350.170 2511.620 1350.490 2511.680 ;
        RECT 1352.010 2511.620 1352.330 2511.680 ;
      LAYER met1 ;
        RECT 1502.830 2504.460 1885.870 2889.200 ;
      LAYER met1 ;
        RECT 2093.990 2781.440 2094.310 2781.500 ;
        RECT 2556.290 2781.440 2556.610 2781.500 ;
        RECT 2093.990 2781.300 2556.610 2781.440 ;
        RECT 2093.990 2781.240 2094.310 2781.300 ;
        RECT 2556.290 2781.240 2556.610 2781.300 ;
        RECT 1893.890 2781.100 1894.210 2781.160 ;
        RECT 2421.970 2781.100 2422.290 2781.160 ;
        RECT 1893.890 2780.960 2422.290 2781.100 ;
        RECT 1893.890 2780.900 1894.210 2780.960 ;
        RECT 2421.970 2780.900 2422.290 2780.960 ;
      LAYER met1 ;
        RECT 2400.000 2610.640 2556.720 2760.720 ;
      LAYER met1 ;
        RECT 2528.690 2587.640 2529.010 2587.700 ;
        RECT 2534.210 2587.640 2534.530 2587.700 ;
        RECT 2528.690 2587.500 2534.530 2587.640 ;
        RECT 2528.690 2587.440 2529.010 2587.500 ;
        RECT 2534.210 2587.440 2534.530 2587.500 ;
        RECT 1621.110 2495.500 1621.430 2495.560 ;
        RECT 1895.270 2495.500 1895.590 2495.560 ;
        RECT 1621.110 2495.360 1895.590 2495.500 ;
        RECT 1621.110 2495.300 1621.430 2495.360 ;
        RECT 1895.270 2495.300 1895.590 2495.360 ;
        RECT 1495.530 2495.160 1495.850 2495.220 ;
        RECT 1552.570 2495.160 1552.890 2495.220 ;
        RECT 1495.530 2495.020 1552.890 2495.160 ;
        RECT 1495.530 2494.960 1495.850 2495.020 ;
        RECT 1552.570 2494.960 1552.890 2495.020 ;
        RECT 1600.410 2495.160 1600.730 2495.220 ;
        RECT 1887.910 2495.160 1888.230 2495.220 ;
        RECT 1600.410 2495.020 1888.230 2495.160 ;
        RECT 1600.410 2494.960 1600.730 2495.020 ;
        RECT 1887.910 2494.960 1888.230 2495.020 ;
        RECT 1501.970 2494.820 1502.290 2494.880 ;
        RECT 1559.470 2494.820 1559.790 2494.880 ;
        RECT 1501.970 2494.680 1559.790 2494.820 ;
        RECT 1501.970 2494.620 1502.290 2494.680 ;
        RECT 1559.470 2494.620 1559.790 2494.680 ;
        RECT 1586.610 2494.820 1586.930 2494.880 ;
        RECT 1887.450 2494.820 1887.770 2494.880 ;
        RECT 1586.610 2494.680 1887.770 2494.820 ;
        RECT 1586.610 2494.620 1586.930 2494.680 ;
        RECT 1887.450 2494.620 1887.770 2494.680 ;
        RECT 1495.070 2494.480 1495.390 2494.540 ;
        RECT 1514.850 2494.480 1515.170 2494.540 ;
        RECT 1495.070 2494.340 1515.170 2494.480 ;
        RECT 1495.070 2494.280 1495.390 2494.340 ;
        RECT 1514.850 2494.280 1515.170 2494.340 ;
        RECT 1544.290 2494.480 1544.610 2494.540 ;
        RECT 1894.810 2494.480 1895.130 2494.540 ;
        RECT 1544.290 2494.340 1895.130 2494.480 ;
        RECT 1544.290 2494.280 1544.610 2494.340 ;
        RECT 1894.810 2494.280 1895.130 2494.340 ;
        RECT 1494.610 2494.140 1494.930 2494.200 ;
        RECT 1573.730 2494.140 1574.050 2494.200 ;
        RECT 1494.610 2494.000 1574.050 2494.140 ;
        RECT 1494.610 2493.940 1494.930 2494.000 ;
        RECT 1573.730 2493.940 1574.050 2494.000 ;
        RECT 1869.510 2494.140 1869.830 2494.200 ;
        RECT 2394.370 2494.140 2394.690 2494.200 ;
        RECT 1869.510 2494.000 2394.690 2494.140 ;
        RECT 1869.510 2493.940 1869.830 2494.000 ;
        RECT 2394.370 2493.940 2394.690 2494.000 ;
        RECT 1501.510 2491.420 1501.830 2491.480 ;
        RECT 1504.270 2491.420 1504.590 2491.480 ;
        RECT 1501.510 2491.280 1504.590 2491.420 ;
        RECT 1501.510 2491.220 1501.830 2491.280 ;
        RECT 1504.270 2491.220 1504.590 2491.280 ;
        RECT 1679.530 2489.720 1679.850 2489.780 ;
        RECT 1683.210 2489.720 1683.530 2489.780 ;
        RECT 1679.530 2489.580 1683.530 2489.720 ;
        RECT 1679.530 2489.520 1679.850 2489.580 ;
        RECT 1683.210 2489.520 1683.530 2489.580 ;
        RECT 1593.510 2489.380 1593.830 2489.440 ;
        RECT 1778.890 2489.380 1779.210 2489.440 ;
        RECT 1593.510 2489.240 1779.210 2489.380 ;
        RECT 1593.510 2489.180 1593.830 2489.240 ;
        RECT 1778.890 2489.180 1779.210 2489.240 ;
        RECT 1645.490 2489.040 1645.810 2489.100 ;
        RECT 1789.930 2489.040 1790.250 2489.100 ;
        RECT 1645.490 2488.900 1790.250 2489.040 ;
        RECT 1645.490 2488.840 1645.810 2488.900 ;
        RECT 1789.930 2488.840 1790.250 2488.900 ;
        RECT 1421.010 2488.700 1421.330 2488.760 ;
        RECT 1842.370 2488.700 1842.690 2488.760 ;
        RECT 1421.010 2488.560 1842.690 2488.700 ;
        RECT 1421.010 2488.500 1421.330 2488.560 ;
        RECT 1842.370 2488.500 1842.690 2488.560 ;
        RECT 1455.050 2488.360 1455.370 2488.420 ;
        RECT 1885.610 2488.360 1885.930 2488.420 ;
        RECT 1455.050 2488.220 1885.930 2488.360 ;
        RECT 1455.050 2488.160 1455.370 2488.220 ;
        RECT 1885.610 2488.160 1885.930 2488.220 ;
        RECT 1420.550 2488.020 1420.870 2488.080 ;
        RECT 1874.570 2488.020 1874.890 2488.080 ;
        RECT 1420.550 2487.880 1874.890 2488.020 ;
        RECT 1420.550 2487.820 1420.870 2487.880 ;
        RECT 1874.570 2487.820 1874.890 2487.880 ;
        RECT 1448.610 2487.000 1448.930 2487.060 ;
        RECT 1832.250 2487.000 1832.570 2487.060 ;
        RECT 1448.610 2486.860 1832.570 2487.000 ;
        RECT 1448.610 2486.800 1448.930 2486.860 ;
        RECT 1832.250 2486.800 1832.570 2486.860 ;
        RECT 1454.590 2486.660 1454.910 2486.720 ;
        RECT 1757.730 2486.660 1758.050 2486.720 ;
        RECT 1454.590 2486.520 1758.050 2486.660 ;
        RECT 1454.590 2486.460 1454.910 2486.520 ;
        RECT 1757.730 2486.460 1758.050 2486.520 ;
        RECT 1427.910 2486.320 1428.230 2486.380 ;
        RECT 1725.530 2486.320 1725.850 2486.380 ;
        RECT 1427.910 2486.180 1725.850 2486.320 ;
        RECT 1427.910 2486.120 1428.230 2486.180 ;
        RECT 1725.530 2486.120 1725.850 2486.180 ;
        RECT 1528.190 2485.980 1528.510 2486.040 ;
        RECT 1811.090 2485.980 1811.410 2486.040 ;
        RECT 1528.190 2485.840 1811.410 2485.980 ;
        RECT 1528.190 2485.780 1528.510 2485.840 ;
        RECT 1811.090 2485.780 1811.410 2485.840 ;
        RECT 1386.510 2485.640 1386.830 2485.700 ;
        RECT 1587.530 2485.640 1587.850 2485.700 ;
        RECT 1386.510 2485.500 1587.850 2485.640 ;
        RECT 1386.510 2485.440 1386.830 2485.500 ;
        RECT 1587.530 2485.440 1587.850 2485.500 ;
        RECT 1397.090 2485.300 1397.410 2485.360 ;
        RECT 1534.170 2485.300 1534.490 2485.360 ;
        RECT 1397.090 2485.160 1534.490 2485.300 ;
        RECT 1397.090 2485.100 1397.410 2485.160 ;
        RECT 1534.170 2485.100 1534.490 2485.160 ;
        RECT 1572.350 2485.300 1572.670 2485.360 ;
        RECT 1746.690 2485.300 1747.010 2485.360 ;
        RECT 1572.350 2485.160 1747.010 2485.300 ;
        RECT 1572.350 2485.100 1572.670 2485.160 ;
        RECT 1746.690 2485.100 1747.010 2485.160 ;
        RECT 1441.710 2484.960 1442.030 2485.020 ;
        RECT 1608.690 2484.960 1609.010 2485.020 ;
        RECT 1441.710 2484.820 1609.010 2484.960 ;
        RECT 1441.710 2484.760 1442.030 2484.820 ;
        RECT 1608.690 2484.760 1609.010 2484.820 ;
        RECT 1535.090 2484.620 1535.410 2484.680 ;
        RECT 1576.490 2484.620 1576.810 2484.680 ;
        RECT 1535.090 2484.480 1576.810 2484.620 ;
        RECT 1535.090 2484.420 1535.410 2484.480 ;
        RECT 1576.490 2484.420 1576.810 2484.480 ;
        RECT 1545.210 2484.280 1545.530 2484.340 ;
        RECT 1548.890 2484.280 1549.210 2484.340 ;
        RECT 1545.210 2484.140 1549.210 2484.280 ;
        RECT 1545.210 2484.080 1545.530 2484.140 ;
        RECT 1548.890 2484.080 1549.210 2484.140 ;
        RECT 1610.990 2484.280 1611.310 2484.340 ;
        RECT 1619.730 2484.280 1620.050 2484.340 ;
        RECT 1610.990 2484.140 1620.050 2484.280 ;
        RECT 1610.990 2484.080 1611.310 2484.140 ;
        RECT 1619.730 2484.080 1620.050 2484.140 ;
        RECT 1673.090 2484.280 1673.410 2484.340 ;
        RECT 1679.530 2484.280 1679.850 2484.340 ;
        RECT 1673.090 2484.140 1679.850 2484.280 ;
        RECT 1673.090 2484.080 1673.410 2484.140 ;
        RECT 1679.530 2484.080 1679.850 2484.140 ;
        RECT 1679.990 2484.280 1680.310 2484.340 ;
        RECT 1715.410 2484.280 1715.730 2484.340 ;
        RECT 1679.990 2484.140 1715.730 2484.280 ;
        RECT 1679.990 2484.080 1680.310 2484.140 ;
        RECT 1715.410 2484.080 1715.730 2484.140 ;
        RECT 1351.090 2429.340 1351.410 2429.600 ;
        RECT 1351.180 2428.920 1351.320 2429.340 ;
        RECT 1532.330 2429.000 1532.650 2429.260 ;
        RECT 1351.090 2428.660 1351.410 2428.920 ;
        RECT 1532.420 2428.520 1532.560 2429.000 ;
        RECT 1532.790 2428.520 1533.110 2428.580 ;
        RECT 1532.420 2428.380 1533.110 2428.520 ;
        RECT 1532.790 2428.320 1533.110 2428.380 ;
        RECT 1544.290 2414.920 1544.610 2414.980 ;
        RECT 1545.210 2414.920 1545.530 2414.980 ;
        RECT 1544.290 2414.780 1545.530 2414.920 ;
        RECT 1544.290 2414.720 1544.610 2414.780 ;
        RECT 1545.210 2414.720 1545.530 2414.780 ;
        RECT 1351.090 2380.580 1351.410 2380.640 ;
        RECT 1351.550 2380.580 1351.870 2380.640 ;
        RECT 1351.090 2380.440 1351.870 2380.580 ;
        RECT 1351.090 2380.380 1351.410 2380.440 ;
        RECT 1351.550 2380.380 1351.870 2380.440 ;
        RECT 1545.210 2380.380 1545.530 2380.640 ;
        RECT 1544.750 2380.240 1545.070 2380.300 ;
        RECT 1545.300 2380.240 1545.440 2380.380 ;
        RECT 1544.750 2380.100 1545.440 2380.240 ;
        RECT 1544.750 2380.040 1545.070 2380.100 ;
        RECT 1351.090 2366.980 1351.410 2367.040 ;
        RECT 1351.550 2366.980 1351.870 2367.040 ;
        RECT 1351.090 2366.840 1351.870 2366.980 ;
        RECT 1351.090 2366.780 1351.410 2366.840 ;
        RECT 1351.550 2366.780 1351.870 2366.840 ;
        RECT 1531.870 2366.980 1532.190 2367.040 ;
        RECT 1533.250 2366.980 1533.570 2367.040 ;
        RECT 1531.870 2366.840 1533.570 2366.980 ;
        RECT 1531.870 2366.780 1532.190 2366.840 ;
        RECT 1533.250 2366.780 1533.570 2366.840 ;
        RECT 1532.330 2359.840 1532.650 2359.900 ;
        RECT 1533.250 2359.840 1533.570 2359.900 ;
        RECT 1532.330 2359.700 1533.570 2359.840 ;
        RECT 1532.330 2359.640 1532.650 2359.700 ;
        RECT 1533.250 2359.640 1533.570 2359.700 ;
        RECT 1351.090 2332.440 1351.410 2332.700 ;
        RECT 1351.180 2332.020 1351.320 2332.440 ;
        RECT 1544.290 2332.300 1544.610 2332.360 ;
        RECT 1545.210 2332.300 1545.530 2332.360 ;
        RECT 1544.290 2332.160 1545.530 2332.300 ;
        RECT 1544.290 2332.100 1544.610 2332.160 ;
        RECT 1545.210 2332.100 1545.530 2332.160 ;
        RECT 1351.090 2331.760 1351.410 2332.020 ;
        RECT 1533.250 2318.700 1533.570 2318.760 ;
        RECT 1532.880 2318.560 1533.570 2318.700 ;
        RECT 1532.880 2318.420 1533.020 2318.560 ;
        RECT 1533.250 2318.500 1533.570 2318.560 ;
        RECT 1532.790 2318.160 1533.110 2318.420 ;
        RECT 1543.830 2318.360 1544.150 2318.420 ;
        RECT 1544.290 2318.360 1544.610 2318.420 ;
        RECT 1543.830 2318.220 1544.610 2318.360 ;
        RECT 1543.830 2318.160 1544.150 2318.220 ;
        RECT 1544.290 2318.160 1544.610 2318.220 ;
        RECT 1559.010 2318.360 1559.330 2318.420 ;
        RECT 1559.470 2318.360 1559.790 2318.420 ;
        RECT 1559.010 2318.220 1559.790 2318.360 ;
        RECT 1559.010 2318.160 1559.330 2318.220 ;
        RECT 1559.470 2318.160 1559.790 2318.220 ;
        RECT 1350.170 2294.220 1350.490 2294.280 ;
        RECT 1351.090 2294.220 1351.410 2294.280 ;
        RECT 1350.170 2294.080 1351.410 2294.220 ;
        RECT 1350.170 2294.020 1350.490 2294.080 ;
        RECT 1351.090 2294.020 1351.410 2294.080 ;
        RECT 1543.830 2283.680 1544.150 2283.740 ;
        RECT 1544.750 2283.680 1545.070 2283.740 ;
        RECT 1543.830 2283.540 1545.070 2283.680 ;
        RECT 1543.830 2283.480 1544.150 2283.540 ;
        RECT 1544.750 2283.480 1545.070 2283.540 ;
        RECT 1559.010 2270.420 1559.330 2270.480 ;
        RECT 1559.470 2270.420 1559.790 2270.480 ;
        RECT 1559.010 2270.280 1559.790 2270.420 ;
        RECT 1559.010 2270.220 1559.330 2270.280 ;
        RECT 1559.470 2270.220 1559.790 2270.280 ;
        RECT 1543.830 2269.740 1544.150 2269.800 ;
        RECT 1545.210 2269.740 1545.530 2269.800 ;
        RECT 1543.830 2269.600 1545.530 2269.740 ;
        RECT 1543.830 2269.540 1544.150 2269.600 ;
        RECT 1545.210 2269.540 1545.530 2269.600 ;
        RECT 1531.410 2262.940 1531.730 2263.000 ;
        RECT 1532.330 2262.940 1532.650 2263.000 ;
        RECT 1531.410 2262.800 1532.650 2262.940 ;
        RECT 1531.410 2262.740 1531.730 2262.800 ;
        RECT 1532.330 2262.740 1532.650 2262.800 ;
        RECT 1559.470 2262.940 1559.790 2263.000 ;
        RECT 1560.390 2262.940 1560.710 2263.000 ;
        RECT 1559.470 2262.800 1560.710 2262.940 ;
        RECT 1559.470 2262.740 1559.790 2262.800 ;
        RECT 1560.390 2262.740 1560.710 2262.800 ;
        RECT 1351.090 2235.880 1351.410 2236.140 ;
        RECT 1351.180 2235.460 1351.320 2235.880 ;
        RECT 1351.090 2235.200 1351.410 2235.460 ;
        RECT 1531.410 2215.000 1531.730 2215.060 ;
        RECT 1532.790 2215.000 1533.110 2215.060 ;
        RECT 1531.410 2214.860 1533.110 2215.000 ;
        RECT 1531.410 2214.800 1531.730 2214.860 ;
        RECT 1532.790 2214.800 1533.110 2214.860 ;
        RECT 1559.470 2215.000 1559.790 2215.060 ;
        RECT 1560.390 2215.000 1560.710 2215.060 ;
        RECT 1559.470 2214.860 1560.710 2215.000 ;
        RECT 1559.470 2214.800 1559.790 2214.860 ;
        RECT 1560.390 2214.800 1560.710 2214.860 ;
        RECT 1350.170 2197.660 1350.490 2197.720 ;
        RECT 1351.090 2197.660 1351.410 2197.720 ;
        RECT 1350.170 2197.520 1351.410 2197.660 ;
        RECT 1350.170 2197.460 1350.490 2197.520 ;
        RECT 1351.090 2197.460 1351.410 2197.520 ;
        RECT 1532.790 2187.800 1533.110 2187.860 ;
        RECT 1532.420 2187.660 1533.110 2187.800 ;
        RECT 1532.420 2187.180 1532.560 2187.660 ;
        RECT 1532.790 2187.600 1533.110 2187.660 ;
        RECT 1532.330 2186.920 1532.650 2187.180 ;
        RECT 1531.870 2173.180 1532.190 2173.240 ;
        RECT 1532.330 2173.180 1532.650 2173.240 ;
        RECT 1531.870 2173.040 1532.650 2173.180 ;
        RECT 1531.870 2172.980 1532.190 2173.040 ;
        RECT 1532.330 2172.980 1532.650 2173.040 ;
        RECT 1531.410 2166.380 1531.730 2166.440 ;
        RECT 1531.870 2166.380 1532.190 2166.440 ;
        RECT 1531.410 2166.240 1532.190 2166.380 ;
        RECT 1531.410 2166.180 1531.730 2166.240 ;
        RECT 1531.870 2166.180 1532.190 2166.240 ;
        RECT 1559.470 2166.380 1559.790 2166.440 ;
        RECT 1560.390 2166.380 1560.710 2166.440 ;
        RECT 1559.470 2166.240 1560.710 2166.380 ;
        RECT 1559.470 2166.180 1559.790 2166.240 ;
        RECT 1560.390 2166.180 1560.710 2166.240 ;
        RECT 1351.090 2139.320 1351.410 2139.580 ;
        RECT 1351.180 2138.900 1351.320 2139.320 ;
        RECT 1351.090 2138.640 1351.410 2138.900 ;
        RECT 1350.630 2125.240 1350.950 2125.300 ;
        RECT 1351.090 2125.240 1351.410 2125.300 ;
        RECT 1350.630 2125.100 1351.410 2125.240 ;
        RECT 1350.630 2125.040 1350.950 2125.100 ;
        RECT 1351.090 2125.040 1351.410 2125.100 ;
        RECT 1531.410 2124.900 1531.730 2124.960 ;
        RECT 1532.790 2124.900 1533.110 2124.960 ;
        RECT 1531.410 2124.760 1533.110 2124.900 ;
        RECT 1531.410 2124.700 1531.730 2124.760 ;
        RECT 1532.790 2124.700 1533.110 2124.760 ;
        RECT 1559.470 2118.440 1559.790 2118.500 ;
        RECT 1560.390 2118.440 1560.710 2118.500 ;
        RECT 1559.470 2118.300 1560.710 2118.440 ;
        RECT 1559.470 2118.240 1559.790 2118.300 ;
        RECT 1560.390 2118.240 1560.710 2118.300 ;
        RECT 1532.790 2111.300 1533.110 2111.360 ;
        RECT 1533.710 2111.300 1534.030 2111.360 ;
        RECT 1532.790 2111.160 1534.030 2111.300 ;
        RECT 1532.790 2111.100 1533.110 2111.160 ;
        RECT 1533.710 2111.100 1534.030 2111.160 ;
        RECT 1350.630 2090.560 1350.950 2090.620 ;
        RECT 1351.550 2090.560 1351.870 2090.620 ;
        RECT 1350.630 2090.420 1351.870 2090.560 ;
        RECT 1350.630 2090.360 1350.950 2090.420 ;
        RECT 1351.550 2090.360 1351.870 2090.420 ;
        RECT 1559.470 2069.820 1559.790 2069.880 ;
        RECT 1560.390 2069.820 1560.710 2069.880 ;
        RECT 1559.470 2069.680 1560.710 2069.820 ;
        RECT 1559.470 2069.620 1559.790 2069.680 ;
        RECT 1560.390 2069.620 1560.710 2069.680 ;
        RECT 1532.330 2063.360 1532.650 2063.420 ;
        RECT 1533.710 2063.360 1534.030 2063.420 ;
        RECT 1532.330 2063.220 1534.030 2063.360 ;
        RECT 1532.330 2063.160 1532.650 2063.220 ;
        RECT 1533.710 2063.160 1534.030 2063.220 ;
        RECT 1244.830 2055.540 1245.150 2055.600 ;
        RECT 1346.030 2055.540 1346.350 2055.600 ;
        RECT 1244.830 2055.400 1346.350 2055.540 ;
        RECT 1244.830 2055.340 1245.150 2055.400 ;
        RECT 1346.030 2055.340 1346.350 2055.400 ;
        RECT 1287.150 2055.200 1287.470 2055.260 ;
        RECT 1346.490 2055.200 1346.810 2055.260 ;
        RECT 1287.150 2055.060 1346.810 2055.200 ;
        RECT 1287.150 2055.000 1287.470 2055.060 ;
        RECT 1346.490 2055.000 1346.810 2055.060 ;
        RECT 1230.110 2054.860 1230.430 2054.920 ;
        RECT 1335.450 2054.860 1335.770 2054.920 ;
        RECT 1230.110 2054.720 1335.770 2054.860 ;
        RECT 1230.110 2054.660 1230.430 2054.720 ;
        RECT 1335.450 2054.660 1335.770 2054.720 ;
        RECT 1116.950 2054.520 1117.270 2054.580 ;
        RECT 1332.690 2054.520 1333.010 2054.580 ;
        RECT 1116.950 2054.380 1333.010 2054.520 ;
        RECT 1116.950 2054.320 1117.270 2054.380 ;
        RECT 1332.690 2054.320 1333.010 2054.380 ;
        RECT 1130.750 2054.180 1131.070 2054.240 ;
        RECT 1352.930 2054.180 1353.250 2054.240 ;
        RECT 1130.750 2054.040 1353.250 2054.180 ;
        RECT 1130.750 2053.980 1131.070 2054.040 ;
        RECT 1352.930 2053.980 1353.250 2054.040 ;
        RECT 1216.310 2053.840 1216.630 2053.900 ;
        RECT 1346.950 2053.840 1347.270 2053.900 ;
        RECT 1216.310 2053.700 1347.270 2053.840 ;
        RECT 1216.310 2053.640 1216.630 2053.700 ;
        RECT 1346.950 2053.640 1347.270 2053.700 ;
        RECT 1059.910 2053.500 1060.230 2053.560 ;
        RECT 1334.990 2053.500 1335.310 2053.560 ;
        RECT 1059.910 2053.360 1335.310 2053.500 ;
        RECT 1059.910 2053.300 1060.230 2053.360 ;
        RECT 1334.990 2053.300 1335.310 2053.360 ;
        RECT 1031.390 2053.160 1031.710 2053.220 ;
        RECT 1353.850 2053.160 1354.170 2053.220 ;
        RECT 1031.390 2053.020 1354.170 2053.160 ;
        RECT 1031.390 2052.960 1031.710 2053.020 ;
        RECT 1353.850 2052.960 1354.170 2053.020 ;
        RECT 1016.670 2052.820 1016.990 2052.880 ;
        RECT 1347.410 2052.820 1347.730 2052.880 ;
        RECT 1016.670 2052.680 1347.730 2052.820 ;
        RECT 1016.670 2052.620 1016.990 2052.680 ;
        RECT 1347.410 2052.620 1347.730 2052.680 ;
        RECT 1350.170 2052.820 1350.490 2052.880 ;
        RECT 1352.010 2052.820 1352.330 2052.880 ;
        RECT 1350.170 2052.680 1352.330 2052.820 ;
        RECT 1350.170 2052.620 1350.490 2052.680 ;
        RECT 1352.010 2052.620 1352.330 2052.680 ;
        RECT 1201.590 2052.480 1201.910 2052.540 ;
        RECT 1333.150 2052.480 1333.470 2052.540 ;
        RECT 1201.590 2052.340 1333.470 2052.480 ;
        RECT 1201.590 2052.280 1201.910 2052.340 ;
        RECT 1333.150 2052.280 1333.470 2052.340 ;
        RECT 1187.790 2052.140 1188.110 2052.200 ;
        RECT 1335.910 2052.140 1336.230 2052.200 ;
        RECT 1187.790 2052.000 1336.230 2052.140 ;
        RECT 1187.790 2051.940 1188.110 2052.000 ;
        RECT 1335.910 2051.940 1336.230 2052.000 ;
        RECT 1173.070 2051.800 1173.390 2051.860 ;
        RECT 1345.570 2051.800 1345.890 2051.860 ;
        RECT 1173.070 2051.660 1345.890 2051.800 ;
        RECT 1173.070 2051.600 1173.390 2051.660 ;
        RECT 1345.570 2051.600 1345.890 2051.660 ;
        RECT 1159.270 2051.460 1159.590 2051.520 ;
        RECT 1352.470 2051.460 1352.790 2051.520 ;
        RECT 1159.270 2051.320 1352.790 2051.460 ;
        RECT 1159.270 2051.260 1159.590 2051.320 ;
        RECT 1352.470 2051.260 1352.790 2051.320 ;
        RECT 1144.550 2051.120 1144.870 2051.180 ;
        RECT 1353.390 2051.120 1353.710 2051.180 ;
        RECT 1144.550 2050.980 1353.710 2051.120 ;
        RECT 1144.550 2050.920 1144.870 2050.980 ;
        RECT 1353.390 2050.920 1353.710 2050.980 ;
        RECT 977.110 2050.780 977.430 2050.840 ;
        RECT 1088.430 2050.780 1088.750 2050.840 ;
        RECT 977.110 2050.640 1088.750 2050.780 ;
        RECT 977.110 2050.580 977.430 2050.640 ;
        RECT 1088.430 2050.580 1088.750 2050.640 ;
        RECT 1273.350 2050.780 1273.670 2050.840 ;
        RECT 1333.610 2050.780 1333.930 2050.840 ;
        RECT 1273.350 2050.640 1333.930 2050.780 ;
        RECT 1273.350 2050.580 1273.670 2050.640 ;
        RECT 1333.610 2050.580 1333.930 2050.640 ;
        RECT 977.570 2050.440 977.890 2050.500 ;
        RECT 1102.230 2050.440 1102.550 2050.500 ;
        RECT 977.570 2050.300 1102.550 2050.440 ;
        RECT 977.570 2050.240 977.890 2050.300 ;
        RECT 1102.230 2050.240 1102.550 2050.300 ;
        RECT 1258.630 2050.440 1258.950 2050.500 ;
        RECT 1337.750 2050.440 1338.070 2050.500 ;
        RECT 1258.630 2050.300 1338.070 2050.440 ;
        RECT 1258.630 2050.240 1258.950 2050.300 ;
        RECT 1337.750 2050.240 1338.070 2050.300 ;
        RECT 984.010 2050.100 984.330 2050.160 ;
        RECT 1073.710 2050.100 1074.030 2050.160 ;
        RECT 984.010 2049.960 1074.030 2050.100 ;
        RECT 984.010 2049.900 984.330 2049.960 ;
        RECT 1073.710 2049.900 1074.030 2049.960 ;
        RECT 1000.110 2049.760 1000.430 2049.820 ;
        RECT 1045.190 2049.760 1045.510 2049.820 ;
        RECT 1000.110 2049.620 1045.510 2049.760 ;
        RECT 1000.110 2049.560 1000.430 2049.620 ;
        RECT 1045.190 2049.560 1045.510 2049.620 ;
        RECT 1301.870 2049.760 1302.190 2049.820 ;
        RECT 1347.870 2049.760 1348.190 2049.820 ;
        RECT 1301.870 2049.620 1348.190 2049.760 ;
        RECT 1301.870 2049.560 1302.190 2049.620 ;
        RECT 1347.870 2049.560 1348.190 2049.620 ;
        RECT 984.470 2049.420 984.790 2049.480 ;
        RECT 1002.870 2049.420 1003.190 2049.480 ;
        RECT 984.470 2049.280 1003.190 2049.420 ;
        RECT 984.470 2049.220 984.790 2049.280 ;
        RECT 1002.870 2049.220 1003.190 2049.280 ;
        RECT 1315.670 2049.420 1315.990 2049.480 ;
        RECT 1336.370 2049.420 1336.690 2049.480 ;
        RECT 1315.670 2049.280 1336.690 2049.420 ;
        RECT 1315.670 2049.220 1315.990 2049.280 ;
        RECT 1336.370 2049.220 1336.690 2049.280 ;
        RECT 976.190 2048.060 976.510 2048.120 ;
        RECT 1014.370 2048.060 1014.690 2048.120 ;
        RECT 976.190 2047.920 1014.690 2048.060 ;
        RECT 976.190 2047.860 976.510 2047.920 ;
        RECT 1014.370 2047.860 1014.690 2047.920 ;
        RECT 983.090 2047.720 983.410 2047.780 ;
        RECT 1028.170 2047.720 1028.490 2047.780 ;
        RECT 983.090 2047.580 1028.490 2047.720 ;
        RECT 983.090 2047.520 983.410 2047.580 ;
        RECT 1028.170 2047.520 1028.490 2047.580 ;
        RECT 982.630 2047.380 982.950 2047.440 ;
        RECT 1062.670 2047.380 1062.990 2047.440 ;
        RECT 982.630 2047.240 1062.990 2047.380 ;
        RECT 982.630 2047.180 982.950 2047.240 ;
        RECT 1062.670 2047.180 1062.990 2047.240 ;
        RECT 975.730 2047.040 976.050 2047.100 ;
        RECT 1076.470 2047.040 1076.790 2047.100 ;
        RECT 975.730 2046.900 1076.790 2047.040 ;
        RECT 975.730 2046.840 976.050 2046.900 ;
        RECT 1076.470 2046.840 1076.790 2046.900 ;
        RECT 983.550 2046.700 983.870 2046.760 ;
        RECT 1097.630 2046.700 1097.950 2046.760 ;
        RECT 983.550 2046.560 1097.950 2046.700 ;
        RECT 983.550 2046.500 983.870 2046.560 ;
        RECT 1097.630 2046.500 1097.950 2046.560 ;
        RECT 976.650 2046.360 976.970 2046.420 ;
        RECT 1097.170 2046.360 1097.490 2046.420 ;
        RECT 976.650 2046.220 1097.490 2046.360 ;
        RECT 976.650 2046.160 976.970 2046.220 ;
        RECT 1097.170 2046.160 1097.490 2046.220 ;
        RECT 972.510 2046.020 972.830 2046.080 ;
        RECT 1111.430 2046.020 1111.750 2046.080 ;
        RECT 972.510 2045.880 1111.750 2046.020 ;
        RECT 972.510 2045.820 972.830 2045.880 ;
        RECT 1111.430 2045.820 1111.750 2045.880 ;
        RECT 965.610 2045.680 965.930 2045.740 ;
        RECT 1110.970 2045.680 1111.290 2045.740 ;
        RECT 965.610 2045.540 1111.290 2045.680 ;
        RECT 965.610 2045.480 965.930 2045.540 ;
        RECT 1110.970 2045.480 1111.290 2045.540 ;
        RECT 1330.850 2036.500 1331.170 2036.560 ;
        RECT 1343.730 2036.500 1344.050 2036.560 ;
        RECT 1330.850 2036.360 1344.050 2036.500 ;
        RECT 1330.850 2036.300 1331.170 2036.360 ;
        RECT 1343.730 2036.300 1344.050 2036.360 ;
        RECT 529.990 1988.560 530.310 1988.620 ;
        RECT 650.510 1988.560 650.830 1988.620 ;
        RECT 529.990 1988.420 650.830 1988.560 ;
        RECT 529.990 1988.360 530.310 1988.420 ;
        RECT 650.510 1988.360 650.830 1988.420 ;
        RECT 579.210 1987.540 579.530 1987.600 ;
        RECT 638.090 1987.540 638.410 1987.600 ;
        RECT 579.210 1987.400 638.410 1987.540 ;
        RECT 579.210 1987.340 579.530 1987.400 ;
        RECT 638.090 1987.340 638.410 1987.400 ;
        RECT 420.510 1978.700 420.830 1978.760 ;
        RECT 419.680 1978.560 420.830 1978.700 ;
        RECT 419.680 1977.680 419.820 1978.560 ;
        RECT 420.510 1978.500 420.830 1978.560 ;
        RECT 420.050 1978.160 420.370 1978.420 ;
        RECT 420.140 1978.020 420.280 1978.160 ;
        RECT 842.790 1978.020 843.110 1978.080 ;
        RECT 420.140 1977.880 843.110 1978.020 ;
        RECT 842.790 1977.820 843.110 1977.880 ;
        RECT 897.530 1977.680 897.850 1977.740 ;
        RECT 419.680 1977.540 897.850 1977.680 ;
        RECT 897.530 1977.480 897.850 1977.540 ;
      LAYER met1 ;
        RECT 362.830 1710.640 628.110 1977.400 ;
      LAYER met1 ;
        RECT 998.730 1713.500 999.050 1713.560 ;
        RECT 1001.030 1713.500 1001.350 1713.560 ;
        RECT 998.730 1713.360 1001.350 1713.500 ;
        RECT 998.730 1713.300 999.050 1713.360 ;
        RECT 1001.030 1713.300 1001.350 1713.360 ;
      LAYER met1 ;
        RECT 1002.830 1710.640 1329.750 2032.080 ;
      LAYER met1 ;
        RECT 1350.170 2029.020 1350.490 2029.080 ;
        RECT 1352.010 2029.020 1352.330 2029.080 ;
        RECT 1350.170 2028.880 1352.330 2029.020 ;
        RECT 1350.170 2028.820 1350.490 2028.880 ;
        RECT 1352.010 2028.820 1352.330 2028.880 ;
        RECT 1350.170 2028.340 1350.490 2028.400 ;
        RECT 1351.550 2028.340 1351.870 2028.400 ;
        RECT 1350.170 2028.200 1351.870 2028.340 ;
        RECT 1350.170 2028.140 1350.490 2028.200 ;
        RECT 1351.550 2028.140 1351.870 2028.200 ;
        RECT 1559.470 2021.880 1559.790 2021.940 ;
        RECT 1560.390 2021.880 1560.710 2021.940 ;
        RECT 1559.470 2021.740 1560.710 2021.880 ;
        RECT 1559.470 2021.680 1559.790 2021.740 ;
        RECT 1560.390 2021.680 1560.710 2021.740 ;
        RECT 1543.370 2004.540 1543.690 2004.600 ;
        RECT 1544.290 2004.540 1544.610 2004.600 ;
        RECT 1543.370 2004.400 1544.610 2004.540 ;
        RECT 1543.370 2004.340 1543.690 2004.400 ;
        RECT 1544.290 2004.340 1544.610 2004.400 ;
        RECT 1350.170 1980.740 1350.490 1980.800 ;
        RECT 1350.630 1980.740 1350.950 1980.800 ;
        RECT 1532.790 1980.740 1533.110 1980.800 ;
        RECT 1350.170 1980.600 1350.950 1980.740 ;
        RECT 1350.170 1980.540 1350.490 1980.600 ;
        RECT 1350.630 1980.540 1350.950 1980.600 ;
        RECT 1532.420 1980.600 1533.110 1980.740 ;
        RECT 1532.420 1980.120 1532.560 1980.600 ;
        RECT 1532.790 1980.540 1533.110 1980.600 ;
        RECT 1543.370 1980.400 1543.690 1980.460 ;
        RECT 1543.830 1980.400 1544.150 1980.460 ;
        RECT 1543.370 1980.260 1544.150 1980.400 ;
        RECT 1543.370 1980.200 1543.690 1980.260 ;
        RECT 1543.830 1980.200 1544.150 1980.260 ;
        RECT 1350.170 1980.060 1350.490 1980.120 ;
        RECT 1350.630 1980.060 1350.950 1980.120 ;
        RECT 1350.170 1979.920 1350.950 1980.060 ;
        RECT 1350.170 1979.860 1350.490 1979.920 ;
        RECT 1350.630 1979.860 1350.950 1979.920 ;
        RECT 1532.330 1979.860 1532.650 1980.120 ;
        RECT 1559.470 1973.260 1559.790 1973.320 ;
        RECT 1560.390 1973.260 1560.710 1973.320 ;
        RECT 1559.470 1973.120 1560.710 1973.260 ;
        RECT 1559.470 1973.060 1559.790 1973.120 ;
        RECT 1560.390 1973.060 1560.710 1973.120 ;
        RECT 1543.830 1956.260 1544.150 1956.320 ;
        RECT 1544.750 1956.260 1545.070 1956.320 ;
        RECT 1543.830 1956.120 1545.070 1956.260 ;
        RECT 1543.830 1956.060 1544.150 1956.120 ;
        RECT 1544.750 1956.060 1545.070 1956.120 ;
        RECT 2294.090 1947.080 2294.410 1947.140 ;
        RECT 2380.110 1947.080 2380.430 1947.140 ;
        RECT 2294.090 1946.940 2380.430 1947.080 ;
        RECT 2294.090 1946.880 2294.410 1946.940 ;
        RECT 2380.110 1946.880 2380.430 1946.940 ;
        RECT 2076.510 1946.740 2076.830 1946.800 ;
        RECT 2321.230 1946.740 2321.550 1946.800 ;
        RECT 2076.510 1946.600 2321.550 1946.740 ;
        RECT 2076.510 1946.540 2076.830 1946.600 ;
        RECT 2321.230 1946.540 2321.550 1946.600 ;
        RECT 2082.950 1946.400 2083.270 1946.460 ;
        RECT 2438.070 1946.400 2438.390 1946.460 ;
        RECT 2082.950 1946.260 2438.390 1946.400 ;
        RECT 2082.950 1946.200 2083.270 1946.260 ;
        RECT 2438.070 1946.200 2438.390 1946.260 ;
        RECT 2083.410 1946.060 2083.730 1946.120 ;
        RECT 2496.950 1946.060 2497.270 1946.120 ;
        RECT 2083.410 1945.920 2497.270 1946.060 ;
        RECT 2083.410 1945.860 2083.730 1945.920 ;
        RECT 2496.950 1945.860 2497.270 1945.920 ;
        RECT 1350.170 1932.120 1350.490 1932.180 ;
        RECT 1351.090 1932.120 1351.410 1932.180 ;
        RECT 1350.170 1931.980 1351.410 1932.120 ;
        RECT 1350.170 1931.920 1350.490 1931.980 ;
        RECT 1351.090 1931.920 1351.410 1931.980 ;
        RECT 1532.330 1931.920 1532.650 1932.180 ;
        RECT 1532.420 1931.500 1532.560 1931.920 ;
        RECT 1545.210 1931.580 1545.530 1931.840 ;
        RECT 1532.330 1931.240 1532.650 1931.500 ;
        RECT 1544.290 1931.440 1544.610 1931.500 ;
        RECT 1545.300 1931.440 1545.440 1931.580 ;
        RECT 1544.290 1931.300 1545.440 1931.440 ;
        RECT 1544.290 1931.240 1544.610 1931.300 ;
        RECT 1724.610 1928.720 1724.930 1928.780 ;
        RECT 2044.310 1928.720 2044.630 1928.780 ;
        RECT 1724.610 1928.580 2044.630 1928.720 ;
        RECT 1724.610 1928.520 1724.930 1928.580 ;
        RECT 2044.310 1928.520 2044.630 1928.580 ;
        RECT 1828.110 1928.040 1828.430 1928.100 ;
        RECT 1964.270 1928.040 1964.590 1928.100 ;
        RECT 1828.110 1927.900 1964.590 1928.040 ;
        RECT 1828.110 1927.840 1828.430 1927.900 ;
        RECT 1964.270 1927.840 1964.590 1927.900 ;
        RECT 1745.310 1927.700 1745.630 1927.760 ;
        RECT 1929.310 1927.700 1929.630 1927.760 ;
        RECT 1745.310 1927.560 1929.630 1927.700 ;
        RECT 1745.310 1927.500 1745.630 1927.560 ;
        RECT 1929.310 1927.500 1929.630 1927.560 ;
        RECT 1779.810 1927.360 1780.130 1927.420 ;
        RECT 1998.310 1927.360 1998.630 1927.420 ;
        RECT 1779.810 1927.220 1998.630 1927.360 ;
        RECT 1779.810 1927.160 1780.130 1927.220 ;
        RECT 1998.310 1927.160 1998.630 1927.220 ;
        RECT 1786.710 1927.020 1787.030 1927.080 ;
        RECT 2033.270 1927.020 2033.590 1927.080 ;
        RECT 1786.710 1926.880 2033.590 1927.020 ;
        RECT 1786.710 1926.820 1787.030 1926.880 ;
        RECT 2033.270 1926.820 2033.590 1926.880 ;
        RECT 1759.110 1926.680 1759.430 1926.740 ;
        RECT 2010.270 1926.680 2010.590 1926.740 ;
        RECT 1759.110 1926.540 2010.590 1926.680 ;
        RECT 1759.110 1926.480 1759.430 1926.540 ;
        RECT 2010.270 1926.480 2010.590 1926.540 ;
        RECT 1738.410 1926.340 1738.730 1926.400 ;
        RECT 1987.270 1926.340 1987.590 1926.400 ;
        RECT 1738.410 1926.200 1987.590 1926.340 ;
        RECT 1738.410 1926.140 1738.730 1926.200 ;
        RECT 1987.270 1926.140 1987.590 1926.200 ;
        RECT 1717.250 1926.000 1717.570 1926.060 ;
        RECT 1975.310 1926.000 1975.630 1926.060 ;
        RECT 1717.250 1925.860 1975.630 1926.000 ;
        RECT 1717.250 1925.800 1717.570 1925.860 ;
        RECT 1975.310 1925.800 1975.630 1925.860 ;
        RECT 1772.910 1925.660 1773.230 1925.720 ;
        RECT 2067.310 1925.660 2067.630 1925.720 ;
        RECT 1772.910 1925.520 2067.630 1925.660 ;
        RECT 1772.910 1925.460 1773.230 1925.520 ;
        RECT 2067.310 1925.460 2067.630 1925.520 ;
        RECT 1559.470 1925.320 1559.790 1925.380 ;
        RECT 1560.390 1925.320 1560.710 1925.380 ;
        RECT 1559.470 1925.180 1560.710 1925.320 ;
        RECT 1559.470 1925.120 1559.790 1925.180 ;
        RECT 1560.390 1925.120 1560.710 1925.180 ;
        RECT 1827.650 1925.320 1827.970 1925.380 ;
        RECT 1952.310 1925.320 1952.630 1925.380 ;
        RECT 1827.650 1925.180 1952.630 1925.320 ;
        RECT 1827.650 1925.120 1827.970 1925.180 ;
        RECT 1952.310 1925.120 1952.630 1925.180 ;
        RECT 1351.090 1907.980 1351.410 1908.040 ;
        RECT 1352.010 1907.980 1352.330 1908.040 ;
        RECT 1351.090 1907.840 1352.330 1907.980 ;
        RECT 1351.090 1907.780 1351.410 1907.840 ;
        RECT 1352.010 1907.780 1352.330 1907.840 ;
        RECT 1544.290 1897.440 1544.610 1897.500 ;
        RECT 1545.210 1897.440 1545.530 1897.500 ;
        RECT 1544.290 1897.300 1545.530 1897.440 ;
        RECT 1544.290 1897.240 1544.610 1897.300 ;
        RECT 1545.210 1897.240 1545.530 1897.300 ;
        RECT 1531.870 1883.840 1532.190 1883.900 ;
        RECT 1532.330 1883.840 1532.650 1883.900 ;
        RECT 1531.870 1883.700 1532.650 1883.840 ;
        RECT 1531.870 1883.640 1532.190 1883.700 ;
        RECT 1532.330 1883.640 1532.650 1883.700 ;
        RECT 1752.210 1883.840 1752.530 1883.900 ;
        RECT 1904.470 1883.840 1904.790 1883.900 ;
        RECT 1752.210 1883.700 1904.790 1883.840 ;
        RECT 1752.210 1883.640 1752.530 1883.700 ;
        RECT 1904.470 1883.640 1904.790 1883.700 ;
        RECT 1573.730 1883.500 1574.050 1883.560 ;
        RECT 1574.650 1883.500 1574.970 1883.560 ;
        RECT 1573.730 1883.360 1574.970 1883.500 ;
        RECT 1573.730 1883.300 1574.050 1883.360 ;
        RECT 1574.650 1883.300 1574.970 1883.360 ;
        RECT 1558.550 1876.700 1558.870 1876.760 ;
        RECT 1559.470 1876.700 1559.790 1876.760 ;
        RECT 1558.550 1876.560 1559.790 1876.700 ;
        RECT 1558.550 1876.500 1558.870 1876.560 ;
        RECT 1559.470 1876.500 1559.790 1876.560 ;
        RECT 1821.210 1870.240 1821.530 1870.300 ;
        RECT 1904.470 1870.240 1904.790 1870.300 ;
        RECT 1821.210 1870.100 1904.790 1870.240 ;
        RECT 1821.210 1870.040 1821.530 1870.100 ;
        RECT 1904.470 1870.040 1904.790 1870.100 ;
        RECT 1544.290 1859.700 1544.610 1859.760 ;
        RECT 1545.210 1859.700 1545.530 1859.760 ;
        RECT 1544.290 1859.560 1545.530 1859.700 ;
        RECT 1544.290 1859.500 1544.610 1859.560 ;
        RECT 1545.210 1859.500 1545.530 1859.560 ;
        RECT 1731.510 1849.500 1731.830 1849.560 ;
        RECT 1904.470 1849.500 1904.790 1849.560 ;
        RECT 1731.510 1849.360 1904.790 1849.500 ;
        RECT 1731.510 1849.300 1731.830 1849.360 ;
        RECT 1904.470 1849.300 1904.790 1849.360 ;
        RECT 1350.170 1835.560 1350.490 1835.620 ;
        RECT 1351.090 1835.560 1351.410 1835.620 ;
        RECT 1350.170 1835.420 1351.410 1835.560 ;
        RECT 1350.170 1835.360 1350.490 1835.420 ;
        RECT 1351.090 1835.360 1351.410 1835.420 ;
        RECT 1531.870 1835.560 1532.190 1835.620 ;
        RECT 1532.790 1835.560 1533.110 1835.620 ;
        RECT 1531.870 1835.420 1533.110 1835.560 ;
        RECT 1531.870 1835.360 1532.190 1835.420 ;
        RECT 1532.790 1835.360 1533.110 1835.420 ;
        RECT 1558.550 1828.760 1558.870 1828.820 ;
        RECT 1559.930 1828.760 1560.250 1828.820 ;
        RECT 1558.550 1828.620 1560.250 1828.760 ;
        RECT 1558.550 1828.560 1558.870 1828.620 ;
        RECT 1559.930 1828.560 1560.250 1828.620 ;
        RECT 1544.290 1821.960 1544.610 1822.020 ;
        RECT 1545.210 1821.960 1545.530 1822.020 ;
        RECT 1544.290 1821.820 1545.530 1821.960 ;
        RECT 1544.290 1821.760 1544.610 1821.820 ;
        RECT 1545.210 1821.760 1545.530 1821.820 ;
        RECT 1662.510 1814.820 1662.830 1814.880 ;
        RECT 1904.470 1814.820 1904.790 1814.880 ;
        RECT 1662.510 1814.680 1904.790 1814.820 ;
        RECT 1662.510 1814.620 1662.830 1814.680 ;
        RECT 1904.470 1814.620 1904.790 1814.680 ;
        RECT 1351.090 1801.020 1351.410 1801.280 ;
        RECT 1351.180 1800.880 1351.320 1801.020 ;
        RECT 1351.550 1800.880 1351.870 1800.940 ;
        RECT 1351.180 1800.740 1351.870 1800.880 ;
        RECT 1351.550 1800.680 1351.870 1800.740 ;
        RECT 1350.170 1786.940 1350.490 1787.000 ;
        RECT 1351.550 1786.940 1351.870 1787.000 ;
        RECT 1350.170 1786.800 1351.870 1786.940 ;
        RECT 1350.170 1786.740 1350.490 1786.800 ;
        RECT 1351.550 1786.740 1351.870 1786.800 ;
        RECT 1573.730 1786.940 1574.050 1787.000 ;
        RECT 1574.650 1786.940 1574.970 1787.000 ;
        RECT 1573.730 1786.800 1574.970 1786.940 ;
        RECT 1573.730 1786.740 1574.050 1786.800 ;
        RECT 1574.650 1786.740 1574.970 1786.800 ;
        RECT 1532.790 1786.600 1533.110 1786.660 ;
        RECT 1534.170 1786.600 1534.490 1786.660 ;
        RECT 1532.790 1786.460 1534.490 1786.600 ;
        RECT 1532.790 1786.400 1533.110 1786.460 ;
        RECT 1534.170 1786.400 1534.490 1786.460 ;
        RECT 1350.170 1780.140 1350.490 1780.200 ;
        RECT 1350.630 1780.140 1350.950 1780.200 ;
        RECT 1350.170 1780.000 1350.950 1780.140 ;
        RECT 1350.170 1779.940 1350.490 1780.000 ;
        RECT 1350.630 1779.940 1350.950 1780.000 ;
        RECT 1559.470 1780.140 1559.790 1780.200 ;
        RECT 1560.390 1780.140 1560.710 1780.200 ;
        RECT 1559.470 1780.000 1560.710 1780.140 ;
        RECT 1559.470 1779.940 1559.790 1780.000 ;
        RECT 1560.390 1779.940 1560.710 1780.000 ;
        RECT 1766.010 1766.540 1766.330 1766.600 ;
        RECT 1904.470 1766.540 1904.790 1766.600 ;
        RECT 1766.010 1766.400 1904.790 1766.540 ;
        RECT 1766.010 1766.340 1766.330 1766.400 ;
        RECT 1904.470 1766.340 1904.790 1766.400 ;
      LAYER met1 ;
        RECT 1922.830 1760.240 2072.190 1905.280 ;
      LAYER met1 ;
        RECT 1533.250 1739.340 1533.570 1739.400 ;
        RECT 1534.170 1739.340 1534.490 1739.400 ;
        RECT 1533.250 1739.200 1534.490 1739.340 ;
        RECT 1533.250 1739.140 1533.570 1739.200 ;
        RECT 1534.170 1739.140 1534.490 1739.200 ;
        RECT 1532.790 1738.660 1533.110 1738.720 ;
        RECT 1533.710 1738.660 1534.030 1738.720 ;
        RECT 1532.790 1738.520 1534.030 1738.660 ;
        RECT 1532.790 1738.460 1533.110 1738.520 ;
        RECT 1533.710 1738.460 1534.030 1738.520 ;
        RECT 1820.750 1738.660 1821.070 1738.720 ;
        RECT 1933.910 1738.660 1934.230 1738.720 ;
        RECT 1820.750 1738.520 1934.230 1738.660 ;
        RECT 1820.750 1738.460 1821.070 1738.520 ;
        RECT 1933.910 1738.460 1934.230 1738.520 ;
        RECT 1800.510 1738.320 1800.830 1738.380 ;
        RECT 1956.910 1738.320 1957.230 1738.380 ;
        RECT 1800.510 1738.180 1957.230 1738.320 ;
        RECT 1800.510 1738.120 1800.830 1738.180 ;
        RECT 1956.910 1738.120 1957.230 1738.180 ;
        RECT 1814.310 1737.980 1814.630 1738.040 ;
        RECT 1990.950 1737.980 1991.270 1738.040 ;
        RECT 1814.310 1737.840 1991.270 1737.980 ;
        RECT 1814.310 1737.780 1814.630 1737.840 ;
        RECT 1990.950 1737.780 1991.270 1737.840 ;
        RECT 1793.610 1737.640 1793.930 1737.700 ;
        RECT 1967.950 1737.640 1968.270 1737.700 ;
        RECT 1793.610 1737.500 1968.270 1737.640 ;
        RECT 1793.610 1737.440 1793.930 1737.500 ;
        RECT 1967.950 1737.440 1968.270 1737.500 ;
        RECT 1807.410 1737.300 1807.730 1737.360 ;
        RECT 2013.950 1737.300 2014.270 1737.360 ;
        RECT 1807.410 1737.160 2014.270 1737.300 ;
        RECT 1807.410 1737.100 1807.730 1737.160 ;
        RECT 2013.950 1737.100 2014.270 1737.160 ;
        RECT 1751.750 1736.960 1752.070 1737.020 ;
        RECT 1979.910 1736.960 1980.230 1737.020 ;
        RECT 1751.750 1736.820 1980.230 1736.960 ;
        RECT 1751.750 1736.760 1752.070 1736.820 ;
        RECT 1979.910 1736.760 1980.230 1736.820 ;
        RECT 1772.450 1736.620 1772.770 1736.680 ;
        RECT 2002.910 1736.620 2003.230 1736.680 ;
        RECT 1772.450 1736.480 2003.230 1736.620 ;
        RECT 1772.450 1736.420 1772.770 1736.480 ;
        RECT 2002.910 1736.420 2003.230 1736.480 ;
        RECT 1806.950 1736.280 1807.270 1736.340 ;
        RECT 2036.950 1736.280 2037.270 1736.340 ;
        RECT 1806.950 1736.140 2037.270 1736.280 ;
        RECT 1806.950 1736.080 1807.270 1736.140 ;
        RECT 2036.950 1736.080 2037.270 1736.140 ;
        RECT 1703.910 1735.940 1704.230 1736.000 ;
        RECT 1944.950 1735.940 1945.270 1736.000 ;
        RECT 1703.910 1735.800 1945.270 1735.940 ;
        RECT 1703.910 1735.740 1704.230 1735.800 ;
        RECT 1944.950 1735.740 1945.270 1735.800 ;
        RECT 1800.050 1735.600 1800.370 1735.660 ;
        RECT 2071.910 1735.600 2072.230 1735.660 ;
        RECT 1800.050 1735.460 2072.230 1735.600 ;
        RECT 1800.050 1735.400 1800.370 1735.460 ;
        RECT 2071.910 1735.400 2072.230 1735.460 ;
        RECT 1365.810 1735.260 1366.130 1735.320 ;
        RECT 1553.030 1735.260 1553.350 1735.320 ;
        RECT 1365.810 1735.120 1553.350 1735.260 ;
        RECT 1365.810 1735.060 1366.130 1735.120 ;
        RECT 1553.030 1735.060 1553.350 1735.120 ;
        RECT 1669.410 1735.260 1669.730 1735.320 ;
        RECT 2059.950 1735.260 2060.270 1735.320 ;
        RECT 1669.410 1735.120 2060.270 1735.260 ;
        RECT 1669.410 1735.060 1669.730 1735.120 ;
        RECT 2059.950 1735.060 2060.270 1735.120 ;
        RECT 1350.630 1732.200 1350.950 1732.260 ;
        RECT 1352.010 1732.200 1352.330 1732.260 ;
        RECT 1350.630 1732.060 1352.330 1732.200 ;
        RECT 1350.630 1732.000 1350.950 1732.060 ;
        RECT 1352.010 1732.000 1352.330 1732.060 ;
        RECT 1559.470 1732.200 1559.790 1732.260 ;
        RECT 1560.390 1732.200 1560.710 1732.260 ;
        RECT 1559.470 1732.060 1560.710 1732.200 ;
        RECT 1559.470 1732.000 1559.790 1732.060 ;
        RECT 1560.390 1732.000 1560.710 1732.060 ;
        RECT 1544.290 1725.400 1544.610 1725.460 ;
        RECT 1545.210 1725.400 1545.530 1725.460 ;
        RECT 1544.290 1725.260 1545.530 1725.400 ;
        RECT 1544.290 1725.200 1544.610 1725.260 ;
        RECT 1545.210 1725.200 1545.530 1725.260 ;
        RECT 1350.630 1725.060 1350.950 1725.120 ;
        RECT 1352.010 1725.060 1352.330 1725.120 ;
        RECT 1350.630 1724.920 1352.330 1725.060 ;
        RECT 1350.630 1724.860 1350.950 1724.920 ;
        RECT 1352.010 1724.860 1352.330 1724.920 ;
      LAYER met1 ;
        RECT 2302.830 1710.640 2522.640 1926.000 ;
      LAYER met1 ;
        RECT 1559.010 1700.920 1559.330 1700.980 ;
        RECT 1560.390 1700.920 1560.710 1700.980 ;
        RECT 1559.010 1700.780 1560.710 1700.920 ;
        RECT 1559.010 1700.720 1559.330 1700.780 ;
        RECT 1560.390 1700.720 1560.710 1700.780 ;
        RECT 999.190 1695.140 999.510 1695.200 ;
        RECT 1070.490 1695.140 1070.810 1695.200 ;
        RECT 999.190 1695.000 1070.810 1695.140 ;
        RECT 999.190 1694.940 999.510 1695.000 ;
        RECT 1070.490 1694.940 1070.810 1695.000 ;
        RECT 974.810 1694.800 975.130 1694.860 ;
        RECT 1048.870 1694.800 1049.190 1694.860 ;
        RECT 974.810 1694.660 1049.190 1694.800 ;
        RECT 974.810 1694.600 975.130 1694.660 ;
        RECT 1048.870 1694.600 1049.190 1694.660 ;
        RECT 1289.910 1694.800 1290.230 1694.860 ;
        RECT 1347.870 1694.800 1348.190 1694.860 ;
        RECT 1289.910 1694.660 1348.190 1694.800 ;
        RECT 1289.910 1694.600 1290.230 1694.660 ;
        RECT 1347.870 1694.600 1348.190 1694.660 ;
        RECT 999.650 1694.460 999.970 1694.520 ;
        RECT 1076.470 1694.460 1076.790 1694.520 ;
        RECT 999.650 1694.320 1076.790 1694.460 ;
        RECT 999.650 1694.260 999.970 1694.320 ;
        RECT 1076.470 1694.260 1076.790 1694.320 ;
        RECT 1234.710 1694.460 1235.030 1694.520 ;
        RECT 1335.450 1694.460 1335.770 1694.520 ;
        RECT 1234.710 1694.320 1335.770 1694.460 ;
        RECT 1234.710 1694.260 1235.030 1694.320 ;
        RECT 1335.450 1694.260 1335.770 1694.320 ;
        RECT 982.170 1694.120 982.490 1694.180 ;
        RECT 1104.990 1694.120 1105.310 1694.180 ;
        RECT 982.170 1693.980 1105.310 1694.120 ;
        RECT 982.170 1693.920 982.490 1693.980 ;
        RECT 1104.990 1693.920 1105.310 1693.980 ;
        RECT 1186.410 1694.120 1186.730 1694.180 ;
        RECT 1335.910 1694.120 1336.230 1694.180 ;
        RECT 1186.410 1693.980 1336.230 1694.120 ;
        RECT 1186.410 1693.920 1186.730 1693.980 ;
        RECT 1335.910 1693.920 1336.230 1693.980 ;
        RECT 975.270 1693.780 975.590 1693.840 ;
        RECT 1110.970 1693.780 1111.290 1693.840 ;
        RECT 975.270 1693.640 1111.290 1693.780 ;
        RECT 975.270 1693.580 975.590 1693.640 ;
        RECT 1110.970 1693.580 1111.290 1693.640 ;
        RECT 1185.950 1693.780 1186.270 1693.840 ;
        RECT 1336.370 1693.780 1336.690 1693.840 ;
        RECT 1185.950 1693.640 1336.690 1693.780 ;
        RECT 1185.950 1693.580 1186.270 1693.640 ;
        RECT 1336.370 1693.580 1336.690 1693.640 ;
        RECT 1310.610 1692.420 1310.930 1692.480 ;
        RECT 1343.730 1692.420 1344.050 1692.480 ;
        RECT 1310.610 1692.280 1344.050 1692.420 ;
        RECT 1310.610 1692.220 1310.930 1692.280 ;
        RECT 1343.730 1692.220 1344.050 1692.280 ;
        RECT 1573.730 1690.860 1574.050 1691.120 ;
        RECT 1532.790 1690.720 1533.110 1690.780 ;
        RECT 1533.710 1690.720 1534.030 1690.780 ;
        RECT 1532.790 1690.580 1534.030 1690.720 ;
        RECT 1573.820 1690.720 1573.960 1690.860 ;
        RECT 1574.190 1690.720 1574.510 1690.780 ;
        RECT 1573.820 1690.580 1574.510 1690.720 ;
        RECT 1532.790 1690.520 1533.110 1690.580 ;
        RECT 1533.710 1690.520 1534.030 1690.580 ;
        RECT 1574.190 1690.520 1574.510 1690.580 ;
        RECT 1116.030 1690.040 1116.350 1690.100 ;
        RECT 1186.870 1690.040 1187.190 1690.100 ;
        RECT 1116.030 1689.900 1187.190 1690.040 ;
        RECT 1116.030 1689.840 1116.350 1689.900 ;
        RECT 1186.870 1689.840 1187.190 1689.900 ;
        RECT 1159.270 1689.700 1159.590 1689.760 ;
        RECT 1221.370 1689.700 1221.690 1689.760 ;
        RECT 1159.270 1689.560 1221.690 1689.700 ;
        RECT 1159.270 1689.500 1159.590 1689.560 ;
        RECT 1221.370 1689.500 1221.690 1689.560 ;
        RECT 1268.750 1689.700 1269.070 1689.760 ;
        RECT 1315.670 1689.700 1315.990 1689.760 ;
        RECT 1268.750 1689.560 1315.990 1689.700 ;
        RECT 1268.750 1689.500 1269.070 1689.560 ;
        RECT 1315.670 1689.500 1315.990 1689.560 ;
        RECT 1102.230 1689.360 1102.550 1689.420 ;
        RECT 1203.890 1689.360 1204.210 1689.420 ;
        RECT 1102.230 1689.220 1204.210 1689.360 ;
        RECT 1102.230 1689.160 1102.550 1689.220 ;
        RECT 1203.890 1689.160 1204.210 1689.220 ;
        RECT 1214.010 1689.360 1214.330 1689.420 ;
        RECT 1287.150 1689.360 1287.470 1689.420 ;
        RECT 1214.010 1689.220 1287.470 1689.360 ;
        RECT 1214.010 1689.160 1214.330 1689.220 ;
        RECT 1287.150 1689.160 1287.470 1689.220 ;
        RECT 1130.750 1689.020 1131.070 1689.080 ;
        RECT 1196.990 1689.020 1197.310 1689.080 ;
        RECT 1130.750 1688.880 1197.310 1689.020 ;
        RECT 1130.750 1688.820 1131.070 1688.880 ;
        RECT 1196.990 1688.820 1197.310 1688.880 ;
        RECT 1217.690 1689.020 1218.010 1689.080 ;
        RECT 1230.110 1689.020 1230.430 1689.080 ;
        RECT 1217.690 1688.880 1230.430 1689.020 ;
        RECT 1217.690 1688.820 1218.010 1688.880 ;
        RECT 1230.110 1688.820 1230.430 1688.880 ;
        RECT 1248.050 1689.020 1248.370 1689.080 ;
        RECT 1300.950 1689.020 1301.270 1689.080 ;
        RECT 1248.050 1688.880 1301.270 1689.020 ;
        RECT 1248.050 1688.820 1248.370 1688.880 ;
        RECT 1300.950 1688.820 1301.270 1688.880 ;
        RECT 463.750 1688.680 464.070 1688.740 ;
        RECT 468.810 1688.680 469.130 1688.740 ;
        RECT 463.750 1688.540 469.130 1688.680 ;
        RECT 463.750 1688.480 464.070 1688.540 ;
        RECT 468.810 1688.480 469.130 1688.540 ;
        RECT 514.350 1688.680 514.670 1688.740 ;
        RECT 517.110 1688.680 517.430 1688.740 ;
        RECT 514.350 1688.540 517.430 1688.680 ;
        RECT 514.350 1688.480 514.670 1688.540 ;
        RECT 517.110 1688.480 517.430 1688.540 ;
        RECT 1073.710 1688.680 1074.030 1688.740 ;
        RECT 1293.590 1688.680 1293.910 1688.740 ;
        RECT 1073.710 1688.540 1293.910 1688.680 ;
        RECT 1073.710 1688.480 1074.030 1688.540 ;
        RECT 1293.590 1688.480 1293.910 1688.540 ;
        RECT 1030.470 1688.340 1030.790 1688.400 ;
        RECT 1264.150 1688.340 1264.470 1688.400 ;
        RECT 1030.470 1688.200 1264.470 1688.340 ;
        RECT 1030.470 1688.140 1030.790 1688.200 ;
        RECT 1264.150 1688.140 1264.470 1688.200 ;
        RECT 2000.610 1688.000 2000.930 1688.060 ;
        RECT 2302.830 1688.000 2303.150 1688.060 ;
        RECT 2000.610 1687.860 2303.150 1688.000 ;
        RECT 2000.610 1687.800 2000.930 1687.860 ;
        RECT 2302.830 1687.800 2303.150 1687.860 ;
        RECT 2048.910 1687.660 2049.230 1687.720 ;
        RECT 2360.790 1687.660 2361.110 1687.720 ;
        RECT 2048.910 1687.520 2361.110 1687.660 ;
        RECT 2048.910 1687.460 2049.230 1687.520 ;
        RECT 2360.790 1687.460 2361.110 1687.520 ;
        RECT 2042.010 1687.320 2042.330 1687.380 ;
        RECT 2419.670 1687.320 2419.990 1687.380 ;
        RECT 2042.010 1687.180 2419.990 1687.320 ;
        RECT 2042.010 1687.120 2042.330 1687.180 ;
        RECT 2419.670 1687.120 2419.990 1687.180 ;
        RECT 2069.610 1686.980 2069.930 1687.040 ;
        RECT 2477.630 1686.980 2477.950 1687.040 ;
        RECT 2069.610 1686.840 2477.950 1686.980 ;
        RECT 2069.610 1686.780 2069.930 1686.840 ;
        RECT 2477.630 1686.780 2477.950 1686.840 ;
        RECT 1144.550 1686.640 1144.870 1686.700 ;
        RECT 1180.890 1686.640 1181.210 1686.700 ;
        RECT 1144.550 1686.500 1181.210 1686.640 ;
        RECT 1144.550 1686.440 1144.870 1686.500 ;
        RECT 1180.890 1686.440 1181.210 1686.500 ;
        RECT 1196.990 1686.640 1197.310 1686.700 ;
        RECT 1237.010 1686.640 1237.330 1686.700 ;
        RECT 1196.990 1686.500 1237.330 1686.640 ;
        RECT 1196.990 1686.440 1197.310 1686.500 ;
        RECT 1237.010 1686.440 1237.330 1686.500 ;
        RECT 1002.870 1685.620 1003.190 1685.680 ;
        RECT 1038.290 1685.620 1038.610 1685.680 ;
        RECT 1002.870 1685.480 1038.610 1685.620 ;
        RECT 1002.870 1685.420 1003.190 1685.480 ;
        RECT 1038.290 1685.420 1038.610 1685.480 ;
        RECT 1173.070 1684.600 1173.390 1684.660 ;
        RECT 1188.250 1684.600 1188.570 1684.660 ;
        RECT 1173.070 1684.460 1188.570 1684.600 ;
        RECT 1173.070 1684.400 1173.390 1684.460 ;
        RECT 1188.250 1684.400 1188.570 1684.460 ;
        RECT 1193.310 1684.600 1193.630 1684.660 ;
        RECT 1215.390 1684.600 1215.710 1684.660 ;
        RECT 1193.310 1684.460 1215.710 1684.600 ;
        RECT 1193.310 1684.400 1193.630 1684.460 ;
        RECT 1215.390 1684.400 1215.710 1684.460 ;
        RECT 1016.670 1684.260 1016.990 1684.320 ;
        RECT 1020.810 1684.260 1021.130 1684.320 ;
        RECT 1016.670 1684.120 1021.130 1684.260 ;
        RECT 1016.670 1684.060 1016.990 1684.120 ;
        RECT 1020.810 1684.060 1021.130 1684.120 ;
        RECT 1187.790 1684.260 1188.110 1684.320 ;
        RECT 1196.990 1684.260 1197.310 1684.320 ;
        RECT 1187.790 1684.120 1197.310 1684.260 ;
        RECT 1187.790 1684.060 1188.110 1684.120 ;
        RECT 1196.990 1684.060 1197.310 1684.120 ;
        RECT 1238.390 1684.260 1238.710 1684.320 ;
        RECT 1243.910 1684.260 1244.230 1684.320 ;
        RECT 1238.390 1684.120 1244.230 1684.260 ;
        RECT 1238.390 1684.060 1238.710 1684.120 ;
        RECT 1243.910 1684.060 1244.230 1684.120 ;
        RECT 1272.430 1684.260 1272.750 1684.320 ;
        RECT 1291.290 1684.260 1291.610 1684.320 ;
        RECT 1272.430 1684.120 1291.610 1684.260 ;
        RECT 1272.430 1684.060 1272.750 1684.120 ;
        RECT 1291.290 1684.060 1291.610 1684.120 ;
        RECT 1531.410 1683.580 1531.730 1683.640 ;
        RECT 1532.330 1683.580 1532.650 1683.640 ;
        RECT 1531.410 1683.440 1532.650 1683.580 ;
        RECT 1531.410 1683.380 1531.730 1683.440 ;
        RECT 1532.330 1683.380 1532.650 1683.440 ;
        RECT 1572.810 1683.580 1573.130 1683.640 ;
        RECT 1574.190 1683.580 1574.510 1683.640 ;
        RECT 1572.810 1683.440 1574.510 1683.580 ;
        RECT 1572.810 1683.380 1573.130 1683.440 ;
        RECT 1574.190 1683.380 1574.510 1683.440 ;
        RECT 1350.630 1676.780 1350.950 1676.840 ;
        RECT 1351.090 1676.780 1351.410 1676.840 ;
        RECT 1350.630 1676.640 1351.410 1676.780 ;
        RECT 1350.630 1676.580 1350.950 1676.640 ;
        RECT 1351.090 1676.580 1351.410 1676.640 ;
        RECT 1069.570 1642.440 1069.890 1642.500 ;
        RECT 1070.030 1642.440 1070.350 1642.500 ;
        RECT 1069.570 1642.300 1070.350 1642.440 ;
        RECT 1069.570 1642.240 1069.890 1642.300 ;
        RECT 1070.030 1642.240 1070.350 1642.300 ;
        RECT 1104.070 1642.440 1104.390 1642.500 ;
        RECT 1104.990 1642.440 1105.310 1642.500 ;
        RECT 1104.070 1642.300 1105.310 1642.440 ;
        RECT 1104.070 1642.240 1104.390 1642.300 ;
        RECT 1104.990 1642.240 1105.310 1642.300 ;
        RECT 1221.370 1642.440 1221.690 1642.500 ;
        RECT 1243.910 1642.440 1244.230 1642.500 ;
        RECT 1221.370 1642.300 1244.230 1642.440 ;
        RECT 1221.370 1642.240 1221.690 1642.300 ;
        RECT 1243.910 1642.240 1244.230 1642.300 ;
        RECT 1264.150 1642.440 1264.470 1642.500 ;
        RECT 1276.570 1642.440 1276.890 1642.500 ;
        RECT 1264.150 1642.300 1276.890 1642.440 ;
        RECT 1264.150 1642.240 1264.470 1642.300 ;
        RECT 1276.570 1642.240 1276.890 1642.300 ;
        RECT 1351.090 1642.440 1351.410 1642.500 ;
        RECT 1351.550 1642.440 1351.870 1642.500 ;
        RECT 1351.090 1642.300 1351.870 1642.440 ;
        RECT 1351.090 1642.240 1351.410 1642.300 ;
        RECT 1351.550 1642.240 1351.870 1642.300 ;
        RECT 1544.290 1642.440 1544.610 1642.500 ;
        RECT 1545.210 1642.440 1545.530 1642.500 ;
        RECT 1544.290 1642.300 1545.530 1642.440 ;
        RECT 1544.290 1642.240 1544.610 1642.300 ;
        RECT 1545.210 1642.240 1545.530 1642.300 ;
        RECT 1572.810 1635.640 1573.130 1635.700 ;
        RECT 1573.730 1635.640 1574.050 1635.700 ;
        RECT 1572.810 1635.500 1574.050 1635.640 ;
        RECT 1572.810 1635.440 1573.130 1635.500 ;
        RECT 1573.730 1635.440 1574.050 1635.500 ;
        RECT 1532.790 1635.300 1533.110 1635.360 ;
        RECT 1533.710 1635.300 1534.030 1635.360 ;
        RECT 1532.790 1635.160 1534.030 1635.300 ;
        RECT 1532.790 1635.100 1533.110 1635.160 ;
        RECT 1533.710 1635.100 1534.030 1635.160 ;
        RECT 1350.170 1593.820 1350.490 1593.880 ;
        RECT 1351.550 1593.820 1351.870 1593.880 ;
        RECT 1350.170 1593.680 1351.870 1593.820 ;
        RECT 1350.170 1593.620 1350.490 1593.680 ;
        RECT 1351.550 1593.620 1351.870 1593.680 ;
        RECT 1543.830 1593.820 1544.150 1593.880 ;
        RECT 1544.750 1593.820 1545.070 1593.880 ;
        RECT 1543.830 1593.680 1545.070 1593.820 ;
        RECT 1543.830 1593.620 1544.150 1593.680 ;
        RECT 1544.750 1593.620 1545.070 1593.680 ;
        RECT 1559.470 1593.820 1559.790 1593.880 ;
        RECT 1560.390 1593.820 1560.710 1593.880 ;
        RECT 1559.470 1593.680 1560.710 1593.820 ;
        RECT 1559.470 1593.620 1559.790 1593.680 ;
        RECT 1560.390 1593.620 1560.710 1593.680 ;
        RECT 1533.710 1587.020 1534.030 1587.080 ;
        RECT 1534.170 1587.020 1534.490 1587.080 ;
        RECT 1533.710 1586.880 1534.490 1587.020 ;
        RECT 1533.710 1586.820 1534.030 1586.880 ;
        RECT 1534.170 1586.820 1534.490 1586.880 ;
        RECT 1543.830 1587.020 1544.150 1587.080 ;
        RECT 1545.210 1587.020 1545.530 1587.080 ;
        RECT 1543.830 1586.880 1545.530 1587.020 ;
        RECT 1543.830 1586.820 1544.150 1586.880 ;
        RECT 1545.210 1586.820 1545.530 1586.880 ;
        RECT 1350.170 1546.220 1350.490 1546.280 ;
        RECT 1351.550 1546.220 1351.870 1546.280 ;
        RECT 1350.170 1546.080 1351.870 1546.220 ;
        RECT 1350.170 1546.020 1350.490 1546.080 ;
        RECT 1351.550 1546.020 1351.870 1546.080 ;
        RECT 1534.170 1545.680 1534.490 1545.940 ;
        RECT 1559.470 1545.880 1559.790 1545.940 ;
        RECT 1560.390 1545.880 1560.710 1545.940 ;
        RECT 1559.470 1545.740 1560.710 1545.880 ;
        RECT 1559.470 1545.680 1559.790 1545.740 ;
        RECT 1560.390 1545.680 1560.710 1545.740 ;
        RECT 1573.730 1545.880 1574.050 1545.940 ;
        RECT 1574.190 1545.880 1574.510 1545.940 ;
        RECT 1573.730 1545.740 1574.510 1545.880 ;
        RECT 1573.730 1545.680 1574.050 1545.740 ;
        RECT 1574.190 1545.680 1574.510 1545.740 ;
        RECT 1350.630 1545.540 1350.950 1545.600 ;
        RECT 1351.550 1545.540 1351.870 1545.600 ;
        RECT 1350.630 1545.400 1351.870 1545.540 ;
        RECT 1350.630 1545.340 1350.950 1545.400 ;
        RECT 1351.550 1545.340 1351.870 1545.400 ;
        RECT 1534.260 1545.260 1534.400 1545.680 ;
        RECT 1534.170 1545.000 1534.490 1545.260 ;
        RECT 1350.630 1510.860 1350.950 1510.920 ;
        RECT 1351.550 1510.860 1351.870 1510.920 ;
        RECT 1350.630 1510.720 1351.870 1510.860 ;
        RECT 1350.630 1510.660 1350.950 1510.720 ;
        RECT 1351.550 1510.660 1351.870 1510.720 ;
        RECT 1532.790 1497.600 1533.110 1497.660 ;
        RECT 1534.170 1497.600 1534.490 1497.660 ;
        RECT 1532.790 1497.460 1534.490 1497.600 ;
        RECT 1532.790 1497.400 1533.110 1497.460 ;
        RECT 1534.170 1497.400 1534.490 1497.460 ;
        RECT 1350.170 1497.260 1350.490 1497.320 ;
        RECT 1351.550 1497.260 1351.870 1497.320 ;
        RECT 1350.170 1497.120 1351.870 1497.260 ;
        RECT 1350.170 1497.060 1350.490 1497.120 ;
        RECT 1351.550 1497.060 1351.870 1497.120 ;
        RECT 1559.470 1497.260 1559.790 1497.320 ;
        RECT 1560.390 1497.260 1560.710 1497.320 ;
        RECT 1559.470 1497.120 1560.710 1497.260 ;
        RECT 1559.470 1497.060 1559.790 1497.120 ;
        RECT 1560.390 1497.060 1560.710 1497.120 ;
        RECT 1487.250 1461.220 1487.570 1461.280 ;
        RECT 1518.990 1461.220 1519.310 1461.280 ;
        RECT 1487.250 1461.080 1519.310 1461.220 ;
        RECT 1487.250 1461.020 1487.570 1461.080 ;
        RECT 1518.990 1461.020 1519.310 1461.080 ;
        RECT 1486.790 1460.880 1487.110 1460.940 ;
        RECT 1526.350 1460.880 1526.670 1460.940 ;
        RECT 1486.790 1460.740 1526.670 1460.880 ;
        RECT 1486.790 1460.680 1487.110 1460.740 ;
        RECT 1526.350 1460.680 1526.670 1460.740 ;
        RECT 1614.210 1459.520 1614.530 1459.580 ;
        RECT 1893.430 1459.520 1893.750 1459.580 ;
        RECT 1614.210 1459.380 1893.750 1459.520 ;
        RECT 1614.210 1459.320 1614.530 1459.380 ;
        RECT 1893.430 1459.320 1893.750 1459.380 ;
        RECT 1495.530 1459.180 1495.850 1459.240 ;
        RECT 1894.350 1459.180 1894.670 1459.240 ;
        RECT 1495.530 1459.040 1894.670 1459.180 ;
        RECT 1495.530 1458.980 1495.850 1459.040 ;
        RECT 1894.350 1458.980 1894.670 1459.040 ;
        RECT 1350.170 1449.660 1350.490 1449.720 ;
        RECT 1351.550 1449.660 1351.870 1449.720 ;
        RECT 1350.170 1449.520 1351.870 1449.660 ;
        RECT 1350.170 1449.460 1350.490 1449.520 ;
        RECT 1351.550 1449.460 1351.870 1449.520 ;
        RECT 1544.290 1449.320 1544.610 1449.380 ;
        RECT 1545.210 1449.320 1545.530 1449.380 ;
        RECT 1544.290 1449.180 1545.530 1449.320 ;
        RECT 1544.290 1449.120 1544.610 1449.180 ;
        RECT 1545.210 1449.120 1545.530 1449.180 ;
        RECT 1559.470 1449.320 1559.790 1449.380 ;
        RECT 1560.390 1449.320 1560.710 1449.380 ;
        RECT 1559.470 1449.180 1560.710 1449.320 ;
        RECT 1559.470 1449.120 1559.790 1449.180 ;
        RECT 1560.390 1449.120 1560.710 1449.180 ;
        RECT 1573.730 1449.320 1574.050 1449.380 ;
        RECT 1574.190 1449.320 1574.510 1449.380 ;
        RECT 1573.730 1449.180 1574.510 1449.320 ;
        RECT 1573.730 1449.120 1574.050 1449.180 ;
        RECT 1574.190 1449.120 1574.510 1449.180 ;
        RECT 1350.630 1448.980 1350.950 1449.040 ;
        RECT 1351.550 1448.980 1351.870 1449.040 ;
        RECT 1350.630 1448.840 1351.870 1448.980 ;
        RECT 1350.630 1448.780 1350.950 1448.840 ;
        RECT 1351.550 1448.780 1351.870 1448.840 ;
        RECT 1544.290 1435.380 1544.610 1435.440 ;
        RECT 1545.210 1435.380 1545.530 1435.440 ;
        RECT 1544.290 1435.240 1545.530 1435.380 ;
        RECT 1544.290 1435.180 1544.610 1435.240 ;
        RECT 1545.210 1435.180 1545.530 1435.240 ;
        RECT 1350.630 1414.300 1350.950 1414.360 ;
        RECT 1351.550 1414.300 1351.870 1414.360 ;
        RECT 1350.630 1414.160 1351.870 1414.300 ;
        RECT 1350.630 1414.100 1350.950 1414.160 ;
        RECT 1351.550 1414.100 1351.870 1414.160 ;
        RECT 1104.070 1400.700 1104.390 1400.760 ;
        RECT 1104.990 1400.700 1105.310 1400.760 ;
        RECT 1104.070 1400.560 1105.310 1400.700 ;
        RECT 1104.070 1400.500 1104.390 1400.560 ;
        RECT 1104.990 1400.500 1105.310 1400.560 ;
        RECT 1350.170 1400.700 1350.490 1400.760 ;
        RECT 1351.550 1400.700 1351.870 1400.760 ;
        RECT 1350.170 1400.560 1351.870 1400.700 ;
        RECT 1350.170 1400.500 1350.490 1400.560 ;
        RECT 1351.550 1400.500 1351.870 1400.560 ;
        RECT 1543.370 1400.700 1543.690 1400.760 ;
        RECT 1544.750 1400.700 1545.070 1400.760 ;
        RECT 1543.370 1400.560 1545.070 1400.700 ;
        RECT 1543.370 1400.500 1543.690 1400.560 ;
        RECT 1544.750 1400.500 1545.070 1400.560 ;
        RECT 1559.470 1400.700 1559.790 1400.760 ;
        RECT 1560.390 1400.700 1560.710 1400.760 ;
        RECT 1559.470 1400.560 1560.710 1400.700 ;
        RECT 1559.470 1400.500 1559.790 1400.560 ;
        RECT 1560.390 1400.500 1560.710 1400.560 ;
        RECT 1069.110 1353.100 1069.430 1353.160 ;
        RECT 1069.110 1352.960 1069.800 1353.100 ;
        RECT 1069.110 1352.900 1069.430 1352.960 ;
        RECT 1069.660 1352.820 1069.800 1352.960 ;
        RECT 1069.570 1352.560 1069.890 1352.820 ;
        RECT 1104.070 1352.760 1104.390 1352.820 ;
        RECT 1104.990 1352.760 1105.310 1352.820 ;
        RECT 1104.070 1352.620 1105.310 1352.760 ;
        RECT 1104.070 1352.560 1104.390 1352.620 ;
        RECT 1104.990 1352.560 1105.310 1352.620 ;
        RECT 1350.170 1352.760 1350.490 1352.820 ;
        RECT 1351.090 1352.760 1351.410 1352.820 ;
        RECT 1350.170 1352.620 1351.410 1352.760 ;
        RECT 1350.170 1352.560 1350.490 1352.620 ;
        RECT 1351.090 1352.560 1351.410 1352.620 ;
        RECT 1543.370 1352.760 1543.690 1352.820 ;
        RECT 1544.290 1352.760 1544.610 1352.820 ;
        RECT 1543.370 1352.620 1544.610 1352.760 ;
        RECT 1543.370 1352.560 1543.690 1352.620 ;
        RECT 1544.290 1352.560 1544.610 1352.620 ;
        RECT 1559.470 1352.760 1559.790 1352.820 ;
        RECT 1560.390 1352.760 1560.710 1352.820 ;
        RECT 1559.470 1352.620 1560.710 1352.760 ;
        RECT 1559.470 1352.560 1559.790 1352.620 ;
        RECT 1560.390 1352.560 1560.710 1352.620 ;
        RECT 1573.730 1352.760 1574.050 1352.820 ;
        RECT 1574.190 1352.760 1574.510 1352.820 ;
        RECT 1573.730 1352.620 1574.510 1352.760 ;
        RECT 1573.730 1352.560 1574.050 1352.620 ;
        RECT 1574.190 1352.560 1574.510 1352.620 ;
        RECT 1532.790 1338.820 1533.110 1338.880 ;
        RECT 1533.710 1338.820 1534.030 1338.880 ;
        RECT 1532.790 1338.680 1534.030 1338.820 ;
        RECT 1532.790 1338.620 1533.110 1338.680 ;
        RECT 1533.710 1338.620 1534.030 1338.680 ;
        RECT 1350.630 1317.740 1350.950 1317.800 ;
        RECT 1351.550 1317.740 1351.870 1317.800 ;
        RECT 1350.630 1317.600 1351.870 1317.740 ;
        RECT 1350.630 1317.540 1350.950 1317.600 ;
        RECT 1351.550 1317.540 1351.870 1317.600 ;
        RECT 1104.070 1304.140 1104.390 1304.200 ;
        RECT 1104.990 1304.140 1105.310 1304.200 ;
        RECT 1104.070 1304.000 1105.310 1304.140 ;
        RECT 1104.070 1303.940 1104.390 1304.000 ;
        RECT 1104.990 1303.940 1105.310 1304.000 ;
        RECT 1350.170 1304.140 1350.490 1304.200 ;
        RECT 1351.550 1304.140 1351.870 1304.200 ;
        RECT 1350.170 1304.000 1351.870 1304.140 ;
        RECT 1350.170 1303.940 1350.490 1304.000 ;
        RECT 1351.550 1303.940 1351.870 1304.000 ;
        RECT 1069.110 1303.800 1069.430 1303.860 ;
        RECT 1069.570 1303.800 1069.890 1303.860 ;
        RECT 1069.110 1303.660 1069.890 1303.800 ;
        RECT 1069.110 1303.600 1069.430 1303.660 ;
        RECT 1069.570 1303.600 1069.890 1303.660 ;
        RECT 1543.370 1297.340 1543.690 1297.400 ;
        RECT 1545.210 1297.340 1545.530 1297.400 ;
        RECT 1543.370 1297.200 1545.530 1297.340 ;
        RECT 1543.370 1297.140 1543.690 1297.200 ;
        RECT 1545.210 1297.140 1545.530 1297.200 ;
        RECT 1545.210 1270.140 1545.530 1270.200 ;
        RECT 1544.380 1270.000 1545.530 1270.140 ;
        RECT 1544.380 1269.520 1544.520 1270.000 ;
        RECT 1545.210 1269.940 1545.530 1270.000 ;
        RECT 1544.290 1269.260 1544.610 1269.520 ;
        RECT 1104.070 1256.540 1104.390 1256.600 ;
        RECT 1104.990 1256.540 1105.310 1256.600 ;
        RECT 1104.070 1256.400 1105.310 1256.540 ;
        RECT 1104.070 1256.340 1104.390 1256.400 ;
        RECT 1104.990 1256.340 1105.310 1256.400 ;
        RECT 1350.170 1256.540 1350.490 1256.600 ;
        RECT 1350.170 1256.400 1351.780 1256.540 ;
        RECT 1350.170 1256.340 1350.490 1256.400 ;
        RECT 1351.640 1256.260 1351.780 1256.400 ;
        RECT 1351.550 1256.000 1351.870 1256.260 ;
        RECT 1544.290 1220.980 1544.610 1221.240 ;
        RECT 1544.380 1220.560 1544.520 1220.980 ;
        RECT 1544.290 1220.300 1544.610 1220.560 ;
        RECT 1350.630 1207.580 1350.950 1207.640 ;
        RECT 1351.550 1207.580 1351.870 1207.640 ;
        RECT 1350.630 1207.440 1351.870 1207.580 ;
        RECT 1350.630 1207.380 1350.950 1207.440 ;
        RECT 1351.550 1207.380 1351.870 1207.440 ;
        RECT 1350.170 1159.300 1350.490 1159.360 ;
        RECT 1352.010 1159.300 1352.330 1159.360 ;
        RECT 1350.170 1159.160 1352.330 1159.300 ;
        RECT 1350.170 1159.100 1350.490 1159.160 ;
        RECT 1352.010 1159.100 1352.330 1159.160 ;
        RECT 1543.830 1159.300 1544.150 1159.360 ;
        RECT 1544.290 1159.300 1544.610 1159.360 ;
        RECT 1543.830 1159.160 1544.610 1159.300 ;
        RECT 1543.830 1159.100 1544.150 1159.160 ;
        RECT 1544.290 1159.100 1544.610 1159.160 ;
        RECT 1351.090 1111.020 1351.410 1111.080 ;
        RECT 1352.010 1111.020 1352.330 1111.080 ;
        RECT 1351.090 1110.880 1352.330 1111.020 ;
        RECT 1351.090 1110.820 1351.410 1110.880 ;
        RECT 1352.010 1110.820 1352.330 1110.880 ;
        RECT 1530.950 1111.020 1531.270 1111.080 ;
        RECT 1532.790 1111.020 1533.110 1111.080 ;
        RECT 1530.950 1110.880 1533.110 1111.020 ;
        RECT 1530.950 1110.820 1531.270 1110.880 ;
        RECT 1532.790 1110.820 1533.110 1110.880 ;
        RECT 1351.090 1076.820 1351.410 1077.080 ;
        RECT 1351.180 1076.060 1351.320 1076.820 ;
        RECT 1351.090 1075.800 1351.410 1076.060 ;
        RECT 1530.950 1076.000 1531.270 1076.060 ;
        RECT 1532.790 1076.000 1533.110 1076.060 ;
        RECT 1530.950 1075.860 1533.110 1076.000 ;
        RECT 1530.950 1075.800 1531.270 1075.860 ;
        RECT 1532.790 1075.800 1533.110 1075.860 ;
        RECT 1730.590 1062.740 1730.910 1062.800 ;
        RECT 1731.510 1062.740 1731.830 1062.800 ;
        RECT 1730.590 1062.600 1731.830 1062.740 ;
        RECT 1730.590 1062.540 1730.910 1062.600 ;
        RECT 1731.510 1062.540 1731.830 1062.600 ;
        RECT 1489.550 1055.600 1489.870 1055.660 ;
        RECT 1519.450 1055.600 1519.770 1055.660 ;
        RECT 1489.550 1055.460 1519.770 1055.600 ;
        RECT 1489.550 1055.400 1489.870 1055.460 ;
        RECT 1519.450 1055.400 1519.770 1055.460 ;
        RECT 993.670 1052.200 993.990 1052.260 ;
        RECT 1062.670 1052.200 1062.990 1052.260 ;
        RECT 993.670 1052.060 1062.990 1052.200 ;
        RECT 993.670 1052.000 993.990 1052.060 ;
        RECT 1062.670 1052.000 1062.990 1052.060 ;
        RECT 1237.010 1048.800 1237.330 1048.860 ;
        RECT 1239.310 1048.800 1239.630 1048.860 ;
        RECT 1237.010 1048.660 1239.630 1048.800 ;
        RECT 1237.010 1048.600 1237.330 1048.660 ;
        RECT 1239.310 1048.600 1239.630 1048.660 ;
        RECT 982.630 1025.680 982.950 1025.740 ;
        RECT 1146.390 1025.680 1146.710 1025.740 ;
        RECT 982.630 1025.540 1146.710 1025.680 ;
        RECT 982.630 1025.480 982.950 1025.540 ;
        RECT 1146.390 1025.480 1146.710 1025.540 ;
        RECT 975.730 1025.340 976.050 1025.400 ;
        RECT 1152.370 1025.340 1152.690 1025.400 ;
        RECT 975.730 1025.200 1152.690 1025.340 ;
        RECT 975.730 1025.140 976.050 1025.200 ;
        RECT 1152.370 1025.140 1152.690 1025.200 ;
        RECT 972.510 1025.000 972.830 1025.060 ;
        RECT 1154.670 1025.000 1154.990 1025.060 ;
        RECT 972.510 1024.860 1154.990 1025.000 ;
        RECT 972.510 1024.800 972.830 1024.860 ;
        RECT 1154.670 1024.800 1154.990 1024.860 ;
        RECT 1472.070 1025.000 1472.390 1025.060 ;
        RECT 1891.590 1025.000 1891.910 1025.060 ;
        RECT 1472.070 1024.860 1891.910 1025.000 ;
        RECT 1472.070 1024.800 1472.390 1024.860 ;
        RECT 1891.590 1024.800 1891.910 1024.860 ;
        RECT 965.610 1024.660 965.930 1024.720 ;
        RECT 1163.410 1024.660 1163.730 1024.720 ;
        RECT 965.610 1024.520 1163.730 1024.660 ;
        RECT 965.610 1024.460 965.930 1024.520 ;
        RECT 1163.410 1024.460 1163.730 1024.520 ;
        RECT 1385.590 1024.660 1385.910 1024.720 ;
        RECT 1892.050 1024.660 1892.370 1024.720 ;
        RECT 1385.590 1024.520 1892.370 1024.660 ;
        RECT 1385.590 1024.460 1385.910 1024.520 ;
        RECT 1892.050 1024.460 1892.370 1024.520 ;
        RECT 997.350 1021.260 997.670 1021.320 ;
        RECT 1223.210 1021.260 1223.530 1021.320 ;
        RECT 997.350 1021.120 1223.530 1021.260 ;
        RECT 997.350 1021.060 997.670 1021.120 ;
        RECT 1223.210 1021.060 1223.530 1021.120 ;
        RECT 1250.810 1021.260 1251.130 1021.320 ;
        RECT 1339.130 1021.260 1339.450 1021.320 ;
        RECT 1250.810 1021.120 1339.450 1021.260 ;
        RECT 1250.810 1021.060 1251.130 1021.120 ;
        RECT 1339.130 1021.060 1339.450 1021.120 ;
        RECT 1571.890 1021.260 1572.210 1021.320 ;
        RECT 1900.790 1021.260 1901.110 1021.320 ;
        RECT 1571.890 1021.120 1901.110 1021.260 ;
        RECT 1571.890 1021.060 1572.210 1021.120 ;
        RECT 1900.790 1021.060 1901.110 1021.120 ;
        RECT 988.610 1020.920 988.930 1020.980 ;
        RECT 1228.270 1020.920 1228.590 1020.980 ;
        RECT 988.610 1020.780 1228.590 1020.920 ;
        RECT 988.610 1020.720 988.930 1020.780 ;
        RECT 1228.270 1020.720 1228.590 1020.780 ;
        RECT 1243.450 1020.920 1243.770 1020.980 ;
        RECT 1340.970 1020.920 1341.290 1020.980 ;
        RECT 1243.450 1020.780 1341.290 1020.920 ;
        RECT 1243.450 1020.720 1243.770 1020.780 ;
        RECT 1340.970 1020.720 1341.290 1020.780 ;
        RECT 1469.310 1020.920 1469.630 1020.980 ;
        RECT 1704.370 1020.920 1704.690 1020.980 ;
        RECT 1469.310 1020.780 1704.690 1020.920 ;
        RECT 1469.310 1020.720 1469.630 1020.780 ;
        RECT 1704.370 1020.720 1704.690 1020.780 ;
        RECT 1716.790 1020.920 1717.110 1020.980 ;
        RECT 2084.330 1020.920 2084.650 1020.980 ;
        RECT 1716.790 1020.780 2084.650 1020.920 ;
        RECT 1716.790 1020.720 1717.110 1020.780 ;
        RECT 2084.330 1020.720 2084.650 1020.780 ;
        RECT 996.890 1020.580 997.210 1020.640 ;
        RECT 1265.990 1020.580 1266.310 1020.640 ;
        RECT 1337.290 1020.580 1337.610 1020.640 ;
        RECT 996.890 1020.440 1258.860 1020.580 ;
        RECT 996.890 1020.380 997.210 1020.440 ;
        RECT 987.690 1020.240 988.010 1020.300 ;
        RECT 1258.170 1020.240 1258.490 1020.300 ;
        RECT 987.690 1020.100 1258.490 1020.240 ;
        RECT 1258.720 1020.240 1258.860 1020.440 ;
        RECT 1265.990 1020.440 1337.610 1020.580 ;
        RECT 1265.990 1020.380 1266.310 1020.440 ;
        RECT 1337.290 1020.380 1337.610 1020.440 ;
        RECT 1530.490 1020.580 1530.810 1020.640 ;
        RECT 1903.550 1020.580 1903.870 1020.640 ;
        RECT 1530.490 1020.440 1903.870 1020.580 ;
        RECT 1530.490 1020.380 1530.810 1020.440 ;
        RECT 1903.550 1020.380 1903.870 1020.440 ;
        RECT 1268.290 1020.240 1268.610 1020.300 ;
        RECT 1258.720 1020.100 1268.610 1020.240 ;
        RECT 987.690 1020.040 988.010 1020.100 ;
        RECT 1258.170 1020.040 1258.490 1020.100 ;
        RECT 1268.290 1020.040 1268.610 1020.100 ;
        RECT 1286.230 1020.240 1286.550 1020.300 ;
        RECT 1338.670 1020.240 1338.990 1020.300 ;
        RECT 1286.230 1020.100 1338.990 1020.240 ;
        RECT 1286.230 1020.040 1286.550 1020.100 ;
        RECT 1338.670 1020.040 1338.990 1020.100 ;
        RECT 1503.810 1020.240 1504.130 1020.300 ;
        RECT 1897.570 1020.240 1897.890 1020.300 ;
        RECT 1503.810 1020.100 1897.890 1020.240 ;
        RECT 1503.810 1020.040 1504.130 1020.100 ;
        RECT 1897.570 1020.040 1897.890 1020.100 ;
        RECT 996.430 1019.900 996.750 1019.960 ;
        RECT 1290.370 1019.900 1290.690 1019.960 ;
        RECT 996.430 1019.760 1290.690 1019.900 ;
        RECT 996.430 1019.700 996.750 1019.760 ;
        RECT 1290.370 1019.700 1290.690 1019.760 ;
        RECT 1495.070 1019.900 1495.390 1019.960 ;
        RECT 1901.250 1019.900 1901.570 1019.960 ;
        RECT 1495.070 1019.760 1901.570 1019.900 ;
        RECT 1495.070 1019.700 1495.390 1019.760 ;
        RECT 1901.250 1019.700 1901.570 1019.760 ;
        RECT 989.070 1019.560 989.390 1019.620 ;
        RECT 1283.470 1019.560 1283.790 1019.620 ;
        RECT 989.070 1019.420 1283.790 1019.560 ;
        RECT 989.070 1019.360 989.390 1019.420 ;
        RECT 1283.470 1019.360 1283.790 1019.420 ;
        RECT 1462.410 1019.560 1462.730 1019.620 ;
        RECT 1898.490 1019.560 1898.810 1019.620 ;
        RECT 1462.410 1019.420 1898.810 1019.560 ;
        RECT 1462.410 1019.360 1462.730 1019.420 ;
        RECT 1898.490 1019.360 1898.810 1019.420 ;
        RECT 990.450 1019.220 990.770 1019.280 ;
        RECT 1300.030 1019.220 1300.350 1019.280 ;
        RECT 990.450 1019.080 1300.350 1019.220 ;
        RECT 990.450 1019.020 990.770 1019.080 ;
        RECT 1300.030 1019.020 1300.350 1019.080 ;
        RECT 1461.950 1019.220 1462.270 1019.280 ;
        RECT 1898.030 1019.220 1898.350 1019.280 ;
        RECT 1461.950 1019.080 1898.350 1019.220 ;
        RECT 1461.950 1019.020 1462.270 1019.080 ;
        RECT 1898.030 1019.020 1898.350 1019.080 ;
        RECT 988.150 1018.880 988.470 1018.940 ;
        RECT 1312.910 1018.880 1313.230 1018.940 ;
        RECT 988.150 1018.740 1313.230 1018.880 ;
        RECT 988.150 1018.680 988.470 1018.740 ;
        RECT 1312.910 1018.680 1313.230 1018.740 ;
        RECT 1434.810 1018.880 1435.130 1018.940 ;
        RECT 1892.970 1018.880 1893.290 1018.940 ;
        RECT 1434.810 1018.740 1893.290 1018.880 ;
        RECT 1434.810 1018.680 1435.130 1018.740 ;
        RECT 1892.970 1018.680 1893.290 1018.740 ;
        RECT 989.530 1018.540 989.850 1018.600 ;
        RECT 1324.870 1018.540 1325.190 1018.600 ;
        RECT 989.530 1018.400 1325.190 1018.540 ;
        RECT 989.530 1018.340 989.850 1018.400 ;
        RECT 1324.870 1018.340 1325.190 1018.400 ;
        RECT 1357.070 1018.540 1357.390 1018.600 ;
        RECT 1849.270 1018.540 1849.590 1018.600 ;
        RECT 1357.070 1018.400 1849.590 1018.540 ;
        RECT 1357.070 1018.340 1357.390 1018.400 ;
        RECT 1849.270 1018.340 1849.590 1018.400 ;
        RECT 990.910 1018.200 991.230 1018.260 ;
        RECT 1335.450 1018.200 1335.770 1018.260 ;
        RECT 990.910 1018.060 1335.770 1018.200 ;
        RECT 990.910 1018.000 991.230 1018.060 ;
        RECT 1335.450 1018.000 1335.770 1018.060 ;
        RECT 1400.310 1018.200 1400.630 1018.260 ;
        RECT 1898.950 1018.200 1899.270 1018.260 ;
        RECT 1400.310 1018.060 1899.270 1018.200 ;
        RECT 1400.310 1018.000 1400.630 1018.060 ;
        RECT 1898.950 1018.000 1899.270 1018.060 ;
        RECT 989.990 1017.860 990.310 1017.920 ;
        RECT 1347.870 1017.860 1348.190 1017.920 ;
        RECT 989.990 1017.720 1348.190 1017.860 ;
        RECT 989.990 1017.660 990.310 1017.720 ;
        RECT 1347.870 1017.660 1348.190 1017.720 ;
        RECT 1352.010 1017.860 1352.330 1017.920 ;
        RECT 1899.410 1017.860 1899.730 1017.920 ;
        RECT 1352.010 1017.720 1899.730 1017.860 ;
        RECT 1352.010 1017.660 1352.330 1017.720 ;
        RECT 1899.410 1017.660 1899.730 1017.720 ;
        RECT 991.370 1017.520 991.690 1017.580 ;
        RECT 1197.910 1017.520 1198.230 1017.580 ;
        RECT 991.370 1017.380 1198.230 1017.520 ;
        RECT 991.370 1017.320 991.690 1017.380 ;
        RECT 1197.910 1017.320 1198.230 1017.380 ;
        RECT 1203.430 1017.520 1203.750 1017.580 ;
        RECT 1343.270 1017.520 1343.590 1017.580 ;
        RECT 1203.430 1017.380 1343.590 1017.520 ;
        RECT 1203.430 1017.320 1203.750 1017.380 ;
        RECT 1343.270 1017.320 1343.590 1017.380 ;
        RECT 1565.450 1017.520 1565.770 1017.580 ;
        RECT 1890.670 1017.520 1890.990 1017.580 ;
        RECT 1565.450 1017.380 1890.990 1017.520 ;
        RECT 1565.450 1017.320 1565.770 1017.380 ;
        RECT 1890.670 1017.320 1890.990 1017.380 ;
        RECT 992.750 1017.180 993.070 1017.240 ;
        RECT 1159.730 1017.180 1160.050 1017.240 ;
        RECT 992.750 1017.040 1160.050 1017.180 ;
        RECT 992.750 1016.980 993.070 1017.040 ;
        RECT 1159.730 1016.980 1160.050 1017.040 ;
        RECT 1276.110 1017.180 1276.430 1017.240 ;
        RECT 1340.510 1017.180 1340.830 1017.240 ;
        RECT 1276.110 1017.040 1340.830 1017.180 ;
        RECT 1276.110 1016.980 1276.430 1017.040 ;
        RECT 1340.510 1016.980 1340.830 1017.040 ;
        RECT 1478.510 1017.180 1478.830 1017.240 ;
        RECT 1766.470 1017.180 1766.790 1017.240 ;
        RECT 1478.510 1017.040 1766.790 1017.180 ;
        RECT 1478.510 1016.980 1478.830 1017.040 ;
        RECT 1766.470 1016.980 1766.790 1017.040 ;
        RECT 1257.710 1016.840 1258.030 1016.900 ;
        RECT 1286.230 1016.840 1286.550 1016.900 ;
        RECT 1257.710 1016.700 1286.550 1016.840 ;
        RECT 1257.710 1016.640 1258.030 1016.700 ;
        RECT 1286.230 1016.640 1286.550 1016.700 ;
        RECT 1297.270 1016.840 1297.590 1016.900 ;
        RECT 1336.830 1016.840 1337.150 1016.900 ;
        RECT 1297.270 1016.700 1337.150 1016.840 ;
        RECT 1297.270 1016.640 1297.590 1016.700 ;
        RECT 1336.830 1016.640 1337.150 1016.700 ;
        RECT 1512.090 1016.840 1512.410 1016.900 ;
        RECT 1656.070 1016.840 1656.390 1016.900 ;
        RECT 1512.090 1016.700 1656.390 1016.840 ;
        RECT 1512.090 1016.640 1512.410 1016.700 ;
        RECT 1656.070 1016.640 1656.390 1016.700 ;
        RECT 1490.010 1016.500 1490.330 1016.560 ;
        RECT 1622.950 1016.500 1623.270 1016.560 ;
        RECT 1490.010 1016.360 1623.270 1016.500 ;
        RECT 1490.010 1016.300 1490.330 1016.360 ;
        RECT 1622.950 1016.300 1623.270 1016.360 ;
        RECT 1869.970 1014.800 1870.290 1014.860 ;
        RECT 1886.530 1014.800 1886.850 1014.860 ;
        RECT 1869.970 1014.660 1886.850 1014.800 ;
        RECT 1869.970 1014.600 1870.290 1014.660 ;
        RECT 1886.530 1014.600 1886.850 1014.660 ;
        RECT 1333.150 1014.460 1333.470 1014.520 ;
        RECT 1330.940 1014.320 1333.470 1014.460 ;
        RECT 1048.410 1014.120 1048.730 1014.180 ;
        RECT 1214.470 1014.120 1214.790 1014.180 ;
        RECT 1238.390 1014.120 1238.710 1014.180 ;
        RECT 1048.410 1013.980 1214.790 1014.120 ;
        RECT 1048.410 1013.920 1048.730 1013.980 ;
        RECT 1214.470 1013.920 1214.790 1013.980 ;
        RECT 1229.740 1013.980 1238.710 1014.120 ;
        RECT 977.110 1013.780 977.430 1013.840 ;
        RECT 1189.630 1013.780 1189.950 1013.840 ;
        RECT 977.110 1013.640 1189.950 1013.780 ;
        RECT 977.110 1013.580 977.430 1013.640 ;
        RECT 1189.630 1013.580 1189.950 1013.640 ;
        RECT 984.470 1013.440 984.790 1013.500 ;
        RECT 1145.470 1013.440 1145.790 1013.500 ;
        RECT 984.470 1013.300 1145.790 1013.440 ;
        RECT 984.470 1013.240 984.790 1013.300 ;
        RECT 1145.470 1013.240 1145.790 1013.300 ;
        RECT 1173.070 1013.440 1173.390 1013.500 ;
        RECT 1218.610 1013.440 1218.930 1013.500 ;
        RECT 1173.070 1013.300 1218.930 1013.440 ;
        RECT 1173.070 1013.240 1173.390 1013.300 ;
        RECT 1218.610 1013.240 1218.930 1013.300 ;
        RECT 789.890 1013.100 790.210 1013.160 ;
        RECT 888.330 1013.100 888.650 1013.160 ;
        RECT 789.890 1012.960 888.650 1013.100 ;
        RECT 789.890 1012.900 790.210 1012.960 ;
        RECT 888.330 1012.900 888.650 1012.960 ;
        RECT 983.090 1013.100 983.410 1013.160 ;
        RECT 1012.530 1013.100 1012.850 1013.160 ;
        RECT 983.090 1012.960 1012.850 1013.100 ;
        RECT 983.090 1012.900 983.410 1012.960 ;
        RECT 1012.530 1012.900 1012.850 1012.960 ;
        RECT 1020.810 1013.100 1021.130 1013.160 ;
        RECT 1196.070 1013.100 1196.390 1013.160 ;
        RECT 1204.350 1013.100 1204.670 1013.160 ;
        RECT 1020.810 1012.960 1196.390 1013.100 ;
        RECT 1020.810 1012.900 1021.130 1012.960 ;
        RECT 1196.070 1012.900 1196.390 1012.960 ;
        RECT 1196.620 1012.960 1204.670 1013.100 ;
        RECT 796.790 1012.760 797.110 1012.820 ;
        RECT 844.630 1012.760 844.950 1012.820 ;
        RECT 796.790 1012.620 844.950 1012.760 ;
        RECT 796.790 1012.560 797.110 1012.620 ;
        RECT 844.630 1012.560 844.950 1012.620 ;
        RECT 977.570 1012.760 977.890 1012.820 ;
        RECT 1196.620 1012.760 1196.760 1012.960 ;
        RECT 1204.350 1012.900 1204.670 1012.960 ;
        RECT 1213.550 1013.100 1213.870 1013.160 ;
        RECT 1229.740 1013.100 1229.880 1013.980 ;
        RECT 1238.390 1013.920 1238.710 1013.980 ;
        RECT 1255.410 1014.120 1255.730 1014.180 ;
        RECT 1330.940 1014.120 1331.080 1014.320 ;
        RECT 1333.150 1014.260 1333.470 1014.320 ;
        RECT 1790.390 1014.460 1790.710 1014.520 ;
        RECT 1790.390 1014.320 1828.340 1014.460 ;
        RECT 1790.390 1014.260 1790.710 1014.320 ;
        RECT 1255.410 1013.980 1331.080 1014.120 ;
        RECT 1331.310 1014.120 1331.630 1014.180 ;
        RECT 1334.530 1014.120 1334.850 1014.180 ;
        RECT 1331.310 1013.980 1334.850 1014.120 ;
        RECT 1255.410 1013.920 1255.730 1013.980 ;
        RECT 1331.310 1013.920 1331.630 1013.980 ;
        RECT 1334.530 1013.920 1334.850 1013.980 ;
        RECT 1338.670 1014.120 1338.990 1014.180 ;
        RECT 1353.390 1014.120 1353.710 1014.180 ;
        RECT 1338.670 1013.980 1353.710 1014.120 ;
        RECT 1338.670 1013.920 1338.990 1013.980 ;
        RECT 1353.390 1013.920 1353.710 1013.980 ;
        RECT 1355.230 1014.120 1355.550 1014.180 ;
        RECT 1357.990 1014.120 1358.310 1014.180 ;
        RECT 1513.010 1014.120 1513.330 1014.180 ;
        RECT 1355.230 1013.980 1358.310 1014.120 ;
        RECT 1355.230 1013.920 1355.550 1013.980 ;
        RECT 1357.990 1013.920 1358.310 1013.980 ;
        RECT 1511.720 1013.980 1513.330 1014.120 ;
        RECT 1261.390 1013.780 1261.710 1013.840 ;
        RECT 1341.430 1013.780 1341.750 1013.840 ;
        RECT 1261.390 1013.640 1341.750 1013.780 ;
        RECT 1261.390 1013.580 1261.710 1013.640 ;
        RECT 1341.430 1013.580 1341.750 1013.640 ;
        RECT 1488.630 1013.780 1488.950 1013.840 ;
        RECT 1511.720 1013.780 1511.860 1013.980 ;
        RECT 1513.010 1013.920 1513.330 1013.980 ;
        RECT 1538.310 1014.120 1538.630 1014.180 ;
        RECT 1550.270 1014.120 1550.590 1014.180 ;
        RECT 1762.790 1014.120 1763.110 1014.180 ;
        RECT 1538.310 1013.980 1546.820 1014.120 ;
        RECT 1538.310 1013.920 1538.630 1013.980 ;
        RECT 1528.190 1013.780 1528.510 1013.840 ;
        RECT 1488.630 1013.640 1511.860 1013.780 ;
        RECT 1512.180 1013.640 1528.510 1013.780 ;
        RECT 1488.630 1013.580 1488.950 1013.640 ;
        RECT 1286.690 1013.440 1287.010 1013.500 ;
        RECT 1213.550 1012.960 1229.880 1013.100 ;
        RECT 1231.580 1013.300 1287.010 1013.440 ;
        RECT 1213.550 1012.900 1213.870 1012.960 ;
        RECT 977.570 1012.620 1196.760 1012.760 ;
        RECT 1203.890 1012.760 1204.210 1012.820 ;
        RECT 1231.580 1012.760 1231.720 1013.300 ;
        RECT 1286.690 1013.240 1287.010 1013.300 ;
        RECT 1287.610 1013.440 1287.930 1013.500 ;
        RECT 1289.910 1013.440 1290.230 1013.500 ;
        RECT 1287.610 1013.300 1290.230 1013.440 ;
        RECT 1287.610 1013.240 1287.930 1013.300 ;
        RECT 1289.910 1013.240 1290.230 1013.300 ;
        RECT 1293.590 1013.440 1293.910 1013.500 ;
        RECT 1317.970 1013.440 1318.290 1013.500 ;
        RECT 1293.590 1013.300 1318.290 1013.440 ;
        RECT 1293.590 1013.240 1293.910 1013.300 ;
        RECT 1317.970 1013.240 1318.290 1013.300 ;
        RECT 1487.710 1013.440 1488.030 1013.500 ;
        RECT 1509.330 1013.440 1509.650 1013.500 ;
        RECT 1487.710 1013.300 1509.650 1013.440 ;
        RECT 1487.710 1013.240 1488.030 1013.300 ;
        RECT 1509.330 1013.240 1509.650 1013.300 ;
        RECT 1253.110 1013.100 1253.430 1013.160 ;
        RECT 1345.570 1013.100 1345.890 1013.160 ;
        RECT 1253.110 1012.960 1345.890 1013.100 ;
        RECT 1253.110 1012.900 1253.430 1012.960 ;
        RECT 1345.570 1012.900 1345.890 1012.960 ;
        RECT 1496.910 1013.100 1497.230 1013.160 ;
        RECT 1511.630 1013.100 1511.950 1013.160 ;
        RECT 1496.910 1012.960 1511.950 1013.100 ;
        RECT 1496.910 1012.900 1497.230 1012.960 ;
        RECT 1511.630 1012.900 1511.950 1012.960 ;
        RECT 1346.490 1012.760 1346.810 1012.820 ;
        RECT 1203.890 1012.620 1231.720 1012.760 ;
        RECT 1236.640 1012.620 1346.810 1012.760 ;
        RECT 977.570 1012.560 977.890 1012.620 ;
        RECT 1203.890 1012.560 1204.210 1012.620 ;
        RECT 782.990 1012.420 783.310 1012.480 ;
        RECT 884.190 1012.420 884.510 1012.480 ;
        RECT 782.990 1012.280 884.510 1012.420 ;
        RECT 782.990 1012.220 783.310 1012.280 ;
        RECT 884.190 1012.220 884.510 1012.280 ;
        RECT 1000.110 1012.420 1000.430 1012.480 ;
        RECT 1179.970 1012.420 1180.290 1012.480 ;
        RECT 1000.110 1012.280 1180.290 1012.420 ;
        RECT 1000.110 1012.220 1000.430 1012.280 ;
        RECT 1179.970 1012.220 1180.290 1012.280 ;
        RECT 1180.430 1012.420 1180.750 1012.480 ;
        RECT 1186.410 1012.420 1186.730 1012.480 ;
        RECT 1180.430 1012.280 1186.730 1012.420 ;
        RECT 1180.430 1012.220 1180.750 1012.280 ;
        RECT 1186.410 1012.220 1186.730 1012.280 ;
        RECT 1196.990 1012.420 1197.310 1012.480 ;
        RECT 1218.150 1012.420 1218.470 1012.480 ;
        RECT 1196.990 1012.280 1218.470 1012.420 ;
        RECT 1196.990 1012.220 1197.310 1012.280 ;
        RECT 1218.150 1012.220 1218.470 1012.280 ;
        RECT 1218.610 1012.420 1218.930 1012.480 ;
        RECT 1221.370 1012.420 1221.690 1012.480 ;
        RECT 1218.610 1012.280 1221.690 1012.420 ;
        RECT 1218.610 1012.220 1218.930 1012.280 ;
        RECT 1221.370 1012.220 1221.690 1012.280 ;
        RECT 707.090 1012.080 707.410 1012.140 ;
        RECT 841.870 1012.080 842.190 1012.140 ;
        RECT 707.090 1011.940 842.190 1012.080 ;
        RECT 707.090 1011.880 707.410 1011.940 ;
        RECT 841.870 1011.880 842.190 1011.940 ;
        RECT 984.010 1012.080 984.330 1012.140 ;
        RECT 1173.070 1012.080 1173.390 1012.140 ;
        RECT 984.010 1011.940 1173.390 1012.080 ;
        RECT 984.010 1011.880 984.330 1011.940 ;
        RECT 1173.070 1011.880 1173.390 1011.940 ;
        RECT 769.190 1011.740 769.510 1011.800 ;
        RECT 910.870 1011.740 911.190 1011.800 ;
        RECT 769.190 1011.600 911.190 1011.740 ;
        RECT 769.190 1011.540 769.510 1011.600 ;
        RECT 910.870 1011.540 911.190 1011.600 ;
        RECT 976.190 1011.740 976.510 1011.800 ;
        RECT 1003.790 1011.740 1004.110 1011.800 ;
        RECT 976.190 1011.600 1004.110 1011.740 ;
        RECT 976.190 1011.540 976.510 1011.600 ;
        RECT 1003.790 1011.540 1004.110 1011.600 ;
        RECT 1038.290 1011.740 1038.610 1011.800 ;
        RECT 1093.030 1011.740 1093.350 1011.800 ;
        RECT 1038.290 1011.600 1093.350 1011.740 ;
        RECT 1038.290 1011.540 1038.610 1011.600 ;
        RECT 1093.030 1011.540 1093.350 1011.600 ;
        RECT 1104.070 1011.740 1104.390 1011.800 ;
        RECT 1105.450 1011.740 1105.770 1011.800 ;
        RECT 1104.070 1011.600 1105.770 1011.740 ;
        RECT 1104.070 1011.540 1104.390 1011.600 ;
        RECT 1105.450 1011.540 1105.770 1011.600 ;
        RECT 1145.010 1011.740 1145.330 1011.800 ;
        RECT 1197.450 1011.740 1197.770 1011.800 ;
        RECT 1145.010 1011.600 1197.770 1011.740 ;
        RECT 1145.010 1011.540 1145.330 1011.600 ;
        RECT 1197.450 1011.540 1197.770 1011.600 ;
        RECT 1217.230 1011.740 1217.550 1011.800 ;
        RECT 1236.640 1011.740 1236.780 1012.620 ;
        RECT 1346.490 1012.560 1346.810 1012.620 ;
        RECT 1489.550 1012.760 1489.870 1012.820 ;
        RECT 1512.180 1012.760 1512.320 1013.640 ;
        RECT 1528.190 1013.580 1528.510 1013.640 ;
        RECT 1530.950 1013.780 1531.270 1013.840 ;
        RECT 1546.680 1013.780 1546.820 1013.980 ;
        RECT 1550.270 1013.980 1763.110 1014.120 ;
        RECT 1550.270 1013.920 1550.590 1013.980 ;
        RECT 1762.790 1013.920 1763.110 1013.980 ;
        RECT 1777.510 1014.120 1777.830 1014.180 ;
        RECT 1779.810 1014.120 1780.130 1014.180 ;
        RECT 1777.510 1013.980 1780.130 1014.120 ;
        RECT 1828.200 1014.120 1828.340 1014.320 ;
        RECT 1869.970 1014.120 1870.290 1014.180 ;
        RECT 1828.200 1013.980 1870.290 1014.120 ;
        RECT 1777.510 1013.920 1777.830 1013.980 ;
        RECT 1779.810 1013.920 1780.130 1013.980 ;
        RECT 1869.970 1013.920 1870.290 1013.980 ;
        RECT 2061.790 1014.120 2062.110 1014.180 ;
        RECT 2287.190 1014.120 2287.510 1014.180 ;
        RECT 2061.790 1013.980 2287.510 1014.120 ;
        RECT 2061.790 1013.920 2062.110 1013.980 ;
        RECT 2287.190 1013.920 2287.510 1013.980 ;
        RECT 1886.070 1013.780 1886.390 1013.840 ;
        RECT 1530.950 1013.640 1546.360 1013.780 ;
        RECT 1546.680 1013.640 1886.390 1013.780 ;
        RECT 1530.950 1013.580 1531.270 1013.640 ;
        RECT 1512.550 1013.440 1512.870 1013.500 ;
        RECT 1512.550 1013.300 1545.900 1013.440 ;
        RECT 1512.550 1013.240 1512.870 1013.300 ;
        RECT 1524.510 1013.100 1524.830 1013.160 ;
        RECT 1542.910 1013.100 1543.230 1013.160 ;
        RECT 1524.510 1012.960 1543.230 1013.100 ;
        RECT 1524.510 1012.900 1524.830 1012.960 ;
        RECT 1542.910 1012.900 1543.230 1012.960 ;
        RECT 1489.550 1012.620 1512.320 1012.760 ;
        RECT 1518.990 1012.760 1519.310 1012.820 ;
        RECT 1521.290 1012.760 1521.610 1012.820 ;
        RECT 1518.990 1012.620 1521.610 1012.760 ;
        RECT 1489.550 1012.560 1489.870 1012.620 ;
        RECT 1518.990 1012.560 1519.310 1012.620 ;
        RECT 1521.290 1012.560 1521.610 1012.620 ;
        RECT 1541.530 1012.760 1541.850 1012.820 ;
        RECT 1545.210 1012.760 1545.530 1012.820 ;
        RECT 1541.530 1012.620 1545.530 1012.760 ;
        RECT 1545.760 1012.760 1545.900 1013.300 ;
        RECT 1546.220 1013.100 1546.360 1013.640 ;
        RECT 1886.070 1013.580 1886.390 1013.640 ;
        RECT 1998.310 1013.780 1998.630 1013.840 ;
        RECT 2000.610 1013.780 2000.930 1013.840 ;
        RECT 1998.310 1013.640 2000.930 1013.780 ;
        RECT 1998.310 1013.580 1998.630 1013.640 ;
        RECT 2000.610 1013.580 2000.930 1013.640 ;
        RECT 2057.190 1013.780 2057.510 1013.840 ;
        RECT 2287.650 1013.780 2287.970 1013.840 ;
        RECT 2057.190 1013.640 2287.970 1013.780 ;
        RECT 2057.190 1013.580 2057.510 1013.640 ;
        RECT 2287.650 1013.580 2287.970 1013.640 ;
        RECT 1553.030 1013.440 1553.350 1013.500 ;
        RECT 1673.090 1013.440 1673.410 1013.500 ;
        RECT 1553.030 1013.300 1673.410 1013.440 ;
        RECT 1553.030 1013.240 1553.350 1013.300 ;
        RECT 1673.090 1013.240 1673.410 1013.300 ;
        RECT 1708.510 1013.440 1708.830 1013.500 ;
        RECT 1762.790 1013.440 1763.110 1013.500 ;
        RECT 1790.390 1013.440 1790.710 1013.500 ;
        RECT 1708.510 1013.300 1752.900 1013.440 ;
        RECT 1708.510 1013.240 1708.830 1013.300 ;
        RECT 1625.250 1013.100 1625.570 1013.160 ;
        RECT 1546.220 1012.960 1625.570 1013.100 ;
        RECT 1625.250 1012.900 1625.570 1012.960 ;
        RECT 1724.150 1013.100 1724.470 1013.160 ;
        RECT 1751.290 1013.100 1751.610 1013.160 ;
        RECT 1724.150 1012.960 1751.610 1013.100 ;
        RECT 1724.150 1012.900 1724.470 1012.960 ;
        RECT 1751.290 1012.900 1751.610 1012.960 ;
        RECT 1628.470 1012.760 1628.790 1012.820 ;
        RECT 1545.760 1012.620 1628.790 1012.760 ;
        RECT 1541.530 1012.560 1541.850 1012.620 ;
        RECT 1545.210 1012.560 1545.530 1012.620 ;
        RECT 1628.470 1012.560 1628.790 1012.620 ;
        RECT 1721.390 1012.760 1721.710 1012.820 ;
        RECT 1724.610 1012.760 1724.930 1012.820 ;
        RECT 1721.390 1012.620 1724.930 1012.760 ;
        RECT 1721.390 1012.560 1721.710 1012.620 ;
        RECT 1724.610 1012.560 1724.930 1012.620 ;
        RECT 1743.010 1012.760 1743.330 1012.820 ;
        RECT 1745.310 1012.760 1745.630 1012.820 ;
        RECT 1743.010 1012.620 1745.630 1012.760 ;
        RECT 1743.010 1012.560 1743.330 1012.620 ;
        RECT 1745.310 1012.560 1745.630 1012.620 ;
        RECT 1747.610 1012.760 1747.930 1012.820 ;
        RECT 1751.750 1012.760 1752.070 1012.820 ;
        RECT 1747.610 1012.620 1752.070 1012.760 ;
        RECT 1752.760 1012.760 1752.900 1013.300 ;
        RECT 1762.790 1013.300 1790.710 1013.440 ;
        RECT 1762.790 1013.240 1763.110 1013.300 ;
        RECT 1790.390 1013.240 1790.710 1013.300 ;
        RECT 1790.850 1013.440 1791.170 1013.500 ;
        RECT 1793.610 1013.440 1793.930 1013.500 ;
        RECT 1790.850 1013.300 1793.930 1013.440 ;
        RECT 1790.850 1013.240 1791.170 1013.300 ;
        RECT 1793.610 1013.240 1793.930 1013.300 ;
        RECT 1794.070 1013.440 1794.390 1013.500 ;
        RECT 2086.170 1013.440 2086.490 1013.500 ;
        RECT 1794.070 1013.300 2086.490 1013.440 ;
        RECT 1794.070 1013.240 1794.390 1013.300 ;
        RECT 2086.170 1013.240 2086.490 1013.300 ;
        RECT 1753.130 1013.100 1753.450 1013.160 ;
        RECT 2085.710 1013.100 2086.030 1013.160 ;
        RECT 1753.130 1012.960 2086.030 1013.100 ;
        RECT 1753.130 1012.900 1753.450 1012.960 ;
        RECT 2085.710 1012.900 2086.030 1012.960 ;
        RECT 2085.250 1012.760 2085.570 1012.820 ;
        RECT 1752.760 1012.620 2085.570 1012.760 ;
        RECT 1747.610 1012.560 1747.930 1012.620 ;
        RECT 1751.750 1012.560 1752.070 1012.620 ;
        RECT 2085.250 1012.560 2085.570 1012.620 ;
        RECT 1237.010 1012.420 1237.330 1012.480 ;
        RECT 1340.050 1012.420 1340.370 1012.480 ;
        RECT 1237.010 1012.280 1340.370 1012.420 ;
        RECT 1237.010 1012.220 1237.330 1012.280 ;
        RECT 1340.050 1012.220 1340.370 1012.280 ;
        RECT 1411.350 1012.420 1411.670 1012.480 ;
        RECT 1414.110 1012.420 1414.430 1012.480 ;
        RECT 1411.350 1012.280 1414.430 1012.420 ;
        RECT 1411.350 1012.220 1411.670 1012.280 ;
        RECT 1414.110 1012.220 1414.430 1012.280 ;
        RECT 1467.470 1012.420 1467.790 1012.480 ;
        RECT 1468.850 1012.420 1469.170 1012.480 ;
        RECT 1467.470 1012.280 1469.170 1012.420 ;
        RECT 1467.470 1012.220 1467.790 1012.280 ;
        RECT 1468.850 1012.220 1469.170 1012.280 ;
        RECT 1480.350 1012.420 1480.670 1012.480 ;
        RECT 1482.650 1012.420 1482.970 1012.480 ;
        RECT 1480.350 1012.280 1482.970 1012.420 ;
        RECT 1480.350 1012.220 1480.670 1012.280 ;
        RECT 1482.650 1012.220 1482.970 1012.280 ;
        RECT 1501.970 1012.420 1502.290 1012.480 ;
        RECT 1875.490 1012.420 1875.810 1012.480 ;
        RECT 1893.890 1012.420 1894.210 1012.480 ;
        RECT 1501.970 1012.280 1873.880 1012.420 ;
        RECT 1501.970 1012.220 1502.290 1012.280 ;
        RECT 1297.730 1012.080 1298.050 1012.140 ;
        RECT 1217.230 1011.600 1236.780 1011.740 ;
        RECT 1244.460 1011.940 1298.050 1012.080 ;
        RECT 1217.230 1011.540 1217.550 1011.600 ;
        RECT 762.290 1011.400 762.610 1011.460 ;
        RECT 905.350 1011.400 905.670 1011.460 ;
        RECT 762.290 1011.260 905.670 1011.400 ;
        RECT 762.290 1011.200 762.610 1011.260 ;
        RECT 905.350 1011.200 905.670 1011.260 ;
        RECT 995.970 1011.400 996.290 1011.460 ;
        RECT 1053.470 1011.400 1053.790 1011.460 ;
        RECT 995.970 1011.260 1053.790 1011.400 ;
        RECT 995.970 1011.200 996.290 1011.260 ;
        RECT 1053.470 1011.200 1053.790 1011.260 ;
        RECT 1100.390 1011.400 1100.710 1011.460 ;
        RECT 1145.470 1011.400 1145.790 1011.460 ;
        RECT 1100.390 1011.260 1145.790 1011.400 ;
        RECT 1100.390 1011.200 1100.710 1011.260 ;
        RECT 1145.470 1011.200 1145.790 1011.260 ;
        RECT 1196.530 1011.400 1196.850 1011.460 ;
        RECT 1244.460 1011.400 1244.600 1011.940 ;
        RECT 1297.730 1011.880 1298.050 1011.940 ;
        RECT 1324.410 1012.080 1324.730 1012.140 ;
        RECT 1334.070 1012.080 1334.390 1012.140 ;
        RECT 1324.410 1011.940 1334.390 1012.080 ;
        RECT 1324.410 1011.880 1324.730 1011.940 ;
        RECT 1334.070 1011.880 1334.390 1011.940 ;
        RECT 1334.530 1012.080 1334.850 1012.140 ;
        RECT 1352.930 1012.080 1353.250 1012.140 ;
        RECT 1334.530 1011.940 1353.250 1012.080 ;
        RECT 1334.530 1011.880 1334.850 1011.940 ;
        RECT 1352.930 1011.880 1353.250 1011.940 ;
        RECT 1441.250 1012.080 1441.570 1012.140 ;
        RECT 1610.990 1012.080 1611.310 1012.140 ;
        RECT 1441.250 1011.940 1611.310 1012.080 ;
        RECT 1441.250 1011.880 1441.570 1011.940 ;
        RECT 1610.990 1011.880 1611.310 1011.940 ;
        RECT 1665.270 1012.080 1665.590 1012.140 ;
        RECT 1669.410 1012.080 1669.730 1012.140 ;
        RECT 1665.270 1011.940 1669.730 1012.080 ;
        RECT 1665.270 1011.880 1665.590 1011.940 ;
        RECT 1669.410 1011.880 1669.730 1011.940 ;
        RECT 1669.870 1012.080 1670.190 1012.140 ;
        RECT 1872.730 1012.080 1873.050 1012.140 ;
        RECT 1669.870 1011.940 1873.050 1012.080 ;
        RECT 1669.870 1011.880 1670.190 1011.940 ;
        RECT 1872.730 1011.880 1873.050 1011.940 ;
        RECT 1286.690 1011.740 1287.010 1011.800 ;
        RECT 1304.170 1011.740 1304.490 1011.800 ;
        RECT 1286.690 1011.600 1304.490 1011.740 ;
        RECT 1286.690 1011.540 1287.010 1011.600 ;
        RECT 1304.170 1011.540 1304.490 1011.600 ;
        RECT 1304.630 1011.740 1304.950 1011.800 ;
        RECT 1332.690 1011.740 1333.010 1011.800 ;
        RECT 1304.630 1011.600 1333.010 1011.740 ;
        RECT 1304.630 1011.540 1304.950 1011.600 ;
        RECT 1332.690 1011.540 1333.010 1011.600 ;
        RECT 1333.150 1011.740 1333.470 1011.800 ;
        RECT 1353.850 1011.740 1354.170 1011.800 ;
        RECT 1333.150 1011.600 1354.170 1011.740 ;
        RECT 1333.150 1011.540 1333.470 1011.600 ;
        RECT 1353.850 1011.540 1354.170 1011.600 ;
        RECT 1506.570 1011.740 1506.890 1011.800 ;
        RECT 1873.190 1011.740 1873.510 1011.800 ;
        RECT 1506.570 1011.600 1873.510 1011.740 ;
        RECT 1873.740 1011.740 1873.880 1012.280 ;
        RECT 1875.490 1012.280 1894.210 1012.420 ;
        RECT 1875.490 1012.220 1875.810 1012.280 ;
        RECT 1893.890 1012.220 1894.210 1012.280 ;
        RECT 2000.610 1012.420 2000.930 1012.480 ;
        RECT 2294.090 1012.420 2294.410 1012.480 ;
        RECT 2000.610 1012.280 2294.410 1012.420 ;
        RECT 2000.610 1012.220 2000.930 1012.280 ;
        RECT 2294.090 1012.220 2294.410 1012.280 ;
        RECT 1874.110 1012.080 1874.430 1012.140 ;
        RECT 2046.610 1012.080 2046.930 1012.140 ;
        RECT 2048.910 1012.080 2049.230 1012.140 ;
        RECT 2087.090 1012.080 2087.410 1012.140 ;
        RECT 1874.110 1011.940 2046.380 1012.080 ;
        RECT 1874.110 1011.880 1874.430 1011.940 ;
        RECT 1892.510 1011.740 1892.830 1011.800 ;
        RECT 1873.740 1011.600 1892.830 1011.740 ;
        RECT 1506.570 1011.540 1506.890 1011.600 ;
        RECT 1873.190 1011.540 1873.510 1011.600 ;
        RECT 1892.510 1011.540 1892.830 1011.600 ;
        RECT 1196.530 1011.260 1244.600 1011.400 ;
        RECT 1245.290 1011.400 1245.610 1011.460 ;
        RECT 1294.050 1011.400 1294.370 1011.460 ;
        RECT 1346.950 1011.400 1347.270 1011.460 ;
        RECT 1245.290 1011.260 1294.370 1011.400 ;
        RECT 1196.530 1011.200 1196.850 1011.260 ;
        RECT 1245.290 1011.200 1245.610 1011.260 ;
        RECT 1294.050 1011.200 1294.370 1011.260 ;
        RECT 1294.600 1011.260 1347.270 1011.400 ;
        RECT 517.110 1011.060 517.430 1011.120 ;
        RECT 712.610 1011.060 712.930 1011.120 ;
        RECT 517.110 1010.920 712.930 1011.060 ;
        RECT 517.110 1010.860 517.430 1010.920 ;
        RECT 712.610 1010.860 712.930 1010.920 ;
        RECT 755.390 1011.060 755.710 1011.120 ;
        RECT 901.210 1011.060 901.530 1011.120 ;
        RECT 755.390 1010.920 901.530 1011.060 ;
        RECT 755.390 1010.860 755.710 1010.920 ;
        RECT 901.210 1010.860 901.530 1010.920 ;
        RECT 995.050 1011.060 995.370 1011.120 ;
        RECT 1289.910 1011.060 1290.230 1011.120 ;
        RECT 1294.600 1011.060 1294.740 1011.260 ;
        RECT 1346.950 1011.200 1347.270 1011.260 ;
        RECT 1444.010 1011.400 1444.330 1011.460 ;
        RECT 1479.890 1011.400 1480.210 1011.460 ;
        RECT 1444.010 1011.260 1480.210 1011.400 ;
        RECT 1444.010 1011.200 1444.330 1011.260 ;
        RECT 1479.890 1011.200 1480.210 1011.260 ;
        RECT 1484.950 1011.400 1485.270 1011.460 ;
        RECT 1899.870 1011.400 1900.190 1011.460 ;
        RECT 1484.950 1011.260 1900.190 1011.400 ;
        RECT 2046.240 1011.400 2046.380 1011.940 ;
        RECT 2046.610 1011.940 2049.230 1012.080 ;
        RECT 2046.610 1011.880 2046.930 1011.940 ;
        RECT 2048.910 1011.880 2049.230 1011.940 ;
        RECT 2049.920 1011.940 2087.410 1012.080 ;
        RECT 2049.920 1011.400 2050.060 1011.940 ;
        RECT 2087.090 1011.880 2087.410 1011.940 ;
        RECT 2069.150 1011.740 2069.470 1011.800 ;
        RECT 2540.190 1011.740 2540.510 1011.800 ;
        RECT 2069.150 1011.600 2540.510 1011.740 ;
        RECT 2069.150 1011.540 2069.470 1011.600 ;
        RECT 2540.190 1011.540 2540.510 1011.600 ;
        RECT 2046.240 1011.260 2050.060 1011.400 ;
        RECT 2053.050 1011.400 2053.370 1011.460 ;
        RECT 2539.730 1011.400 2540.050 1011.460 ;
        RECT 2053.050 1011.260 2540.050 1011.400 ;
        RECT 1484.950 1011.200 1485.270 1011.260 ;
        RECT 1899.870 1011.200 1900.190 1011.260 ;
        RECT 2053.050 1011.200 2053.370 1011.260 ;
        RECT 2539.730 1011.200 2540.050 1011.260 ;
        RECT 995.050 1010.920 1288.990 1011.060 ;
        RECT 995.050 1010.860 995.370 1010.920 ;
        RECT 468.810 1010.720 469.130 1010.780 ;
        RECT 673.510 1010.720 673.830 1010.780 ;
        RECT 468.810 1010.580 673.830 1010.720 ;
        RECT 468.810 1010.520 469.130 1010.580 ;
        RECT 673.510 1010.520 673.830 1010.580 ;
        RECT 720.890 1010.720 721.210 1010.780 ;
        RECT 892.470 1010.720 892.790 1010.780 ;
        RECT 720.890 1010.580 892.790 1010.720 ;
        RECT 720.890 1010.520 721.210 1010.580 ;
        RECT 892.470 1010.520 892.790 1010.580 ;
        RECT 995.510 1010.720 995.830 1010.780 ;
        RECT 1288.850 1010.720 1288.990 1010.920 ;
        RECT 1289.910 1010.920 1294.740 1011.060 ;
        RECT 1322.570 1011.060 1322.890 1011.120 ;
        RECT 1346.030 1011.060 1346.350 1011.120 ;
        RECT 1322.570 1010.920 1346.350 1011.060 ;
        RECT 1289.910 1010.860 1290.230 1010.920 ;
        RECT 1322.570 1010.860 1322.890 1010.920 ;
        RECT 1346.030 1010.860 1346.350 1010.920 ;
        RECT 1427.910 1011.060 1428.230 1011.120 ;
        RECT 1891.130 1011.060 1891.450 1011.120 ;
        RECT 1427.910 1010.920 1891.450 1011.060 ;
        RECT 1427.910 1010.860 1428.230 1010.920 ;
        RECT 1891.130 1010.860 1891.450 1010.920 ;
        RECT 2041.550 1011.060 2041.870 1011.120 ;
        RECT 2539.270 1011.060 2539.590 1011.120 ;
        RECT 2041.550 1010.920 2539.590 1011.060 ;
        RECT 2041.550 1010.860 2041.870 1010.920 ;
        RECT 2539.270 1010.860 2539.590 1010.920 ;
        RECT 1307.850 1010.720 1308.170 1010.780 ;
        RECT 995.510 1010.580 1282.780 1010.720 ;
        RECT 1288.850 1010.580 1308.170 1010.720 ;
        RECT 995.510 1010.520 995.830 1010.580 ;
        RECT 983.550 1010.380 983.870 1010.440 ;
        RECT 1138.570 1010.380 1138.890 1010.440 ;
        RECT 983.550 1010.240 1138.890 1010.380 ;
        RECT 983.550 1010.180 983.870 1010.240 ;
        RECT 1138.570 1010.180 1138.890 1010.240 ;
        RECT 1145.470 1010.380 1145.790 1010.440 ;
        RECT 1196.530 1010.380 1196.850 1010.440 ;
        RECT 1145.470 1010.240 1196.850 1010.380 ;
        RECT 1145.470 1010.180 1145.790 1010.240 ;
        RECT 1196.530 1010.180 1196.850 1010.240 ;
        RECT 1196.990 1010.380 1197.310 1010.440 ;
        RECT 1200.210 1010.380 1200.530 1010.440 ;
        RECT 1196.990 1010.240 1200.530 1010.380 ;
        RECT 1196.990 1010.180 1197.310 1010.240 ;
        RECT 1200.210 1010.180 1200.530 1010.240 ;
        RECT 1221.370 1010.380 1221.690 1010.440 ;
        RECT 1224.130 1010.380 1224.450 1010.440 ;
        RECT 1221.370 1010.240 1224.450 1010.380 ;
        RECT 1221.370 1010.180 1221.690 1010.240 ;
        RECT 1224.130 1010.180 1224.450 1010.240 ;
        RECT 976.650 1010.040 976.970 1010.100 ;
        RECT 1133.050 1010.040 1133.370 1010.100 ;
        RECT 976.650 1009.900 1133.370 1010.040 ;
        RECT 976.650 1009.840 976.970 1009.900 ;
        RECT 1133.050 1009.840 1133.370 1009.900 ;
        RECT 1145.930 1010.040 1146.250 1010.100 ;
        RECT 1179.510 1010.040 1179.830 1010.100 ;
        RECT 1145.930 1009.900 1179.830 1010.040 ;
        RECT 1145.930 1009.840 1146.250 1009.900 ;
        RECT 1179.510 1009.840 1179.830 1009.900 ;
        RECT 1179.970 1010.040 1180.290 1010.100 ;
        RECT 1230.570 1010.040 1230.890 1010.100 ;
        RECT 1179.970 1009.900 1230.890 1010.040 ;
        RECT 1282.640 1010.040 1282.780 1010.580 ;
        RECT 1307.850 1010.520 1308.170 1010.580 ;
        RECT 1328.090 1010.720 1328.410 1010.780 ;
        RECT 1347.410 1010.720 1347.730 1010.780 ;
        RECT 1328.090 1010.580 1347.730 1010.720 ;
        RECT 1328.090 1010.520 1328.410 1010.580 ;
        RECT 1347.410 1010.520 1347.730 1010.580 ;
        RECT 1376.850 1010.720 1377.170 1010.780 ;
        RECT 1379.610 1010.720 1379.930 1010.780 ;
        RECT 1376.850 1010.580 1379.930 1010.720 ;
        RECT 1376.850 1010.520 1377.170 1010.580 ;
        RECT 1379.610 1010.520 1379.930 1010.580 ;
        RECT 1409.050 1010.720 1409.370 1010.780 ;
        RECT 1413.650 1010.720 1413.970 1010.780 ;
        RECT 1409.050 1010.580 1413.970 1010.720 ;
        RECT 1409.050 1010.520 1409.370 1010.580 ;
        RECT 1413.650 1010.520 1413.970 1010.580 ;
        RECT 1415.950 1010.720 1416.270 1010.780 ;
        RECT 1679.990 1010.720 1680.310 1010.780 ;
        RECT 1415.950 1010.580 1680.310 1010.720 ;
        RECT 1415.950 1010.520 1416.270 1010.580 ;
        RECT 1679.990 1010.520 1680.310 1010.580 ;
        RECT 1737.950 1010.720 1738.270 1010.780 ;
        RECT 1794.070 1010.720 1794.390 1010.780 ;
        RECT 1737.950 1010.580 1794.390 1010.720 ;
        RECT 1737.950 1010.520 1738.270 1010.580 ;
        RECT 1794.070 1010.520 1794.390 1010.580 ;
        RECT 1794.990 1010.720 1795.310 1010.780 ;
        RECT 1800.510 1010.720 1800.830 1010.780 ;
        RECT 1794.990 1010.580 1800.830 1010.720 ;
        RECT 1794.990 1010.520 1795.310 1010.580 ;
        RECT 1800.510 1010.520 1800.830 1010.580 ;
        RECT 1823.510 1010.720 1823.830 1010.780 ;
        RECT 1828.110 1010.720 1828.430 1010.780 ;
        RECT 1823.510 1010.580 1828.430 1010.720 ;
        RECT 1823.510 1010.520 1823.830 1010.580 ;
        RECT 1828.110 1010.520 1828.430 1010.580 ;
        RECT 1867.670 1010.720 1867.990 1010.780 ;
        RECT 1869.510 1010.720 1869.830 1010.780 ;
        RECT 1867.670 1010.580 1869.830 1010.720 ;
        RECT 1867.670 1010.520 1867.990 1010.580 ;
        RECT 1869.510 1010.520 1869.830 1010.580 ;
        RECT 1879.630 1010.720 1879.950 1010.780 ;
        RECT 2528.690 1010.720 2529.010 1010.780 ;
        RECT 1879.630 1010.580 2529.010 1010.720 ;
        RECT 1879.630 1010.520 1879.950 1010.580 ;
        RECT 2528.690 1010.520 2529.010 1010.580 ;
        RECT 1283.010 1010.380 1283.330 1010.440 ;
        RECT 1352.470 1010.380 1352.790 1010.440 ;
        RECT 1283.010 1010.240 1352.790 1010.380 ;
        RECT 1283.010 1010.180 1283.330 1010.240 ;
        RECT 1352.470 1010.180 1352.790 1010.240 ;
        RECT 1504.270 1010.380 1504.590 1010.440 ;
        RECT 1507.950 1010.380 1508.270 1010.440 ;
        RECT 1512.550 1010.380 1512.870 1010.440 ;
        RECT 1582.470 1010.380 1582.790 1010.440 ;
        RECT 1586.610 1010.380 1586.930 1010.440 ;
        RECT 1504.270 1010.240 1508.270 1010.380 ;
        RECT 1504.270 1010.180 1504.590 1010.240 ;
        RECT 1507.950 1010.180 1508.270 1010.240 ;
        RECT 1508.500 1010.240 1512.870 1010.380 ;
        RECT 1311.070 1010.040 1311.390 1010.100 ;
        RECT 1282.640 1009.900 1311.390 1010.040 ;
        RECT 1179.970 1009.840 1180.290 1009.900 ;
        RECT 1230.570 1009.840 1230.890 1009.900 ;
        RECT 1311.070 1009.840 1311.390 1009.900 ;
        RECT 1311.530 1010.040 1311.850 1010.100 ;
        RECT 1341.890 1010.040 1342.210 1010.100 ;
        RECT 1311.530 1009.900 1342.210 1010.040 ;
        RECT 1311.530 1009.840 1311.850 1009.900 ;
        RECT 1341.890 1009.840 1342.210 1009.900 ;
        RECT 1374.550 1010.040 1374.870 1010.100 ;
        RECT 1397.090 1010.040 1397.410 1010.100 ;
        RECT 1374.550 1009.900 1397.410 1010.040 ;
        RECT 1374.550 1009.840 1374.870 1009.900 ;
        RECT 1397.090 1009.840 1397.410 1009.900 ;
        RECT 1402.610 1010.040 1402.930 1010.100 ;
        RECT 1407.210 1010.040 1407.530 1010.100 ;
        RECT 1402.610 1009.900 1407.530 1010.040 ;
        RECT 1402.610 1009.840 1402.930 1009.900 ;
        RECT 1407.210 1009.840 1407.530 1009.900 ;
        RECT 1493.230 1010.040 1493.550 1010.100 ;
        RECT 1508.500 1010.040 1508.640 1010.240 ;
        RECT 1512.550 1010.180 1512.870 1010.240 ;
        RECT 1513.100 1010.240 1579.940 1010.380 ;
        RECT 1493.230 1009.900 1508.640 1010.040 ;
        RECT 1508.870 1010.040 1509.190 1010.100 ;
        RECT 1513.100 1010.040 1513.240 1010.240 ;
        RECT 1508.870 1009.900 1513.240 1010.040 ;
        RECT 1534.630 1010.040 1534.950 1010.100 ;
        RECT 1573.270 1010.040 1573.590 1010.100 ;
        RECT 1534.630 1009.900 1573.590 1010.040 ;
        RECT 1579.800 1010.040 1579.940 1010.240 ;
        RECT 1582.470 1010.240 1586.930 1010.380 ;
        RECT 1582.470 1010.180 1582.790 1010.240 ;
        RECT 1586.610 1010.180 1586.930 1010.240 ;
        RECT 1591.210 1010.380 1591.530 1010.440 ;
        RECT 1593.510 1010.380 1593.830 1010.440 ;
        RECT 1591.210 1010.240 1593.830 1010.380 ;
        RECT 1591.210 1010.180 1591.530 1010.240 ;
        RECT 1593.510 1010.180 1593.830 1010.240 ;
        RECT 1599.030 1010.380 1599.350 1010.440 ;
        RECT 1600.410 1010.380 1600.730 1010.440 ;
        RECT 1599.030 1010.240 1600.730 1010.380 ;
        RECT 1599.030 1010.180 1599.350 1010.240 ;
        RECT 1600.410 1010.180 1600.730 1010.240 ;
        RECT 1660.670 1010.380 1660.990 1010.440 ;
        RECT 1669.870 1010.380 1670.190 1010.440 ;
        RECT 1660.670 1010.240 1670.190 1010.380 ;
        RECT 1660.670 1010.180 1660.990 1010.240 ;
        RECT 1669.870 1010.180 1670.190 1010.240 ;
        RECT 1755.890 1010.380 1756.210 1010.440 ;
        RECT 2086.630 1010.380 2086.950 1010.440 ;
        RECT 1755.890 1010.240 2086.950 1010.380 ;
        RECT 1755.890 1010.180 1756.210 1010.240 ;
        RECT 2086.630 1010.180 2086.950 1010.240 ;
        RECT 1593.050 1010.040 1593.370 1010.100 ;
        RECT 1645.490 1010.040 1645.810 1010.100 ;
        RECT 1579.800 1009.900 1583.620 1010.040 ;
        RECT 1493.230 1009.840 1493.550 1009.900 ;
        RECT 1508.870 1009.840 1509.190 1009.900 ;
        RECT 1534.630 1009.840 1534.950 1009.900 ;
        RECT 1573.270 1009.840 1573.590 1009.900 ;
        RECT 978.030 1009.700 978.350 1009.760 ;
        RECT 1057.150 1009.700 1057.470 1009.760 ;
        RECT 978.030 1009.560 1057.470 1009.700 ;
        RECT 978.030 1009.500 978.350 1009.560 ;
        RECT 1057.150 1009.500 1057.470 1009.560 ;
        RECT 1062.210 1009.700 1062.530 1009.760 ;
        RECT 1191.470 1009.700 1191.790 1009.760 ;
        RECT 1062.210 1009.560 1191.790 1009.700 ;
        RECT 1062.210 1009.500 1062.530 1009.560 ;
        RECT 1191.470 1009.500 1191.790 1009.560 ;
        RECT 1200.210 1009.700 1200.530 1009.760 ;
        RECT 1217.690 1009.700 1218.010 1009.760 ;
        RECT 1200.210 1009.560 1218.010 1009.700 ;
        RECT 1200.210 1009.500 1200.530 1009.560 ;
        RECT 1217.690 1009.500 1218.010 1009.560 ;
        RECT 1267.830 1009.700 1268.150 1009.760 ;
        RECT 1293.590 1009.700 1293.910 1009.760 ;
        RECT 1267.830 1009.560 1293.910 1009.700 ;
        RECT 1267.830 1009.500 1268.150 1009.560 ;
        RECT 1293.590 1009.500 1293.910 1009.560 ;
        RECT 1307.390 1009.700 1307.710 1009.760 ;
        RECT 1310.610 1009.700 1310.930 1009.760 ;
        RECT 1334.530 1009.700 1334.850 1009.760 ;
        RECT 1307.390 1009.560 1310.930 1009.700 ;
        RECT 1307.390 1009.500 1307.710 1009.560 ;
        RECT 1310.610 1009.500 1310.930 1009.560 ;
        RECT 1311.160 1009.560 1334.850 1009.700 ;
        RECT 984.930 1009.360 985.250 1009.420 ;
        RECT 1012.530 1009.360 1012.850 1009.420 ;
        RECT 1083.370 1009.360 1083.690 1009.420 ;
        RECT 984.930 1009.220 1012.300 1009.360 ;
        RECT 984.930 1009.160 985.250 1009.220 ;
        RECT 991.830 1009.020 992.150 1009.080 ;
        RECT 1011.610 1009.020 1011.930 1009.080 ;
        RECT 991.830 1008.880 1011.930 1009.020 ;
        RECT 1012.160 1009.020 1012.300 1009.220 ;
        RECT 1012.530 1009.220 1083.690 1009.360 ;
        RECT 1012.530 1009.160 1012.850 1009.220 ;
        RECT 1083.370 1009.160 1083.690 1009.220 ;
        RECT 1089.810 1009.360 1090.130 1009.420 ;
        RECT 1228.730 1009.360 1229.050 1009.420 ;
        RECT 1089.810 1009.220 1229.050 1009.360 ;
        RECT 1089.810 1009.160 1090.130 1009.220 ;
        RECT 1228.730 1009.160 1229.050 1009.220 ;
        RECT 1272.890 1009.360 1273.210 1009.420 ;
        RECT 1304.630 1009.360 1304.950 1009.420 ;
        RECT 1272.890 1009.220 1304.950 1009.360 ;
        RECT 1272.890 1009.160 1273.210 1009.220 ;
        RECT 1304.630 1009.160 1304.950 1009.220 ;
        RECT 1310.150 1009.360 1310.470 1009.420 ;
        RECT 1311.160 1009.360 1311.300 1009.560 ;
        RECT 1334.530 1009.500 1334.850 1009.560 ;
        RECT 1487.250 1009.700 1487.570 1009.760 ;
        RECT 1493.690 1009.700 1494.010 1009.760 ;
        RECT 1487.250 1009.560 1494.010 1009.700 ;
        RECT 1487.250 1009.500 1487.570 1009.560 ;
        RECT 1493.690 1009.500 1494.010 1009.560 ;
        RECT 1502.430 1009.700 1502.750 1009.760 ;
        RECT 1582.930 1009.700 1583.250 1009.760 ;
        RECT 1502.430 1009.560 1583.250 1009.700 ;
        RECT 1583.480 1009.700 1583.620 1009.900 ;
        RECT 1593.050 1009.900 1645.810 1010.040 ;
        RECT 1593.050 1009.840 1593.370 1009.900 ;
        RECT 1645.490 1009.840 1645.810 1009.900 ;
        RECT 1712.650 1010.040 1712.970 1010.100 ;
        RECT 1717.250 1010.040 1717.570 1010.100 ;
        RECT 1712.650 1009.900 1717.570 1010.040 ;
        RECT 1712.650 1009.840 1712.970 1009.900 ;
        RECT 1717.250 1009.840 1717.570 1009.900 ;
        RECT 1734.270 1010.040 1734.590 1010.100 ;
        RECT 1738.410 1010.040 1738.730 1010.100 ;
        RECT 1734.270 1009.900 1738.730 1010.040 ;
        RECT 1734.270 1009.840 1734.590 1009.900 ;
        RECT 1738.410 1009.840 1738.730 1009.900 ;
        RECT 1786.250 1010.040 1786.570 1010.100 ;
        RECT 2084.790 1010.040 2085.110 1010.100 ;
        RECT 1786.250 1009.900 2085.110 1010.040 ;
        RECT 1786.250 1009.840 1786.570 1009.900 ;
        RECT 2084.790 1009.840 2085.110 1009.900 ;
        RECT 1600.870 1009.700 1601.190 1009.760 ;
        RECT 1583.480 1009.560 1601.190 1009.700 ;
        RECT 1502.430 1009.500 1502.750 1009.560 ;
        RECT 1582.930 1009.500 1583.250 1009.560 ;
        RECT 1600.870 1009.500 1601.190 1009.560 ;
        RECT 1831.790 1009.700 1832.110 1009.760 ;
        RECT 1831.790 1009.560 2042.700 1009.700 ;
        RECT 1831.790 1009.500 1832.110 1009.560 ;
        RECT 1342.350 1009.360 1342.670 1009.420 ;
        RECT 1310.150 1009.220 1311.300 1009.360 ;
        RECT 1311.620 1009.220 1342.670 1009.360 ;
        RECT 1310.150 1009.160 1310.470 1009.220 ;
        RECT 1113.730 1009.020 1114.050 1009.080 ;
        RECT 1012.160 1008.880 1114.050 1009.020 ;
        RECT 991.830 1008.820 992.150 1008.880 ;
        RECT 1011.610 1008.820 1011.930 1008.880 ;
        RECT 1113.730 1008.820 1114.050 1008.880 ;
        RECT 1196.070 1009.020 1196.390 1009.080 ;
        RECT 1237.010 1009.020 1237.330 1009.080 ;
        RECT 1196.070 1008.880 1237.330 1009.020 ;
        RECT 1196.070 1008.820 1196.390 1008.880 ;
        RECT 1237.010 1008.820 1237.330 1008.880 ;
        RECT 1278.410 1009.020 1278.730 1009.080 ;
        RECT 1311.620 1009.020 1311.760 1009.220 ;
        RECT 1342.350 1009.160 1342.670 1009.220 ;
        RECT 1496.450 1009.360 1496.770 1009.420 ;
        RECT 1508.870 1009.360 1509.190 1009.420 ;
        RECT 1496.450 1009.220 1509.190 1009.360 ;
        RECT 1496.450 1009.160 1496.770 1009.220 ;
        RECT 1508.870 1009.160 1509.190 1009.220 ;
        RECT 1509.330 1009.360 1509.650 1009.420 ;
        RECT 1530.950 1009.360 1531.270 1009.420 ;
        RECT 1509.330 1009.220 1531.270 1009.360 ;
        RECT 1509.330 1009.160 1509.650 1009.220 ;
        RECT 1530.950 1009.160 1531.270 1009.220 ;
        RECT 1531.410 1009.360 1531.730 1009.420 ;
        RECT 1535.090 1009.360 1535.410 1009.420 ;
        RECT 1566.370 1009.360 1566.690 1009.420 ;
        RECT 1531.410 1009.220 1535.410 1009.360 ;
        RECT 1531.410 1009.160 1531.730 1009.220 ;
        RECT 1535.090 1009.160 1535.410 1009.220 ;
        RECT 1535.640 1009.220 1566.690 1009.360 ;
        RECT 1278.410 1008.880 1311.760 1009.020 ;
        RECT 1497.370 1009.020 1497.690 1009.080 ;
        RECT 1535.640 1009.020 1535.780 1009.220 ;
        RECT 1566.370 1009.160 1566.690 1009.220 ;
        RECT 1873.190 1009.360 1873.510 1009.420 ;
        RECT 1900.330 1009.360 1900.650 1009.420 ;
        RECT 1873.190 1009.220 1900.650 1009.360 ;
        RECT 1873.190 1009.160 1873.510 1009.220 ;
        RECT 1900.330 1009.160 1900.650 1009.220 ;
        RECT 2037.870 1009.360 2038.190 1009.420 ;
        RECT 2042.010 1009.360 2042.330 1009.420 ;
        RECT 2037.870 1009.220 2042.330 1009.360 ;
        RECT 2037.870 1009.160 2038.190 1009.220 ;
        RECT 2042.010 1009.160 2042.330 1009.220 ;
        RECT 1497.370 1008.880 1535.780 1009.020 ;
        RECT 1548.890 1009.020 1549.210 1009.080 ;
        RECT 1605.930 1009.020 1606.250 1009.080 ;
        RECT 1548.890 1008.880 1606.250 1009.020 ;
        RECT 2042.560 1009.020 2042.700 1009.560 ;
        RECT 2065.930 1009.360 2066.250 1009.420 ;
        RECT 2069.610 1009.360 2069.930 1009.420 ;
        RECT 2065.930 1009.220 2069.930 1009.360 ;
        RECT 2065.930 1009.160 2066.250 1009.220 ;
        RECT 2069.610 1009.160 2069.930 1009.220 ;
        RECT 2079.270 1009.360 2079.590 1009.420 ;
        RECT 2083.410 1009.360 2083.730 1009.420 ;
        RECT 2079.270 1009.220 2083.730 1009.360 ;
        RECT 2079.270 1009.160 2079.590 1009.220 ;
        RECT 2083.410 1009.160 2083.730 1009.220 ;
        RECT 2093.990 1009.020 2094.310 1009.080 ;
        RECT 2042.560 1008.880 2094.310 1009.020 ;
        RECT 1278.410 1008.820 1278.730 1008.880 ;
        RECT 1497.370 1008.820 1497.690 1008.880 ;
        RECT 1548.890 1008.820 1549.210 1008.880 ;
        RECT 1605.930 1008.820 1606.250 1008.880 ;
        RECT 2093.990 1008.820 2094.310 1008.880 ;
        RECT 1003.790 1008.680 1004.110 1008.740 ;
        RECT 1092.110 1008.680 1092.430 1008.740 ;
        RECT 1003.790 1008.540 1092.430 1008.680 ;
        RECT 1003.790 1008.480 1004.110 1008.540 ;
        RECT 1092.110 1008.480 1092.430 1008.540 ;
        RECT 1093.030 1008.680 1093.350 1008.740 ;
        RECT 1145.010 1008.680 1145.330 1008.740 ;
        RECT 1093.030 1008.540 1145.330 1008.680 ;
        RECT 1093.030 1008.480 1093.350 1008.540 ;
        RECT 1145.010 1008.480 1145.330 1008.540 ;
        RECT 1197.450 1008.680 1197.770 1008.740 ;
        RECT 1245.290 1008.680 1245.610 1008.740 ;
        RECT 1197.450 1008.540 1245.610 1008.680 ;
        RECT 1197.450 1008.480 1197.770 1008.540 ;
        RECT 1245.290 1008.480 1245.610 1008.540 ;
        RECT 1264.150 1008.680 1264.470 1008.740 ;
        RECT 1268.750 1008.680 1269.070 1008.740 ;
        RECT 1264.150 1008.540 1269.070 1008.680 ;
        RECT 1264.150 1008.480 1264.470 1008.540 ;
        RECT 1268.750 1008.480 1269.070 1008.540 ;
        RECT 1274.730 1008.680 1275.050 1008.740 ;
        RECT 1311.530 1008.680 1311.850 1008.740 ;
        RECT 1339.590 1008.680 1339.910 1008.740 ;
        RECT 1274.730 1008.540 1311.850 1008.680 ;
        RECT 1274.730 1008.480 1275.050 1008.540 ;
        RECT 1311.530 1008.480 1311.850 1008.540 ;
        RECT 1315.760 1008.540 1339.910 1008.680 ;
        RECT 998.730 1008.340 999.050 1008.400 ;
        RECT 1097.170 1008.340 1097.490 1008.400 ;
        RECT 998.730 1008.200 1097.490 1008.340 ;
        RECT 998.730 1008.140 999.050 1008.200 ;
        RECT 1097.170 1008.140 1097.490 1008.200 ;
        RECT 1179.510 1008.340 1179.830 1008.400 ;
        RECT 1204.810 1008.340 1205.130 1008.400 ;
        RECT 1179.510 1008.200 1205.130 1008.340 ;
        RECT 1179.510 1008.140 1179.830 1008.200 ;
        RECT 1204.810 1008.140 1205.130 1008.200 ;
        RECT 1261.850 1008.340 1262.170 1008.400 ;
        RECT 1315.210 1008.340 1315.530 1008.400 ;
        RECT 1261.850 1008.200 1315.530 1008.340 ;
        RECT 1261.850 1008.140 1262.170 1008.200 ;
        RECT 1315.210 1008.140 1315.530 1008.200 ;
        RECT 638.090 1008.000 638.410 1008.060 ;
        RECT 669.830 1008.000 670.150 1008.060 ;
        RECT 638.090 1007.860 670.150 1008.000 ;
        RECT 638.090 1007.800 638.410 1007.860 ;
        RECT 669.830 1007.800 670.150 1007.860 ;
        RECT 994.590 1008.000 994.910 1008.060 ;
        RECT 1078.770 1008.000 1079.090 1008.060 ;
        RECT 994.590 1007.860 1079.090 1008.000 ;
        RECT 994.590 1007.800 994.910 1007.860 ;
        RECT 1078.770 1007.800 1079.090 1007.860 ;
        RECT 1209.870 1008.000 1210.190 1008.060 ;
        RECT 1214.010 1008.000 1214.330 1008.060 ;
        RECT 1209.870 1007.860 1214.330 1008.000 ;
        RECT 1209.870 1007.800 1210.190 1007.860 ;
        RECT 1214.010 1007.800 1214.330 1007.860 ;
        RECT 1222.750 1008.000 1223.070 1008.060 ;
        RECT 1315.760 1008.000 1315.900 1008.540 ;
        RECT 1339.590 1008.480 1339.910 1008.540 ;
        RECT 1368.110 1008.680 1368.430 1008.740 ;
        RECT 1372.710 1008.680 1373.030 1008.740 ;
        RECT 1368.110 1008.540 1373.030 1008.680 ;
        RECT 1368.110 1008.480 1368.430 1008.540 ;
        RECT 1372.710 1008.480 1373.030 1008.540 ;
        RECT 1383.290 1008.680 1383.610 1008.740 ;
        RECT 1386.510 1008.680 1386.830 1008.740 ;
        RECT 1383.290 1008.540 1386.830 1008.680 ;
        RECT 1383.290 1008.480 1383.610 1008.540 ;
        RECT 1386.510 1008.480 1386.830 1008.540 ;
        RECT 1489.090 1008.680 1489.410 1008.740 ;
        RECT 1534.630 1008.680 1534.950 1008.740 ;
        RECT 1489.090 1008.540 1534.950 1008.680 ;
        RECT 1489.090 1008.480 1489.410 1008.540 ;
        RECT 1534.630 1008.480 1534.950 1008.540 ;
        RECT 1552.570 1008.680 1552.890 1008.740 ;
        RECT 1554.410 1008.680 1554.730 1008.740 ;
        RECT 1552.570 1008.540 1554.730 1008.680 ;
        RECT 1552.570 1008.480 1552.890 1008.540 ;
        RECT 1554.410 1008.480 1554.730 1008.540 ;
        RECT 1769.230 1008.680 1769.550 1008.740 ;
        RECT 1772.450 1008.680 1772.770 1008.740 ;
        RECT 1769.230 1008.540 1772.770 1008.680 ;
        RECT 1769.230 1008.480 1769.550 1008.540 ;
        RECT 1772.450 1008.480 1772.770 1008.540 ;
        RECT 1782.110 1008.680 1782.430 1008.740 ;
        RECT 1786.710 1008.680 1787.030 1008.740 ;
        RECT 1782.110 1008.540 1787.030 1008.680 ;
        RECT 1782.110 1008.480 1782.430 1008.540 ;
        RECT 1786.710 1008.480 1787.030 1008.540 ;
        RECT 1330.390 1008.340 1330.710 1008.400 ;
        RECT 1343.270 1008.340 1343.590 1008.400 ;
        RECT 1330.390 1008.200 1343.590 1008.340 ;
        RECT 1330.390 1008.140 1330.710 1008.200 ;
        RECT 1343.270 1008.140 1343.590 1008.200 ;
        RECT 1495.990 1008.340 1496.310 1008.400 ;
        RECT 1555.790 1008.340 1556.110 1008.400 ;
        RECT 1495.990 1008.200 1556.110 1008.340 ;
        RECT 1495.990 1008.140 1496.310 1008.200 ;
        RECT 1555.790 1008.140 1556.110 1008.200 ;
        RECT 1222.750 1007.860 1315.900 1008.000 ;
        RECT 1450.450 1008.000 1450.770 1008.060 ;
        RECT 1455.050 1008.000 1455.370 1008.060 ;
        RECT 1450.450 1007.860 1455.370 1008.000 ;
        RECT 1222.750 1007.800 1223.070 1007.860 ;
        RECT 1450.450 1007.800 1450.770 1007.860 ;
        RECT 1455.050 1007.800 1455.370 1007.860 ;
        RECT 1461.030 1008.000 1461.350 1008.060 ;
        RECT 1462.410 1008.000 1462.730 1008.060 ;
        RECT 1461.030 1007.860 1462.730 1008.000 ;
        RECT 1461.030 1007.800 1461.350 1007.860 ;
        RECT 1462.410 1007.800 1462.730 1007.860 ;
        RECT 1488.170 1008.000 1488.490 1008.060 ;
        RECT 1518.070 1008.000 1518.390 1008.060 ;
        RECT 1488.170 1007.860 1518.390 1008.000 ;
        RECT 1488.170 1007.800 1488.490 1007.860 ;
        RECT 1518.070 1007.800 1518.390 1007.860 ;
        RECT 650.510 1007.660 650.830 1007.720 ;
        RECT 671.670 1007.660 671.990 1007.720 ;
        RECT 650.510 1007.520 671.990 1007.660 ;
        RECT 650.510 1007.460 650.830 1007.520 ;
        RECT 671.670 1007.460 671.990 1007.520 ;
        RECT 992.290 1007.660 992.610 1007.720 ;
        RECT 1053.010 1007.660 1053.330 1007.720 ;
        RECT 992.290 1007.520 1053.330 1007.660 ;
        RECT 992.290 1007.460 992.610 1007.520 ;
        RECT 1053.010 1007.460 1053.330 1007.520 ;
        RECT 1053.470 1007.660 1053.790 1007.720 ;
        RECT 1100.390 1007.660 1100.710 1007.720 ;
        RECT 1053.470 1007.520 1100.710 1007.660 ;
        RECT 1053.470 1007.460 1053.790 1007.520 ;
        RECT 1100.390 1007.460 1100.710 1007.520 ;
        RECT 1191.470 1007.660 1191.790 1007.720 ;
        RECT 1210.330 1007.660 1210.650 1007.720 ;
        RECT 1191.470 1007.520 1210.650 1007.660 ;
        RECT 1191.470 1007.460 1191.790 1007.520 ;
        RECT 1210.330 1007.460 1210.650 1007.520 ;
        RECT 1293.590 1007.660 1293.910 1007.720 ;
        RECT 1333.610 1007.660 1333.930 1007.720 ;
        RECT 1293.590 1007.520 1333.930 1007.660 ;
        RECT 1293.590 1007.460 1293.910 1007.520 ;
        RECT 1333.610 1007.460 1333.930 1007.520 ;
        RECT 1334.990 1007.660 1335.310 1007.720 ;
        RECT 1340.510 1007.660 1340.830 1007.720 ;
        RECT 1334.990 1007.520 1340.830 1007.660 ;
        RECT 1334.990 1007.460 1335.310 1007.520 ;
        RECT 1340.510 1007.460 1340.830 1007.520 ;
        RECT 1417.790 1007.660 1418.110 1007.720 ;
        RECT 1421.010 1007.660 1421.330 1007.720 ;
        RECT 1417.790 1007.520 1421.330 1007.660 ;
        RECT 1417.790 1007.460 1418.110 1007.520 ;
        RECT 1421.010 1007.460 1421.330 1007.520 ;
        RECT 1437.570 1007.660 1437.890 1007.720 ;
        RECT 1441.710 1007.660 1442.030 1007.720 ;
        RECT 1437.570 1007.520 1442.030 1007.660 ;
        RECT 1437.570 1007.460 1437.890 1007.520 ;
        RECT 1441.710 1007.460 1442.030 1007.520 ;
        RECT 1446.310 1007.660 1446.630 1007.720 ;
        RECT 1448.610 1007.660 1448.930 1007.720 ;
        RECT 1446.310 1007.520 1448.930 1007.660 ;
        RECT 1446.310 1007.460 1446.630 1007.520 ;
        RECT 1448.610 1007.460 1448.930 1007.520 ;
        RECT 1452.750 1007.660 1453.070 1007.720 ;
        RECT 1455.510 1007.660 1455.830 1007.720 ;
        RECT 1452.750 1007.520 1455.830 1007.660 ;
        RECT 1452.750 1007.460 1453.070 1007.520 ;
        RECT 1455.510 1007.460 1455.830 1007.520 ;
        RECT 1459.190 1007.660 1459.510 1007.720 ;
        RECT 1461.950 1007.660 1462.270 1007.720 ;
        RECT 1459.190 1007.520 1462.270 1007.660 ;
        RECT 1459.190 1007.460 1459.510 1007.520 ;
        RECT 1461.950 1007.460 1462.270 1007.520 ;
        RECT 1511.630 1007.660 1511.950 1007.720 ;
        RECT 1545.670 1007.660 1545.990 1007.720 ;
        RECT 1511.630 1007.520 1545.990 1007.660 ;
        RECT 1511.630 1007.460 1511.950 1007.520 ;
        RECT 1545.670 1007.460 1545.990 1007.520 ;
        RECT 1610.990 1007.660 1611.310 1007.720 ;
        RECT 1614.210 1007.660 1614.530 1007.720 ;
        RECT 1610.990 1007.520 1614.530 1007.660 ;
        RECT 1610.990 1007.460 1611.310 1007.520 ;
        RECT 1614.210 1007.460 1614.530 1007.520 ;
        RECT 1617.430 1007.660 1617.750 1007.720 ;
        RECT 1635.370 1007.660 1635.690 1007.720 ;
        RECT 1617.430 1007.520 1635.690 1007.660 ;
        RECT 1617.430 1007.460 1617.750 1007.520 ;
        RECT 1635.370 1007.460 1635.690 1007.520 ;
        RECT 1803.730 1007.660 1804.050 1007.720 ;
        RECT 1806.950 1007.660 1807.270 1007.720 ;
        RECT 1803.730 1007.520 1807.270 1007.660 ;
        RECT 1803.730 1007.460 1804.050 1007.520 ;
        RECT 1806.950 1007.460 1807.270 1007.520 ;
        RECT 910.870 1001.880 911.190 1001.940 ;
        RECT 912.250 1001.880 912.570 1001.940 ;
        RECT 910.870 1001.740 912.570 1001.880 ;
        RECT 910.870 1001.680 911.190 1001.740 ;
        RECT 912.250 1001.680 912.570 1001.740 ;
        RECT 1532.790 1001.200 1533.110 1001.260 ;
        RECT 1535.780 1001.200 1536.100 1001.260 ;
        RECT 1532.790 1001.060 1536.100 1001.200 ;
        RECT 1532.790 1001.000 1533.110 1001.060 ;
        RECT 1535.780 1001.000 1536.100 1001.060 ;
        RECT 1559.470 1001.200 1559.790 1001.260 ;
        RECT 1561.540 1001.200 1561.860 1001.260 ;
        RECT 1559.470 1001.060 1561.860 1001.200 ;
        RECT 1559.470 1001.000 1559.790 1001.060 ;
        RECT 1561.540 1001.000 1561.860 1001.060 ;
        RECT 1815.460 1001.200 1815.780 1001.260 ;
        RECT 1821.210 1001.200 1821.530 1001.260 ;
        RECT 1815.460 1001.060 1821.530 1001.200 ;
        RECT 1815.460 1001.000 1815.780 1001.060 ;
        RECT 1821.210 1001.000 1821.530 1001.060 ;
      LAYER met1 ;
        RECT 670.070 604.460 2164.080 998.440 ;
      LAYER via ;
        RECT 1351.120 2917.580 1351.380 2917.840 ;
        RECT 1535.120 2917.580 1535.380 2917.840 ;
        RECT 1501.540 2917.240 1501.800 2917.500 ;
        RECT 1546.160 2917.240 1546.420 2917.500 ;
        RECT 1414.140 2916.900 1414.400 2917.160 ;
        RECT 1567.320 2916.900 1567.580 2917.160 ;
        RECT 1479.920 2915.540 1480.180 2915.800 ;
        RECT 1641.840 2915.540 1642.100 2915.800 ;
        RECT 1495.560 2915.200 1495.820 2915.460 ;
        RECT 1705.320 2915.200 1705.580 2915.460 ;
        RECT 1379.640 2914.860 1379.900 2915.120 ;
        RECT 1598.600 2914.860 1598.860 2915.120 ;
        RECT 1407.240 2914.520 1407.500 2914.780 ;
        RECT 1630.800 2914.520 1631.060 2914.780 ;
        RECT 1461.520 2914.180 1461.780 2914.440 ;
        RECT 1694.280 2914.180 1694.540 2914.440 ;
        RECT 1494.640 2913.840 1494.900 2914.100 ;
        RECT 1768.800 2913.840 1769.060 2914.100 ;
        RECT 1789.960 2913.840 1790.220 2914.100 ;
        RECT 1895.300 2913.840 1895.560 2914.100 ;
        RECT 1502.000 2913.500 1502.260 2913.760 ;
        RECT 1812.040 2913.500 1812.300 2913.760 ;
        RECT 1372.740 2913.160 1373.000 2913.420 ;
        RECT 1843.320 2913.160 1843.580 2913.420 ;
        RECT 1493.720 2912.820 1493.980 2913.080 ;
        RECT 1801.000 2912.820 1801.260 2913.080 ;
        RECT 1833.200 2912.820 1833.460 2913.080 ;
        RECT 1887.480 2912.820 1887.740 2913.080 ;
        RECT 1496.940 2912.480 1497.200 2912.740 ;
        RECT 1663.000 2912.480 1663.260 2912.740 ;
        RECT 1854.360 2912.480 1854.620 2912.740 ;
        RECT 1886.560 2912.480 1886.820 2912.740 ;
        RECT 1495.100 2912.140 1495.360 2912.400 ;
        RECT 1609.640 2912.140 1609.900 2912.400 ;
        RECT 1351.120 2911.800 1351.380 2912.060 ;
        RECT 1502.460 2911.800 1502.720 2912.060 ;
        RECT 1779.840 2911.800 1780.100 2912.060 ;
        RECT 1864.480 2911.800 1864.740 2912.060 ;
        RECT 1894.840 2911.800 1895.100 2912.060 ;
        RECT 1351.120 2911.120 1351.380 2911.380 ;
        RECT 1455.540 2900.920 1455.800 2901.180 ;
        RECT 1758.680 2900.920 1758.940 2901.180 ;
        RECT 1496.480 2898.200 1496.740 2898.460 ;
        RECT 1524.080 2898.200 1524.340 2898.460 ;
        RECT 1497.400 2896.500 1497.660 2896.760 ;
        RECT 1503.380 2896.500 1503.640 2896.760 ;
        RECT 1876.900 2896.500 1877.160 2896.760 ;
        RECT 1887.940 2896.500 1888.200 2896.760 ;
        RECT 1351.120 2849.920 1351.380 2850.180 ;
        RECT 1358.020 2849.580 1358.280 2849.840 ;
        RECT 1490.040 2849.580 1490.300 2849.840 ;
        RECT 1351.120 2849.240 1351.380 2849.500 ;
        RECT 1350.660 2842.780 1350.920 2843.040 ;
        RECT 1351.120 2842.780 1351.380 2843.040 ;
        RECT 1476.240 2829.180 1476.500 2829.440 ;
        RECT 1490.040 2829.180 1490.300 2829.440 ;
        RECT 1000.600 2810.480 1000.860 2810.740 ;
        RECT 1048.440 2810.480 1048.700 2810.740 ;
        RECT 985.420 2810.140 985.680 2810.400 ;
        RECT 1073.740 2810.140 1074.000 2810.400 ;
        RECT 978.520 2809.800 978.780 2810.060 ;
        RECT 1027.740 2809.800 1028.000 2810.060 ;
        RECT 978.980 2809.460 979.240 2809.720 ;
        RECT 1043.380 2809.460 1043.640 2809.720 ;
        RECT 985.880 2809.120 986.140 2809.380 ;
        RECT 1058.100 2809.120 1058.360 2809.380 ;
        RECT 979.440 2808.780 979.700 2809.040 ;
        RECT 1000.600 2808.780 1000.860 2809.040 ;
        RECT 1048.440 2808.440 1048.700 2808.700 ;
        RECT 1089.380 2808.440 1089.640 2808.700 ;
        RECT 986.340 2800.960 986.600 2801.220 ;
        RECT 1010.260 2800.960 1010.520 2801.220 ;
        RECT 1351.580 2794.840 1351.840 2795.100 ;
        RECT 1352.960 2794.840 1353.220 2795.100 ;
        RECT 445.840 2769.340 446.100 2769.600 ;
        RECT 796.820 2769.340 797.080 2769.600 ;
        RECT 532.320 2767.980 532.580 2768.240 ;
        RECT 707.120 2767.980 707.380 2768.240 ;
        RECT 518.520 2767.640 518.780 2767.900 ;
        RECT 755.420 2767.640 755.680 2767.900 ;
        RECT 489.080 2767.300 489.340 2767.560 ;
        RECT 769.220 2767.300 769.480 2767.560 ;
        RECT 588.900 2684.000 589.160 2684.260 ;
        RECT 720.920 2684.000 721.180 2684.260 ;
        RECT 588.900 2663.600 589.160 2663.860 ;
        RECT 789.920 2663.600 790.180 2663.860 ;
        RECT 978.060 2643.880 978.320 2644.140 ;
        RECT 987.260 2643.880 987.520 2644.140 ;
        RECT 1358.480 2780.900 1358.740 2781.160 ;
        RECT 1485.440 2780.900 1485.700 2781.160 ;
        RECT 1351.580 2767.300 1351.840 2767.560 ;
        RECT 1351.120 2766.620 1351.380 2766.880 ;
        RECT 1350.660 2739.080 1350.920 2739.340 ;
        RECT 1351.120 2739.080 1351.380 2739.340 ;
        RECT 1350.200 2691.140 1350.460 2691.400 ;
        RECT 1350.660 2691.140 1350.920 2691.400 ;
        RECT 1434.380 2691.140 1434.640 2691.400 ;
        RECT 1489.120 2691.140 1489.380 2691.400 ;
        RECT 1350.200 2670.060 1350.460 2670.320 ;
        RECT 1351.120 2670.060 1351.380 2670.320 ;
        RECT 1351.120 2622.460 1351.380 2622.720 ;
        RECT 1351.120 2621.780 1351.380 2622.040 ;
        RECT 1393.440 2608.180 1393.700 2608.440 ;
        RECT 1488.660 2608.180 1488.920 2608.440 ;
        RECT 999.220 2605.460 999.480 2605.720 ;
        RECT 1111.920 2605.460 1112.180 2605.720 ;
        RECT 999.680 2605.120 999.940 2605.380 ;
        RECT 1112.840 2605.120 1113.100 2605.380 ;
        RECT 982.200 2604.780 982.460 2605.040 ;
        RECT 1113.300 2604.780 1113.560 2605.040 ;
        RECT 975.300 2604.440 975.560 2604.700 ;
        RECT 1112.380 2604.440 1112.640 2604.700 ;
        RECT 1392.980 2594.580 1393.240 2594.840 ;
        RECT 1488.200 2594.580 1488.460 2594.840 ;
        RECT 533.240 2591.520 533.500 2591.780 ;
        RECT 762.320 2591.520 762.580 2591.780 ;
        RECT 984.960 2591.520 985.220 2591.780 ;
        RECT 1048.900 2591.520 1049.160 2591.780 ;
        RECT 504.720 2591.180 504.980 2591.440 ;
        RECT 783.020 2591.180 783.280 2591.440 ;
        RECT 974.840 2591.180 975.100 2591.440 ;
        RECT 1094.900 2591.180 1095.160 2591.440 ;
        RECT 1028.200 2587.440 1028.460 2587.700 ;
        RECT 1033.260 2587.440 1033.520 2587.700 ;
        RECT 1413.680 2580.640 1413.940 2580.900 ;
        RECT 1488.200 2580.640 1488.460 2580.900 ;
        RECT 1468.880 2546.300 1469.140 2546.560 ;
        RECT 1484.520 2546.300 1484.780 2546.560 ;
        RECT 1350.200 2511.620 1350.460 2511.880 ;
        RECT 1352.040 2511.620 1352.300 2511.880 ;
        RECT 2094.020 2781.240 2094.280 2781.500 ;
        RECT 2556.320 2781.240 2556.580 2781.500 ;
        RECT 1893.920 2780.900 1894.180 2781.160 ;
        RECT 2422.000 2780.900 2422.260 2781.160 ;
        RECT 2528.720 2587.440 2528.980 2587.700 ;
        RECT 2534.240 2587.440 2534.500 2587.700 ;
        RECT 1621.140 2495.300 1621.400 2495.560 ;
        RECT 1895.300 2495.300 1895.560 2495.560 ;
        RECT 1495.560 2494.960 1495.820 2495.220 ;
        RECT 1552.600 2494.960 1552.860 2495.220 ;
        RECT 1600.440 2494.960 1600.700 2495.220 ;
        RECT 1887.940 2494.960 1888.200 2495.220 ;
        RECT 1502.000 2494.620 1502.260 2494.880 ;
        RECT 1559.500 2494.620 1559.760 2494.880 ;
        RECT 1586.640 2494.620 1586.900 2494.880 ;
        RECT 1887.480 2494.620 1887.740 2494.880 ;
        RECT 1495.100 2494.280 1495.360 2494.540 ;
        RECT 1514.880 2494.280 1515.140 2494.540 ;
        RECT 1544.320 2494.280 1544.580 2494.540 ;
        RECT 1894.840 2494.280 1895.100 2494.540 ;
        RECT 1494.640 2493.940 1494.900 2494.200 ;
        RECT 1573.760 2493.940 1574.020 2494.200 ;
        RECT 1869.540 2493.940 1869.800 2494.200 ;
        RECT 2394.400 2493.940 2394.660 2494.200 ;
        RECT 1501.540 2491.220 1501.800 2491.480 ;
        RECT 1504.300 2491.220 1504.560 2491.480 ;
        RECT 1679.560 2489.520 1679.820 2489.780 ;
        RECT 1683.240 2489.520 1683.500 2489.780 ;
        RECT 1593.540 2489.180 1593.800 2489.440 ;
        RECT 1778.920 2489.180 1779.180 2489.440 ;
        RECT 1645.520 2488.840 1645.780 2489.100 ;
        RECT 1789.960 2488.840 1790.220 2489.100 ;
        RECT 1421.040 2488.500 1421.300 2488.760 ;
        RECT 1842.400 2488.500 1842.660 2488.760 ;
        RECT 1455.080 2488.160 1455.340 2488.420 ;
        RECT 1885.640 2488.160 1885.900 2488.420 ;
        RECT 1420.580 2487.820 1420.840 2488.080 ;
        RECT 1874.600 2487.820 1874.860 2488.080 ;
        RECT 1448.640 2486.800 1448.900 2487.060 ;
        RECT 1832.280 2486.800 1832.540 2487.060 ;
        RECT 1454.620 2486.460 1454.880 2486.720 ;
        RECT 1757.760 2486.460 1758.020 2486.720 ;
        RECT 1427.940 2486.120 1428.200 2486.380 ;
        RECT 1725.560 2486.120 1725.820 2486.380 ;
        RECT 1528.220 2485.780 1528.480 2486.040 ;
        RECT 1811.120 2485.780 1811.380 2486.040 ;
        RECT 1386.540 2485.440 1386.800 2485.700 ;
        RECT 1587.560 2485.440 1587.820 2485.700 ;
        RECT 1397.120 2485.100 1397.380 2485.360 ;
        RECT 1534.200 2485.100 1534.460 2485.360 ;
        RECT 1572.380 2485.100 1572.640 2485.360 ;
        RECT 1746.720 2485.100 1746.980 2485.360 ;
        RECT 1441.740 2484.760 1442.000 2485.020 ;
        RECT 1608.720 2484.760 1608.980 2485.020 ;
        RECT 1535.120 2484.420 1535.380 2484.680 ;
        RECT 1576.520 2484.420 1576.780 2484.680 ;
        RECT 1545.240 2484.080 1545.500 2484.340 ;
        RECT 1548.920 2484.080 1549.180 2484.340 ;
        RECT 1611.020 2484.080 1611.280 2484.340 ;
        RECT 1619.760 2484.080 1620.020 2484.340 ;
        RECT 1673.120 2484.080 1673.380 2484.340 ;
        RECT 1679.560 2484.080 1679.820 2484.340 ;
        RECT 1680.020 2484.080 1680.280 2484.340 ;
        RECT 1715.440 2484.080 1715.700 2484.340 ;
        RECT 1351.120 2429.340 1351.380 2429.600 ;
        RECT 1532.360 2429.000 1532.620 2429.260 ;
        RECT 1351.120 2428.660 1351.380 2428.920 ;
        RECT 1532.820 2428.320 1533.080 2428.580 ;
        RECT 1544.320 2414.720 1544.580 2414.980 ;
        RECT 1545.240 2414.720 1545.500 2414.980 ;
        RECT 1351.120 2380.380 1351.380 2380.640 ;
        RECT 1351.580 2380.380 1351.840 2380.640 ;
        RECT 1545.240 2380.380 1545.500 2380.640 ;
        RECT 1544.780 2380.040 1545.040 2380.300 ;
        RECT 1351.120 2366.780 1351.380 2367.040 ;
        RECT 1351.580 2366.780 1351.840 2367.040 ;
        RECT 1531.900 2366.780 1532.160 2367.040 ;
        RECT 1533.280 2366.780 1533.540 2367.040 ;
        RECT 1532.360 2359.640 1532.620 2359.900 ;
        RECT 1533.280 2359.640 1533.540 2359.900 ;
        RECT 1351.120 2332.440 1351.380 2332.700 ;
        RECT 1544.320 2332.100 1544.580 2332.360 ;
        RECT 1545.240 2332.100 1545.500 2332.360 ;
        RECT 1351.120 2331.760 1351.380 2332.020 ;
        RECT 1533.280 2318.500 1533.540 2318.760 ;
        RECT 1532.820 2318.160 1533.080 2318.420 ;
        RECT 1543.860 2318.160 1544.120 2318.420 ;
        RECT 1544.320 2318.160 1544.580 2318.420 ;
        RECT 1559.040 2318.160 1559.300 2318.420 ;
        RECT 1559.500 2318.160 1559.760 2318.420 ;
        RECT 1350.200 2294.020 1350.460 2294.280 ;
        RECT 1351.120 2294.020 1351.380 2294.280 ;
        RECT 1543.860 2283.480 1544.120 2283.740 ;
        RECT 1544.780 2283.480 1545.040 2283.740 ;
        RECT 1559.040 2270.220 1559.300 2270.480 ;
        RECT 1559.500 2270.220 1559.760 2270.480 ;
        RECT 1543.860 2269.540 1544.120 2269.800 ;
        RECT 1545.240 2269.540 1545.500 2269.800 ;
        RECT 1531.440 2262.740 1531.700 2263.000 ;
        RECT 1532.360 2262.740 1532.620 2263.000 ;
        RECT 1559.500 2262.740 1559.760 2263.000 ;
        RECT 1560.420 2262.740 1560.680 2263.000 ;
        RECT 1351.120 2235.880 1351.380 2236.140 ;
        RECT 1351.120 2235.200 1351.380 2235.460 ;
        RECT 1531.440 2214.800 1531.700 2215.060 ;
        RECT 1532.820 2214.800 1533.080 2215.060 ;
        RECT 1559.500 2214.800 1559.760 2215.060 ;
        RECT 1560.420 2214.800 1560.680 2215.060 ;
        RECT 1350.200 2197.460 1350.460 2197.720 ;
        RECT 1351.120 2197.460 1351.380 2197.720 ;
        RECT 1532.820 2187.600 1533.080 2187.860 ;
        RECT 1532.360 2186.920 1532.620 2187.180 ;
        RECT 1531.900 2172.980 1532.160 2173.240 ;
        RECT 1532.360 2172.980 1532.620 2173.240 ;
        RECT 1531.440 2166.180 1531.700 2166.440 ;
        RECT 1531.900 2166.180 1532.160 2166.440 ;
        RECT 1559.500 2166.180 1559.760 2166.440 ;
        RECT 1560.420 2166.180 1560.680 2166.440 ;
        RECT 1351.120 2139.320 1351.380 2139.580 ;
        RECT 1351.120 2138.640 1351.380 2138.900 ;
        RECT 1350.660 2125.040 1350.920 2125.300 ;
        RECT 1351.120 2125.040 1351.380 2125.300 ;
        RECT 1531.440 2124.700 1531.700 2124.960 ;
        RECT 1532.820 2124.700 1533.080 2124.960 ;
        RECT 1559.500 2118.240 1559.760 2118.500 ;
        RECT 1560.420 2118.240 1560.680 2118.500 ;
        RECT 1532.820 2111.100 1533.080 2111.360 ;
        RECT 1533.740 2111.100 1534.000 2111.360 ;
        RECT 1350.660 2090.360 1350.920 2090.620 ;
        RECT 1351.580 2090.360 1351.840 2090.620 ;
        RECT 1559.500 2069.620 1559.760 2069.880 ;
        RECT 1560.420 2069.620 1560.680 2069.880 ;
        RECT 1532.360 2063.160 1532.620 2063.420 ;
        RECT 1533.740 2063.160 1534.000 2063.420 ;
        RECT 1244.860 2055.340 1245.120 2055.600 ;
        RECT 1346.060 2055.340 1346.320 2055.600 ;
        RECT 1287.180 2055.000 1287.440 2055.260 ;
        RECT 1346.520 2055.000 1346.780 2055.260 ;
        RECT 1230.140 2054.660 1230.400 2054.920 ;
        RECT 1335.480 2054.660 1335.740 2054.920 ;
        RECT 1116.980 2054.320 1117.240 2054.580 ;
        RECT 1332.720 2054.320 1332.980 2054.580 ;
        RECT 1130.780 2053.980 1131.040 2054.240 ;
        RECT 1352.960 2053.980 1353.220 2054.240 ;
        RECT 1216.340 2053.640 1216.600 2053.900 ;
        RECT 1346.980 2053.640 1347.240 2053.900 ;
        RECT 1059.940 2053.300 1060.200 2053.560 ;
        RECT 1335.020 2053.300 1335.280 2053.560 ;
        RECT 1031.420 2052.960 1031.680 2053.220 ;
        RECT 1353.880 2052.960 1354.140 2053.220 ;
        RECT 1016.700 2052.620 1016.960 2052.880 ;
        RECT 1347.440 2052.620 1347.700 2052.880 ;
        RECT 1350.200 2052.620 1350.460 2052.880 ;
        RECT 1352.040 2052.620 1352.300 2052.880 ;
        RECT 1201.620 2052.280 1201.880 2052.540 ;
        RECT 1333.180 2052.280 1333.440 2052.540 ;
        RECT 1187.820 2051.940 1188.080 2052.200 ;
        RECT 1335.940 2051.940 1336.200 2052.200 ;
        RECT 1173.100 2051.600 1173.360 2051.860 ;
        RECT 1345.600 2051.600 1345.860 2051.860 ;
        RECT 1159.300 2051.260 1159.560 2051.520 ;
        RECT 1352.500 2051.260 1352.760 2051.520 ;
        RECT 1144.580 2050.920 1144.840 2051.180 ;
        RECT 1353.420 2050.920 1353.680 2051.180 ;
        RECT 977.140 2050.580 977.400 2050.840 ;
        RECT 1088.460 2050.580 1088.720 2050.840 ;
        RECT 1273.380 2050.580 1273.640 2050.840 ;
        RECT 1333.640 2050.580 1333.900 2050.840 ;
        RECT 977.600 2050.240 977.860 2050.500 ;
        RECT 1102.260 2050.240 1102.520 2050.500 ;
        RECT 1258.660 2050.240 1258.920 2050.500 ;
        RECT 1337.780 2050.240 1338.040 2050.500 ;
        RECT 984.040 2049.900 984.300 2050.160 ;
        RECT 1073.740 2049.900 1074.000 2050.160 ;
        RECT 1000.140 2049.560 1000.400 2049.820 ;
        RECT 1045.220 2049.560 1045.480 2049.820 ;
        RECT 1301.900 2049.560 1302.160 2049.820 ;
        RECT 1347.900 2049.560 1348.160 2049.820 ;
        RECT 984.500 2049.220 984.760 2049.480 ;
        RECT 1002.900 2049.220 1003.160 2049.480 ;
        RECT 1315.700 2049.220 1315.960 2049.480 ;
        RECT 1336.400 2049.220 1336.660 2049.480 ;
        RECT 976.220 2047.860 976.480 2048.120 ;
        RECT 1014.400 2047.860 1014.660 2048.120 ;
        RECT 983.120 2047.520 983.380 2047.780 ;
        RECT 1028.200 2047.520 1028.460 2047.780 ;
        RECT 982.660 2047.180 982.920 2047.440 ;
        RECT 1062.700 2047.180 1062.960 2047.440 ;
        RECT 975.760 2046.840 976.020 2047.100 ;
        RECT 1076.500 2046.840 1076.760 2047.100 ;
        RECT 983.580 2046.500 983.840 2046.760 ;
        RECT 1097.660 2046.500 1097.920 2046.760 ;
        RECT 976.680 2046.160 976.940 2046.420 ;
        RECT 1097.200 2046.160 1097.460 2046.420 ;
        RECT 972.540 2045.820 972.800 2046.080 ;
        RECT 1111.460 2045.820 1111.720 2046.080 ;
        RECT 965.640 2045.480 965.900 2045.740 ;
        RECT 1111.000 2045.480 1111.260 2045.740 ;
        RECT 1330.880 2036.300 1331.140 2036.560 ;
        RECT 1343.760 2036.300 1344.020 2036.560 ;
        RECT 530.020 1988.360 530.280 1988.620 ;
        RECT 650.540 1988.360 650.800 1988.620 ;
        RECT 579.240 1987.340 579.500 1987.600 ;
        RECT 638.120 1987.340 638.380 1987.600 ;
        RECT 420.540 1978.500 420.800 1978.760 ;
        RECT 420.080 1978.160 420.340 1978.420 ;
        RECT 842.820 1977.820 843.080 1978.080 ;
        RECT 897.560 1977.480 897.820 1977.740 ;
        RECT 998.760 1713.300 999.020 1713.560 ;
        RECT 1001.060 1713.300 1001.320 1713.560 ;
        RECT 1350.200 2028.820 1350.460 2029.080 ;
        RECT 1352.040 2028.820 1352.300 2029.080 ;
        RECT 1350.200 2028.140 1350.460 2028.400 ;
        RECT 1351.580 2028.140 1351.840 2028.400 ;
        RECT 1559.500 2021.680 1559.760 2021.940 ;
        RECT 1560.420 2021.680 1560.680 2021.940 ;
        RECT 1543.400 2004.340 1543.660 2004.600 ;
        RECT 1544.320 2004.340 1544.580 2004.600 ;
        RECT 1350.200 1980.540 1350.460 1980.800 ;
        RECT 1350.660 1980.540 1350.920 1980.800 ;
        RECT 1532.820 1980.540 1533.080 1980.800 ;
        RECT 1543.400 1980.200 1543.660 1980.460 ;
        RECT 1543.860 1980.200 1544.120 1980.460 ;
        RECT 1350.200 1979.860 1350.460 1980.120 ;
        RECT 1350.660 1979.860 1350.920 1980.120 ;
        RECT 1532.360 1979.860 1532.620 1980.120 ;
        RECT 1559.500 1973.060 1559.760 1973.320 ;
        RECT 1560.420 1973.060 1560.680 1973.320 ;
        RECT 1543.860 1956.060 1544.120 1956.320 ;
        RECT 1544.780 1956.060 1545.040 1956.320 ;
        RECT 2294.120 1946.880 2294.380 1947.140 ;
        RECT 2380.140 1946.880 2380.400 1947.140 ;
        RECT 2076.540 1946.540 2076.800 1946.800 ;
        RECT 2321.260 1946.540 2321.520 1946.800 ;
        RECT 2082.980 1946.200 2083.240 1946.460 ;
        RECT 2438.100 1946.200 2438.360 1946.460 ;
        RECT 2083.440 1945.860 2083.700 1946.120 ;
        RECT 2496.980 1945.860 2497.240 1946.120 ;
        RECT 1350.200 1931.920 1350.460 1932.180 ;
        RECT 1351.120 1931.920 1351.380 1932.180 ;
        RECT 1532.360 1931.920 1532.620 1932.180 ;
        RECT 1545.240 1931.580 1545.500 1931.840 ;
        RECT 1532.360 1931.240 1532.620 1931.500 ;
        RECT 1544.320 1931.240 1544.580 1931.500 ;
        RECT 1724.640 1928.520 1724.900 1928.780 ;
        RECT 2044.340 1928.520 2044.600 1928.780 ;
        RECT 1828.140 1927.840 1828.400 1928.100 ;
        RECT 1964.300 1927.840 1964.560 1928.100 ;
        RECT 1745.340 1927.500 1745.600 1927.760 ;
        RECT 1929.340 1927.500 1929.600 1927.760 ;
        RECT 1779.840 1927.160 1780.100 1927.420 ;
        RECT 1998.340 1927.160 1998.600 1927.420 ;
        RECT 1786.740 1926.820 1787.000 1927.080 ;
        RECT 2033.300 1926.820 2033.560 1927.080 ;
        RECT 1759.140 1926.480 1759.400 1926.740 ;
        RECT 2010.300 1926.480 2010.560 1926.740 ;
        RECT 1738.440 1926.140 1738.700 1926.400 ;
        RECT 1987.300 1926.140 1987.560 1926.400 ;
        RECT 1717.280 1925.800 1717.540 1926.060 ;
        RECT 1975.340 1925.800 1975.600 1926.060 ;
        RECT 1772.940 1925.460 1773.200 1925.720 ;
        RECT 2067.340 1925.460 2067.600 1925.720 ;
        RECT 1559.500 1925.120 1559.760 1925.380 ;
        RECT 1560.420 1925.120 1560.680 1925.380 ;
        RECT 1827.680 1925.120 1827.940 1925.380 ;
        RECT 1952.340 1925.120 1952.600 1925.380 ;
        RECT 1351.120 1907.780 1351.380 1908.040 ;
        RECT 1352.040 1907.780 1352.300 1908.040 ;
        RECT 1544.320 1897.240 1544.580 1897.500 ;
        RECT 1545.240 1897.240 1545.500 1897.500 ;
        RECT 1531.900 1883.640 1532.160 1883.900 ;
        RECT 1532.360 1883.640 1532.620 1883.900 ;
        RECT 1752.240 1883.640 1752.500 1883.900 ;
        RECT 1904.500 1883.640 1904.760 1883.900 ;
        RECT 1573.760 1883.300 1574.020 1883.560 ;
        RECT 1574.680 1883.300 1574.940 1883.560 ;
        RECT 1558.580 1876.500 1558.840 1876.760 ;
        RECT 1559.500 1876.500 1559.760 1876.760 ;
        RECT 1821.240 1870.040 1821.500 1870.300 ;
        RECT 1904.500 1870.040 1904.760 1870.300 ;
        RECT 1544.320 1859.500 1544.580 1859.760 ;
        RECT 1545.240 1859.500 1545.500 1859.760 ;
        RECT 1731.540 1849.300 1731.800 1849.560 ;
        RECT 1904.500 1849.300 1904.760 1849.560 ;
        RECT 1350.200 1835.360 1350.460 1835.620 ;
        RECT 1351.120 1835.360 1351.380 1835.620 ;
        RECT 1531.900 1835.360 1532.160 1835.620 ;
        RECT 1532.820 1835.360 1533.080 1835.620 ;
        RECT 1558.580 1828.560 1558.840 1828.820 ;
        RECT 1559.960 1828.560 1560.220 1828.820 ;
        RECT 1544.320 1821.760 1544.580 1822.020 ;
        RECT 1545.240 1821.760 1545.500 1822.020 ;
        RECT 1662.540 1814.620 1662.800 1814.880 ;
        RECT 1904.500 1814.620 1904.760 1814.880 ;
        RECT 1351.120 1801.020 1351.380 1801.280 ;
        RECT 1351.580 1800.680 1351.840 1800.940 ;
        RECT 1350.200 1786.740 1350.460 1787.000 ;
        RECT 1351.580 1786.740 1351.840 1787.000 ;
        RECT 1573.760 1786.740 1574.020 1787.000 ;
        RECT 1574.680 1786.740 1574.940 1787.000 ;
        RECT 1532.820 1786.400 1533.080 1786.660 ;
        RECT 1534.200 1786.400 1534.460 1786.660 ;
        RECT 1350.200 1779.940 1350.460 1780.200 ;
        RECT 1350.660 1779.940 1350.920 1780.200 ;
        RECT 1559.500 1779.940 1559.760 1780.200 ;
        RECT 1560.420 1779.940 1560.680 1780.200 ;
        RECT 1766.040 1766.340 1766.300 1766.600 ;
        RECT 1904.500 1766.340 1904.760 1766.600 ;
        RECT 1533.280 1739.140 1533.540 1739.400 ;
        RECT 1534.200 1739.140 1534.460 1739.400 ;
        RECT 1532.820 1738.460 1533.080 1738.720 ;
        RECT 1533.740 1738.460 1534.000 1738.720 ;
        RECT 1820.780 1738.460 1821.040 1738.720 ;
        RECT 1933.940 1738.460 1934.200 1738.720 ;
        RECT 1800.540 1738.120 1800.800 1738.380 ;
        RECT 1956.940 1738.120 1957.200 1738.380 ;
        RECT 1814.340 1737.780 1814.600 1738.040 ;
        RECT 1990.980 1737.780 1991.240 1738.040 ;
        RECT 1793.640 1737.440 1793.900 1737.700 ;
        RECT 1967.980 1737.440 1968.240 1737.700 ;
        RECT 1807.440 1737.100 1807.700 1737.360 ;
        RECT 2013.980 1737.100 2014.240 1737.360 ;
        RECT 1751.780 1736.760 1752.040 1737.020 ;
        RECT 1979.940 1736.760 1980.200 1737.020 ;
        RECT 1772.480 1736.420 1772.740 1736.680 ;
        RECT 2002.940 1736.420 2003.200 1736.680 ;
        RECT 1806.980 1736.080 1807.240 1736.340 ;
        RECT 2036.980 1736.080 2037.240 1736.340 ;
        RECT 1703.940 1735.740 1704.200 1736.000 ;
        RECT 1944.980 1735.740 1945.240 1736.000 ;
        RECT 1800.080 1735.400 1800.340 1735.660 ;
        RECT 2071.940 1735.400 2072.200 1735.660 ;
        RECT 1365.840 1735.060 1366.100 1735.320 ;
        RECT 1553.060 1735.060 1553.320 1735.320 ;
        RECT 1669.440 1735.060 1669.700 1735.320 ;
        RECT 2059.980 1735.060 2060.240 1735.320 ;
        RECT 1350.660 1732.000 1350.920 1732.260 ;
        RECT 1352.040 1732.000 1352.300 1732.260 ;
        RECT 1559.500 1732.000 1559.760 1732.260 ;
        RECT 1560.420 1732.000 1560.680 1732.260 ;
        RECT 1544.320 1725.200 1544.580 1725.460 ;
        RECT 1545.240 1725.200 1545.500 1725.460 ;
        RECT 1350.660 1724.860 1350.920 1725.120 ;
        RECT 1352.040 1724.860 1352.300 1725.120 ;
        RECT 1559.040 1700.720 1559.300 1700.980 ;
        RECT 1560.420 1700.720 1560.680 1700.980 ;
        RECT 999.220 1694.940 999.480 1695.200 ;
        RECT 1070.520 1694.940 1070.780 1695.200 ;
        RECT 974.840 1694.600 975.100 1694.860 ;
        RECT 1048.900 1694.600 1049.160 1694.860 ;
        RECT 1289.940 1694.600 1290.200 1694.860 ;
        RECT 1347.900 1694.600 1348.160 1694.860 ;
        RECT 999.680 1694.260 999.940 1694.520 ;
        RECT 1076.500 1694.260 1076.760 1694.520 ;
        RECT 1234.740 1694.260 1235.000 1694.520 ;
        RECT 1335.480 1694.260 1335.740 1694.520 ;
        RECT 982.200 1693.920 982.460 1694.180 ;
        RECT 1105.020 1693.920 1105.280 1694.180 ;
        RECT 1186.440 1693.920 1186.700 1694.180 ;
        RECT 1335.940 1693.920 1336.200 1694.180 ;
        RECT 975.300 1693.580 975.560 1693.840 ;
        RECT 1111.000 1693.580 1111.260 1693.840 ;
        RECT 1185.980 1693.580 1186.240 1693.840 ;
        RECT 1336.400 1693.580 1336.660 1693.840 ;
        RECT 1310.640 1692.220 1310.900 1692.480 ;
        RECT 1343.760 1692.220 1344.020 1692.480 ;
        RECT 1573.760 1690.860 1574.020 1691.120 ;
        RECT 1532.820 1690.520 1533.080 1690.780 ;
        RECT 1533.740 1690.520 1534.000 1690.780 ;
        RECT 1574.220 1690.520 1574.480 1690.780 ;
        RECT 1116.060 1689.840 1116.320 1690.100 ;
        RECT 1186.900 1689.840 1187.160 1690.100 ;
        RECT 1159.300 1689.500 1159.560 1689.760 ;
        RECT 1221.400 1689.500 1221.660 1689.760 ;
        RECT 1268.780 1689.500 1269.040 1689.760 ;
        RECT 1315.700 1689.500 1315.960 1689.760 ;
        RECT 1102.260 1689.160 1102.520 1689.420 ;
        RECT 1203.920 1689.160 1204.180 1689.420 ;
        RECT 1214.040 1689.160 1214.300 1689.420 ;
        RECT 1287.180 1689.160 1287.440 1689.420 ;
        RECT 1130.780 1688.820 1131.040 1689.080 ;
        RECT 1197.020 1688.820 1197.280 1689.080 ;
        RECT 1217.720 1688.820 1217.980 1689.080 ;
        RECT 1230.140 1688.820 1230.400 1689.080 ;
        RECT 1248.080 1688.820 1248.340 1689.080 ;
        RECT 1300.980 1688.820 1301.240 1689.080 ;
        RECT 463.780 1688.480 464.040 1688.740 ;
        RECT 468.840 1688.480 469.100 1688.740 ;
        RECT 514.380 1688.480 514.640 1688.740 ;
        RECT 517.140 1688.480 517.400 1688.740 ;
        RECT 1073.740 1688.480 1074.000 1688.740 ;
        RECT 1293.620 1688.480 1293.880 1688.740 ;
        RECT 1030.500 1688.140 1030.760 1688.400 ;
        RECT 1264.180 1688.140 1264.440 1688.400 ;
        RECT 2000.640 1687.800 2000.900 1688.060 ;
        RECT 2302.860 1687.800 2303.120 1688.060 ;
        RECT 2048.940 1687.460 2049.200 1687.720 ;
        RECT 2360.820 1687.460 2361.080 1687.720 ;
        RECT 2042.040 1687.120 2042.300 1687.380 ;
        RECT 2419.700 1687.120 2419.960 1687.380 ;
        RECT 2069.640 1686.780 2069.900 1687.040 ;
        RECT 2477.660 1686.780 2477.920 1687.040 ;
        RECT 1144.580 1686.440 1144.840 1686.700 ;
        RECT 1180.920 1686.440 1181.180 1686.700 ;
        RECT 1197.020 1686.440 1197.280 1686.700 ;
        RECT 1237.040 1686.440 1237.300 1686.700 ;
        RECT 1002.900 1685.420 1003.160 1685.680 ;
        RECT 1038.320 1685.420 1038.580 1685.680 ;
        RECT 1173.100 1684.400 1173.360 1684.660 ;
        RECT 1188.280 1684.400 1188.540 1684.660 ;
        RECT 1193.340 1684.400 1193.600 1684.660 ;
        RECT 1215.420 1684.400 1215.680 1684.660 ;
        RECT 1016.700 1684.060 1016.960 1684.320 ;
        RECT 1020.840 1684.060 1021.100 1684.320 ;
        RECT 1187.820 1684.060 1188.080 1684.320 ;
        RECT 1197.020 1684.060 1197.280 1684.320 ;
        RECT 1238.420 1684.060 1238.680 1684.320 ;
        RECT 1243.940 1684.060 1244.200 1684.320 ;
        RECT 1272.460 1684.060 1272.720 1684.320 ;
        RECT 1291.320 1684.060 1291.580 1684.320 ;
        RECT 1531.440 1683.380 1531.700 1683.640 ;
        RECT 1532.360 1683.380 1532.620 1683.640 ;
        RECT 1572.840 1683.380 1573.100 1683.640 ;
        RECT 1574.220 1683.380 1574.480 1683.640 ;
        RECT 1350.660 1676.580 1350.920 1676.840 ;
        RECT 1351.120 1676.580 1351.380 1676.840 ;
        RECT 1069.600 1642.240 1069.860 1642.500 ;
        RECT 1070.060 1642.240 1070.320 1642.500 ;
        RECT 1104.100 1642.240 1104.360 1642.500 ;
        RECT 1105.020 1642.240 1105.280 1642.500 ;
        RECT 1221.400 1642.240 1221.660 1642.500 ;
        RECT 1243.940 1642.240 1244.200 1642.500 ;
        RECT 1264.180 1642.240 1264.440 1642.500 ;
        RECT 1276.600 1642.240 1276.860 1642.500 ;
        RECT 1351.120 1642.240 1351.380 1642.500 ;
        RECT 1351.580 1642.240 1351.840 1642.500 ;
        RECT 1544.320 1642.240 1544.580 1642.500 ;
        RECT 1545.240 1642.240 1545.500 1642.500 ;
        RECT 1572.840 1635.440 1573.100 1635.700 ;
        RECT 1573.760 1635.440 1574.020 1635.700 ;
        RECT 1532.820 1635.100 1533.080 1635.360 ;
        RECT 1533.740 1635.100 1534.000 1635.360 ;
        RECT 1350.200 1593.620 1350.460 1593.880 ;
        RECT 1351.580 1593.620 1351.840 1593.880 ;
        RECT 1543.860 1593.620 1544.120 1593.880 ;
        RECT 1544.780 1593.620 1545.040 1593.880 ;
        RECT 1559.500 1593.620 1559.760 1593.880 ;
        RECT 1560.420 1593.620 1560.680 1593.880 ;
        RECT 1533.740 1586.820 1534.000 1587.080 ;
        RECT 1534.200 1586.820 1534.460 1587.080 ;
        RECT 1543.860 1586.820 1544.120 1587.080 ;
        RECT 1545.240 1586.820 1545.500 1587.080 ;
        RECT 1350.200 1546.020 1350.460 1546.280 ;
        RECT 1351.580 1546.020 1351.840 1546.280 ;
        RECT 1534.200 1545.680 1534.460 1545.940 ;
        RECT 1559.500 1545.680 1559.760 1545.940 ;
        RECT 1560.420 1545.680 1560.680 1545.940 ;
        RECT 1573.760 1545.680 1574.020 1545.940 ;
        RECT 1574.220 1545.680 1574.480 1545.940 ;
        RECT 1350.660 1545.340 1350.920 1545.600 ;
        RECT 1351.580 1545.340 1351.840 1545.600 ;
        RECT 1534.200 1545.000 1534.460 1545.260 ;
        RECT 1350.660 1510.660 1350.920 1510.920 ;
        RECT 1351.580 1510.660 1351.840 1510.920 ;
        RECT 1532.820 1497.400 1533.080 1497.660 ;
        RECT 1534.200 1497.400 1534.460 1497.660 ;
        RECT 1350.200 1497.060 1350.460 1497.320 ;
        RECT 1351.580 1497.060 1351.840 1497.320 ;
        RECT 1559.500 1497.060 1559.760 1497.320 ;
        RECT 1560.420 1497.060 1560.680 1497.320 ;
        RECT 1487.280 1461.020 1487.540 1461.280 ;
        RECT 1519.020 1461.020 1519.280 1461.280 ;
        RECT 1486.820 1460.680 1487.080 1460.940 ;
        RECT 1526.380 1460.680 1526.640 1460.940 ;
        RECT 1614.240 1459.320 1614.500 1459.580 ;
        RECT 1893.460 1459.320 1893.720 1459.580 ;
        RECT 1495.560 1458.980 1495.820 1459.240 ;
        RECT 1894.380 1458.980 1894.640 1459.240 ;
        RECT 1350.200 1449.460 1350.460 1449.720 ;
        RECT 1351.580 1449.460 1351.840 1449.720 ;
        RECT 1544.320 1449.120 1544.580 1449.380 ;
        RECT 1545.240 1449.120 1545.500 1449.380 ;
        RECT 1559.500 1449.120 1559.760 1449.380 ;
        RECT 1560.420 1449.120 1560.680 1449.380 ;
        RECT 1573.760 1449.120 1574.020 1449.380 ;
        RECT 1574.220 1449.120 1574.480 1449.380 ;
        RECT 1350.660 1448.780 1350.920 1449.040 ;
        RECT 1351.580 1448.780 1351.840 1449.040 ;
        RECT 1544.320 1435.180 1544.580 1435.440 ;
        RECT 1545.240 1435.180 1545.500 1435.440 ;
        RECT 1350.660 1414.100 1350.920 1414.360 ;
        RECT 1351.580 1414.100 1351.840 1414.360 ;
        RECT 1104.100 1400.500 1104.360 1400.760 ;
        RECT 1105.020 1400.500 1105.280 1400.760 ;
        RECT 1350.200 1400.500 1350.460 1400.760 ;
        RECT 1351.580 1400.500 1351.840 1400.760 ;
        RECT 1543.400 1400.500 1543.660 1400.760 ;
        RECT 1544.780 1400.500 1545.040 1400.760 ;
        RECT 1559.500 1400.500 1559.760 1400.760 ;
        RECT 1560.420 1400.500 1560.680 1400.760 ;
        RECT 1069.140 1352.900 1069.400 1353.160 ;
        RECT 1069.600 1352.560 1069.860 1352.820 ;
        RECT 1104.100 1352.560 1104.360 1352.820 ;
        RECT 1105.020 1352.560 1105.280 1352.820 ;
        RECT 1350.200 1352.560 1350.460 1352.820 ;
        RECT 1351.120 1352.560 1351.380 1352.820 ;
        RECT 1543.400 1352.560 1543.660 1352.820 ;
        RECT 1544.320 1352.560 1544.580 1352.820 ;
        RECT 1559.500 1352.560 1559.760 1352.820 ;
        RECT 1560.420 1352.560 1560.680 1352.820 ;
        RECT 1573.760 1352.560 1574.020 1352.820 ;
        RECT 1574.220 1352.560 1574.480 1352.820 ;
        RECT 1532.820 1338.620 1533.080 1338.880 ;
        RECT 1533.740 1338.620 1534.000 1338.880 ;
        RECT 1350.660 1317.540 1350.920 1317.800 ;
        RECT 1351.580 1317.540 1351.840 1317.800 ;
        RECT 1104.100 1303.940 1104.360 1304.200 ;
        RECT 1105.020 1303.940 1105.280 1304.200 ;
        RECT 1350.200 1303.940 1350.460 1304.200 ;
        RECT 1351.580 1303.940 1351.840 1304.200 ;
        RECT 1069.140 1303.600 1069.400 1303.860 ;
        RECT 1069.600 1303.600 1069.860 1303.860 ;
        RECT 1543.400 1297.140 1543.660 1297.400 ;
        RECT 1545.240 1297.140 1545.500 1297.400 ;
        RECT 1545.240 1269.940 1545.500 1270.200 ;
        RECT 1544.320 1269.260 1544.580 1269.520 ;
        RECT 1104.100 1256.340 1104.360 1256.600 ;
        RECT 1105.020 1256.340 1105.280 1256.600 ;
        RECT 1350.200 1256.340 1350.460 1256.600 ;
        RECT 1351.580 1256.000 1351.840 1256.260 ;
        RECT 1544.320 1220.980 1544.580 1221.240 ;
        RECT 1544.320 1220.300 1544.580 1220.560 ;
        RECT 1350.660 1207.380 1350.920 1207.640 ;
        RECT 1351.580 1207.380 1351.840 1207.640 ;
        RECT 1350.200 1159.100 1350.460 1159.360 ;
        RECT 1352.040 1159.100 1352.300 1159.360 ;
        RECT 1543.860 1159.100 1544.120 1159.360 ;
        RECT 1544.320 1159.100 1544.580 1159.360 ;
        RECT 1351.120 1110.820 1351.380 1111.080 ;
        RECT 1352.040 1110.820 1352.300 1111.080 ;
        RECT 1530.980 1110.820 1531.240 1111.080 ;
        RECT 1532.820 1110.820 1533.080 1111.080 ;
        RECT 1351.120 1076.820 1351.380 1077.080 ;
        RECT 1351.120 1075.800 1351.380 1076.060 ;
        RECT 1530.980 1075.800 1531.240 1076.060 ;
        RECT 1532.820 1075.800 1533.080 1076.060 ;
        RECT 1730.620 1062.540 1730.880 1062.800 ;
        RECT 1731.540 1062.540 1731.800 1062.800 ;
        RECT 1489.580 1055.400 1489.840 1055.660 ;
        RECT 1519.480 1055.400 1519.740 1055.660 ;
        RECT 993.700 1052.000 993.960 1052.260 ;
        RECT 1062.700 1052.000 1062.960 1052.260 ;
        RECT 1237.040 1048.600 1237.300 1048.860 ;
        RECT 1239.340 1048.600 1239.600 1048.860 ;
        RECT 982.660 1025.480 982.920 1025.740 ;
        RECT 1146.420 1025.480 1146.680 1025.740 ;
        RECT 975.760 1025.140 976.020 1025.400 ;
        RECT 1152.400 1025.140 1152.660 1025.400 ;
        RECT 972.540 1024.800 972.800 1025.060 ;
        RECT 1154.700 1024.800 1154.960 1025.060 ;
        RECT 1472.100 1024.800 1472.360 1025.060 ;
        RECT 1891.620 1024.800 1891.880 1025.060 ;
        RECT 965.640 1024.460 965.900 1024.720 ;
        RECT 1163.440 1024.460 1163.700 1024.720 ;
        RECT 1385.620 1024.460 1385.880 1024.720 ;
        RECT 1892.080 1024.460 1892.340 1024.720 ;
        RECT 997.380 1021.060 997.640 1021.320 ;
        RECT 1223.240 1021.060 1223.500 1021.320 ;
        RECT 1250.840 1021.060 1251.100 1021.320 ;
        RECT 1339.160 1021.060 1339.420 1021.320 ;
        RECT 1571.920 1021.060 1572.180 1021.320 ;
        RECT 1900.820 1021.060 1901.080 1021.320 ;
        RECT 988.640 1020.720 988.900 1020.980 ;
        RECT 1228.300 1020.720 1228.560 1020.980 ;
        RECT 1243.480 1020.720 1243.740 1020.980 ;
        RECT 1341.000 1020.720 1341.260 1020.980 ;
        RECT 1469.340 1020.720 1469.600 1020.980 ;
        RECT 1704.400 1020.720 1704.660 1020.980 ;
        RECT 1716.820 1020.720 1717.080 1020.980 ;
        RECT 2084.360 1020.720 2084.620 1020.980 ;
        RECT 996.920 1020.380 997.180 1020.640 ;
        RECT 987.720 1020.040 987.980 1020.300 ;
        RECT 1258.200 1020.040 1258.460 1020.300 ;
        RECT 1266.020 1020.380 1266.280 1020.640 ;
        RECT 1337.320 1020.380 1337.580 1020.640 ;
        RECT 1530.520 1020.380 1530.780 1020.640 ;
        RECT 1903.580 1020.380 1903.840 1020.640 ;
        RECT 1268.320 1020.040 1268.580 1020.300 ;
        RECT 1286.260 1020.040 1286.520 1020.300 ;
        RECT 1338.700 1020.040 1338.960 1020.300 ;
        RECT 1503.840 1020.040 1504.100 1020.300 ;
        RECT 1897.600 1020.040 1897.860 1020.300 ;
        RECT 996.460 1019.700 996.720 1019.960 ;
        RECT 1290.400 1019.700 1290.660 1019.960 ;
        RECT 1495.100 1019.700 1495.360 1019.960 ;
        RECT 1901.280 1019.700 1901.540 1019.960 ;
        RECT 989.100 1019.360 989.360 1019.620 ;
        RECT 1283.500 1019.360 1283.760 1019.620 ;
        RECT 1462.440 1019.360 1462.700 1019.620 ;
        RECT 1898.520 1019.360 1898.780 1019.620 ;
        RECT 990.480 1019.020 990.740 1019.280 ;
        RECT 1300.060 1019.020 1300.320 1019.280 ;
        RECT 1461.980 1019.020 1462.240 1019.280 ;
        RECT 1898.060 1019.020 1898.320 1019.280 ;
        RECT 988.180 1018.680 988.440 1018.940 ;
        RECT 1312.940 1018.680 1313.200 1018.940 ;
        RECT 1434.840 1018.680 1435.100 1018.940 ;
        RECT 1893.000 1018.680 1893.260 1018.940 ;
        RECT 989.560 1018.340 989.820 1018.600 ;
        RECT 1324.900 1018.340 1325.160 1018.600 ;
        RECT 1357.100 1018.340 1357.360 1018.600 ;
        RECT 1849.300 1018.340 1849.560 1018.600 ;
        RECT 990.940 1018.000 991.200 1018.260 ;
        RECT 1335.480 1018.000 1335.740 1018.260 ;
        RECT 1400.340 1018.000 1400.600 1018.260 ;
        RECT 1898.980 1018.000 1899.240 1018.260 ;
        RECT 990.020 1017.660 990.280 1017.920 ;
        RECT 1347.900 1017.660 1348.160 1017.920 ;
        RECT 1352.040 1017.660 1352.300 1017.920 ;
        RECT 1899.440 1017.660 1899.700 1017.920 ;
        RECT 991.400 1017.320 991.660 1017.580 ;
        RECT 1197.940 1017.320 1198.200 1017.580 ;
        RECT 1203.460 1017.320 1203.720 1017.580 ;
        RECT 1343.300 1017.320 1343.560 1017.580 ;
        RECT 1565.480 1017.320 1565.740 1017.580 ;
        RECT 1890.700 1017.320 1890.960 1017.580 ;
        RECT 992.780 1016.980 993.040 1017.240 ;
        RECT 1159.760 1016.980 1160.020 1017.240 ;
        RECT 1276.140 1016.980 1276.400 1017.240 ;
        RECT 1340.540 1016.980 1340.800 1017.240 ;
        RECT 1478.540 1016.980 1478.800 1017.240 ;
        RECT 1766.500 1016.980 1766.760 1017.240 ;
        RECT 1257.740 1016.640 1258.000 1016.900 ;
        RECT 1286.260 1016.640 1286.520 1016.900 ;
        RECT 1297.300 1016.640 1297.560 1016.900 ;
        RECT 1336.860 1016.640 1337.120 1016.900 ;
        RECT 1512.120 1016.640 1512.380 1016.900 ;
        RECT 1656.100 1016.640 1656.360 1016.900 ;
        RECT 1490.040 1016.300 1490.300 1016.560 ;
        RECT 1622.980 1016.300 1623.240 1016.560 ;
        RECT 1870.000 1014.600 1870.260 1014.860 ;
        RECT 1886.560 1014.600 1886.820 1014.860 ;
        RECT 1048.440 1013.920 1048.700 1014.180 ;
        RECT 1214.500 1013.920 1214.760 1014.180 ;
        RECT 977.140 1013.580 977.400 1013.840 ;
        RECT 1189.660 1013.580 1189.920 1013.840 ;
        RECT 984.500 1013.240 984.760 1013.500 ;
        RECT 1145.500 1013.240 1145.760 1013.500 ;
        RECT 1173.100 1013.240 1173.360 1013.500 ;
        RECT 1218.640 1013.240 1218.900 1013.500 ;
        RECT 789.920 1012.900 790.180 1013.160 ;
        RECT 888.360 1012.900 888.620 1013.160 ;
        RECT 983.120 1012.900 983.380 1013.160 ;
        RECT 1012.560 1012.900 1012.820 1013.160 ;
        RECT 1020.840 1012.900 1021.100 1013.160 ;
        RECT 1196.100 1012.900 1196.360 1013.160 ;
        RECT 796.820 1012.560 797.080 1012.820 ;
        RECT 844.660 1012.560 844.920 1012.820 ;
        RECT 977.600 1012.560 977.860 1012.820 ;
        RECT 1204.380 1012.900 1204.640 1013.160 ;
        RECT 1213.580 1012.900 1213.840 1013.160 ;
        RECT 1238.420 1013.920 1238.680 1014.180 ;
        RECT 1255.440 1013.920 1255.700 1014.180 ;
        RECT 1333.180 1014.260 1333.440 1014.520 ;
        RECT 1790.420 1014.260 1790.680 1014.520 ;
        RECT 1331.340 1013.920 1331.600 1014.180 ;
        RECT 1334.560 1013.920 1334.820 1014.180 ;
        RECT 1338.700 1013.920 1338.960 1014.180 ;
        RECT 1353.420 1013.920 1353.680 1014.180 ;
        RECT 1355.260 1013.920 1355.520 1014.180 ;
        RECT 1358.020 1013.920 1358.280 1014.180 ;
        RECT 1261.420 1013.580 1261.680 1013.840 ;
        RECT 1341.460 1013.580 1341.720 1013.840 ;
        RECT 1488.660 1013.580 1488.920 1013.840 ;
        RECT 1513.040 1013.920 1513.300 1014.180 ;
        RECT 1538.340 1013.920 1538.600 1014.180 ;
        RECT 1203.920 1012.560 1204.180 1012.820 ;
        RECT 1286.720 1013.240 1286.980 1013.500 ;
        RECT 1287.640 1013.240 1287.900 1013.500 ;
        RECT 1289.940 1013.240 1290.200 1013.500 ;
        RECT 1293.620 1013.240 1293.880 1013.500 ;
        RECT 1318.000 1013.240 1318.260 1013.500 ;
        RECT 1487.740 1013.240 1488.000 1013.500 ;
        RECT 1509.360 1013.240 1509.620 1013.500 ;
        RECT 1253.140 1012.900 1253.400 1013.160 ;
        RECT 1345.600 1012.900 1345.860 1013.160 ;
        RECT 1496.940 1012.900 1497.200 1013.160 ;
        RECT 1511.660 1012.900 1511.920 1013.160 ;
        RECT 783.020 1012.220 783.280 1012.480 ;
        RECT 884.220 1012.220 884.480 1012.480 ;
        RECT 1000.140 1012.220 1000.400 1012.480 ;
        RECT 1180.000 1012.220 1180.260 1012.480 ;
        RECT 1180.460 1012.220 1180.720 1012.480 ;
        RECT 1186.440 1012.220 1186.700 1012.480 ;
        RECT 1197.020 1012.220 1197.280 1012.480 ;
        RECT 1218.180 1012.220 1218.440 1012.480 ;
        RECT 1218.640 1012.220 1218.900 1012.480 ;
        RECT 1221.400 1012.220 1221.660 1012.480 ;
        RECT 707.120 1011.880 707.380 1012.140 ;
        RECT 841.900 1011.880 842.160 1012.140 ;
        RECT 984.040 1011.880 984.300 1012.140 ;
        RECT 1173.100 1011.880 1173.360 1012.140 ;
        RECT 769.220 1011.540 769.480 1011.800 ;
        RECT 910.900 1011.540 911.160 1011.800 ;
        RECT 976.220 1011.540 976.480 1011.800 ;
        RECT 1003.820 1011.540 1004.080 1011.800 ;
        RECT 1038.320 1011.540 1038.580 1011.800 ;
        RECT 1093.060 1011.540 1093.320 1011.800 ;
        RECT 1104.100 1011.540 1104.360 1011.800 ;
        RECT 1105.480 1011.540 1105.740 1011.800 ;
        RECT 1145.040 1011.540 1145.300 1011.800 ;
        RECT 1197.480 1011.540 1197.740 1011.800 ;
        RECT 1217.260 1011.540 1217.520 1011.800 ;
        RECT 1346.520 1012.560 1346.780 1012.820 ;
        RECT 1489.580 1012.560 1489.840 1012.820 ;
        RECT 1528.220 1013.580 1528.480 1013.840 ;
        RECT 1530.980 1013.580 1531.240 1013.840 ;
        RECT 1550.300 1013.920 1550.560 1014.180 ;
        RECT 1762.820 1013.920 1763.080 1014.180 ;
        RECT 1777.540 1013.920 1777.800 1014.180 ;
        RECT 1779.840 1013.920 1780.100 1014.180 ;
        RECT 1870.000 1013.920 1870.260 1014.180 ;
        RECT 2061.820 1013.920 2062.080 1014.180 ;
        RECT 2287.220 1013.920 2287.480 1014.180 ;
        RECT 1512.580 1013.240 1512.840 1013.500 ;
        RECT 1524.540 1012.900 1524.800 1013.160 ;
        RECT 1542.940 1012.900 1543.200 1013.160 ;
        RECT 1519.020 1012.560 1519.280 1012.820 ;
        RECT 1521.320 1012.560 1521.580 1012.820 ;
        RECT 1541.560 1012.560 1541.820 1012.820 ;
        RECT 1545.240 1012.560 1545.500 1012.820 ;
        RECT 1886.100 1013.580 1886.360 1013.840 ;
        RECT 1998.340 1013.580 1998.600 1013.840 ;
        RECT 2000.640 1013.580 2000.900 1013.840 ;
        RECT 2057.220 1013.580 2057.480 1013.840 ;
        RECT 2287.680 1013.580 2287.940 1013.840 ;
        RECT 1553.060 1013.240 1553.320 1013.500 ;
        RECT 1673.120 1013.240 1673.380 1013.500 ;
        RECT 1708.540 1013.240 1708.800 1013.500 ;
        RECT 1625.280 1012.900 1625.540 1013.160 ;
        RECT 1724.180 1012.900 1724.440 1013.160 ;
        RECT 1751.320 1012.900 1751.580 1013.160 ;
        RECT 1628.500 1012.560 1628.760 1012.820 ;
        RECT 1721.420 1012.560 1721.680 1012.820 ;
        RECT 1724.640 1012.560 1724.900 1012.820 ;
        RECT 1743.040 1012.560 1743.300 1012.820 ;
        RECT 1745.340 1012.560 1745.600 1012.820 ;
        RECT 1747.640 1012.560 1747.900 1012.820 ;
        RECT 1751.780 1012.560 1752.040 1012.820 ;
        RECT 1762.820 1013.240 1763.080 1013.500 ;
        RECT 1790.420 1013.240 1790.680 1013.500 ;
        RECT 1790.880 1013.240 1791.140 1013.500 ;
        RECT 1793.640 1013.240 1793.900 1013.500 ;
        RECT 1794.100 1013.240 1794.360 1013.500 ;
        RECT 2086.200 1013.240 2086.460 1013.500 ;
        RECT 1753.160 1012.900 1753.420 1013.160 ;
        RECT 2085.740 1012.900 2086.000 1013.160 ;
        RECT 2085.280 1012.560 2085.540 1012.820 ;
        RECT 1237.040 1012.220 1237.300 1012.480 ;
        RECT 1340.080 1012.220 1340.340 1012.480 ;
        RECT 1411.380 1012.220 1411.640 1012.480 ;
        RECT 1414.140 1012.220 1414.400 1012.480 ;
        RECT 1467.500 1012.220 1467.760 1012.480 ;
        RECT 1468.880 1012.220 1469.140 1012.480 ;
        RECT 1480.380 1012.220 1480.640 1012.480 ;
        RECT 1482.680 1012.220 1482.940 1012.480 ;
        RECT 1502.000 1012.220 1502.260 1012.480 ;
        RECT 762.320 1011.200 762.580 1011.460 ;
        RECT 905.380 1011.200 905.640 1011.460 ;
        RECT 996.000 1011.200 996.260 1011.460 ;
        RECT 1053.500 1011.200 1053.760 1011.460 ;
        RECT 1100.420 1011.200 1100.680 1011.460 ;
        RECT 1145.500 1011.200 1145.760 1011.460 ;
        RECT 1196.560 1011.200 1196.820 1011.460 ;
        RECT 1297.760 1011.880 1298.020 1012.140 ;
        RECT 1324.440 1011.880 1324.700 1012.140 ;
        RECT 1334.100 1011.880 1334.360 1012.140 ;
        RECT 1334.560 1011.880 1334.820 1012.140 ;
        RECT 1352.960 1011.880 1353.220 1012.140 ;
        RECT 1441.280 1011.880 1441.540 1012.140 ;
        RECT 1611.020 1011.880 1611.280 1012.140 ;
        RECT 1665.300 1011.880 1665.560 1012.140 ;
        RECT 1669.440 1011.880 1669.700 1012.140 ;
        RECT 1669.900 1011.880 1670.160 1012.140 ;
        RECT 1872.760 1011.880 1873.020 1012.140 ;
        RECT 1286.720 1011.540 1286.980 1011.800 ;
        RECT 1304.200 1011.540 1304.460 1011.800 ;
        RECT 1304.660 1011.540 1304.920 1011.800 ;
        RECT 1332.720 1011.540 1332.980 1011.800 ;
        RECT 1333.180 1011.540 1333.440 1011.800 ;
        RECT 1353.880 1011.540 1354.140 1011.800 ;
        RECT 1506.600 1011.540 1506.860 1011.800 ;
        RECT 1873.220 1011.540 1873.480 1011.800 ;
        RECT 1875.520 1012.220 1875.780 1012.480 ;
        RECT 1893.920 1012.220 1894.180 1012.480 ;
        RECT 2000.640 1012.220 2000.900 1012.480 ;
        RECT 2294.120 1012.220 2294.380 1012.480 ;
        RECT 1874.140 1011.880 1874.400 1012.140 ;
        RECT 1892.540 1011.540 1892.800 1011.800 ;
        RECT 1245.320 1011.200 1245.580 1011.460 ;
        RECT 1294.080 1011.200 1294.340 1011.460 ;
        RECT 517.140 1010.860 517.400 1011.120 ;
        RECT 712.640 1010.860 712.900 1011.120 ;
        RECT 755.420 1010.860 755.680 1011.120 ;
        RECT 901.240 1010.860 901.500 1011.120 ;
        RECT 995.080 1010.860 995.340 1011.120 ;
        RECT 468.840 1010.520 469.100 1010.780 ;
        RECT 673.540 1010.520 673.800 1010.780 ;
        RECT 720.920 1010.520 721.180 1010.780 ;
        RECT 892.500 1010.520 892.760 1010.780 ;
        RECT 995.540 1010.520 995.800 1010.780 ;
        RECT 1289.940 1010.860 1290.200 1011.120 ;
        RECT 1346.980 1011.200 1347.240 1011.460 ;
        RECT 1444.040 1011.200 1444.300 1011.460 ;
        RECT 1479.920 1011.200 1480.180 1011.460 ;
        RECT 1484.980 1011.200 1485.240 1011.460 ;
        RECT 1899.900 1011.200 1900.160 1011.460 ;
        RECT 2046.640 1011.880 2046.900 1012.140 ;
        RECT 2048.940 1011.880 2049.200 1012.140 ;
        RECT 2087.120 1011.880 2087.380 1012.140 ;
        RECT 2069.180 1011.540 2069.440 1011.800 ;
        RECT 2540.220 1011.540 2540.480 1011.800 ;
        RECT 2053.080 1011.200 2053.340 1011.460 ;
        RECT 2539.760 1011.200 2540.020 1011.460 ;
        RECT 1322.600 1010.860 1322.860 1011.120 ;
        RECT 1346.060 1010.860 1346.320 1011.120 ;
        RECT 1427.940 1010.860 1428.200 1011.120 ;
        RECT 1891.160 1010.860 1891.420 1011.120 ;
        RECT 2041.580 1010.860 2041.840 1011.120 ;
        RECT 2539.300 1010.860 2539.560 1011.120 ;
        RECT 983.580 1010.180 983.840 1010.440 ;
        RECT 1138.600 1010.180 1138.860 1010.440 ;
        RECT 1145.500 1010.180 1145.760 1010.440 ;
        RECT 1196.560 1010.180 1196.820 1010.440 ;
        RECT 1197.020 1010.180 1197.280 1010.440 ;
        RECT 1200.240 1010.180 1200.500 1010.440 ;
        RECT 1221.400 1010.180 1221.660 1010.440 ;
        RECT 1224.160 1010.180 1224.420 1010.440 ;
        RECT 976.680 1009.840 976.940 1010.100 ;
        RECT 1133.080 1009.840 1133.340 1010.100 ;
        RECT 1145.960 1009.840 1146.220 1010.100 ;
        RECT 1179.540 1009.840 1179.800 1010.100 ;
        RECT 1180.000 1009.840 1180.260 1010.100 ;
        RECT 1230.600 1009.840 1230.860 1010.100 ;
        RECT 1307.880 1010.520 1308.140 1010.780 ;
        RECT 1328.120 1010.520 1328.380 1010.780 ;
        RECT 1347.440 1010.520 1347.700 1010.780 ;
        RECT 1376.880 1010.520 1377.140 1010.780 ;
        RECT 1379.640 1010.520 1379.900 1010.780 ;
        RECT 1409.080 1010.520 1409.340 1010.780 ;
        RECT 1413.680 1010.520 1413.940 1010.780 ;
        RECT 1415.980 1010.520 1416.240 1010.780 ;
        RECT 1680.020 1010.520 1680.280 1010.780 ;
        RECT 1737.980 1010.520 1738.240 1010.780 ;
        RECT 1794.100 1010.520 1794.360 1010.780 ;
        RECT 1795.020 1010.520 1795.280 1010.780 ;
        RECT 1800.540 1010.520 1800.800 1010.780 ;
        RECT 1823.540 1010.520 1823.800 1010.780 ;
        RECT 1828.140 1010.520 1828.400 1010.780 ;
        RECT 1867.700 1010.520 1867.960 1010.780 ;
        RECT 1869.540 1010.520 1869.800 1010.780 ;
        RECT 1879.660 1010.520 1879.920 1010.780 ;
        RECT 2528.720 1010.520 2528.980 1010.780 ;
        RECT 1283.040 1010.180 1283.300 1010.440 ;
        RECT 1352.500 1010.180 1352.760 1010.440 ;
        RECT 1504.300 1010.180 1504.560 1010.440 ;
        RECT 1507.980 1010.180 1508.240 1010.440 ;
        RECT 1311.100 1009.840 1311.360 1010.100 ;
        RECT 1311.560 1009.840 1311.820 1010.100 ;
        RECT 1341.920 1009.840 1342.180 1010.100 ;
        RECT 1374.580 1009.840 1374.840 1010.100 ;
        RECT 1397.120 1009.840 1397.380 1010.100 ;
        RECT 1402.640 1009.840 1402.900 1010.100 ;
        RECT 1407.240 1009.840 1407.500 1010.100 ;
        RECT 1493.260 1009.840 1493.520 1010.100 ;
        RECT 1512.580 1010.180 1512.840 1010.440 ;
        RECT 1508.900 1009.840 1509.160 1010.100 ;
        RECT 1534.660 1009.840 1534.920 1010.100 ;
        RECT 1573.300 1009.840 1573.560 1010.100 ;
        RECT 1582.500 1010.180 1582.760 1010.440 ;
        RECT 1586.640 1010.180 1586.900 1010.440 ;
        RECT 1591.240 1010.180 1591.500 1010.440 ;
        RECT 1593.540 1010.180 1593.800 1010.440 ;
        RECT 1599.060 1010.180 1599.320 1010.440 ;
        RECT 1600.440 1010.180 1600.700 1010.440 ;
        RECT 1660.700 1010.180 1660.960 1010.440 ;
        RECT 1669.900 1010.180 1670.160 1010.440 ;
        RECT 1755.920 1010.180 1756.180 1010.440 ;
        RECT 2086.660 1010.180 2086.920 1010.440 ;
        RECT 978.060 1009.500 978.320 1009.760 ;
        RECT 1057.180 1009.500 1057.440 1009.760 ;
        RECT 1062.240 1009.500 1062.500 1009.760 ;
        RECT 1191.500 1009.500 1191.760 1009.760 ;
        RECT 1200.240 1009.500 1200.500 1009.760 ;
        RECT 1217.720 1009.500 1217.980 1009.760 ;
        RECT 1267.860 1009.500 1268.120 1009.760 ;
        RECT 1293.620 1009.500 1293.880 1009.760 ;
        RECT 1307.420 1009.500 1307.680 1009.760 ;
        RECT 1310.640 1009.500 1310.900 1009.760 ;
        RECT 984.960 1009.160 985.220 1009.420 ;
        RECT 991.860 1008.820 992.120 1009.080 ;
        RECT 1011.640 1008.820 1011.900 1009.080 ;
        RECT 1012.560 1009.160 1012.820 1009.420 ;
        RECT 1083.400 1009.160 1083.660 1009.420 ;
        RECT 1089.840 1009.160 1090.100 1009.420 ;
        RECT 1228.760 1009.160 1229.020 1009.420 ;
        RECT 1272.920 1009.160 1273.180 1009.420 ;
        RECT 1304.660 1009.160 1304.920 1009.420 ;
        RECT 1310.180 1009.160 1310.440 1009.420 ;
        RECT 1334.560 1009.500 1334.820 1009.760 ;
        RECT 1487.280 1009.500 1487.540 1009.760 ;
        RECT 1493.720 1009.500 1493.980 1009.760 ;
        RECT 1502.460 1009.500 1502.720 1009.760 ;
        RECT 1582.960 1009.500 1583.220 1009.760 ;
        RECT 1593.080 1009.840 1593.340 1010.100 ;
        RECT 1645.520 1009.840 1645.780 1010.100 ;
        RECT 1712.680 1009.840 1712.940 1010.100 ;
        RECT 1717.280 1009.840 1717.540 1010.100 ;
        RECT 1734.300 1009.840 1734.560 1010.100 ;
        RECT 1738.440 1009.840 1738.700 1010.100 ;
        RECT 1786.280 1009.840 1786.540 1010.100 ;
        RECT 2084.820 1009.840 2085.080 1010.100 ;
        RECT 1600.900 1009.500 1601.160 1009.760 ;
        RECT 1831.820 1009.500 1832.080 1009.760 ;
        RECT 1113.760 1008.820 1114.020 1009.080 ;
        RECT 1196.100 1008.820 1196.360 1009.080 ;
        RECT 1237.040 1008.820 1237.300 1009.080 ;
        RECT 1278.440 1008.820 1278.700 1009.080 ;
        RECT 1342.380 1009.160 1342.640 1009.420 ;
        RECT 1496.480 1009.160 1496.740 1009.420 ;
        RECT 1508.900 1009.160 1509.160 1009.420 ;
        RECT 1509.360 1009.160 1509.620 1009.420 ;
        RECT 1530.980 1009.160 1531.240 1009.420 ;
        RECT 1531.440 1009.160 1531.700 1009.420 ;
        RECT 1535.120 1009.160 1535.380 1009.420 ;
        RECT 1497.400 1008.820 1497.660 1009.080 ;
        RECT 1566.400 1009.160 1566.660 1009.420 ;
        RECT 1873.220 1009.160 1873.480 1009.420 ;
        RECT 1900.360 1009.160 1900.620 1009.420 ;
        RECT 2037.900 1009.160 2038.160 1009.420 ;
        RECT 2042.040 1009.160 2042.300 1009.420 ;
        RECT 1548.920 1008.820 1549.180 1009.080 ;
        RECT 1605.960 1008.820 1606.220 1009.080 ;
        RECT 2065.960 1009.160 2066.220 1009.420 ;
        RECT 2069.640 1009.160 2069.900 1009.420 ;
        RECT 2079.300 1009.160 2079.560 1009.420 ;
        RECT 2083.440 1009.160 2083.700 1009.420 ;
        RECT 2094.020 1008.820 2094.280 1009.080 ;
        RECT 1003.820 1008.480 1004.080 1008.740 ;
        RECT 1092.140 1008.480 1092.400 1008.740 ;
        RECT 1093.060 1008.480 1093.320 1008.740 ;
        RECT 1145.040 1008.480 1145.300 1008.740 ;
        RECT 1197.480 1008.480 1197.740 1008.740 ;
        RECT 1245.320 1008.480 1245.580 1008.740 ;
        RECT 1264.180 1008.480 1264.440 1008.740 ;
        RECT 1268.780 1008.480 1269.040 1008.740 ;
        RECT 1274.760 1008.480 1275.020 1008.740 ;
        RECT 1311.560 1008.480 1311.820 1008.740 ;
        RECT 998.760 1008.140 999.020 1008.400 ;
        RECT 1097.200 1008.140 1097.460 1008.400 ;
        RECT 1179.540 1008.140 1179.800 1008.400 ;
        RECT 1204.840 1008.140 1205.100 1008.400 ;
        RECT 1261.880 1008.140 1262.140 1008.400 ;
        RECT 1315.240 1008.140 1315.500 1008.400 ;
        RECT 638.120 1007.800 638.380 1008.060 ;
        RECT 669.860 1007.800 670.120 1008.060 ;
        RECT 994.620 1007.800 994.880 1008.060 ;
        RECT 1078.800 1007.800 1079.060 1008.060 ;
        RECT 1209.900 1007.800 1210.160 1008.060 ;
        RECT 1214.040 1007.800 1214.300 1008.060 ;
        RECT 1222.780 1007.800 1223.040 1008.060 ;
        RECT 1339.620 1008.480 1339.880 1008.740 ;
        RECT 1368.140 1008.480 1368.400 1008.740 ;
        RECT 1372.740 1008.480 1373.000 1008.740 ;
        RECT 1383.320 1008.480 1383.580 1008.740 ;
        RECT 1386.540 1008.480 1386.800 1008.740 ;
        RECT 1489.120 1008.480 1489.380 1008.740 ;
        RECT 1534.660 1008.480 1534.920 1008.740 ;
        RECT 1552.600 1008.480 1552.860 1008.740 ;
        RECT 1554.440 1008.480 1554.700 1008.740 ;
        RECT 1769.260 1008.480 1769.520 1008.740 ;
        RECT 1772.480 1008.480 1772.740 1008.740 ;
        RECT 1782.140 1008.480 1782.400 1008.740 ;
        RECT 1786.740 1008.480 1787.000 1008.740 ;
        RECT 1330.420 1008.140 1330.680 1008.400 ;
        RECT 1343.300 1008.140 1343.560 1008.400 ;
        RECT 1496.020 1008.140 1496.280 1008.400 ;
        RECT 1555.820 1008.140 1556.080 1008.400 ;
        RECT 1450.480 1007.800 1450.740 1008.060 ;
        RECT 1455.080 1007.800 1455.340 1008.060 ;
        RECT 1461.060 1007.800 1461.320 1008.060 ;
        RECT 1462.440 1007.800 1462.700 1008.060 ;
        RECT 1488.200 1007.800 1488.460 1008.060 ;
        RECT 1518.100 1007.800 1518.360 1008.060 ;
        RECT 650.540 1007.460 650.800 1007.720 ;
        RECT 671.700 1007.460 671.960 1007.720 ;
        RECT 992.320 1007.460 992.580 1007.720 ;
        RECT 1053.040 1007.460 1053.300 1007.720 ;
        RECT 1053.500 1007.460 1053.760 1007.720 ;
        RECT 1100.420 1007.460 1100.680 1007.720 ;
        RECT 1191.500 1007.460 1191.760 1007.720 ;
        RECT 1210.360 1007.460 1210.620 1007.720 ;
        RECT 1293.620 1007.460 1293.880 1007.720 ;
        RECT 1333.640 1007.460 1333.900 1007.720 ;
        RECT 1335.020 1007.460 1335.280 1007.720 ;
        RECT 1340.540 1007.460 1340.800 1007.720 ;
        RECT 1417.820 1007.460 1418.080 1007.720 ;
        RECT 1421.040 1007.460 1421.300 1007.720 ;
        RECT 1437.600 1007.460 1437.860 1007.720 ;
        RECT 1441.740 1007.460 1442.000 1007.720 ;
        RECT 1446.340 1007.460 1446.600 1007.720 ;
        RECT 1448.640 1007.460 1448.900 1007.720 ;
        RECT 1452.780 1007.460 1453.040 1007.720 ;
        RECT 1455.540 1007.460 1455.800 1007.720 ;
        RECT 1459.220 1007.460 1459.480 1007.720 ;
        RECT 1461.980 1007.460 1462.240 1007.720 ;
        RECT 1511.660 1007.460 1511.920 1007.720 ;
        RECT 1545.700 1007.460 1545.960 1007.720 ;
        RECT 1611.020 1007.460 1611.280 1007.720 ;
        RECT 1614.240 1007.460 1614.500 1007.720 ;
        RECT 1617.460 1007.460 1617.720 1007.720 ;
        RECT 1635.400 1007.460 1635.660 1007.720 ;
        RECT 1803.760 1007.460 1804.020 1007.720 ;
        RECT 1806.980 1007.460 1807.240 1007.720 ;
        RECT 910.900 1001.680 911.160 1001.940 ;
        RECT 912.280 1001.680 912.540 1001.940 ;
        RECT 1532.820 1001.000 1533.080 1001.260 ;
        RECT 1535.810 1001.000 1536.070 1001.260 ;
        RECT 1559.500 1001.000 1559.760 1001.260 ;
        RECT 1561.570 1001.000 1561.830 1001.260 ;
        RECT 1815.490 1001.000 1815.750 1001.260 ;
        RECT 1821.240 1001.000 1821.500 1001.260 ;
      LAYER met2 ;
        RECT 1351.120 2917.550 1351.380 2917.870 ;
        RECT 1535.120 2917.550 1535.380 2917.870 ;
        RECT 1351.180 2912.090 1351.320 2917.550 ;
        RECT 1501.540 2917.210 1501.800 2917.530 ;
        RECT 1414.140 2916.870 1414.400 2917.190 ;
        RECT 1379.640 2914.830 1379.900 2915.150 ;
        RECT 1372.740 2913.130 1373.000 2913.450 ;
        RECT 1351.120 2911.770 1351.380 2912.090 ;
        RECT 1351.120 2911.090 1351.380 2911.410 ;
        RECT 1351.180 2850.210 1351.320 2911.090 ;
        RECT 1351.120 2849.890 1351.380 2850.210 ;
        RECT 1358.020 2849.550 1358.280 2849.870 ;
        RECT 1351.120 2849.210 1351.380 2849.530 ;
        RECT 1350.720 2843.070 1350.860 2843.225 ;
        RECT 1351.180 2843.070 1351.320 2849.210 ;
        RECT 1350.660 2842.810 1350.920 2843.070 ;
        RECT 1351.120 2842.925 1351.380 2843.070 ;
        RECT 1351.110 2842.810 1351.390 2842.925 ;
        RECT 1350.660 2842.750 1351.390 2842.810 ;
        RECT 1350.720 2842.670 1351.390 2842.750 ;
        RECT 1351.110 2842.555 1351.390 2842.670 ;
        RECT 1352.950 2842.555 1353.230 2842.925 ;
        RECT 1000.600 2810.450 1000.860 2810.770 ;
        RECT 1048.440 2810.450 1048.700 2810.770 ;
        RECT 985.420 2810.110 985.680 2810.430 ;
        RECT 978.520 2809.770 978.780 2810.090 ;
        RECT 445.840 2769.310 446.100 2769.630 ;
        RECT 796.820 2769.310 797.080 2769.630 ;
        RECT 445.900 2759.520 446.040 2769.310 ;
        RECT 532.320 2767.950 532.580 2768.270 ;
        RECT 707.120 2767.950 707.380 2768.270 ;
        RECT 518.520 2767.610 518.780 2767.930 ;
        RECT 489.080 2767.270 489.340 2767.590 ;
        RECT 489.140 2759.520 489.280 2767.270 ;
        RECT 518.580 2759.520 518.720 2767.610 ;
        RECT 532.380 2759.520 532.520 2767.950 ;
        RECT 445.730 2759.100 446.040 2759.520 ;
        RECT 488.970 2759.100 489.280 2759.520 ;
        RECT 518.410 2759.100 518.720 2759.520 ;
        RECT 532.210 2759.100 532.520 2759.520 ;
        RECT 445.730 2755.520 446.010 2759.100 ;
        RECT 488.970 2755.520 489.250 2759.100 ;
        RECT 518.410 2755.520 518.690 2759.100 ;
        RECT 532.210 2755.520 532.490 2759.100 ;
      LAYER met2 ;
        RECT 432.860 2755.240 445.450 2755.520 ;
        RECT 446.290 2755.240 460.170 2755.520 ;
        RECT 461.010 2755.240 474.890 2755.520 ;
        RECT 475.730 2755.240 488.690 2755.520 ;
        RECT 489.530 2755.240 503.410 2755.520 ;
        RECT 504.250 2755.240 518.130 2755.520 ;
        RECT 518.970 2755.240 531.930 2755.520 ;
        RECT 532.770 2755.240 546.650 2755.520 ;
        RECT 547.490 2755.240 561.370 2755.520 ;
        RECT 562.210 2755.240 575.170 2755.520 ;
      LAYER met2 ;
        RECT 420.530 2728.995 420.810 2729.365 ;
        RECT 420.070 2707.235 420.350 2707.605 ;
        RECT 420.140 1978.450 420.280 2707.235 ;
        RECT 420.600 1978.790 420.740 2728.995 ;
      LAYER met2 ;
        RECT 432.860 2604.280 575.720 2755.240 ;
      LAYER met2 ;
        RECT 588.890 2686.835 589.170 2687.205 ;
        RECT 588.960 2684.290 589.100 2686.835 ;
        RECT 588.900 2683.970 589.160 2684.290 ;
        RECT 588.890 2666.435 589.170 2666.805 ;
        RECT 588.960 2663.890 589.100 2666.435 ;
        RECT 588.900 2663.570 589.160 2663.890 ;
      LAYER met2 ;
        RECT 433.410 2604.000 446.370 2604.280 ;
        RECT 447.210 2604.000 461.090 2604.280 ;
        RECT 461.930 2604.000 475.810 2604.280 ;
        RECT 476.650 2604.000 489.610 2604.280 ;
        RECT 490.450 2604.000 504.330 2604.280 ;
        RECT 505.170 2604.000 519.050 2604.280 ;
        RECT 519.890 2604.000 532.850 2604.280 ;
        RECT 533.690 2604.000 547.570 2604.280 ;
        RECT 548.410 2604.000 562.290 2604.280 ;
        RECT 563.130 2604.000 575.720 2604.280 ;
      LAYER met2 ;
        RECT 504.610 2600.660 504.890 2604.000 ;
        RECT 533.130 2600.660 533.410 2604.000 ;
        RECT 504.610 2600.000 504.920 2600.660 ;
        RECT 533.130 2600.000 533.440 2600.660 ;
        RECT 504.780 2591.470 504.920 2600.000 ;
        RECT 533.300 2591.810 533.440 2600.000 ;
        RECT 533.240 2591.490 533.500 2591.810 ;
        RECT 504.720 2591.150 504.980 2591.470 ;
        RECT 530.020 1988.330 530.280 1988.650 ;
        RECT 650.540 1988.330 650.800 1988.650 ;
        RECT 528.450 1981.250 528.730 1981.750 ;
        RECT 530.080 1981.250 530.220 1988.330 ;
        RECT 579.240 1987.310 579.500 1987.630 ;
        RECT 638.120 1987.310 638.380 1987.630 ;
        RECT 528.450 1981.110 530.220 1981.250 ;
        RECT 578.130 1981.250 578.410 1981.750 ;
        RECT 579.300 1981.250 579.440 1987.310 ;
        RECT 578.130 1981.110 579.440 1981.250 ;
        RECT 420.540 1978.470 420.800 1978.790 ;
        RECT 420.080 1978.130 420.340 1978.450 ;
        RECT 528.450 1977.750 528.730 1981.110 ;
        RECT 578.130 1977.750 578.410 1981.110 ;
      LAYER met2 ;
        RECT 362.860 1977.470 377.290 1977.750 ;
        RECT 378.130 1977.470 402.130 1977.750 ;
        RECT 402.970 1977.470 427.890 1977.750 ;
        RECT 428.730 1977.470 452.730 1977.750 ;
        RECT 453.570 1977.470 477.570 1977.750 ;
        RECT 478.410 1977.470 502.410 1977.750 ;
        RECT 503.250 1977.470 528.170 1977.750 ;
        RECT 529.010 1977.470 553.010 1977.750 ;
        RECT 553.850 1977.470 577.850 1977.750 ;
        RECT 578.690 1977.470 602.690 1977.750 ;
        RECT 603.530 1977.470 627.530 1977.750 ;
        RECT 362.860 1704.280 628.080 1977.470 ;
        RECT 363.410 1704.000 387.410 1704.280 ;
        RECT 388.250 1704.000 412.250 1704.280 ;
        RECT 413.090 1704.000 437.090 1704.280 ;
        RECT 437.930 1704.000 461.930 1704.280 ;
        RECT 462.770 1704.000 487.690 1704.280 ;
        RECT 488.530 1704.000 512.530 1704.280 ;
        RECT 513.370 1704.000 537.370 1704.280 ;
        RECT 538.210 1704.000 562.210 1704.280 ;
        RECT 563.050 1704.000 587.970 1704.280 ;
        RECT 588.810 1704.000 612.810 1704.280 ;
        RECT 613.650 1704.000 628.080 1704.280 ;
      LAYER met2 ;
        RECT 462.210 1700.410 462.490 1704.000 ;
        RECT 512.810 1700.410 513.090 1704.000 ;
        RECT 462.210 1700.270 463.980 1700.410 ;
        RECT 462.210 1700.000 462.490 1700.270 ;
        RECT 463.840 1688.770 463.980 1700.270 ;
        RECT 512.810 1700.270 514.580 1700.410 ;
        RECT 512.810 1700.000 513.090 1700.270 ;
        RECT 514.440 1688.770 514.580 1700.270 ;
        RECT 463.780 1688.450 464.040 1688.770 ;
        RECT 468.840 1688.450 469.100 1688.770 ;
        RECT 514.380 1688.450 514.640 1688.770 ;
        RECT 517.140 1688.450 517.400 1688.770 ;
        RECT 468.900 1010.810 469.040 1688.450 ;
        RECT 517.200 1011.150 517.340 1688.450 ;
        RECT 517.140 1010.830 517.400 1011.150 ;
        RECT 468.840 1010.490 469.100 1010.810 ;
        RECT 638.180 1008.090 638.320 1987.310 ;
        RECT 638.120 1007.770 638.380 1008.090 ;
        RECT 650.600 1007.750 650.740 1988.330 ;
        RECT 707.180 1012.170 707.320 2767.950 ;
        RECT 755.420 2767.610 755.680 2767.930 ;
        RECT 720.920 2683.970 721.180 2684.290 ;
        RECT 707.120 1011.850 707.380 1012.170 ;
        RECT 712.640 1010.830 712.900 1011.150 ;
        RECT 673.540 1010.490 673.800 1010.810 ;
        RECT 669.860 1007.770 670.120 1008.090 ;
        RECT 650.540 1007.430 650.800 1007.750 ;
        RECT 669.920 1000.010 670.060 1007.770 ;
        RECT 671.700 1007.430 671.960 1007.750 ;
        RECT 671.760 1000.010 671.900 1007.430 ;
        RECT 673.600 1000.010 673.740 1010.490 ;
        RECT 712.700 1000.010 712.840 1010.830 ;
        RECT 720.980 1010.810 721.120 2683.970 ;
        RECT 755.480 1011.150 755.620 2767.610 ;
        RECT 769.220 2767.270 769.480 2767.590 ;
        RECT 762.320 2591.490 762.580 2591.810 ;
        RECT 762.380 1011.490 762.520 2591.490 ;
        RECT 769.280 1011.830 769.420 2767.270 ;
        RECT 789.920 2663.570 790.180 2663.890 ;
        RECT 783.020 2591.150 783.280 2591.470 ;
        RECT 783.080 1012.510 783.220 2591.150 ;
        RECT 789.980 1013.190 790.120 2663.570 ;
        RECT 789.920 1012.870 790.180 1013.190 ;
        RECT 796.880 1012.850 797.020 2769.310 ;
        RECT 978.060 2643.850 978.320 2644.170 ;
        RECT 975.300 2604.410 975.560 2604.730 ;
        RECT 974.840 2591.150 975.100 2591.470 ;
        RECT 972.540 2045.790 972.800 2046.110 ;
        RECT 965.640 2045.450 965.900 2045.770 ;
        RECT 842.820 1977.790 843.080 1978.110 ;
        RECT 796.820 1012.530 797.080 1012.850 ;
        RECT 783.020 1012.190 783.280 1012.510 ;
        RECT 841.900 1011.850 842.160 1012.170 ;
        RECT 769.220 1011.510 769.480 1011.830 ;
        RECT 762.320 1011.170 762.580 1011.490 ;
        RECT 755.420 1010.830 755.680 1011.150 ;
        RECT 720.920 1010.490 721.180 1010.810 ;
        RECT 841.960 1000.010 842.100 1011.850 ;
        RECT 842.880 1000.010 843.020 1977.790 ;
        RECT 897.560 1977.450 897.820 1977.770 ;
        RECT 888.360 1012.870 888.620 1013.190 ;
        RECT 844.660 1012.530 844.920 1012.850 ;
        RECT 844.720 1000.010 844.860 1012.530 ;
        RECT 884.220 1012.190 884.480 1012.510 ;
        RECT 884.280 1000.010 884.420 1012.190 ;
        RECT 888.420 1000.010 888.560 1012.870 ;
        RECT 892.500 1010.490 892.760 1010.810 ;
        RECT 892.560 1000.010 892.700 1010.490 ;
        RECT 897.620 1000.010 897.760 1977.450 ;
        RECT 965.700 1024.750 965.840 2045.450 ;
        RECT 972.600 1025.090 972.740 2045.790 ;
        RECT 974.900 1694.890 975.040 2591.150 ;
        RECT 974.840 1694.570 975.100 1694.890 ;
        RECT 975.360 1693.870 975.500 2604.410 ;
        RECT 977.140 2050.550 977.400 2050.870 ;
        RECT 976.220 2047.830 976.480 2048.150 ;
        RECT 975.760 2046.810 976.020 2047.130 ;
        RECT 975.300 1693.550 975.560 1693.870 ;
        RECT 975.820 1025.430 975.960 2046.810 ;
        RECT 975.760 1025.110 976.020 1025.430 ;
        RECT 972.540 1024.770 972.800 1025.090 ;
        RECT 965.640 1024.430 965.900 1024.750 ;
        RECT 976.280 1011.830 976.420 2047.830 ;
        RECT 976.680 2046.130 976.940 2046.450 ;
        RECT 910.900 1011.510 911.160 1011.830 ;
        RECT 976.220 1011.510 976.480 1011.830 ;
        RECT 905.380 1011.170 905.640 1011.490 ;
        RECT 901.240 1010.830 901.500 1011.150 ;
        RECT 901.300 1000.010 901.440 1010.830 ;
        RECT 905.440 1000.010 905.580 1011.170 ;
        RECT 910.960 1001.970 911.100 1011.510 ;
        RECT 976.740 1010.130 976.880 2046.130 ;
        RECT 977.200 1013.870 977.340 2050.550 ;
        RECT 977.600 2050.210 977.860 2050.530 ;
        RECT 977.140 1013.550 977.400 1013.870 ;
        RECT 977.660 1012.850 977.800 2050.210 ;
        RECT 977.600 1012.530 977.860 1012.850 ;
        RECT 976.680 1009.810 976.940 1010.130 ;
        RECT 978.120 1009.790 978.260 2643.850 ;
        RECT 978.580 1012.365 978.720 2809.770 ;
        RECT 978.980 2809.430 979.240 2809.750 ;
        RECT 979.040 1014.405 979.180 2809.430 ;
        RECT 979.440 2808.750 979.700 2809.070 ;
        RECT 978.970 1014.035 979.250 1014.405 ;
        RECT 978.510 1011.995 978.790 1012.365 ;
        RECT 979.500 1011.685 979.640 2808.750 ;
        RECT 982.200 2604.750 982.460 2605.070 ;
        RECT 982.260 1694.210 982.400 2604.750 ;
        RECT 984.960 2591.490 985.220 2591.810 ;
        RECT 984.040 2049.870 984.300 2050.190 ;
        RECT 983.120 2047.490 983.380 2047.810 ;
        RECT 982.660 2047.150 982.920 2047.470 ;
        RECT 982.200 1693.890 982.460 1694.210 ;
        RECT 982.720 1025.770 982.860 2047.150 ;
        RECT 982.660 1025.450 982.920 1025.770 ;
        RECT 983.180 1013.190 983.320 2047.490 ;
        RECT 983.580 2046.470 983.840 2046.790 ;
        RECT 983.120 1012.870 983.380 1013.190 ;
        RECT 979.430 1011.315 979.710 1011.685 ;
        RECT 983.640 1010.470 983.780 2046.470 ;
        RECT 984.100 1012.170 984.240 2049.870 ;
        RECT 984.500 2049.190 984.760 2049.510 ;
        RECT 984.560 1013.530 984.700 2049.190 ;
        RECT 984.500 1013.210 984.760 1013.530 ;
        RECT 984.040 1011.850 984.300 1012.170 ;
        RECT 983.580 1010.150 983.840 1010.470 ;
        RECT 978.060 1009.470 978.320 1009.790 ;
        RECT 985.020 1009.450 985.160 2591.490 ;
        RECT 985.480 1013.045 985.620 2810.110 ;
        RECT 985.880 2809.090 986.140 2809.410 ;
        RECT 985.410 1012.675 985.690 1013.045 ;
        RECT 985.940 1010.325 986.080 2809.090 ;
        RECT 1000.660 2809.070 1000.800 2810.450 ;
        RECT 1027.740 2809.770 1028.000 2810.090 ;
        RECT 1000.600 2808.750 1000.860 2809.070 ;
        RECT 986.340 2800.930 986.600 2801.250 ;
        RECT 1010.260 2800.930 1010.520 2801.250 ;
        RECT 986.400 1011.005 986.540 2800.930 ;
        RECT 1010.320 2799.970 1010.460 2800.930 ;
        RECT 1027.800 2800.000 1027.940 2809.770 ;
        RECT 1043.380 2809.430 1043.640 2809.750 ;
        RECT 1043.440 2800.000 1043.580 2809.430 ;
        RECT 1048.500 2808.730 1048.640 2810.450 ;
        RECT 1073.740 2810.110 1074.000 2810.430 ;
        RECT 1058.100 2809.090 1058.360 2809.410 ;
        RECT 1048.440 2808.410 1048.700 2808.730 ;
        RECT 1058.160 2800.000 1058.300 2809.090 ;
        RECT 1073.800 2800.000 1073.940 2810.110 ;
        RECT 1089.380 2808.410 1089.640 2808.730 ;
        RECT 1089.440 2800.000 1089.580 2808.410 ;
        RECT 1012.050 2799.970 1012.330 2800.000 ;
        RECT 1010.320 2799.830 1012.330 2799.970 ;
        RECT 1012.050 2796.000 1012.330 2799.830 ;
        RECT 1027.690 2796.000 1027.970 2800.000 ;
        RECT 1043.330 2796.000 1043.610 2800.000 ;
        RECT 1058.050 2796.000 1058.330 2800.000 ;
        RECT 1073.690 2796.000 1073.970 2800.000 ;
        RECT 1089.330 2796.000 1089.610 2800.000 ;
      LAYER met2 ;
        RECT 1002.860 2795.720 1011.770 2796.000 ;
        RECT 1012.610 2795.720 1027.410 2796.000 ;
        RECT 1028.250 2795.720 1043.050 2796.000 ;
        RECT 1043.890 2795.720 1057.770 2796.000 ;
        RECT 1058.610 2795.720 1073.410 2796.000 ;
        RECT 1074.250 2795.720 1089.050 2796.000 ;
        RECT 1089.890 2795.720 1095.120 2796.000 ;
      LAYER met2 ;
        RECT 993.230 2783.395 993.510 2783.765 ;
        RECT 992.770 2739.195 993.050 2739.565 ;
        RECT 992.310 2718.795 992.590 2719.165 ;
        RECT 987.250 2646.035 987.530 2646.405 ;
        RECT 987.320 2644.170 987.460 2646.035 ;
        RECT 987.260 2643.850 987.520 2644.170 ;
        RECT 991.850 2622.915 992.130 2623.285 ;
        RECT 991.390 1955.835 991.670 1956.205 ;
        RECT 990.930 1935.435 991.210 1935.805 ;
        RECT 990.470 1893.275 990.750 1893.645 ;
        RECT 990.010 1871.515 990.290 1871.885 ;
        RECT 989.550 1851.115 989.830 1851.485 ;
        RECT 989.090 1808.955 989.370 1809.325 ;
        RECT 988.630 1787.195 988.910 1787.565 ;
        RECT 988.170 1766.795 988.450 1767.165 ;
        RECT 987.710 1745.035 987.990 1745.405 ;
        RECT 987.780 1020.330 987.920 1745.035 ;
        RECT 987.720 1020.010 987.980 1020.330 ;
        RECT 988.240 1018.970 988.380 1766.795 ;
        RECT 988.700 1021.010 988.840 1787.195 ;
        RECT 988.640 1020.690 988.900 1021.010 ;
        RECT 989.160 1019.650 989.300 1808.955 ;
        RECT 989.100 1019.330 989.360 1019.650 ;
        RECT 988.180 1018.650 988.440 1018.970 ;
        RECT 989.620 1018.630 989.760 1851.115 ;
        RECT 989.560 1018.310 989.820 1018.630 ;
        RECT 990.080 1017.950 990.220 1871.515 ;
        RECT 990.540 1019.310 990.680 1893.275 ;
        RECT 990.480 1018.990 990.740 1019.310 ;
        RECT 991.000 1018.290 991.140 1935.435 ;
        RECT 990.940 1017.970 991.200 1018.290 ;
        RECT 990.020 1017.630 990.280 1017.950 ;
        RECT 991.460 1017.610 991.600 1955.835 ;
        RECT 991.400 1017.290 991.660 1017.610 ;
        RECT 986.330 1010.635 986.610 1011.005 ;
        RECT 985.870 1009.955 986.150 1010.325 ;
        RECT 984.960 1009.130 985.220 1009.450 ;
        RECT 991.920 1009.110 992.060 2622.915 ;
        RECT 991.860 1008.790 992.120 1009.110 ;
        RECT 992.380 1007.750 992.520 2718.795 ;
        RECT 992.840 1017.270 992.980 2739.195 ;
        RECT 992.780 1016.950 993.040 1017.270 ;
        RECT 993.300 1009.645 993.440 2783.395 ;
        RECT 993.690 2760.275 993.970 2760.645 ;
        RECT 993.760 1052.290 993.900 2760.275 ;
        RECT 994.150 2692.275 994.430 2692.645 ;
        RECT 993.700 1051.970 993.960 1052.290 ;
        RECT 994.220 1013.725 994.360 2692.275 ;
        RECT 994.610 2670.515 994.890 2670.885 ;
        RECT 994.150 1013.355 994.430 1013.725 ;
        RECT 993.230 1009.275 993.510 1009.645 ;
        RECT 994.680 1008.090 994.820 2670.515 ;
        RECT 999.220 2605.430 999.480 2605.750 ;
        RECT 995.070 2018.395 995.350 2018.765 ;
        RECT 995.140 1011.150 995.280 2018.395 ;
        RECT 995.530 1997.995 995.810 1998.365 ;
        RECT 995.080 1010.830 995.340 1011.150 ;
        RECT 995.600 1010.810 995.740 1997.995 ;
        RECT 995.990 1976.235 996.270 1976.605 ;
        RECT 996.060 1011.490 996.200 1976.235 ;
        RECT 996.450 1913.675 996.730 1914.045 ;
        RECT 996.520 1019.990 996.660 1913.675 ;
        RECT 996.910 1829.355 997.190 1829.725 ;
        RECT 996.980 1020.670 997.120 1829.355 ;
        RECT 997.370 1724.635 997.650 1725.005 ;
        RECT 997.440 1021.350 997.580 1724.635 ;
        RECT 998.760 1713.270 999.020 1713.590 ;
        RECT 997.380 1021.030 997.640 1021.350 ;
        RECT 996.920 1020.350 997.180 1020.670 ;
        RECT 996.460 1019.670 996.720 1019.990 ;
        RECT 996.000 1011.170 996.260 1011.490 ;
        RECT 995.540 1010.490 995.800 1010.810 ;
        RECT 998.820 1008.430 998.960 1713.270 ;
        RECT 999.280 1695.230 999.420 2605.430 ;
        RECT 999.680 2605.090 999.940 2605.410 ;
        RECT 999.220 1694.910 999.480 1695.230 ;
        RECT 999.740 1694.550 999.880 2605.090 ;
      LAYER met2 ;
        RECT 1002.860 2604.280 1095.120 2795.720 ;
      LAYER met2 ;
        RECT 1353.020 2795.130 1353.160 2842.555 ;
        RECT 1351.580 2794.810 1351.840 2795.130 ;
        RECT 1352.960 2794.810 1353.220 2795.130 ;
        RECT 1110.990 2780.675 1111.270 2781.045 ;
        RECT 1097.190 2644.675 1097.470 2645.045 ;
      LAYER met2 ;
        RECT 1003.410 2604.000 1017.290 2604.280 ;
        RECT 1018.130 2604.000 1032.930 2604.280 ;
        RECT 1033.770 2604.000 1048.570 2604.280 ;
        RECT 1049.410 2604.000 1064.210 2604.280 ;
        RECT 1065.050 2604.000 1079.850 2604.280 ;
        RECT 1080.690 2604.000 1094.570 2604.280 ;
      LAYER met2 ;
        RECT 1002.850 2600.730 1003.130 2604.000 ;
        RECT 1017.570 2600.730 1017.850 2604.000 ;
        RECT 1001.120 2600.590 1003.130 2600.730 ;
        RECT 1000.140 2049.530 1000.400 2049.850 ;
        RECT 999.680 1694.230 999.940 1694.550 ;
        RECT 1000.200 1012.510 1000.340 2049.530 ;
        RECT 1001.120 1713.590 1001.260 2600.590 ;
        RECT 1002.850 2600.000 1003.130 2600.590 ;
        RECT 1014.460 2600.590 1017.850 2600.730 ;
        RECT 1002.900 2049.190 1003.160 2049.510 ;
        RECT 1002.960 2044.110 1003.100 2049.190 ;
        RECT 1014.460 2048.150 1014.600 2600.590 ;
        RECT 1017.570 2600.000 1017.850 2600.590 ;
        RECT 1033.210 2600.000 1033.490 2604.000 ;
        RECT 1048.850 2600.000 1049.130 2604.000 ;
        RECT 1064.490 2600.730 1064.770 2604.000 ;
        RECT 1080.130 2600.730 1080.410 2604.000 ;
        RECT 1062.760 2600.590 1064.770 2600.730 ;
        RECT 1033.320 2587.730 1033.460 2600.000 ;
        RECT 1048.960 2591.810 1049.100 2600.000 ;
        RECT 1048.900 2591.490 1049.160 2591.810 ;
        RECT 1028.200 2587.410 1028.460 2587.730 ;
        RECT 1033.260 2587.410 1033.520 2587.730 ;
        RECT 1016.700 2052.590 1016.960 2052.910 ;
        RECT 1014.400 2047.830 1014.660 2048.150 ;
        RECT 1016.760 2044.110 1016.900 2052.590 ;
        RECT 1028.260 2047.810 1028.400 2587.410 ;
        RECT 1059.940 2053.270 1060.200 2053.590 ;
        RECT 1031.420 2052.930 1031.680 2053.250 ;
        RECT 1028.200 2047.490 1028.460 2047.810 ;
        RECT 1031.480 2044.110 1031.620 2052.930 ;
        RECT 1045.220 2049.530 1045.480 2049.850 ;
        RECT 1045.280 2044.110 1045.420 2049.530 ;
        RECT 1060.000 2044.110 1060.140 2053.270 ;
        RECT 1062.760 2047.470 1062.900 2600.590 ;
        RECT 1064.490 2600.000 1064.770 2600.590 ;
        RECT 1076.560 2600.590 1080.410 2600.730 ;
        RECT 1073.740 2049.870 1074.000 2050.190 ;
        RECT 1062.700 2047.150 1062.960 2047.470 ;
        RECT 1073.800 2044.110 1073.940 2049.870 ;
        RECT 1076.560 2047.130 1076.700 2600.590 ;
        RECT 1080.130 2600.000 1080.410 2600.590 ;
        RECT 1094.850 2600.000 1095.130 2604.000 ;
        RECT 1094.960 2591.470 1095.100 2600.000 ;
        RECT 1094.900 2591.150 1095.160 2591.470 ;
        RECT 1088.460 2050.550 1088.720 2050.870 ;
        RECT 1076.500 2046.810 1076.760 2047.130 ;
        RECT 1088.520 2044.110 1088.660 2050.550 ;
        RECT 1097.260 2046.450 1097.400 2644.675 ;
        RECT 1097.650 2622.235 1097.930 2622.605 ;
        RECT 1097.720 2046.790 1097.860 2622.235 ;
        RECT 1102.260 2050.210 1102.520 2050.530 ;
        RECT 1097.660 2046.470 1097.920 2046.790 ;
        RECT 1097.200 2046.130 1097.460 2046.450 ;
        RECT 1102.320 2044.110 1102.460 2050.210 ;
        RECT 1111.060 2045.770 1111.200 2780.675 ;
        RECT 1351.640 2767.590 1351.780 2794.810 ;
        RECT 1351.580 2767.270 1351.840 2767.590 ;
        RECT 1351.120 2766.590 1351.380 2766.910 ;
        RECT 1111.450 2760.275 1111.730 2760.645 ;
        RECT 1111.520 2046.110 1111.660 2760.275 ;
        RECT 1351.180 2739.370 1351.320 2766.590 ;
        RECT 1350.660 2739.050 1350.920 2739.370 ;
        RECT 1351.120 2739.050 1351.380 2739.370 ;
        RECT 1111.910 2734.435 1112.190 2734.805 ;
        RECT 1111.980 2605.750 1112.120 2734.435 ;
        RECT 1112.370 2712.675 1112.650 2713.045 ;
        RECT 1111.920 2605.430 1112.180 2605.750 ;
        RECT 1112.440 2604.730 1112.580 2712.675 ;
        RECT 1112.830 2691.595 1113.110 2691.965 ;
        RECT 1112.900 2605.410 1113.040 2691.595 ;
        RECT 1350.720 2691.430 1350.860 2739.050 ;
        RECT 1350.200 2691.110 1350.460 2691.430 ;
        RECT 1350.660 2691.110 1350.920 2691.430 ;
        RECT 1350.260 2670.350 1350.400 2691.110 ;
        RECT 1350.200 2670.030 1350.460 2670.350 ;
        RECT 1351.120 2670.030 1351.380 2670.350 ;
        RECT 1113.290 2666.435 1113.570 2666.805 ;
        RECT 1112.840 2605.090 1113.100 2605.410 ;
        RECT 1113.360 2605.070 1113.500 2666.435 ;
        RECT 1351.180 2622.750 1351.320 2670.030 ;
        RECT 1351.120 2622.430 1351.380 2622.750 ;
        RECT 1351.120 2621.750 1351.380 2622.070 ;
        RECT 1113.300 2604.750 1113.560 2605.070 ;
        RECT 1112.380 2604.410 1112.640 2604.730 ;
        RECT 1351.180 2601.525 1351.320 2621.750 ;
        RECT 1350.190 2601.155 1350.470 2601.525 ;
        RECT 1351.110 2601.155 1351.390 2601.525 ;
        RECT 1350.260 2573.530 1350.400 2601.155 ;
        RECT 1350.260 2573.390 1351.780 2573.530 ;
        RECT 1351.640 2560.045 1351.780 2573.390 ;
        RECT 1351.570 2559.675 1351.850 2560.045 ;
        RECT 1350.190 2558.995 1350.470 2559.365 ;
        RECT 1350.260 2511.910 1350.400 2558.995 ;
        RECT 1350.200 2511.590 1350.460 2511.910 ;
        RECT 1352.040 2511.590 1352.300 2511.910 ;
        RECT 1352.100 2463.485 1352.240 2511.590 ;
        RECT 1351.110 2463.115 1351.390 2463.485 ;
        RECT 1352.030 2463.115 1352.310 2463.485 ;
        RECT 1351.180 2429.630 1351.320 2463.115 ;
        RECT 1351.120 2429.310 1351.380 2429.630 ;
        RECT 1351.120 2428.630 1351.380 2428.950 ;
        RECT 1351.180 2380.670 1351.320 2428.630 ;
        RECT 1351.120 2380.350 1351.380 2380.670 ;
        RECT 1351.580 2380.350 1351.840 2380.670 ;
        RECT 1351.640 2367.070 1351.780 2380.350 ;
        RECT 1351.120 2366.750 1351.380 2367.070 ;
        RECT 1351.580 2366.750 1351.840 2367.070 ;
        RECT 1351.180 2332.730 1351.320 2366.750 ;
        RECT 1351.120 2332.410 1351.380 2332.730 ;
        RECT 1351.120 2331.730 1351.380 2332.050 ;
        RECT 1351.180 2294.310 1351.320 2331.730 ;
        RECT 1350.200 2293.990 1350.460 2294.310 ;
        RECT 1351.120 2293.990 1351.380 2294.310 ;
        RECT 1350.260 2270.365 1350.400 2293.990 ;
        RECT 1350.190 2269.995 1350.470 2270.365 ;
        RECT 1351.110 2269.995 1351.390 2270.365 ;
        RECT 1351.180 2236.170 1351.320 2269.995 ;
        RECT 1351.120 2235.850 1351.380 2236.170 ;
        RECT 1351.120 2235.170 1351.380 2235.490 ;
        RECT 1351.180 2197.750 1351.320 2235.170 ;
        RECT 1350.200 2197.430 1350.460 2197.750 ;
        RECT 1351.120 2197.430 1351.380 2197.750 ;
        RECT 1350.260 2173.805 1350.400 2197.430 ;
        RECT 1350.190 2173.435 1350.470 2173.805 ;
        RECT 1351.110 2173.435 1351.390 2173.805 ;
        RECT 1351.180 2139.610 1351.320 2173.435 ;
        RECT 1351.120 2139.290 1351.380 2139.610 ;
        RECT 1351.120 2138.610 1351.380 2138.930 ;
        RECT 1351.180 2125.330 1351.320 2138.610 ;
        RECT 1350.660 2125.010 1350.920 2125.330 ;
        RECT 1351.120 2125.010 1351.380 2125.330 ;
        RECT 1350.720 2090.650 1350.860 2125.010 ;
        RECT 1350.660 2090.330 1350.920 2090.650 ;
        RECT 1351.580 2090.330 1351.840 2090.650 ;
        RECT 1351.640 2077.130 1351.780 2090.330 ;
        RECT 1351.640 2076.990 1352.240 2077.130 ;
        RECT 1244.860 2055.310 1245.120 2055.630 ;
        RECT 1346.060 2055.310 1346.320 2055.630 ;
        RECT 1230.140 2054.630 1230.400 2054.950 ;
        RECT 1116.980 2054.290 1117.240 2054.610 ;
        RECT 1111.460 2045.790 1111.720 2046.110 ;
        RECT 1111.000 2045.450 1111.260 2045.770 ;
        RECT 1117.040 2044.110 1117.180 2054.290 ;
        RECT 1130.780 2053.950 1131.040 2054.270 ;
        RECT 1130.840 2044.110 1130.980 2053.950 ;
        RECT 1216.340 2053.610 1216.600 2053.930 ;
        RECT 1201.620 2052.250 1201.880 2052.570 ;
        RECT 1187.820 2051.910 1188.080 2052.230 ;
        RECT 1173.100 2051.570 1173.360 2051.890 ;
        RECT 1159.300 2051.230 1159.560 2051.550 ;
        RECT 1144.580 2050.890 1144.840 2051.210 ;
        RECT 1144.640 2044.110 1144.780 2050.890 ;
        RECT 1159.360 2044.110 1159.500 2051.230 ;
        RECT 1173.160 2044.110 1173.300 2051.570 ;
        RECT 1187.880 2044.110 1188.020 2051.910 ;
        RECT 1201.680 2044.110 1201.820 2052.250 ;
        RECT 1216.400 2044.110 1216.540 2053.610 ;
        RECT 1230.200 2044.110 1230.340 2054.630 ;
        RECT 1244.920 2044.110 1245.060 2055.310 ;
        RECT 1287.180 2054.970 1287.440 2055.290 ;
        RECT 1273.380 2050.550 1273.640 2050.870 ;
        RECT 1258.660 2050.210 1258.920 2050.530 ;
        RECT 1258.720 2044.110 1258.860 2050.210 ;
        RECT 1273.440 2044.110 1273.580 2050.550 ;
        RECT 1287.240 2044.110 1287.380 2054.970 ;
        RECT 1335.480 2054.630 1335.740 2054.950 ;
        RECT 1332.720 2054.290 1332.980 2054.610 ;
        RECT 1301.900 2049.530 1302.160 2049.850 ;
        RECT 1301.960 2044.110 1302.100 2049.530 ;
        RECT 1315.700 2049.190 1315.960 2049.510 ;
        RECT 1315.760 2044.110 1315.900 2049.190 ;
        RECT 1002.850 2040.110 1003.130 2044.110 ;
        RECT 1016.650 2040.110 1016.930 2044.110 ;
        RECT 1031.370 2040.110 1031.650 2044.110 ;
        RECT 1045.170 2040.110 1045.450 2044.110 ;
        RECT 1059.890 2040.110 1060.170 2044.110 ;
        RECT 1073.690 2040.110 1073.970 2044.110 ;
        RECT 1088.410 2040.110 1088.690 2044.110 ;
        RECT 1102.210 2040.110 1102.490 2044.110 ;
        RECT 1116.930 2040.110 1117.210 2044.110 ;
        RECT 1130.730 2040.110 1131.010 2044.110 ;
        RECT 1144.530 2040.110 1144.810 2044.110 ;
        RECT 1159.250 2040.110 1159.530 2044.110 ;
        RECT 1173.050 2040.110 1173.330 2044.110 ;
        RECT 1187.770 2040.110 1188.050 2044.110 ;
        RECT 1201.570 2040.110 1201.850 2044.110 ;
        RECT 1216.290 2040.110 1216.570 2044.110 ;
        RECT 1230.090 2040.110 1230.370 2044.110 ;
        RECT 1244.810 2040.110 1245.090 2044.110 ;
        RECT 1258.610 2040.110 1258.890 2044.110 ;
        RECT 1273.330 2040.110 1273.610 2044.110 ;
        RECT 1287.130 2040.110 1287.410 2044.110 ;
        RECT 1301.850 2040.110 1302.130 2044.110 ;
        RECT 1315.650 2040.110 1315.930 2044.110 ;
        RECT 1329.450 2040.410 1329.730 2044.110 ;
        RECT 1329.450 2040.270 1331.080 2040.410 ;
        RECT 1329.450 2040.110 1329.730 2040.270 ;
      LAYER met2 ;
        RECT 1003.410 2039.830 1016.370 2040.110 ;
        RECT 1017.210 2039.830 1031.090 2040.110 ;
        RECT 1031.930 2039.830 1044.890 2040.110 ;
        RECT 1045.730 2039.830 1059.610 2040.110 ;
        RECT 1060.450 2039.830 1073.410 2040.110 ;
        RECT 1074.250 2039.830 1088.130 2040.110 ;
        RECT 1088.970 2039.830 1101.930 2040.110 ;
        RECT 1102.770 2039.830 1116.650 2040.110 ;
        RECT 1117.490 2039.830 1130.450 2040.110 ;
        RECT 1131.290 2039.830 1144.250 2040.110 ;
        RECT 1145.090 2039.830 1158.970 2040.110 ;
        RECT 1159.810 2039.830 1172.770 2040.110 ;
        RECT 1173.610 2039.830 1187.490 2040.110 ;
        RECT 1188.330 2039.830 1201.290 2040.110 ;
        RECT 1202.130 2039.830 1216.010 2040.110 ;
        RECT 1216.850 2039.830 1229.810 2040.110 ;
        RECT 1230.650 2039.830 1244.530 2040.110 ;
        RECT 1245.370 2039.830 1258.330 2040.110 ;
        RECT 1259.170 2039.830 1273.050 2040.110 ;
        RECT 1273.890 2039.830 1286.850 2040.110 ;
        RECT 1287.690 2039.830 1301.570 2040.110 ;
        RECT 1302.410 2039.830 1315.370 2040.110 ;
        RECT 1316.210 2039.830 1329.170 2040.110 ;
      LAYER met2 ;
        RECT 1001.060 1713.270 1001.320 1713.590 ;
      LAYER met2 ;
        RECT 1002.860 1704.280 1329.720 2039.830 ;
      LAYER met2 ;
        RECT 1330.940 2036.590 1331.080 2040.270 ;
        RECT 1330.880 2036.270 1331.140 2036.590 ;
      LAYER met2 ;
        RECT 1003.410 1704.000 1016.370 1704.280 ;
        RECT 1017.210 1704.000 1030.170 1704.280 ;
        RECT 1031.010 1704.000 1044.890 1704.280 ;
        RECT 1045.730 1704.000 1058.690 1704.280 ;
        RECT 1059.530 1704.000 1073.410 1704.280 ;
        RECT 1074.250 1704.000 1087.210 1704.280 ;
        RECT 1088.050 1704.000 1101.930 1704.280 ;
        RECT 1102.770 1704.000 1115.730 1704.280 ;
        RECT 1116.570 1704.000 1130.450 1704.280 ;
        RECT 1131.290 1704.000 1144.250 1704.280 ;
        RECT 1145.090 1704.000 1158.970 1704.280 ;
        RECT 1159.810 1704.000 1172.770 1704.280 ;
        RECT 1173.610 1704.000 1187.490 1704.280 ;
        RECT 1188.330 1704.000 1201.290 1704.280 ;
        RECT 1202.130 1704.000 1215.090 1704.280 ;
        RECT 1215.930 1704.000 1229.810 1704.280 ;
        RECT 1230.650 1704.000 1243.610 1704.280 ;
        RECT 1244.450 1704.000 1258.330 1704.280 ;
        RECT 1259.170 1704.000 1272.130 1704.280 ;
        RECT 1272.970 1704.000 1286.850 1704.280 ;
        RECT 1287.690 1704.000 1300.650 1704.280 ;
        RECT 1301.490 1704.000 1315.370 1704.280 ;
        RECT 1316.210 1704.000 1329.170 1704.280 ;
      LAYER met2 ;
        RECT 1002.850 1700.000 1003.130 1704.000 ;
        RECT 1016.650 1700.000 1016.930 1704.000 ;
        RECT 1030.450 1700.000 1030.730 1704.000 ;
        RECT 1045.170 1700.410 1045.450 1704.000 ;
        RECT 1058.970 1700.410 1059.250 1704.000 ;
        RECT 1045.170 1700.270 1048.640 1700.410 ;
        RECT 1045.170 1700.000 1045.450 1700.270 ;
        RECT 1002.960 1685.710 1003.100 1700.000 ;
        RECT 1002.900 1685.390 1003.160 1685.710 ;
        RECT 1016.760 1684.350 1016.900 1700.000 ;
        RECT 1030.560 1688.430 1030.700 1700.000 ;
        RECT 1030.500 1688.110 1030.760 1688.430 ;
        RECT 1038.320 1685.390 1038.580 1685.710 ;
        RECT 1016.700 1684.030 1016.960 1684.350 ;
        RECT 1020.840 1684.030 1021.100 1684.350 ;
        RECT 1020.900 1013.190 1021.040 1684.030 ;
        RECT 1012.560 1012.870 1012.820 1013.190 ;
        RECT 1020.840 1012.870 1021.100 1013.190 ;
        RECT 1000.140 1012.190 1000.400 1012.510 ;
        RECT 1003.820 1011.510 1004.080 1011.830 ;
        RECT 1003.880 1008.770 1004.020 1011.510 ;
        RECT 1012.620 1009.450 1012.760 1012.870 ;
        RECT 1038.380 1011.830 1038.520 1685.390 ;
        RECT 1048.500 1014.210 1048.640 1700.270 ;
        RECT 1058.970 1700.270 1062.440 1700.410 ;
        RECT 1058.970 1700.000 1059.250 1700.270 ;
        RECT 1048.900 1694.570 1049.160 1694.890 ;
        RECT 1048.440 1013.890 1048.700 1014.210 ;
        RECT 1038.320 1011.510 1038.580 1011.830 ;
        RECT 1012.560 1009.130 1012.820 1009.450 ;
        RECT 1011.640 1008.790 1011.900 1009.110 ;
        RECT 1003.820 1008.450 1004.080 1008.770 ;
        RECT 998.760 1008.110 999.020 1008.430 ;
        RECT 994.620 1007.770 994.880 1008.090 ;
        RECT 992.320 1007.430 992.580 1007.750 ;
        RECT 910.900 1001.650 911.160 1001.970 ;
        RECT 912.280 1001.650 912.540 1001.970 ;
        RECT 669.920 1000.000 671.140 1000.010 ;
        RECT 671.760 1000.000 672.980 1000.010 ;
        RECT 673.600 1000.000 675.280 1000.010 ;
        RECT 712.700 1000.000 714.380 1000.010 ;
        RECT 841.960 1000.000 842.260 1000.010 ;
        RECT 842.880 1000.000 844.100 1000.010 ;
        RECT 844.720 1000.000 846.400 1000.010 ;
        RECT 884.280 1000.000 885.500 1000.010 ;
        RECT 888.420 1000.000 889.640 1000.010 ;
        RECT 892.560 1000.000 894.240 1000.010 ;
        RECT 897.620 1000.000 898.380 1000.010 ;
        RECT 901.300 1000.000 902.980 1000.010 ;
        RECT 905.440 1000.000 907.120 1000.010 ;
        RECT 669.920 999.870 671.290 1000.000 ;
        RECT 671.760 999.870 673.130 1000.000 ;
        RECT 673.600 999.870 675.430 1000.000 ;
      LAYER met2 ;
        RECT 670.100 995.720 670.730 998.470 ;
      LAYER met2 ;
        RECT 671.010 996.000 671.290 999.870 ;
      LAYER met2 ;
        RECT 671.570 995.720 672.570 998.470 ;
      LAYER met2 ;
        RECT 672.850 996.000 673.130 999.870 ;
      LAYER met2 ;
        RECT 673.410 995.720 674.870 998.470 ;
      LAYER met2 ;
        RECT 675.150 996.000 675.430 999.870 ;
      LAYER met2 ;
        RECT 675.710 995.720 677.170 998.470 ;
      LAYER met2 ;
        RECT 677.450 996.000 677.730 1000.000 ;
      LAYER met2 ;
        RECT 678.010 995.720 679.010 998.470 ;
      LAYER met2 ;
        RECT 679.290 996.000 679.570 1000.000 ;
      LAYER met2 ;
        RECT 679.850 995.720 681.310 998.470 ;
      LAYER met2 ;
        RECT 681.590 996.000 681.870 1000.000 ;
      LAYER met2 ;
        RECT 682.150 995.720 683.610 998.470 ;
      LAYER met2 ;
        RECT 683.890 996.000 684.170 1000.000 ;
      LAYER met2 ;
        RECT 684.450 995.720 685.450 998.470 ;
      LAYER met2 ;
        RECT 685.730 996.000 686.010 1000.000 ;
      LAYER met2 ;
        RECT 686.290 995.720 687.750 998.470 ;
      LAYER met2 ;
        RECT 688.030 996.000 688.310 1000.000 ;
      LAYER met2 ;
        RECT 688.590 995.720 690.050 998.470 ;
      LAYER met2 ;
        RECT 690.330 996.000 690.610 1000.000 ;
      LAYER met2 ;
        RECT 690.890 995.720 692.350 998.470 ;
      LAYER met2 ;
        RECT 692.630 996.000 692.910 1000.000 ;
      LAYER met2 ;
        RECT 693.190 995.720 694.190 998.470 ;
      LAYER met2 ;
        RECT 694.470 996.000 694.750 1000.000 ;
      LAYER met2 ;
        RECT 695.030 995.720 696.490 998.470 ;
      LAYER met2 ;
        RECT 696.770 996.000 697.050 1000.000 ;
      LAYER met2 ;
        RECT 697.330 995.720 698.790 998.470 ;
      LAYER met2 ;
        RECT 699.070 996.000 699.350 1000.000 ;
      LAYER met2 ;
        RECT 699.630 995.720 700.630 998.470 ;
      LAYER met2 ;
        RECT 700.910 996.000 701.190 1000.000 ;
      LAYER met2 ;
        RECT 701.470 995.720 702.930 998.470 ;
      LAYER met2 ;
        RECT 703.210 996.000 703.490 1000.000 ;
      LAYER met2 ;
        RECT 703.770 995.720 705.230 998.470 ;
      LAYER met2 ;
        RECT 705.510 996.000 705.790 1000.000 ;
      LAYER met2 ;
        RECT 706.070 995.720 707.530 998.470 ;
      LAYER met2 ;
        RECT 707.810 996.000 708.090 1000.000 ;
      LAYER met2 ;
        RECT 708.370 995.720 709.370 998.470 ;
      LAYER met2 ;
        RECT 709.650 996.000 709.930 1000.000 ;
      LAYER met2 ;
        RECT 710.210 995.720 711.670 998.470 ;
      LAYER met2 ;
        RECT 711.950 996.000 712.230 1000.000 ;
        RECT 712.700 999.870 714.530 1000.000 ;
      LAYER met2 ;
        RECT 712.510 995.720 713.970 998.470 ;
      LAYER met2 ;
        RECT 714.250 996.000 714.530 999.870 ;
      LAYER met2 ;
        RECT 714.810 995.720 715.810 998.470 ;
      LAYER met2 ;
        RECT 716.090 996.000 716.370 1000.000 ;
      LAYER met2 ;
        RECT 716.650 995.720 718.110 998.470 ;
      LAYER met2 ;
        RECT 718.390 996.000 718.670 1000.000 ;
      LAYER met2 ;
        RECT 718.950 995.720 720.410 998.470 ;
      LAYER met2 ;
        RECT 720.690 996.000 720.970 1000.000 ;
      LAYER met2 ;
        RECT 721.250 995.720 722.710 998.470 ;
      LAYER met2 ;
        RECT 722.990 996.000 723.270 1000.000 ;
      LAYER met2 ;
        RECT 723.550 995.720 724.550 998.470 ;
      LAYER met2 ;
        RECT 724.830 996.000 725.110 1000.000 ;
      LAYER met2 ;
        RECT 725.390 995.720 726.850 998.470 ;
      LAYER met2 ;
        RECT 727.130 996.000 727.410 1000.000 ;
      LAYER met2 ;
        RECT 727.690 995.720 729.150 998.470 ;
      LAYER met2 ;
        RECT 729.430 996.000 729.710 1000.000 ;
      LAYER met2 ;
        RECT 729.990 995.720 730.990 998.470 ;
      LAYER met2 ;
        RECT 731.270 996.000 731.550 1000.000 ;
      LAYER met2 ;
        RECT 731.830 995.720 733.290 998.470 ;
      LAYER met2 ;
        RECT 733.570 996.000 733.850 1000.000 ;
      LAYER met2 ;
        RECT 734.130 995.720 735.590 998.470 ;
      LAYER met2 ;
        RECT 735.870 996.000 736.150 1000.000 ;
      LAYER met2 ;
        RECT 736.430 995.720 737.890 998.470 ;
      LAYER met2 ;
        RECT 738.170 996.000 738.450 1000.000 ;
      LAYER met2 ;
        RECT 738.730 995.720 739.730 998.470 ;
      LAYER met2 ;
        RECT 740.010 996.000 740.290 1000.000 ;
      LAYER met2 ;
        RECT 740.570 995.720 742.030 998.470 ;
      LAYER met2 ;
        RECT 742.310 996.000 742.590 1000.000 ;
      LAYER met2 ;
        RECT 742.870 995.720 744.330 998.470 ;
      LAYER met2 ;
        RECT 744.610 996.000 744.890 1000.000 ;
      LAYER met2 ;
        RECT 745.170 995.720 746.170 998.470 ;
      LAYER met2 ;
        RECT 746.450 996.000 746.730 1000.000 ;
      LAYER met2 ;
        RECT 747.010 995.720 748.470 998.470 ;
      LAYER met2 ;
        RECT 748.750 996.000 749.030 1000.000 ;
      LAYER met2 ;
        RECT 749.310 995.720 750.770 998.470 ;
      LAYER met2 ;
        RECT 751.050 996.000 751.330 1000.000 ;
      LAYER met2 ;
        RECT 751.610 995.720 753.070 998.470 ;
      LAYER met2 ;
        RECT 753.350 996.000 753.630 1000.000 ;
      LAYER met2 ;
        RECT 753.910 995.720 754.910 998.470 ;
      LAYER met2 ;
        RECT 755.190 996.000 755.470 1000.000 ;
      LAYER met2 ;
        RECT 755.750 995.720 757.210 998.470 ;
      LAYER met2 ;
        RECT 757.490 996.000 757.770 1000.000 ;
      LAYER met2 ;
        RECT 758.050 995.720 759.510 998.470 ;
      LAYER met2 ;
        RECT 759.790 996.000 760.070 1000.000 ;
      LAYER met2 ;
        RECT 760.350 995.720 761.350 998.470 ;
      LAYER met2 ;
        RECT 761.630 996.000 761.910 1000.000 ;
      LAYER met2 ;
        RECT 762.190 995.720 763.650 998.470 ;
      LAYER met2 ;
        RECT 763.930 996.000 764.210 1000.000 ;
      LAYER met2 ;
        RECT 764.490 995.720 765.950 998.470 ;
      LAYER met2 ;
        RECT 766.230 996.000 766.510 1000.000 ;
      LAYER met2 ;
        RECT 766.790 995.720 768.250 998.470 ;
      LAYER met2 ;
        RECT 768.530 996.000 768.810 1000.000 ;
      LAYER met2 ;
        RECT 769.090 995.720 770.090 998.470 ;
      LAYER met2 ;
        RECT 770.370 996.000 770.650 1000.000 ;
      LAYER met2 ;
        RECT 770.930 995.720 772.390 998.470 ;
      LAYER met2 ;
        RECT 772.670 996.000 772.950 1000.000 ;
      LAYER met2 ;
        RECT 773.230 995.720 774.690 998.470 ;
      LAYER met2 ;
        RECT 774.970 996.000 775.250 1000.000 ;
      LAYER met2 ;
        RECT 775.530 995.720 776.530 998.470 ;
      LAYER met2 ;
        RECT 776.810 996.000 777.090 1000.000 ;
      LAYER met2 ;
        RECT 777.370 995.720 778.830 998.470 ;
      LAYER met2 ;
        RECT 779.110 996.000 779.390 1000.000 ;
      LAYER met2 ;
        RECT 779.670 995.720 781.130 998.470 ;
      LAYER met2 ;
        RECT 781.410 996.000 781.690 1000.000 ;
      LAYER met2 ;
        RECT 781.970 995.720 783.430 998.470 ;
      LAYER met2 ;
        RECT 783.710 996.000 783.990 1000.000 ;
      LAYER met2 ;
        RECT 784.270 995.720 785.270 998.470 ;
      LAYER met2 ;
        RECT 785.550 996.000 785.830 1000.000 ;
      LAYER met2 ;
        RECT 786.110 995.720 787.570 998.470 ;
      LAYER met2 ;
        RECT 787.850 996.000 788.130 1000.000 ;
      LAYER met2 ;
        RECT 788.410 995.720 789.870 998.470 ;
      LAYER met2 ;
        RECT 790.150 996.000 790.430 1000.000 ;
      LAYER met2 ;
        RECT 790.710 995.720 791.710 998.470 ;
      LAYER met2 ;
        RECT 791.990 996.000 792.270 1000.000 ;
      LAYER met2 ;
        RECT 792.550 995.720 794.010 998.470 ;
      LAYER met2 ;
        RECT 794.290 996.000 794.570 1000.000 ;
      LAYER met2 ;
        RECT 794.850 995.720 796.310 998.470 ;
      LAYER met2 ;
        RECT 796.590 996.000 796.870 1000.000 ;
      LAYER met2 ;
        RECT 797.150 995.720 798.610 998.470 ;
      LAYER met2 ;
        RECT 798.890 996.000 799.170 1000.000 ;
      LAYER met2 ;
        RECT 799.450 995.720 800.450 998.470 ;
      LAYER met2 ;
        RECT 800.730 996.000 801.010 1000.000 ;
      LAYER met2 ;
        RECT 801.290 995.720 802.750 998.470 ;
      LAYER met2 ;
        RECT 803.030 996.000 803.310 1000.000 ;
      LAYER met2 ;
        RECT 803.590 995.720 805.050 998.470 ;
      LAYER met2 ;
        RECT 805.330 996.000 805.610 1000.000 ;
      LAYER met2 ;
        RECT 805.890 995.720 806.890 998.470 ;
      LAYER met2 ;
        RECT 807.170 996.000 807.450 1000.000 ;
      LAYER met2 ;
        RECT 807.730 995.720 809.190 998.470 ;
      LAYER met2 ;
        RECT 809.470 996.000 809.750 1000.000 ;
      LAYER met2 ;
        RECT 810.030 995.720 811.490 998.470 ;
      LAYER met2 ;
        RECT 811.770 996.000 812.050 1000.000 ;
      LAYER met2 ;
        RECT 812.330 995.720 813.790 998.470 ;
      LAYER met2 ;
        RECT 814.070 996.000 814.350 1000.000 ;
      LAYER met2 ;
        RECT 814.630 995.720 815.630 998.470 ;
      LAYER met2 ;
        RECT 815.910 996.000 816.190 1000.000 ;
      LAYER met2 ;
        RECT 816.470 995.720 817.930 998.470 ;
      LAYER met2 ;
        RECT 818.210 996.000 818.490 1000.000 ;
      LAYER met2 ;
        RECT 818.770 995.720 820.230 998.470 ;
      LAYER met2 ;
        RECT 820.510 996.000 820.790 1000.000 ;
      LAYER met2 ;
        RECT 821.070 995.720 822.070 998.470 ;
      LAYER met2 ;
        RECT 822.350 996.000 822.630 1000.000 ;
      LAYER met2 ;
        RECT 822.910 995.720 824.370 998.470 ;
      LAYER met2 ;
        RECT 824.650 996.000 824.930 1000.000 ;
      LAYER met2 ;
        RECT 825.210 995.720 826.670 998.470 ;
      LAYER met2 ;
        RECT 826.950 996.000 827.230 1000.000 ;
      LAYER met2 ;
        RECT 827.510 995.720 828.970 998.470 ;
      LAYER met2 ;
        RECT 829.250 996.000 829.530 1000.000 ;
      LAYER met2 ;
        RECT 829.810 995.720 830.810 998.470 ;
      LAYER met2 ;
        RECT 831.090 996.000 831.370 1000.000 ;
      LAYER met2 ;
        RECT 831.650 995.720 833.110 998.470 ;
      LAYER met2 ;
        RECT 833.390 996.000 833.670 1000.000 ;
      LAYER met2 ;
        RECT 833.950 995.720 835.410 998.470 ;
      LAYER met2 ;
        RECT 835.690 996.000 835.970 1000.000 ;
      LAYER met2 ;
        RECT 836.250 995.720 837.250 998.470 ;
      LAYER met2 ;
        RECT 837.530 996.000 837.810 1000.000 ;
      LAYER met2 ;
        RECT 838.090 995.720 839.550 998.470 ;
      LAYER met2 ;
        RECT 839.830 996.000 840.110 1000.000 ;
        RECT 841.960 999.870 842.410 1000.000 ;
        RECT 842.880 999.870 844.250 1000.000 ;
        RECT 844.720 999.870 846.550 1000.000 ;
      LAYER met2 ;
        RECT 840.390 995.720 841.850 998.470 ;
      LAYER met2 ;
        RECT 842.130 996.000 842.410 999.870 ;
      LAYER met2 ;
        RECT 842.690 995.720 843.690 998.470 ;
      LAYER met2 ;
        RECT 843.970 996.000 844.250 999.870 ;
      LAYER met2 ;
        RECT 844.530 995.720 845.990 998.470 ;
      LAYER met2 ;
        RECT 846.270 996.000 846.550 999.870 ;
      LAYER met2 ;
        RECT 846.830 995.720 848.290 998.470 ;
      LAYER met2 ;
        RECT 848.570 996.000 848.850 1000.000 ;
      LAYER met2 ;
        RECT 849.130 995.720 850.590 998.470 ;
      LAYER met2 ;
        RECT 850.870 996.000 851.150 1000.000 ;
      LAYER met2 ;
        RECT 851.430 995.720 852.430 998.470 ;
      LAYER met2 ;
        RECT 852.710 996.000 852.990 1000.000 ;
      LAYER met2 ;
        RECT 853.270 995.720 854.730 998.470 ;
      LAYER met2 ;
        RECT 855.010 996.000 855.290 1000.000 ;
      LAYER met2 ;
        RECT 855.570 995.720 857.030 998.470 ;
      LAYER met2 ;
        RECT 857.310 996.000 857.590 1000.000 ;
      LAYER met2 ;
        RECT 857.870 995.720 858.870 998.470 ;
      LAYER met2 ;
        RECT 859.150 996.000 859.430 1000.000 ;
      LAYER met2 ;
        RECT 859.710 995.720 861.170 998.470 ;
      LAYER met2 ;
        RECT 861.450 996.000 861.730 1000.000 ;
      LAYER met2 ;
        RECT 862.010 995.720 863.470 998.470 ;
      LAYER met2 ;
        RECT 863.750 996.000 864.030 1000.000 ;
      LAYER met2 ;
        RECT 864.310 995.720 865.770 998.470 ;
      LAYER met2 ;
        RECT 866.050 996.000 866.330 1000.000 ;
      LAYER met2 ;
        RECT 866.610 995.720 867.610 998.470 ;
      LAYER met2 ;
        RECT 867.890 996.000 868.170 1000.000 ;
      LAYER met2 ;
        RECT 868.450 995.720 869.910 998.470 ;
      LAYER met2 ;
        RECT 870.190 996.000 870.470 1000.000 ;
      LAYER met2 ;
        RECT 870.750 995.720 872.210 998.470 ;
      LAYER met2 ;
        RECT 872.490 996.000 872.770 1000.000 ;
      LAYER met2 ;
        RECT 873.050 995.720 874.050 998.470 ;
      LAYER met2 ;
        RECT 874.330 996.000 874.610 1000.000 ;
      LAYER met2 ;
        RECT 874.890 995.720 876.350 998.470 ;
      LAYER met2 ;
        RECT 876.630 996.000 876.910 1000.000 ;
      LAYER met2 ;
        RECT 877.190 995.720 878.650 998.470 ;
      LAYER met2 ;
        RECT 878.930 996.000 879.210 1000.000 ;
      LAYER met2 ;
        RECT 879.490 995.720 880.950 998.470 ;
      LAYER met2 ;
        RECT 881.230 996.000 881.510 1000.000 ;
      LAYER met2 ;
        RECT 881.790 995.720 882.790 998.470 ;
      LAYER met2 ;
        RECT 883.070 996.000 883.350 1000.000 ;
        RECT 884.280 999.870 885.650 1000.000 ;
      LAYER met2 ;
        RECT 883.630 995.720 885.090 998.470 ;
      LAYER met2 ;
        RECT 885.370 996.000 885.650 999.870 ;
      LAYER met2 ;
        RECT 885.930 995.720 887.390 998.470 ;
      LAYER met2 ;
        RECT 887.670 996.000 887.950 1000.000 ;
        RECT 888.420 999.870 889.790 1000.000 ;
      LAYER met2 ;
        RECT 888.230 995.720 889.230 998.470 ;
      LAYER met2 ;
        RECT 889.510 996.000 889.790 999.870 ;
      LAYER met2 ;
        RECT 890.070 995.720 891.530 998.470 ;
      LAYER met2 ;
        RECT 891.810 996.000 892.090 1000.000 ;
        RECT 892.560 999.870 894.390 1000.000 ;
      LAYER met2 ;
        RECT 892.370 995.720 893.830 998.470 ;
      LAYER met2 ;
        RECT 894.110 996.000 894.390 999.870 ;
      LAYER met2 ;
        RECT 894.670 995.720 896.130 998.470 ;
      LAYER met2 ;
        RECT 896.410 996.000 896.690 1000.000 ;
        RECT 897.620 999.870 898.530 1000.000 ;
      LAYER met2 ;
        RECT 896.970 995.720 897.970 998.470 ;
      LAYER met2 ;
        RECT 898.250 996.000 898.530 999.870 ;
      LAYER met2 ;
        RECT 898.810 995.720 900.270 998.470 ;
      LAYER met2 ;
        RECT 900.550 996.000 900.830 1000.000 ;
        RECT 901.300 999.870 903.130 1000.000 ;
      LAYER met2 ;
        RECT 901.110 995.720 902.570 998.470 ;
      LAYER met2 ;
        RECT 902.850 996.000 903.130 999.870 ;
      LAYER met2 ;
        RECT 903.410 995.720 904.410 998.470 ;
      LAYER met2 ;
        RECT 904.690 996.000 904.970 1000.000 ;
        RECT 905.440 999.870 907.270 1000.000 ;
      LAYER met2 ;
        RECT 905.250 995.720 906.710 998.470 ;
      LAYER met2 ;
        RECT 906.990 996.000 907.270 999.870 ;
      LAYER met2 ;
        RECT 907.550 995.720 909.010 998.470 ;
      LAYER met2 ;
        RECT 909.290 996.000 909.570 1000.000 ;
        RECT 911.590 999.160 911.870 1000.000 ;
        RECT 912.340 999.160 912.480 1001.650 ;
        RECT 1011.700 1000.010 1011.840 1008.790 ;
        RECT 1048.960 1000.010 1049.100 1694.570 ;
        RECT 1053.500 1011.170 1053.760 1011.490 ;
        RECT 1053.560 1007.750 1053.700 1011.170 ;
        RECT 1062.300 1009.790 1062.440 1700.270 ;
        RECT 1073.690 1700.000 1073.970 1704.000 ;
        RECT 1087.490 1700.410 1087.770 1704.000 ;
        RECT 1087.490 1700.270 1090.040 1700.410 ;
        RECT 1087.490 1700.000 1087.770 1700.270 ;
        RECT 1070.520 1694.910 1070.780 1695.230 ;
        RECT 1070.580 1690.210 1070.720 1694.910 ;
        RECT 1070.120 1690.070 1070.720 1690.210 ;
        RECT 1070.120 1642.530 1070.260 1690.070 ;
        RECT 1073.800 1688.770 1073.940 1700.000 ;
        RECT 1076.500 1694.230 1076.760 1694.550 ;
        RECT 1073.740 1688.450 1074.000 1688.770 ;
        RECT 1069.600 1642.210 1069.860 1642.530 ;
        RECT 1070.060 1642.210 1070.320 1642.530 ;
        RECT 1069.660 1400.530 1069.800 1642.210 ;
        RECT 1069.200 1400.390 1069.800 1400.530 ;
        RECT 1069.200 1353.190 1069.340 1400.390 ;
        RECT 1069.140 1352.870 1069.400 1353.190 ;
        RECT 1069.600 1352.530 1069.860 1352.850 ;
        RECT 1069.660 1303.890 1069.800 1352.530 ;
        RECT 1069.140 1303.570 1069.400 1303.890 ;
        RECT 1069.600 1303.570 1069.860 1303.890 ;
        RECT 1069.200 1256.370 1069.340 1303.570 ;
        RECT 1069.200 1256.230 1069.800 1256.370 ;
        RECT 1062.700 1051.970 1062.960 1052.290 ;
        RECT 1057.180 1009.470 1057.440 1009.790 ;
        RECT 1062.240 1009.470 1062.500 1009.790 ;
        RECT 1053.040 1007.430 1053.300 1007.750 ;
        RECT 1053.500 1007.430 1053.760 1007.750 ;
        RECT 1053.100 1000.010 1053.240 1007.430 ;
        RECT 1057.240 1000.010 1057.380 1009.470 ;
        RECT 1062.760 1000.010 1062.900 1051.970 ;
        RECT 1065.910 1009.275 1066.190 1009.645 ;
        RECT 1065.980 1000.010 1066.120 1009.275 ;
        RECT 1069.660 1000.690 1069.800 1256.230 ;
        RECT 1069.660 1000.550 1071.180 1000.690 ;
        RECT 1071.040 1000.010 1071.180 1000.550 ;
        RECT 1076.560 1000.010 1076.700 1694.230 ;
        RECT 1087.530 1009.955 1087.810 1010.325 ;
        RECT 1083.400 1009.130 1083.660 1009.450 ;
        RECT 1078.800 1007.770 1079.060 1008.090 ;
        RECT 1011.700 1000.000 1013.380 1000.010 ;
        RECT 1048.960 1000.000 1050.180 1000.010 ;
        RECT 1053.100 1000.000 1054.780 1000.010 ;
        RECT 1057.240 1000.000 1058.920 1000.010 ;
        RECT 1062.760 1000.000 1063.060 1000.010 ;
        RECT 1065.980 1000.000 1067.660 1000.010 ;
        RECT 1071.040 1000.000 1071.800 1000.010 ;
        RECT 1076.400 1000.000 1076.700 1000.010 ;
        RECT 1078.860 1000.010 1079.000 1007.770 ;
        RECT 1083.460 1000.010 1083.600 1009.130 ;
        RECT 1087.600 1000.010 1087.740 1009.955 ;
        RECT 1089.900 1009.450 1090.040 1700.270 ;
        RECT 1102.210 1700.000 1102.490 1704.000 ;
        RECT 1116.010 1700.000 1116.290 1704.000 ;
        RECT 1130.730 1700.000 1131.010 1704.000 ;
        RECT 1144.530 1700.000 1144.810 1704.000 ;
        RECT 1159.250 1700.000 1159.530 1704.000 ;
        RECT 1173.050 1700.000 1173.330 1704.000 ;
        RECT 1187.770 1700.000 1188.050 1704.000 ;
        RECT 1201.570 1700.410 1201.850 1704.000 ;
        RECT 1200.760 1700.270 1201.850 1700.410 ;
        RECT 1102.320 1689.450 1102.460 1700.000 ;
        RECT 1105.020 1693.890 1105.280 1694.210 ;
        RECT 1102.260 1689.130 1102.520 1689.450 ;
        RECT 1105.080 1642.530 1105.220 1693.890 ;
        RECT 1111.000 1693.550 1111.260 1693.870 ;
        RECT 1104.100 1642.210 1104.360 1642.530 ;
        RECT 1105.020 1642.210 1105.280 1642.530 ;
        RECT 1104.160 1400.790 1104.300 1642.210 ;
        RECT 1104.100 1400.470 1104.360 1400.790 ;
        RECT 1105.020 1400.470 1105.280 1400.790 ;
        RECT 1105.080 1352.850 1105.220 1400.470 ;
        RECT 1104.100 1352.530 1104.360 1352.850 ;
        RECT 1105.020 1352.530 1105.280 1352.850 ;
        RECT 1104.160 1304.230 1104.300 1352.530 ;
        RECT 1104.100 1303.910 1104.360 1304.230 ;
        RECT 1105.020 1303.910 1105.280 1304.230 ;
        RECT 1105.080 1256.630 1105.220 1303.910 ;
        RECT 1104.100 1256.310 1104.360 1256.630 ;
        RECT 1105.020 1256.310 1105.280 1256.630 ;
        RECT 1100.870 1014.035 1101.150 1014.405 ;
        RECT 1093.060 1011.510 1093.320 1011.830 ;
        RECT 1089.840 1009.130 1090.100 1009.450 ;
        RECT 1093.120 1008.770 1093.260 1011.510 ;
        RECT 1100.420 1011.170 1100.680 1011.490 ;
        RECT 1092.140 1008.450 1092.400 1008.770 ;
        RECT 1093.060 1008.450 1093.320 1008.770 ;
        RECT 1092.200 1000.010 1092.340 1008.450 ;
        RECT 1097.200 1008.110 1097.460 1008.430 ;
        RECT 1097.260 1000.010 1097.400 1008.110 ;
        RECT 1100.480 1007.750 1100.620 1011.170 ;
        RECT 1100.420 1007.430 1100.680 1007.750 ;
        RECT 1100.940 1000.010 1101.080 1014.035 ;
        RECT 1104.160 1011.830 1104.300 1256.310 ;
        RECT 1104.100 1011.510 1104.360 1011.830 ;
        RECT 1105.480 1011.510 1105.740 1011.830 ;
        RECT 1105.540 1000.010 1105.680 1011.510 ;
        RECT 1111.060 1000.010 1111.200 1693.550 ;
        RECT 1116.120 1690.130 1116.260 1700.000 ;
        RECT 1116.060 1689.810 1116.320 1690.130 ;
        RECT 1130.840 1689.110 1130.980 1700.000 ;
        RECT 1130.780 1688.790 1131.040 1689.110 ;
        RECT 1144.640 1686.730 1144.780 1700.000 ;
        RECT 1159.360 1689.790 1159.500 1700.000 ;
        RECT 1159.300 1689.470 1159.560 1689.790 ;
        RECT 1144.580 1686.410 1144.840 1686.730 ;
        RECT 1173.160 1684.690 1173.300 1700.000 ;
        RECT 1186.440 1693.890 1186.700 1694.210 ;
        RECT 1185.980 1693.550 1186.240 1693.870 ;
        RECT 1180.920 1686.410 1181.180 1686.730 ;
        RECT 1173.100 1684.370 1173.360 1684.690 ;
        RECT 1146.420 1025.450 1146.680 1025.770 ;
        RECT 1124.790 1013.355 1125.070 1013.725 ;
        RECT 1117.890 1011.995 1118.170 1012.365 ;
        RECT 1113.760 1008.790 1114.020 1009.110 ;
        RECT 1078.860 1000.000 1080.540 1000.010 ;
        RECT 1083.460 1000.000 1085.140 1000.010 ;
        RECT 1087.600 1000.000 1089.280 1000.010 ;
        RECT 1092.200 1000.000 1093.420 1000.010 ;
        RECT 1097.260 1000.000 1098.020 1000.010 ;
        RECT 1100.940 1000.000 1102.160 1000.010 ;
        RECT 1105.540 1000.000 1106.760 1000.010 ;
        RECT 1110.900 1000.000 1111.200 1000.010 ;
        RECT 1113.820 1000.010 1113.960 1008.790 ;
        RECT 1117.960 1000.010 1118.100 1011.995 ;
        RECT 1124.860 1000.010 1125.000 1013.355 ;
        RECT 1145.500 1013.210 1145.760 1013.530 ;
        RECT 1128.930 1012.675 1129.210 1013.045 ;
        RECT 1145.560 1012.930 1145.700 1013.210 ;
        RECT 1145.560 1012.790 1146.160 1012.930 ;
        RECT 1129.000 1000.010 1129.140 1012.675 ;
        RECT 1141.810 1011.315 1142.090 1011.685 ;
        RECT 1145.040 1011.510 1145.300 1011.830 ;
        RECT 1138.600 1010.150 1138.860 1010.470 ;
        RECT 1133.080 1009.810 1133.340 1010.130 ;
        RECT 1133.140 1000.010 1133.280 1009.810 ;
        RECT 1138.660 1000.010 1138.800 1010.150 ;
        RECT 1141.880 1000.010 1142.020 1011.315 ;
        RECT 1145.100 1008.770 1145.240 1011.510 ;
        RECT 1145.500 1011.170 1145.760 1011.490 ;
        RECT 1145.560 1010.470 1145.700 1011.170 ;
        RECT 1145.500 1010.150 1145.760 1010.470 ;
        RECT 1146.020 1010.130 1146.160 1012.790 ;
        RECT 1145.960 1009.810 1146.220 1010.130 ;
        RECT 1145.040 1008.450 1145.300 1008.770 ;
        RECT 1146.480 1000.010 1146.620 1025.450 ;
        RECT 1152.400 1025.110 1152.660 1025.430 ;
        RECT 1152.460 1000.010 1152.600 1025.110 ;
        RECT 1154.700 1024.770 1154.960 1025.090 ;
        RECT 1113.820 1000.000 1115.500 1000.010 ;
        RECT 1117.960 1000.000 1119.640 1000.010 ;
        RECT 1124.860 1000.000 1126.080 1000.010 ;
        RECT 1129.000 1000.000 1130.680 1000.010 ;
        RECT 1133.140 1000.000 1134.820 1000.010 ;
        RECT 1138.660 1000.000 1138.960 1000.010 ;
        RECT 1141.880 1000.000 1143.560 1000.010 ;
        RECT 1146.480 1000.000 1147.700 1000.010 ;
        RECT 1152.300 1000.000 1152.600 1000.010 ;
        RECT 1154.760 1000.010 1154.900 1024.770 ;
        RECT 1163.440 1024.430 1163.700 1024.750 ;
        RECT 1159.760 1016.950 1160.020 1017.270 ;
        RECT 1159.820 1000.010 1159.960 1016.950 ;
        RECT 1163.500 1000.010 1163.640 1024.430 ;
        RECT 1173.100 1013.210 1173.360 1013.530 ;
        RECT 1173.160 1012.170 1173.300 1013.210 ;
        RECT 1180.000 1012.190 1180.260 1012.510 ;
        RECT 1180.460 1012.190 1180.720 1012.510 ;
        RECT 1173.100 1011.850 1173.360 1012.170 ;
        RECT 1166.190 1010.635 1166.470 1011.005 ;
        RECT 1166.260 1000.010 1166.400 1010.635 ;
        RECT 1180.060 1010.130 1180.200 1012.190 ;
        RECT 1179.540 1009.810 1179.800 1010.130 ;
        RECT 1180.000 1009.810 1180.260 1010.130 ;
        RECT 1179.600 1008.430 1179.740 1009.810 ;
        RECT 1179.540 1008.110 1179.800 1008.430 ;
        RECT 1180.520 1000.010 1180.660 1012.190 ;
        RECT 1154.760 1000.000 1156.440 1000.010 ;
        RECT 1159.820 1000.000 1161.040 1000.010 ;
        RECT 1163.500 1000.000 1165.180 1000.010 ;
        RECT 1166.260 1000.000 1167.480 1000.010 ;
        RECT 1180.360 1000.000 1180.660 1000.010 ;
        RECT 911.590 999.020 912.480 999.160 ;
      LAYER met2 ;
        RECT 909.850 995.720 911.310 998.470 ;
      LAYER met2 ;
        RECT 911.590 996.000 911.870 999.020 ;
      LAYER met2 ;
        RECT 912.150 995.720 913.150 998.470 ;
      LAYER met2 ;
        RECT 913.430 996.000 913.710 1000.000 ;
      LAYER met2 ;
        RECT 913.990 995.720 915.450 998.470 ;
      LAYER met2 ;
        RECT 915.730 996.000 916.010 1000.000 ;
      LAYER met2 ;
        RECT 916.290 995.720 917.750 998.470 ;
      LAYER met2 ;
        RECT 918.030 996.000 918.310 1000.000 ;
      LAYER met2 ;
        RECT 918.590 995.720 919.590 998.470 ;
      LAYER met2 ;
        RECT 919.870 996.000 920.150 1000.000 ;
      LAYER met2 ;
        RECT 920.430 995.720 921.890 998.470 ;
      LAYER met2 ;
        RECT 922.170 996.000 922.450 1000.000 ;
      LAYER met2 ;
        RECT 922.730 995.720 924.190 998.470 ;
      LAYER met2 ;
        RECT 924.470 996.000 924.750 1000.000 ;
      LAYER met2 ;
        RECT 925.030 995.720 926.490 998.470 ;
      LAYER met2 ;
        RECT 926.770 996.000 927.050 1000.000 ;
      LAYER met2 ;
        RECT 927.330 995.720 928.330 998.470 ;
      LAYER met2 ;
        RECT 928.610 996.000 928.890 1000.000 ;
      LAYER met2 ;
        RECT 929.170 995.720 930.630 998.470 ;
      LAYER met2 ;
        RECT 930.910 996.000 931.190 1000.000 ;
      LAYER met2 ;
        RECT 931.470 995.720 932.930 998.470 ;
      LAYER met2 ;
        RECT 933.210 996.000 933.490 1000.000 ;
      LAYER met2 ;
        RECT 933.770 995.720 934.770 998.470 ;
      LAYER met2 ;
        RECT 935.050 996.000 935.330 1000.000 ;
      LAYER met2 ;
        RECT 935.610 995.720 937.070 998.470 ;
      LAYER met2 ;
        RECT 937.350 996.000 937.630 1000.000 ;
      LAYER met2 ;
        RECT 937.910 995.720 939.370 998.470 ;
      LAYER met2 ;
        RECT 939.650 996.000 939.930 1000.000 ;
      LAYER met2 ;
        RECT 940.210 995.720 941.670 998.470 ;
      LAYER met2 ;
        RECT 941.950 996.000 942.230 1000.000 ;
      LAYER met2 ;
        RECT 942.510 995.720 943.510 998.470 ;
      LAYER met2 ;
        RECT 943.790 996.000 944.070 1000.000 ;
      LAYER met2 ;
        RECT 944.350 995.720 945.810 998.470 ;
      LAYER met2 ;
        RECT 946.090 996.000 946.370 1000.000 ;
      LAYER met2 ;
        RECT 946.650 995.720 948.110 998.470 ;
      LAYER met2 ;
        RECT 948.390 996.000 948.670 1000.000 ;
      LAYER met2 ;
        RECT 948.950 995.720 949.950 998.470 ;
      LAYER met2 ;
        RECT 950.230 996.000 950.510 1000.000 ;
      LAYER met2 ;
        RECT 950.790 995.720 952.250 998.470 ;
      LAYER met2 ;
        RECT 952.530 996.000 952.810 1000.000 ;
      LAYER met2 ;
        RECT 953.090 995.720 954.550 998.470 ;
      LAYER met2 ;
        RECT 954.830 996.000 955.110 1000.000 ;
      LAYER met2 ;
        RECT 955.390 995.720 956.850 998.470 ;
      LAYER met2 ;
        RECT 957.130 996.000 957.410 1000.000 ;
      LAYER met2 ;
        RECT 957.690 995.720 958.690 998.470 ;
      LAYER met2 ;
        RECT 958.970 996.000 959.250 1000.000 ;
      LAYER met2 ;
        RECT 959.530 995.720 960.990 998.470 ;
      LAYER met2 ;
        RECT 961.270 996.000 961.550 1000.000 ;
      LAYER met2 ;
        RECT 961.830 995.720 963.290 998.470 ;
      LAYER met2 ;
        RECT 963.570 996.000 963.850 1000.000 ;
      LAYER met2 ;
        RECT 964.130 995.720 965.130 998.470 ;
      LAYER met2 ;
        RECT 965.410 996.000 965.690 1000.000 ;
      LAYER met2 ;
        RECT 965.970 995.720 967.430 998.470 ;
      LAYER met2 ;
        RECT 967.710 996.000 967.990 1000.000 ;
      LAYER met2 ;
        RECT 968.270 995.720 969.730 998.470 ;
      LAYER met2 ;
        RECT 970.010 996.000 970.290 1000.000 ;
      LAYER met2 ;
        RECT 970.570 995.720 972.030 998.470 ;
      LAYER met2 ;
        RECT 972.310 996.000 972.590 1000.000 ;
      LAYER met2 ;
        RECT 972.870 995.720 973.870 998.470 ;
      LAYER met2 ;
        RECT 974.150 996.000 974.430 1000.000 ;
      LAYER met2 ;
        RECT 974.710 995.720 976.170 998.470 ;
      LAYER met2 ;
        RECT 976.450 996.000 976.730 1000.000 ;
      LAYER met2 ;
        RECT 977.010 995.720 978.470 998.470 ;
      LAYER met2 ;
        RECT 978.750 996.000 979.030 1000.000 ;
      LAYER met2 ;
        RECT 979.310 995.720 980.310 998.470 ;
      LAYER met2 ;
        RECT 980.590 996.000 980.870 1000.000 ;
      LAYER met2 ;
        RECT 981.150 995.720 982.610 998.470 ;
      LAYER met2 ;
        RECT 982.890 996.000 983.170 1000.000 ;
      LAYER met2 ;
        RECT 983.450 995.720 984.910 998.470 ;
      LAYER met2 ;
        RECT 985.190 996.000 985.470 1000.000 ;
      LAYER met2 ;
        RECT 985.750 995.720 987.210 998.470 ;
      LAYER met2 ;
        RECT 987.490 996.000 987.770 1000.000 ;
      LAYER met2 ;
        RECT 988.050 995.720 989.050 998.470 ;
      LAYER met2 ;
        RECT 989.330 996.000 989.610 1000.000 ;
      LAYER met2 ;
        RECT 989.890 995.720 991.350 998.470 ;
      LAYER met2 ;
        RECT 991.630 996.000 991.910 1000.000 ;
      LAYER met2 ;
        RECT 992.190 995.720 993.650 998.470 ;
      LAYER met2 ;
        RECT 993.930 996.000 994.210 1000.000 ;
      LAYER met2 ;
        RECT 994.490 995.720 995.490 998.470 ;
      LAYER met2 ;
        RECT 995.770 996.000 996.050 1000.000 ;
      LAYER met2 ;
        RECT 996.330 995.720 997.790 998.470 ;
      LAYER met2 ;
        RECT 998.070 996.000 998.350 1000.000 ;
      LAYER met2 ;
        RECT 998.630 995.720 1000.090 998.470 ;
      LAYER met2 ;
        RECT 1000.370 996.000 1000.650 1000.000 ;
      LAYER met2 ;
        RECT 1000.930 995.720 1002.390 998.470 ;
      LAYER met2 ;
        RECT 1002.670 996.000 1002.950 1000.000 ;
      LAYER met2 ;
        RECT 1003.230 995.720 1004.230 998.470 ;
      LAYER met2 ;
        RECT 1004.510 996.000 1004.790 1000.000 ;
      LAYER met2 ;
        RECT 1005.070 995.720 1006.530 998.470 ;
      LAYER met2 ;
        RECT 1006.810 996.000 1007.090 1000.000 ;
      LAYER met2 ;
        RECT 1007.370 995.720 1008.830 998.470 ;
      LAYER met2 ;
        RECT 1009.110 996.000 1009.390 1000.000 ;
      LAYER met2 ;
        RECT 1009.670 995.720 1010.670 998.470 ;
      LAYER met2 ;
        RECT 1010.950 996.000 1011.230 1000.000 ;
        RECT 1011.700 999.870 1013.530 1000.000 ;
      LAYER met2 ;
        RECT 1011.510 995.720 1012.970 998.470 ;
      LAYER met2 ;
        RECT 1013.250 996.000 1013.530 999.870 ;
      LAYER met2 ;
        RECT 1013.810 995.720 1015.270 998.470 ;
      LAYER met2 ;
        RECT 1015.550 996.000 1015.830 1000.000 ;
      LAYER met2 ;
        RECT 1016.110 995.720 1017.110 998.470 ;
      LAYER met2 ;
        RECT 1017.390 996.000 1017.670 1000.000 ;
      LAYER met2 ;
        RECT 1017.950 995.720 1019.410 998.470 ;
      LAYER met2 ;
        RECT 1019.690 996.000 1019.970 1000.000 ;
      LAYER met2 ;
        RECT 1020.250 995.720 1021.710 998.470 ;
      LAYER met2 ;
        RECT 1021.990 996.000 1022.270 1000.000 ;
      LAYER met2 ;
        RECT 1022.550 995.720 1024.010 998.470 ;
      LAYER met2 ;
        RECT 1024.290 996.000 1024.570 1000.000 ;
      LAYER met2 ;
        RECT 1024.850 995.720 1025.850 998.470 ;
      LAYER met2 ;
        RECT 1026.130 996.000 1026.410 1000.000 ;
      LAYER met2 ;
        RECT 1026.690 995.720 1028.150 998.470 ;
      LAYER met2 ;
        RECT 1028.430 996.000 1028.710 1000.000 ;
      LAYER met2 ;
        RECT 1028.990 995.720 1030.450 998.470 ;
      LAYER met2 ;
        RECT 1030.730 996.000 1031.010 1000.000 ;
      LAYER met2 ;
        RECT 1031.290 995.720 1032.290 998.470 ;
      LAYER met2 ;
        RECT 1032.570 996.000 1032.850 1000.000 ;
      LAYER met2 ;
        RECT 1033.130 995.720 1034.590 998.470 ;
      LAYER met2 ;
        RECT 1034.870 996.000 1035.150 1000.000 ;
      LAYER met2 ;
        RECT 1035.430 995.720 1036.890 998.470 ;
      LAYER met2 ;
        RECT 1037.170 996.000 1037.450 1000.000 ;
      LAYER met2 ;
        RECT 1037.730 995.720 1039.190 998.470 ;
      LAYER met2 ;
        RECT 1039.470 996.000 1039.750 1000.000 ;
      LAYER met2 ;
        RECT 1040.030 995.720 1041.030 998.470 ;
      LAYER met2 ;
        RECT 1041.310 996.000 1041.590 1000.000 ;
      LAYER met2 ;
        RECT 1041.870 995.720 1043.330 998.470 ;
      LAYER met2 ;
        RECT 1043.610 996.000 1043.890 1000.000 ;
      LAYER met2 ;
        RECT 1044.170 995.720 1045.630 998.470 ;
      LAYER met2 ;
        RECT 1045.910 996.000 1046.190 1000.000 ;
      LAYER met2 ;
        RECT 1046.470 995.720 1047.470 998.470 ;
      LAYER met2 ;
        RECT 1047.750 996.000 1048.030 1000.000 ;
        RECT 1048.960 999.870 1050.330 1000.000 ;
      LAYER met2 ;
        RECT 1048.310 995.720 1049.770 998.470 ;
      LAYER met2 ;
        RECT 1050.050 996.000 1050.330 999.870 ;
      LAYER met2 ;
        RECT 1050.610 995.720 1052.070 998.470 ;
      LAYER met2 ;
        RECT 1052.350 996.000 1052.630 1000.000 ;
        RECT 1053.100 999.870 1054.930 1000.000 ;
      LAYER met2 ;
        RECT 1052.910 995.720 1054.370 998.470 ;
      LAYER met2 ;
        RECT 1054.650 996.000 1054.930 999.870 ;
      LAYER met2 ;
        RECT 1055.210 995.720 1056.210 998.470 ;
      LAYER met2 ;
        RECT 1056.490 996.000 1056.770 1000.000 ;
        RECT 1057.240 999.870 1059.070 1000.000 ;
      LAYER met2 ;
        RECT 1057.050 995.720 1058.510 998.470 ;
      LAYER met2 ;
        RECT 1058.790 996.000 1059.070 999.870 ;
      LAYER met2 ;
        RECT 1059.350 995.720 1060.810 998.470 ;
      LAYER met2 ;
        RECT 1061.090 996.000 1061.370 1000.000 ;
        RECT 1062.760 999.870 1063.210 1000.000 ;
      LAYER met2 ;
        RECT 1061.650 995.720 1062.650 998.470 ;
      LAYER met2 ;
        RECT 1062.930 996.000 1063.210 999.870 ;
      LAYER met2 ;
        RECT 1063.490 995.720 1064.950 998.470 ;
      LAYER met2 ;
        RECT 1065.230 996.000 1065.510 1000.000 ;
        RECT 1065.980 999.870 1067.810 1000.000 ;
      LAYER met2 ;
        RECT 1065.790 995.720 1067.250 998.470 ;
      LAYER met2 ;
        RECT 1067.530 996.000 1067.810 999.870 ;
      LAYER met2 ;
        RECT 1068.090 995.720 1069.550 998.470 ;
      LAYER met2 ;
        RECT 1069.830 996.000 1070.110 1000.000 ;
        RECT 1071.040 999.870 1071.950 1000.000 ;
      LAYER met2 ;
        RECT 1070.390 995.720 1071.390 998.470 ;
      LAYER met2 ;
        RECT 1071.670 996.000 1071.950 999.870 ;
      LAYER met2 ;
        RECT 1072.230 995.720 1073.690 998.470 ;
      LAYER met2 ;
        RECT 1073.970 996.000 1074.250 1000.000 ;
        RECT 1076.270 999.870 1076.700 1000.000 ;
      LAYER met2 ;
        RECT 1074.530 995.720 1075.990 998.470 ;
      LAYER met2 ;
        RECT 1076.270 996.000 1076.550 999.870 ;
      LAYER met2 ;
        RECT 1076.830 995.720 1077.830 998.470 ;
      LAYER met2 ;
        RECT 1078.110 996.000 1078.390 1000.000 ;
        RECT 1078.860 999.870 1080.690 1000.000 ;
      LAYER met2 ;
        RECT 1078.670 995.720 1080.130 998.470 ;
      LAYER met2 ;
        RECT 1080.410 996.000 1080.690 999.870 ;
      LAYER met2 ;
        RECT 1080.970 995.720 1082.430 998.470 ;
      LAYER met2 ;
        RECT 1082.710 996.000 1082.990 1000.000 ;
        RECT 1083.460 999.870 1085.290 1000.000 ;
      LAYER met2 ;
        RECT 1083.270 995.720 1084.730 998.470 ;
      LAYER met2 ;
        RECT 1085.010 996.000 1085.290 999.870 ;
      LAYER met2 ;
        RECT 1085.570 995.720 1086.570 998.470 ;
      LAYER met2 ;
        RECT 1086.850 996.000 1087.130 1000.000 ;
        RECT 1087.600 999.870 1089.430 1000.000 ;
      LAYER met2 ;
        RECT 1087.410 995.720 1088.870 998.470 ;
      LAYER met2 ;
        RECT 1089.150 996.000 1089.430 999.870 ;
      LAYER met2 ;
        RECT 1089.710 995.720 1091.170 998.470 ;
      LAYER met2 ;
        RECT 1091.450 996.000 1091.730 1000.000 ;
        RECT 1092.200 999.870 1093.570 1000.000 ;
      LAYER met2 ;
        RECT 1092.010 995.720 1093.010 998.470 ;
      LAYER met2 ;
        RECT 1093.290 996.000 1093.570 999.870 ;
      LAYER met2 ;
        RECT 1093.850 995.720 1095.310 998.470 ;
      LAYER met2 ;
        RECT 1095.590 996.000 1095.870 1000.000 ;
        RECT 1097.260 999.870 1098.170 1000.000 ;
      LAYER met2 ;
        RECT 1096.150 995.720 1097.610 998.470 ;
      LAYER met2 ;
        RECT 1097.890 996.000 1098.170 999.870 ;
      LAYER met2 ;
        RECT 1098.450 995.720 1099.910 998.470 ;
      LAYER met2 ;
        RECT 1100.190 996.000 1100.470 1000.000 ;
        RECT 1100.940 999.870 1102.310 1000.000 ;
      LAYER met2 ;
        RECT 1100.750 995.720 1101.750 998.470 ;
      LAYER met2 ;
        RECT 1102.030 996.000 1102.310 999.870 ;
      LAYER met2 ;
        RECT 1102.590 995.720 1104.050 998.470 ;
      LAYER met2 ;
        RECT 1104.330 996.000 1104.610 1000.000 ;
        RECT 1105.540 999.870 1106.910 1000.000 ;
      LAYER met2 ;
        RECT 1104.890 995.720 1106.350 998.470 ;
      LAYER met2 ;
        RECT 1106.630 996.000 1106.910 999.870 ;
      LAYER met2 ;
        RECT 1107.190 995.720 1108.190 998.470 ;
      LAYER met2 ;
        RECT 1108.470 996.000 1108.750 1000.000 ;
        RECT 1110.770 999.870 1111.200 1000.000 ;
      LAYER met2 ;
        RECT 1109.030 995.720 1110.490 998.470 ;
      LAYER met2 ;
        RECT 1110.770 996.000 1111.050 999.870 ;
      LAYER met2 ;
        RECT 1111.330 995.720 1112.790 998.470 ;
      LAYER met2 ;
        RECT 1113.070 996.000 1113.350 1000.000 ;
        RECT 1113.820 999.870 1115.650 1000.000 ;
      LAYER met2 ;
        RECT 1113.630 995.720 1115.090 998.470 ;
      LAYER met2 ;
        RECT 1115.370 996.000 1115.650 999.870 ;
      LAYER met2 ;
        RECT 1115.930 995.720 1116.930 998.470 ;
      LAYER met2 ;
        RECT 1117.210 996.000 1117.490 1000.000 ;
        RECT 1117.960 999.870 1119.790 1000.000 ;
      LAYER met2 ;
        RECT 1117.770 995.720 1119.230 998.470 ;
      LAYER met2 ;
        RECT 1119.510 996.000 1119.790 999.870 ;
      LAYER met2 ;
        RECT 1120.070 995.720 1121.530 998.470 ;
      LAYER met2 ;
        RECT 1121.810 996.000 1122.090 1000.000 ;
      LAYER met2 ;
        RECT 1122.370 995.720 1123.370 998.470 ;
      LAYER met2 ;
        RECT 1123.650 996.000 1123.930 1000.000 ;
        RECT 1124.860 999.870 1126.230 1000.000 ;
      LAYER met2 ;
        RECT 1124.210 995.720 1125.670 998.470 ;
      LAYER met2 ;
        RECT 1125.950 996.000 1126.230 999.870 ;
      LAYER met2 ;
        RECT 1126.510 995.720 1127.970 998.470 ;
      LAYER met2 ;
        RECT 1128.250 996.000 1128.530 1000.000 ;
        RECT 1129.000 999.870 1130.830 1000.000 ;
      LAYER met2 ;
        RECT 1128.810 995.720 1130.270 998.470 ;
      LAYER met2 ;
        RECT 1130.550 996.000 1130.830 999.870 ;
      LAYER met2 ;
        RECT 1131.110 995.720 1132.110 998.470 ;
      LAYER met2 ;
        RECT 1132.390 996.000 1132.670 1000.000 ;
        RECT 1133.140 999.870 1134.970 1000.000 ;
      LAYER met2 ;
        RECT 1132.950 995.720 1134.410 998.470 ;
      LAYER met2 ;
        RECT 1134.690 996.000 1134.970 999.870 ;
      LAYER met2 ;
        RECT 1135.250 995.720 1136.710 998.470 ;
      LAYER met2 ;
        RECT 1136.990 996.000 1137.270 1000.000 ;
        RECT 1138.660 999.870 1139.110 1000.000 ;
      LAYER met2 ;
        RECT 1137.550 995.720 1138.550 998.470 ;
      LAYER met2 ;
        RECT 1138.830 996.000 1139.110 999.870 ;
      LAYER met2 ;
        RECT 1139.390 995.720 1140.850 998.470 ;
      LAYER met2 ;
        RECT 1141.130 996.000 1141.410 1000.000 ;
        RECT 1141.880 999.870 1143.710 1000.000 ;
      LAYER met2 ;
        RECT 1141.690 995.720 1143.150 998.470 ;
      LAYER met2 ;
        RECT 1143.430 996.000 1143.710 999.870 ;
      LAYER met2 ;
        RECT 1143.990 995.720 1145.450 998.470 ;
      LAYER met2 ;
        RECT 1145.730 996.000 1146.010 1000.000 ;
        RECT 1146.480 999.870 1147.850 1000.000 ;
      LAYER met2 ;
        RECT 1146.290 995.720 1147.290 998.470 ;
      LAYER met2 ;
        RECT 1147.570 996.000 1147.850 999.870 ;
      LAYER met2 ;
        RECT 1148.130 995.720 1149.590 998.470 ;
      LAYER met2 ;
        RECT 1149.870 996.000 1150.150 1000.000 ;
        RECT 1152.170 999.870 1152.600 1000.000 ;
      LAYER met2 ;
        RECT 1150.430 995.720 1151.890 998.470 ;
      LAYER met2 ;
        RECT 1152.170 996.000 1152.450 999.870 ;
      LAYER met2 ;
        RECT 1152.730 995.720 1153.730 998.470 ;
      LAYER met2 ;
        RECT 1154.010 996.000 1154.290 1000.000 ;
        RECT 1154.760 999.870 1156.590 1000.000 ;
      LAYER met2 ;
        RECT 1154.570 995.720 1156.030 998.470 ;
      LAYER met2 ;
        RECT 1156.310 996.000 1156.590 999.870 ;
      LAYER met2 ;
        RECT 1156.870 995.720 1158.330 998.470 ;
      LAYER met2 ;
        RECT 1158.610 996.000 1158.890 1000.000 ;
        RECT 1159.820 999.870 1161.190 1000.000 ;
      LAYER met2 ;
        RECT 1159.170 995.720 1160.630 998.470 ;
      LAYER met2 ;
        RECT 1160.910 996.000 1161.190 999.870 ;
      LAYER met2 ;
        RECT 1161.470 995.720 1162.470 998.470 ;
      LAYER met2 ;
        RECT 1162.750 996.000 1163.030 1000.000 ;
        RECT 1163.500 999.870 1165.330 1000.000 ;
        RECT 1166.260 999.870 1167.630 1000.000 ;
      LAYER met2 ;
        RECT 1163.310 995.720 1164.770 998.470 ;
      LAYER met2 ;
        RECT 1165.050 996.000 1165.330 999.870 ;
      LAYER met2 ;
        RECT 1165.610 995.720 1167.070 998.470 ;
      LAYER met2 ;
        RECT 1167.350 996.000 1167.630 999.870 ;
      LAYER met2 ;
        RECT 1167.910 995.720 1168.910 998.470 ;
      LAYER met2 ;
        RECT 1169.190 996.000 1169.470 1000.000 ;
      LAYER met2 ;
        RECT 1169.750 995.720 1171.210 998.470 ;
      LAYER met2 ;
        RECT 1171.490 996.000 1171.770 1000.000 ;
      LAYER met2 ;
        RECT 1172.050 995.720 1173.510 998.470 ;
      LAYER met2 ;
        RECT 1173.790 996.000 1174.070 1000.000 ;
      LAYER met2 ;
        RECT 1174.350 995.720 1175.350 998.470 ;
      LAYER met2 ;
        RECT 1175.630 996.000 1175.910 1000.000 ;
      LAYER met2 ;
        RECT 1176.190 995.720 1177.650 998.470 ;
      LAYER met2 ;
        RECT 1177.930 996.000 1178.210 1000.000 ;
        RECT 1180.230 999.870 1180.660 1000.000 ;
        RECT 1180.980 1000.010 1181.120 1686.410 ;
        RECT 1186.040 1000.010 1186.180 1693.550 ;
        RECT 1186.500 1012.510 1186.640 1693.890 ;
        RECT 1186.900 1689.810 1187.160 1690.130 ;
        RECT 1186.440 1012.190 1186.700 1012.510 ;
        RECT 1186.960 1000.010 1187.100 1689.810 ;
        RECT 1187.880 1684.350 1188.020 1700.000 ;
        RECT 1197.020 1688.790 1197.280 1689.110 ;
        RECT 1197.080 1686.730 1197.220 1688.790 ;
        RECT 1197.020 1686.410 1197.280 1686.730 ;
        RECT 1188.280 1684.370 1188.540 1684.690 ;
        RECT 1193.340 1684.370 1193.600 1684.690 ;
        RECT 1187.820 1684.030 1188.080 1684.350 ;
        RECT 1180.980 1000.000 1182.660 1000.010 ;
        RECT 1184.500 1000.000 1186.180 1000.010 ;
        RECT 1186.800 1000.000 1187.100 1000.010 ;
        RECT 1180.980 999.870 1182.810 1000.000 ;
      LAYER met2 ;
        RECT 1178.490 995.720 1179.950 998.470 ;
      LAYER met2 ;
        RECT 1180.230 996.000 1180.510 999.870 ;
      LAYER met2 ;
        RECT 1180.790 995.720 1182.250 998.470 ;
      LAYER met2 ;
        RECT 1182.530 996.000 1182.810 999.870 ;
        RECT 1184.370 999.870 1186.180 1000.000 ;
        RECT 1186.670 999.870 1187.100 1000.000 ;
        RECT 1188.340 1000.010 1188.480 1684.370 ;
        RECT 1189.660 1013.550 1189.920 1013.870 ;
        RECT 1189.720 1000.010 1189.860 1013.550 ;
        RECT 1191.500 1009.470 1191.760 1009.790 ;
        RECT 1191.560 1007.750 1191.700 1009.470 ;
        RECT 1191.500 1007.430 1191.760 1007.750 ;
        RECT 1193.400 1000.010 1193.540 1684.370 ;
        RECT 1197.020 1684.030 1197.280 1684.350 ;
        RECT 1200.760 1684.090 1200.900 1700.270 ;
        RECT 1201.570 1700.000 1201.850 1700.270 ;
        RECT 1215.370 1700.000 1215.650 1704.000 ;
        RECT 1230.090 1700.000 1230.370 1704.000 ;
        RECT 1243.890 1700.000 1244.170 1704.000 ;
        RECT 1258.610 1700.410 1258.890 1704.000 ;
        RECT 1258.610 1700.270 1262.080 1700.410 ;
        RECT 1258.610 1700.000 1258.890 1700.270 ;
        RECT 1203.920 1689.130 1204.180 1689.450 ;
        RECT 1214.040 1689.130 1214.300 1689.450 ;
        RECT 1196.100 1012.870 1196.360 1013.190 ;
        RECT 1196.160 1009.110 1196.300 1012.870 ;
        RECT 1197.080 1012.510 1197.220 1684.030 ;
        RECT 1200.300 1683.950 1200.900 1684.090 ;
        RECT 1197.940 1017.290 1198.200 1017.610 ;
        RECT 1197.020 1012.190 1197.280 1012.510 ;
        RECT 1197.480 1011.510 1197.740 1011.830 ;
        RECT 1196.560 1011.170 1196.820 1011.490 ;
        RECT 1196.620 1010.470 1196.760 1011.170 ;
        RECT 1196.560 1010.150 1196.820 1010.470 ;
        RECT 1197.020 1010.150 1197.280 1010.470 ;
        RECT 1196.100 1008.790 1196.360 1009.110 ;
        RECT 1197.080 1000.010 1197.220 1010.150 ;
        RECT 1197.540 1008.770 1197.680 1011.510 ;
        RECT 1197.480 1008.450 1197.740 1008.770 ;
        RECT 1198.000 1000.010 1198.140 1017.290 ;
        RECT 1200.300 1010.470 1200.440 1683.950 ;
        RECT 1203.460 1017.290 1203.720 1017.610 ;
        RECT 1200.240 1010.150 1200.500 1010.470 ;
        RECT 1200.240 1009.470 1200.500 1009.790 ;
        RECT 1200.300 1000.010 1200.440 1009.470 ;
        RECT 1203.520 1000.010 1203.660 1017.290 ;
        RECT 1203.980 1012.850 1204.120 1689.130 ;
        RECT 1204.380 1012.870 1204.640 1013.190 ;
        RECT 1213.580 1012.870 1213.840 1013.190 ;
        RECT 1203.920 1012.530 1204.180 1012.850 ;
        RECT 1204.440 1000.010 1204.580 1012.870 ;
        RECT 1204.840 1008.110 1205.100 1008.430 ;
        RECT 1188.340 1000.000 1189.100 1000.010 ;
        RECT 1189.720 1000.000 1190.940 1000.010 ;
        RECT 1193.240 1000.000 1193.540 1000.010 ;
        RECT 1195.540 1000.000 1197.220 1000.010 ;
        RECT 1197.840 1000.000 1198.140 1000.010 ;
        RECT 1199.680 1000.000 1200.440 1000.010 ;
        RECT 1201.980 1000.000 1203.660 1000.010 ;
        RECT 1204.280 1000.000 1204.580 1000.010 ;
        RECT 1188.340 999.870 1189.250 1000.000 ;
        RECT 1189.720 999.870 1191.090 1000.000 ;
      LAYER met2 ;
        RECT 1183.090 995.720 1184.090 998.470 ;
      LAYER met2 ;
        RECT 1184.370 996.000 1184.650 999.870 ;
      LAYER met2 ;
        RECT 1184.930 995.720 1186.390 998.470 ;
      LAYER met2 ;
        RECT 1186.670 996.000 1186.950 999.870 ;
      LAYER met2 ;
        RECT 1187.230 995.720 1188.690 998.470 ;
      LAYER met2 ;
        RECT 1188.970 996.000 1189.250 999.870 ;
      LAYER met2 ;
        RECT 1189.530 995.720 1190.530 998.470 ;
      LAYER met2 ;
        RECT 1190.810 996.000 1191.090 999.870 ;
        RECT 1193.110 999.870 1193.540 1000.000 ;
        RECT 1195.410 999.870 1197.220 1000.000 ;
        RECT 1197.710 999.870 1198.140 1000.000 ;
        RECT 1199.550 999.870 1200.440 1000.000 ;
        RECT 1201.850 999.870 1203.660 1000.000 ;
        RECT 1204.150 999.870 1204.580 1000.000 ;
        RECT 1204.900 1000.010 1205.040 1008.110 ;
        RECT 1209.900 1007.770 1210.160 1008.090 ;
        RECT 1209.960 1000.010 1210.100 1007.770 ;
        RECT 1210.360 1007.430 1210.620 1007.750 ;
        RECT 1204.900 1000.000 1206.120 1000.010 ;
        RECT 1208.420 1000.000 1210.100 1000.010 ;
        RECT 1204.900 999.870 1206.270 1000.000 ;
      LAYER met2 ;
        RECT 1191.370 995.720 1192.830 998.470 ;
      LAYER met2 ;
        RECT 1193.110 996.000 1193.390 999.870 ;
      LAYER met2 ;
        RECT 1193.670 995.720 1195.130 998.470 ;
      LAYER met2 ;
        RECT 1195.410 996.000 1195.690 999.870 ;
      LAYER met2 ;
        RECT 1195.970 995.720 1197.430 998.470 ;
      LAYER met2 ;
        RECT 1197.710 996.000 1197.990 999.870 ;
      LAYER met2 ;
        RECT 1198.270 995.720 1199.270 998.470 ;
      LAYER met2 ;
        RECT 1199.550 996.000 1199.830 999.870 ;
      LAYER met2 ;
        RECT 1200.110 995.720 1201.570 998.470 ;
      LAYER met2 ;
        RECT 1201.850 996.000 1202.130 999.870 ;
      LAYER met2 ;
        RECT 1202.410 995.720 1203.870 998.470 ;
      LAYER met2 ;
        RECT 1204.150 996.000 1204.430 999.870 ;
      LAYER met2 ;
        RECT 1204.710 995.720 1205.710 998.470 ;
      LAYER met2 ;
        RECT 1205.990 996.000 1206.270 999.870 ;
        RECT 1208.290 999.870 1210.100 1000.000 ;
        RECT 1210.420 1000.010 1210.560 1007.430 ;
        RECT 1213.640 1000.010 1213.780 1012.870 ;
        RECT 1214.100 1008.090 1214.240 1689.130 ;
        RECT 1215.480 1684.690 1215.620 1700.000 ;
        RECT 1221.400 1689.470 1221.660 1689.790 ;
        RECT 1217.720 1688.790 1217.980 1689.110 ;
        RECT 1215.420 1684.370 1215.680 1684.690 ;
        RECT 1214.500 1013.890 1214.760 1014.210 ;
        RECT 1214.040 1007.770 1214.300 1008.090 ;
        RECT 1210.420 1000.000 1210.720 1000.010 ;
        RECT 1213.020 1000.000 1213.780 1000.010 ;
        RECT 1210.420 999.870 1210.870 1000.000 ;
      LAYER met2 ;
        RECT 1206.550 995.720 1208.010 998.470 ;
      LAYER met2 ;
        RECT 1208.290 996.000 1208.570 999.870 ;
      LAYER met2 ;
        RECT 1208.850 995.720 1210.310 998.470 ;
      LAYER met2 ;
        RECT 1210.590 996.000 1210.870 999.870 ;
        RECT 1212.890 999.870 1213.780 1000.000 ;
        RECT 1214.560 1000.010 1214.700 1013.890 ;
        RECT 1217.260 1011.510 1217.520 1011.830 ;
        RECT 1217.320 1000.010 1217.460 1011.510 ;
        RECT 1217.780 1009.790 1217.920 1688.790 ;
        RECT 1221.460 1642.530 1221.600 1689.470 ;
        RECT 1230.200 1689.110 1230.340 1700.000 ;
        RECT 1234.740 1694.230 1235.000 1694.550 ;
        RECT 1230.140 1688.790 1230.400 1689.110 ;
        RECT 1221.400 1642.210 1221.660 1642.530 ;
        RECT 1223.240 1021.030 1223.500 1021.350 ;
        RECT 1218.640 1013.210 1218.900 1013.530 ;
        RECT 1218.700 1012.510 1218.840 1013.210 ;
        RECT 1218.180 1012.190 1218.440 1012.510 ;
        RECT 1218.640 1012.190 1218.900 1012.510 ;
        RECT 1221.400 1012.190 1221.660 1012.510 ;
        RECT 1217.720 1009.470 1217.980 1009.790 ;
        RECT 1214.560 1000.000 1214.860 1000.010 ;
        RECT 1217.160 1000.000 1217.460 1000.010 ;
        RECT 1214.560 999.870 1215.010 1000.000 ;
      LAYER met2 ;
        RECT 1211.150 995.720 1212.610 998.470 ;
      LAYER met2 ;
        RECT 1212.890 996.000 1213.170 999.870 ;
      LAYER met2 ;
        RECT 1213.450 995.720 1214.450 998.470 ;
      LAYER met2 ;
        RECT 1214.730 996.000 1215.010 999.870 ;
        RECT 1217.030 999.870 1217.460 1000.000 ;
        RECT 1218.240 1000.010 1218.380 1012.190 ;
        RECT 1221.460 1010.470 1221.600 1012.190 ;
        RECT 1221.400 1010.150 1221.660 1010.470 ;
        RECT 1222.780 1007.770 1223.040 1008.090 ;
        RECT 1222.840 1000.010 1222.980 1007.770 ;
        RECT 1218.240 1000.000 1219.460 1000.010 ;
        RECT 1221.300 1000.000 1222.980 1000.010 ;
        RECT 1218.240 999.870 1219.610 1000.000 ;
      LAYER met2 ;
        RECT 1215.290 995.720 1216.750 998.470 ;
      LAYER met2 ;
        RECT 1217.030 996.000 1217.310 999.870 ;
      LAYER met2 ;
        RECT 1217.590 995.720 1219.050 998.470 ;
      LAYER met2 ;
        RECT 1219.330 996.000 1219.610 999.870 ;
        RECT 1221.170 999.870 1222.980 1000.000 ;
        RECT 1223.300 1000.010 1223.440 1021.030 ;
        RECT 1228.300 1020.690 1228.560 1021.010 ;
        RECT 1224.160 1010.150 1224.420 1010.470 ;
        RECT 1224.220 1000.010 1224.360 1010.150 ;
        RECT 1228.360 1000.010 1228.500 1020.690 ;
        RECT 1230.600 1009.810 1230.860 1010.130 ;
        RECT 1228.760 1009.130 1229.020 1009.450 ;
        RECT 1223.300 1000.000 1223.600 1000.010 ;
        RECT 1224.220 1000.000 1225.900 1000.010 ;
        RECT 1228.200 1000.000 1228.500 1000.010 ;
        RECT 1223.300 999.870 1223.750 1000.000 ;
        RECT 1224.220 999.870 1226.050 1000.000 ;
      LAYER met2 ;
        RECT 1219.890 995.720 1220.890 998.470 ;
      LAYER met2 ;
        RECT 1221.170 996.000 1221.450 999.870 ;
      LAYER met2 ;
        RECT 1221.730 995.720 1223.190 998.470 ;
      LAYER met2 ;
        RECT 1223.470 996.000 1223.750 999.870 ;
      LAYER met2 ;
        RECT 1224.030 995.720 1225.490 998.470 ;
      LAYER met2 ;
        RECT 1225.770 996.000 1226.050 999.870 ;
        RECT 1228.070 999.870 1228.500 1000.000 ;
        RECT 1228.820 1000.010 1228.960 1009.130 ;
        RECT 1230.660 1000.010 1230.800 1009.810 ;
        RECT 1234.800 1000.010 1234.940 1694.230 ;
        RECT 1237.040 1686.410 1237.300 1686.730 ;
        RECT 1237.100 1048.890 1237.240 1686.410 ;
        RECT 1244.000 1684.350 1244.140 1700.000 ;
        RECT 1248.080 1688.790 1248.340 1689.110 ;
        RECT 1238.420 1684.030 1238.680 1684.350 ;
        RECT 1243.940 1684.030 1244.200 1684.350 ;
        RECT 1237.040 1048.570 1237.300 1048.890 ;
        RECT 1238.480 1014.210 1238.620 1684.030 ;
        RECT 1243.940 1642.210 1244.200 1642.530 ;
        RECT 1239.340 1048.570 1239.600 1048.890 ;
        RECT 1238.420 1013.890 1238.680 1014.210 ;
        RECT 1237.040 1012.190 1237.300 1012.510 ;
        RECT 1237.100 1009.530 1237.240 1012.190 ;
        RECT 1236.640 1009.390 1237.240 1009.530 ;
        RECT 1236.640 1000.010 1236.780 1009.390 ;
        RECT 1237.040 1008.790 1237.300 1009.110 ;
        RECT 1228.820 1000.000 1230.040 1000.010 ;
        RECT 1230.660 1000.000 1232.340 1000.010 ;
        RECT 1234.640 1000.000 1234.940 1000.010 ;
        RECT 1236.480 1000.000 1236.780 1000.010 ;
        RECT 1228.820 999.870 1230.190 1000.000 ;
        RECT 1230.660 999.870 1232.490 1000.000 ;
      LAYER met2 ;
        RECT 1226.330 995.720 1227.790 998.470 ;
      LAYER met2 ;
        RECT 1228.070 996.000 1228.350 999.870 ;
      LAYER met2 ;
        RECT 1228.630 995.720 1229.630 998.470 ;
      LAYER met2 ;
        RECT 1229.910 996.000 1230.190 999.870 ;
      LAYER met2 ;
        RECT 1230.470 995.720 1231.930 998.470 ;
      LAYER met2 ;
        RECT 1232.210 996.000 1232.490 999.870 ;
        RECT 1234.510 999.870 1234.940 1000.000 ;
        RECT 1236.350 999.870 1236.780 1000.000 ;
        RECT 1237.100 1000.010 1237.240 1008.790 ;
        RECT 1239.400 1000.010 1239.540 1048.570 ;
        RECT 1243.480 1020.690 1243.740 1021.010 ;
        RECT 1243.540 1000.010 1243.680 1020.690 ;
        RECT 1244.000 1014.290 1244.140 1642.210 ;
        RECT 1244.000 1014.150 1244.600 1014.290 ;
        RECT 1237.100 1000.000 1238.780 1000.010 ;
        RECT 1239.400 1000.000 1241.080 1000.010 ;
        RECT 1243.380 1000.000 1243.680 1000.010 ;
        RECT 1237.100 999.870 1238.930 1000.000 ;
        RECT 1239.400 999.870 1241.230 1000.000 ;
      LAYER met2 ;
        RECT 1232.770 995.720 1234.230 998.470 ;
      LAYER met2 ;
        RECT 1234.510 996.000 1234.790 999.870 ;
      LAYER met2 ;
        RECT 1235.070 995.720 1236.070 998.470 ;
      LAYER met2 ;
        RECT 1236.350 996.000 1236.630 999.870 ;
      LAYER met2 ;
        RECT 1236.910 995.720 1238.370 998.470 ;
      LAYER met2 ;
        RECT 1238.650 996.000 1238.930 999.870 ;
      LAYER met2 ;
        RECT 1239.210 995.720 1240.670 998.470 ;
      LAYER met2 ;
        RECT 1240.950 996.000 1241.230 999.870 ;
        RECT 1243.250 999.870 1243.680 1000.000 ;
        RECT 1244.460 1000.010 1244.600 1014.150 ;
        RECT 1245.320 1011.170 1245.580 1011.490 ;
        RECT 1245.380 1008.770 1245.520 1011.170 ;
        RECT 1245.320 1008.450 1245.580 1008.770 ;
        RECT 1248.140 1000.010 1248.280 1688.790 ;
        RECT 1250.840 1021.030 1251.100 1021.350 ;
        RECT 1250.900 1000.010 1251.040 1021.030 ;
        RECT 1258.200 1020.010 1258.460 1020.330 ;
        RECT 1257.740 1016.610 1258.000 1016.930 ;
        RECT 1255.440 1013.890 1255.700 1014.210 ;
        RECT 1253.140 1012.870 1253.400 1013.190 ;
        RECT 1253.200 1000.010 1253.340 1012.870 ;
        RECT 1255.500 1000.010 1255.640 1013.890 ;
        RECT 1257.800 1000.010 1257.940 1016.610 ;
        RECT 1244.460 1000.000 1245.220 1000.010 ;
        RECT 1247.520 1000.000 1248.280 1000.010 ;
        RECT 1249.820 1000.000 1251.040 1000.010 ;
        RECT 1251.660 1000.000 1253.340 1000.010 ;
        RECT 1253.960 1000.000 1255.640 1000.010 ;
        RECT 1256.260 1000.000 1257.940 1000.010 ;
        RECT 1244.460 999.870 1245.370 1000.000 ;
      LAYER met2 ;
        RECT 1241.510 995.720 1242.970 998.470 ;
      LAYER met2 ;
        RECT 1243.250 996.000 1243.530 999.870 ;
      LAYER met2 ;
        RECT 1243.810 995.720 1244.810 998.470 ;
      LAYER met2 ;
        RECT 1245.090 996.000 1245.370 999.870 ;
        RECT 1247.390 999.870 1248.280 1000.000 ;
        RECT 1249.690 999.870 1251.040 1000.000 ;
        RECT 1251.530 999.870 1253.340 1000.000 ;
        RECT 1253.830 999.870 1255.640 1000.000 ;
        RECT 1256.130 999.870 1257.940 1000.000 ;
        RECT 1258.260 1000.010 1258.400 1020.010 ;
        RECT 1261.420 1013.550 1261.680 1013.870 ;
        RECT 1261.480 1000.010 1261.620 1013.550 ;
        RECT 1261.940 1008.430 1262.080 1700.270 ;
        RECT 1272.410 1700.000 1272.690 1704.000 ;
        RECT 1287.130 1700.000 1287.410 1704.000 ;
        RECT 1300.930 1700.000 1301.210 1704.000 ;
        RECT 1315.650 1700.000 1315.930 1704.000 ;
        RECT 1329.450 1700.410 1329.730 1704.000 ;
        RECT 1329.450 1700.270 1331.540 1700.410 ;
        RECT 1329.450 1700.000 1329.730 1700.270 ;
        RECT 1268.780 1689.470 1269.040 1689.790 ;
        RECT 1264.180 1688.110 1264.440 1688.430 ;
        RECT 1264.240 1642.530 1264.380 1688.110 ;
        RECT 1264.180 1642.210 1264.440 1642.530 ;
        RECT 1266.020 1020.350 1266.280 1020.670 ;
        RECT 1264.180 1008.450 1264.440 1008.770 ;
        RECT 1261.880 1008.110 1262.140 1008.430 ;
        RECT 1264.240 1000.010 1264.380 1008.450 ;
        RECT 1266.080 1000.010 1266.220 1020.350 ;
        RECT 1268.320 1020.010 1268.580 1020.330 ;
        RECT 1267.860 1009.470 1268.120 1009.790 ;
        RECT 1267.920 1000.010 1268.060 1009.470 ;
        RECT 1258.260 1000.000 1258.560 1000.010 ;
        RECT 1260.400 1000.000 1261.620 1000.010 ;
        RECT 1262.700 1000.000 1264.380 1000.010 ;
        RECT 1265.000 1000.000 1266.220 1000.010 ;
        RECT 1266.840 1000.000 1268.060 1000.010 ;
        RECT 1258.260 999.870 1258.710 1000.000 ;
      LAYER met2 ;
        RECT 1245.650 995.720 1247.110 998.470 ;
      LAYER met2 ;
        RECT 1247.390 996.000 1247.670 999.870 ;
      LAYER met2 ;
        RECT 1247.950 995.720 1249.410 998.470 ;
      LAYER met2 ;
        RECT 1249.690 996.000 1249.970 999.870 ;
      LAYER met2 ;
        RECT 1250.250 995.720 1251.250 998.470 ;
      LAYER met2 ;
        RECT 1251.530 996.000 1251.810 999.870 ;
      LAYER met2 ;
        RECT 1252.090 995.720 1253.550 998.470 ;
      LAYER met2 ;
        RECT 1253.830 996.000 1254.110 999.870 ;
      LAYER met2 ;
        RECT 1254.390 995.720 1255.850 998.470 ;
      LAYER met2 ;
        RECT 1256.130 996.000 1256.410 999.870 ;
      LAYER met2 ;
        RECT 1256.690 995.720 1258.150 998.470 ;
      LAYER met2 ;
        RECT 1258.430 996.000 1258.710 999.870 ;
        RECT 1260.270 999.870 1261.620 1000.000 ;
        RECT 1262.570 999.870 1264.380 1000.000 ;
        RECT 1264.870 999.870 1266.220 1000.000 ;
        RECT 1266.710 999.870 1268.060 1000.000 ;
        RECT 1268.380 1000.010 1268.520 1020.010 ;
        RECT 1268.840 1008.770 1268.980 1689.470 ;
        RECT 1272.520 1684.350 1272.660 1700.000 ;
        RECT 1287.240 1689.450 1287.380 1700.000 ;
        RECT 1289.940 1694.570 1290.200 1694.890 ;
        RECT 1287.180 1689.130 1287.440 1689.450 ;
        RECT 1272.460 1684.030 1272.720 1684.350 ;
        RECT 1276.600 1642.210 1276.860 1642.530 ;
        RECT 1276.140 1016.950 1276.400 1017.270 ;
        RECT 1272.920 1009.130 1273.180 1009.450 ;
        RECT 1268.780 1008.450 1269.040 1008.770 ;
        RECT 1272.980 1000.010 1273.120 1009.130 ;
        RECT 1274.760 1008.450 1275.020 1008.770 ;
        RECT 1274.820 1000.010 1274.960 1008.450 ;
        RECT 1276.200 1000.010 1276.340 1016.950 ;
        RECT 1276.660 1009.700 1276.800 1642.210 ;
        RECT 1286.260 1020.010 1286.520 1020.330 ;
        RECT 1283.500 1019.330 1283.760 1019.650 ;
        RECT 1283.040 1010.150 1283.300 1010.470 ;
        RECT 1276.660 1009.560 1279.100 1009.700 ;
        RECT 1278.440 1008.790 1278.700 1009.110 ;
        RECT 1278.500 1000.010 1278.640 1008.790 ;
        RECT 1268.380 1000.000 1269.140 1000.010 ;
        RECT 1271.440 1000.000 1273.120 1000.010 ;
        RECT 1273.740 1000.000 1274.960 1000.010 ;
        RECT 1275.580 1000.000 1276.340 1000.010 ;
        RECT 1277.880 1000.000 1278.640 1000.010 ;
        RECT 1268.380 999.870 1269.290 1000.000 ;
      LAYER met2 ;
        RECT 1258.990 995.720 1259.990 998.470 ;
      LAYER met2 ;
        RECT 1260.270 996.000 1260.550 999.870 ;
      LAYER met2 ;
        RECT 1260.830 995.720 1262.290 998.470 ;
      LAYER met2 ;
        RECT 1262.570 996.000 1262.850 999.870 ;
      LAYER met2 ;
        RECT 1263.130 995.720 1264.590 998.470 ;
      LAYER met2 ;
        RECT 1264.870 996.000 1265.150 999.870 ;
      LAYER met2 ;
        RECT 1265.430 995.720 1266.430 998.470 ;
      LAYER met2 ;
        RECT 1266.710 996.000 1266.990 999.870 ;
      LAYER met2 ;
        RECT 1267.270 995.720 1268.730 998.470 ;
      LAYER met2 ;
        RECT 1269.010 996.000 1269.290 999.870 ;
        RECT 1271.310 999.870 1273.120 1000.000 ;
        RECT 1273.610 999.870 1274.960 1000.000 ;
        RECT 1275.450 999.870 1276.340 1000.000 ;
        RECT 1277.750 999.870 1278.640 1000.000 ;
        RECT 1278.960 1000.010 1279.100 1009.560 ;
        RECT 1283.100 1000.010 1283.240 1010.150 ;
        RECT 1278.960 1000.000 1280.180 1000.010 ;
        RECT 1282.020 1000.000 1283.240 1000.010 ;
        RECT 1278.960 999.870 1280.330 1000.000 ;
      LAYER met2 ;
        RECT 1269.570 995.720 1271.030 998.470 ;
      LAYER met2 ;
        RECT 1271.310 996.000 1271.590 999.870 ;
      LAYER met2 ;
        RECT 1271.870 995.720 1273.330 998.470 ;
      LAYER met2 ;
        RECT 1273.610 996.000 1273.890 999.870 ;
      LAYER met2 ;
        RECT 1274.170 995.720 1275.170 998.470 ;
      LAYER met2 ;
        RECT 1275.450 996.000 1275.730 999.870 ;
      LAYER met2 ;
        RECT 1276.010 995.720 1277.470 998.470 ;
      LAYER met2 ;
        RECT 1277.750 996.000 1278.030 999.870 ;
      LAYER met2 ;
        RECT 1278.310 995.720 1279.770 998.470 ;
      LAYER met2 ;
        RECT 1280.050 996.000 1280.330 999.870 ;
        RECT 1281.890 999.870 1283.240 1000.000 ;
        RECT 1283.560 1000.010 1283.700 1019.330 ;
        RECT 1286.320 1016.930 1286.460 1020.010 ;
        RECT 1286.260 1016.610 1286.520 1016.930 ;
        RECT 1290.000 1013.530 1290.140 1694.570 ;
        RECT 1301.040 1689.110 1301.180 1700.000 ;
        RECT 1310.640 1692.190 1310.900 1692.510 ;
        RECT 1300.980 1688.790 1301.240 1689.110 ;
        RECT 1293.620 1688.450 1293.880 1688.770 ;
        RECT 1291.320 1684.030 1291.580 1684.350 ;
        RECT 1290.400 1019.670 1290.660 1019.990 ;
        RECT 1286.720 1013.210 1286.980 1013.530 ;
        RECT 1287.640 1013.210 1287.900 1013.530 ;
        RECT 1289.940 1013.210 1290.200 1013.530 ;
        RECT 1286.780 1011.830 1286.920 1013.210 ;
        RECT 1286.720 1011.510 1286.980 1011.830 ;
        RECT 1287.700 1000.010 1287.840 1013.210 ;
        RECT 1289.940 1010.830 1290.200 1011.150 ;
        RECT 1290.000 1000.010 1290.140 1010.830 ;
        RECT 1283.560 1000.000 1284.320 1000.010 ;
        RECT 1286.620 1000.000 1287.840 1000.010 ;
        RECT 1288.920 1000.000 1290.140 1000.010 ;
        RECT 1283.560 999.870 1284.470 1000.000 ;
      LAYER met2 ;
        RECT 1280.610 995.720 1281.610 998.470 ;
      LAYER met2 ;
        RECT 1281.890 996.000 1282.170 999.870 ;
      LAYER met2 ;
        RECT 1282.450 995.720 1283.910 998.470 ;
      LAYER met2 ;
        RECT 1284.190 996.000 1284.470 999.870 ;
        RECT 1286.490 999.870 1287.840 1000.000 ;
        RECT 1288.790 999.870 1290.140 1000.000 ;
        RECT 1290.460 1000.010 1290.600 1019.670 ;
        RECT 1291.380 1000.010 1291.520 1684.030 ;
        RECT 1293.680 1013.530 1293.820 1688.450 ;
        RECT 1300.060 1018.990 1300.320 1019.310 ;
        RECT 1297.300 1016.610 1297.560 1016.930 ;
        RECT 1293.620 1013.210 1293.880 1013.530 ;
        RECT 1294.080 1011.170 1294.340 1011.490 ;
        RECT 1293.620 1009.470 1293.880 1009.790 ;
        RECT 1293.680 1007.750 1293.820 1009.470 ;
        RECT 1293.620 1007.430 1293.880 1007.750 ;
        RECT 1294.140 1000.010 1294.280 1011.170 ;
        RECT 1297.360 1000.010 1297.500 1016.610 ;
        RECT 1297.760 1011.850 1298.020 1012.170 ;
        RECT 1290.460 1000.000 1290.760 1000.010 ;
        RECT 1291.380 1000.000 1293.060 1000.010 ;
        RECT 1294.140 1000.000 1295.360 1000.010 ;
        RECT 1297.200 1000.000 1297.500 1000.010 ;
        RECT 1290.460 999.870 1290.910 1000.000 ;
        RECT 1291.380 999.870 1293.210 1000.000 ;
        RECT 1294.140 999.870 1295.510 1000.000 ;
      LAYER met2 ;
        RECT 1284.750 995.720 1286.210 998.470 ;
      LAYER met2 ;
        RECT 1286.490 996.000 1286.770 999.870 ;
      LAYER met2 ;
        RECT 1287.050 995.720 1288.510 998.470 ;
      LAYER met2 ;
        RECT 1288.790 996.000 1289.070 999.870 ;
      LAYER met2 ;
        RECT 1289.350 995.720 1290.350 998.470 ;
      LAYER met2 ;
        RECT 1290.630 996.000 1290.910 999.870 ;
      LAYER met2 ;
        RECT 1291.190 995.720 1292.650 998.470 ;
      LAYER met2 ;
        RECT 1292.930 996.000 1293.210 999.870 ;
      LAYER met2 ;
        RECT 1293.490 995.720 1294.950 998.470 ;
      LAYER met2 ;
        RECT 1295.230 996.000 1295.510 999.870 ;
        RECT 1297.070 999.870 1297.500 1000.000 ;
        RECT 1297.820 1000.010 1297.960 1011.850 ;
        RECT 1300.120 1000.010 1300.260 1018.990 ;
        RECT 1304.200 1011.510 1304.460 1011.830 ;
        RECT 1304.660 1011.510 1304.920 1011.830 ;
        RECT 1304.260 1000.010 1304.400 1011.510 ;
        RECT 1304.720 1009.450 1304.860 1011.510 ;
        RECT 1307.880 1010.490 1308.140 1010.810 ;
        RECT 1307.420 1009.470 1307.680 1009.790 ;
        RECT 1304.660 1009.130 1304.920 1009.450 ;
        RECT 1307.480 1000.010 1307.620 1009.470 ;
        RECT 1297.820 1000.000 1299.500 1000.010 ;
        RECT 1300.120 1000.000 1301.800 1000.010 ;
        RECT 1304.100 1000.000 1304.400 1000.010 ;
        RECT 1305.940 1000.000 1307.620 1000.010 ;
        RECT 1297.820 999.870 1299.650 1000.000 ;
        RECT 1300.120 999.870 1301.950 1000.000 ;
      LAYER met2 ;
        RECT 1295.790 995.720 1296.790 998.470 ;
      LAYER met2 ;
        RECT 1297.070 996.000 1297.350 999.870 ;
      LAYER met2 ;
        RECT 1297.630 995.720 1299.090 998.470 ;
      LAYER met2 ;
        RECT 1299.370 996.000 1299.650 999.870 ;
      LAYER met2 ;
        RECT 1299.930 995.720 1301.390 998.470 ;
      LAYER met2 ;
        RECT 1301.670 996.000 1301.950 999.870 ;
        RECT 1303.970 999.870 1304.400 1000.000 ;
        RECT 1305.810 999.870 1307.620 1000.000 ;
        RECT 1307.940 1000.010 1308.080 1010.490 ;
        RECT 1310.700 1009.790 1310.840 1692.190 ;
        RECT 1315.760 1689.790 1315.900 1700.000 ;
        RECT 1315.700 1689.470 1315.960 1689.790 ;
        RECT 1331.400 1076.170 1331.540 1700.270 ;
        RECT 1330.940 1076.030 1331.540 1076.170 ;
        RECT 1330.940 1028.570 1331.080 1076.030 ;
        RECT 1330.480 1028.430 1331.080 1028.570 ;
        RECT 1312.940 1018.650 1313.200 1018.970 ;
        RECT 1311.100 1009.810 1311.360 1010.130 ;
        RECT 1311.560 1009.810 1311.820 1010.130 ;
        RECT 1310.640 1009.470 1310.900 1009.790 ;
        RECT 1310.180 1009.130 1310.440 1009.450 ;
        RECT 1310.240 1000.010 1310.380 1009.130 ;
        RECT 1311.160 1000.010 1311.300 1009.810 ;
        RECT 1311.620 1008.770 1311.760 1009.810 ;
        RECT 1311.560 1008.450 1311.820 1008.770 ;
        RECT 1313.000 1000.010 1313.140 1018.650 ;
        RECT 1324.900 1018.310 1325.160 1018.630 ;
        RECT 1318.000 1013.210 1318.260 1013.530 ;
        RECT 1315.240 1008.110 1315.500 1008.430 ;
        RECT 1315.300 1000.010 1315.440 1008.110 ;
        RECT 1318.060 1000.010 1318.200 1013.210 ;
        RECT 1324.440 1011.850 1324.700 1012.170 ;
        RECT 1322.600 1010.830 1322.860 1011.150 ;
        RECT 1322.660 1000.010 1322.800 1010.830 ;
        RECT 1324.500 1000.010 1324.640 1011.850 ;
        RECT 1307.940 1000.000 1308.240 1000.010 ;
        RECT 1310.240 1000.000 1310.540 1000.010 ;
        RECT 1311.160 1000.000 1312.380 1000.010 ;
        RECT 1313.000 1000.000 1314.680 1000.010 ;
        RECT 1315.300 1000.000 1316.980 1000.010 ;
        RECT 1318.060 1000.000 1319.280 1000.010 ;
        RECT 1321.120 1000.000 1322.800 1000.010 ;
        RECT 1323.420 1000.000 1324.640 1000.010 ;
        RECT 1307.940 999.870 1308.390 1000.000 ;
        RECT 1310.240 999.870 1310.690 1000.000 ;
        RECT 1311.160 999.870 1312.530 1000.000 ;
        RECT 1313.000 999.870 1314.830 1000.000 ;
        RECT 1315.300 999.870 1317.130 1000.000 ;
        RECT 1318.060 999.870 1319.430 1000.000 ;
      LAYER met2 ;
        RECT 1302.230 995.720 1303.690 998.470 ;
      LAYER met2 ;
        RECT 1303.970 996.000 1304.250 999.870 ;
      LAYER met2 ;
        RECT 1304.530 995.720 1305.530 998.470 ;
      LAYER met2 ;
        RECT 1305.810 996.000 1306.090 999.870 ;
      LAYER met2 ;
        RECT 1306.370 995.720 1307.830 998.470 ;
      LAYER met2 ;
        RECT 1308.110 996.000 1308.390 999.870 ;
      LAYER met2 ;
        RECT 1308.670 995.720 1310.130 998.470 ;
      LAYER met2 ;
        RECT 1310.410 996.000 1310.690 999.870 ;
      LAYER met2 ;
        RECT 1310.970 995.720 1311.970 998.470 ;
      LAYER met2 ;
        RECT 1312.250 996.000 1312.530 999.870 ;
      LAYER met2 ;
        RECT 1312.810 995.720 1314.270 998.470 ;
      LAYER met2 ;
        RECT 1314.550 996.000 1314.830 999.870 ;
      LAYER met2 ;
        RECT 1315.110 995.720 1316.570 998.470 ;
      LAYER met2 ;
        RECT 1316.850 996.000 1317.130 999.870 ;
      LAYER met2 ;
        RECT 1317.410 995.720 1318.870 998.470 ;
      LAYER met2 ;
        RECT 1319.150 996.000 1319.430 999.870 ;
        RECT 1320.990 999.870 1322.800 1000.000 ;
        RECT 1323.290 999.870 1324.640 1000.000 ;
        RECT 1324.960 1000.010 1325.100 1018.310 ;
        RECT 1328.120 1010.490 1328.380 1010.810 ;
        RECT 1328.180 1000.010 1328.320 1010.490 ;
        RECT 1330.480 1008.430 1330.620 1028.430 ;
        RECT 1331.340 1013.890 1331.600 1014.210 ;
        RECT 1330.420 1008.110 1330.680 1008.430 ;
        RECT 1331.400 1000.010 1331.540 1013.890 ;
        RECT 1332.780 1011.830 1332.920 2054.290 ;
        RECT 1335.020 2053.270 1335.280 2053.590 ;
        RECT 1333.180 2052.250 1333.440 2052.570 ;
        RECT 1333.240 1014.550 1333.380 2052.250 ;
        RECT 1333.640 2050.550 1333.900 2050.870 ;
        RECT 1333.180 1014.230 1333.440 1014.550 ;
        RECT 1332.720 1011.510 1332.980 1011.830 ;
        RECT 1333.180 1011.510 1333.440 1011.830 ;
        RECT 1333.240 1000.010 1333.380 1011.510 ;
        RECT 1333.700 1007.750 1333.840 2050.550 ;
        RECT 1334.090 1997.995 1334.370 1998.365 ;
        RECT 1334.160 1012.170 1334.300 1997.995 ;
        RECT 1334.550 1787.195 1334.830 1787.565 ;
        RECT 1334.620 1014.210 1334.760 1787.195 ;
        RECT 1334.560 1013.890 1334.820 1014.210 ;
        RECT 1334.100 1011.850 1334.360 1012.170 ;
        RECT 1334.560 1011.850 1334.820 1012.170 ;
        RECT 1334.620 1009.790 1334.760 1011.850 ;
        RECT 1334.560 1009.470 1334.820 1009.790 ;
        RECT 1335.080 1007.750 1335.220 2053.270 ;
        RECT 1335.540 1694.550 1335.680 2054.630 ;
        RECT 1335.940 2051.910 1336.200 2052.230 ;
        RECT 1335.480 1694.230 1335.740 1694.550 ;
        RECT 1336.000 1694.210 1336.140 2051.910 ;
        RECT 1345.600 2051.570 1345.860 2051.890 ;
        RECT 1337.780 2050.210 1338.040 2050.530 ;
        RECT 1336.400 2049.190 1336.660 2049.510 ;
        RECT 1335.940 1693.890 1336.200 1694.210 ;
        RECT 1336.460 1693.870 1336.600 2049.190 ;
        RECT 1336.850 1745.035 1337.130 1745.405 ;
        RECT 1336.400 1693.550 1336.660 1693.870 ;
        RECT 1335.480 1017.970 1335.740 1018.290 ;
        RECT 1333.640 1007.430 1333.900 1007.750 ;
        RECT 1335.020 1007.430 1335.280 1007.750 ;
        RECT 1335.540 1000.010 1335.680 1017.970 ;
        RECT 1336.920 1016.930 1337.060 1745.035 ;
        RECT 1337.310 1724.635 1337.590 1725.005 ;
        RECT 1337.380 1020.670 1337.520 1724.635 ;
        RECT 1337.320 1020.350 1337.580 1020.670 ;
        RECT 1336.860 1016.610 1337.120 1016.930 ;
        RECT 1337.840 1000.010 1337.980 2050.210 ;
        RECT 1343.760 2036.270 1344.020 2036.590 ;
        RECT 1338.690 2018.395 1338.970 2018.765 ;
        RECT 1338.760 1020.330 1338.900 2018.395 ;
        RECT 1339.150 1976.235 1339.430 1976.605 ;
        RECT 1339.220 1021.350 1339.360 1976.235 ;
        RECT 1339.610 1955.835 1339.890 1956.205 ;
        RECT 1339.160 1021.030 1339.420 1021.350 ;
        RECT 1338.700 1020.010 1338.960 1020.330 ;
        RECT 1338.700 1013.890 1338.960 1014.210 ;
        RECT 1338.760 1000.010 1338.900 1013.890 ;
        RECT 1339.680 1008.770 1339.820 1955.835 ;
        RECT 1340.070 1934.075 1340.350 1934.445 ;
        RECT 1340.140 1012.510 1340.280 1934.075 ;
        RECT 1340.530 1913.675 1340.810 1914.045 ;
        RECT 1340.600 1017.270 1340.740 1913.675 ;
        RECT 1340.990 1891.915 1341.270 1892.285 ;
        RECT 1341.060 1021.010 1341.200 1891.915 ;
        RECT 1341.450 1871.515 1341.730 1871.885 ;
        RECT 1341.000 1020.690 1341.260 1021.010 ;
        RECT 1340.540 1016.950 1340.800 1017.270 ;
        RECT 1341.520 1013.870 1341.660 1871.515 ;
        RECT 1341.910 1849.755 1342.190 1850.125 ;
        RECT 1341.460 1013.550 1341.720 1013.870 ;
        RECT 1340.080 1012.190 1340.340 1012.510 ;
        RECT 1341.980 1010.130 1342.120 1849.755 ;
        RECT 1342.370 1829.355 1342.650 1829.725 ;
        RECT 1341.920 1009.810 1342.180 1010.130 ;
        RECT 1342.440 1009.450 1342.580 1829.355 ;
        RECT 1342.830 1807.595 1343.110 1807.965 ;
        RECT 1342.380 1009.130 1342.640 1009.450 ;
        RECT 1339.620 1008.450 1339.880 1008.770 ;
        RECT 1340.540 1007.430 1340.800 1007.750 ;
        RECT 1324.960 1000.000 1325.720 1000.010 ;
        RECT 1327.560 1000.000 1328.320 1000.010 ;
        RECT 1329.860 1000.000 1331.540 1000.010 ;
        RECT 1332.160 1000.000 1333.380 1000.010 ;
        RECT 1334.460 1000.000 1335.680 1000.010 ;
        RECT 1336.300 1000.000 1337.980 1000.010 ;
        RECT 1338.600 1000.000 1338.900 1000.010 ;
        RECT 1324.960 999.870 1325.870 1000.000 ;
      LAYER met2 ;
        RECT 1319.710 995.720 1320.710 998.470 ;
      LAYER met2 ;
        RECT 1320.990 996.000 1321.270 999.870 ;
      LAYER met2 ;
        RECT 1321.550 995.720 1323.010 998.470 ;
      LAYER met2 ;
        RECT 1323.290 996.000 1323.570 999.870 ;
      LAYER met2 ;
        RECT 1323.850 995.720 1325.310 998.470 ;
      LAYER met2 ;
        RECT 1325.590 996.000 1325.870 999.870 ;
        RECT 1327.430 999.870 1328.320 1000.000 ;
        RECT 1329.730 999.870 1331.540 1000.000 ;
        RECT 1332.030 999.870 1333.380 1000.000 ;
        RECT 1334.330 999.870 1335.680 1000.000 ;
        RECT 1336.170 999.870 1337.980 1000.000 ;
        RECT 1338.470 999.870 1338.900 1000.000 ;
        RECT 1340.600 1000.010 1340.740 1007.430 ;
        RECT 1342.900 1000.010 1343.040 1807.595 ;
        RECT 1343.290 1766.795 1343.570 1767.165 ;
        RECT 1343.360 1017.610 1343.500 1766.795 ;
        RECT 1343.820 1692.510 1343.960 2036.270 ;
        RECT 1343.760 1692.190 1344.020 1692.510 ;
        RECT 1343.300 1017.290 1343.560 1017.610 ;
        RECT 1345.660 1013.190 1345.800 2051.570 ;
        RECT 1345.600 1012.870 1345.860 1013.190 ;
        RECT 1346.120 1011.150 1346.260 2055.310 ;
        RECT 1346.520 2054.970 1346.780 2055.290 ;
        RECT 1346.580 1012.850 1346.720 2054.970 ;
        RECT 1346.980 2053.610 1347.240 2053.930 ;
        RECT 1346.520 1012.530 1346.780 1012.850 ;
        RECT 1347.040 1011.490 1347.180 2053.610 ;
        RECT 1352.100 2052.910 1352.240 2076.990 ;
        RECT 1352.960 2053.950 1353.220 2054.270 ;
        RECT 1347.440 2052.590 1347.700 2052.910 ;
        RECT 1350.200 2052.590 1350.460 2052.910 ;
        RECT 1352.040 2052.590 1352.300 2052.910 ;
        RECT 1346.980 1011.170 1347.240 1011.490 ;
        RECT 1346.060 1010.830 1346.320 1011.150 ;
        RECT 1347.500 1010.810 1347.640 2052.590 ;
        RECT 1347.900 2049.530 1348.160 2049.850 ;
        RECT 1347.960 1694.890 1348.100 2049.530 ;
        RECT 1350.260 2029.110 1350.400 2052.590 ;
        RECT 1352.500 2051.230 1352.760 2051.550 ;
        RECT 1350.200 2028.790 1350.460 2029.110 ;
        RECT 1352.040 2028.850 1352.300 2029.110 ;
        RECT 1351.640 2028.790 1352.300 2028.850 ;
        RECT 1351.640 2028.710 1352.240 2028.790 ;
        RECT 1351.640 2028.430 1351.780 2028.710 ;
        RECT 1350.200 2028.110 1350.460 2028.430 ;
        RECT 1351.580 2028.110 1351.840 2028.430 ;
        RECT 1350.260 1980.830 1350.400 2028.110 ;
        RECT 1350.200 1980.510 1350.460 1980.830 ;
        RECT 1350.660 1980.510 1350.920 1980.830 ;
        RECT 1350.720 1980.150 1350.860 1980.510 ;
        RECT 1350.200 1979.830 1350.460 1980.150 ;
        RECT 1350.660 1979.830 1350.920 1980.150 ;
        RECT 1350.260 1932.210 1350.400 1979.830 ;
        RECT 1350.200 1931.890 1350.460 1932.210 ;
        RECT 1351.120 1931.890 1351.380 1932.210 ;
        RECT 1351.180 1908.070 1351.320 1931.890 ;
        RECT 1351.120 1907.750 1351.380 1908.070 ;
        RECT 1352.040 1907.750 1352.300 1908.070 ;
        RECT 1352.100 1884.125 1352.240 1907.750 ;
        RECT 1352.030 1883.755 1352.310 1884.125 ;
        RECT 1350.190 1882.395 1350.470 1882.765 ;
        RECT 1350.260 1835.650 1350.400 1882.395 ;
        RECT 1350.200 1835.330 1350.460 1835.650 ;
        RECT 1351.120 1835.330 1351.380 1835.650 ;
        RECT 1351.180 1801.310 1351.320 1835.330 ;
        RECT 1351.120 1800.990 1351.380 1801.310 ;
        RECT 1351.580 1800.650 1351.840 1800.970 ;
        RECT 1351.640 1787.030 1351.780 1800.650 ;
        RECT 1350.200 1786.710 1350.460 1787.030 ;
        RECT 1351.580 1786.710 1351.840 1787.030 ;
        RECT 1350.260 1780.230 1350.400 1786.710 ;
        RECT 1350.200 1779.910 1350.460 1780.230 ;
        RECT 1350.660 1779.910 1350.920 1780.230 ;
        RECT 1350.720 1732.290 1350.860 1779.910 ;
        RECT 1350.660 1731.970 1350.920 1732.290 ;
        RECT 1352.040 1731.970 1352.300 1732.290 ;
        RECT 1352.100 1725.150 1352.240 1731.970 ;
        RECT 1350.660 1724.830 1350.920 1725.150 ;
        RECT 1352.040 1724.830 1352.300 1725.150 ;
        RECT 1347.900 1694.570 1348.160 1694.890 ;
        RECT 1350.720 1676.870 1350.860 1724.830 ;
        RECT 1350.660 1676.550 1350.920 1676.870 ;
        RECT 1351.120 1676.550 1351.380 1676.870 ;
        RECT 1351.180 1642.530 1351.320 1676.550 ;
        RECT 1351.120 1642.210 1351.380 1642.530 ;
        RECT 1351.580 1642.210 1351.840 1642.530 ;
        RECT 1351.640 1641.930 1351.780 1642.210 ;
        RECT 1351.180 1641.790 1351.780 1641.930 ;
        RECT 1351.180 1608.045 1351.320 1641.790 ;
        RECT 1351.110 1607.675 1351.390 1608.045 ;
        RECT 1351.570 1606.995 1351.850 1607.365 ;
        RECT 1351.640 1593.910 1351.780 1606.995 ;
        RECT 1350.200 1593.590 1350.460 1593.910 ;
        RECT 1351.580 1593.590 1351.840 1593.910 ;
        RECT 1350.260 1546.310 1350.400 1593.590 ;
        RECT 1350.200 1545.990 1350.460 1546.310 ;
        RECT 1351.580 1545.990 1351.840 1546.310 ;
        RECT 1351.640 1545.630 1351.780 1545.990 ;
        RECT 1350.660 1545.310 1350.920 1545.630 ;
        RECT 1351.580 1545.310 1351.840 1545.630 ;
        RECT 1350.720 1510.950 1350.860 1545.310 ;
        RECT 1350.660 1510.630 1350.920 1510.950 ;
        RECT 1351.580 1510.630 1351.840 1510.950 ;
        RECT 1351.640 1497.350 1351.780 1510.630 ;
        RECT 1350.200 1497.030 1350.460 1497.350 ;
        RECT 1351.580 1497.030 1351.840 1497.350 ;
        RECT 1350.260 1449.750 1350.400 1497.030 ;
        RECT 1350.200 1449.430 1350.460 1449.750 ;
        RECT 1351.580 1449.430 1351.840 1449.750 ;
        RECT 1351.640 1449.070 1351.780 1449.430 ;
        RECT 1350.660 1448.750 1350.920 1449.070 ;
        RECT 1351.580 1448.750 1351.840 1449.070 ;
        RECT 1350.720 1414.390 1350.860 1448.750 ;
        RECT 1350.660 1414.070 1350.920 1414.390 ;
        RECT 1351.580 1414.070 1351.840 1414.390 ;
        RECT 1351.640 1400.790 1351.780 1414.070 ;
        RECT 1350.200 1400.470 1350.460 1400.790 ;
        RECT 1351.580 1400.470 1351.840 1400.790 ;
        RECT 1350.260 1352.850 1350.400 1400.470 ;
        RECT 1350.200 1352.530 1350.460 1352.850 ;
        RECT 1351.120 1352.530 1351.380 1352.850 ;
        RECT 1351.180 1328.450 1351.320 1352.530 ;
        RECT 1350.720 1328.310 1351.320 1328.450 ;
        RECT 1350.720 1317.830 1350.860 1328.310 ;
        RECT 1350.660 1317.510 1350.920 1317.830 ;
        RECT 1351.580 1317.510 1351.840 1317.830 ;
        RECT 1351.640 1304.230 1351.780 1317.510 ;
        RECT 1350.200 1303.910 1350.460 1304.230 ;
        RECT 1351.580 1303.910 1351.840 1304.230 ;
        RECT 1350.260 1256.630 1350.400 1303.910 ;
        RECT 1350.200 1256.310 1350.460 1256.630 ;
        RECT 1351.580 1255.970 1351.840 1256.290 ;
        RECT 1351.640 1255.805 1351.780 1255.970 ;
        RECT 1350.650 1255.435 1350.930 1255.805 ;
        RECT 1351.570 1255.435 1351.850 1255.805 ;
        RECT 1350.720 1207.670 1350.860 1255.435 ;
        RECT 1350.660 1207.350 1350.920 1207.670 ;
        RECT 1351.580 1207.525 1351.840 1207.670 ;
        RECT 1351.570 1207.155 1351.850 1207.525 ;
        RECT 1350.190 1206.475 1350.470 1206.845 ;
        RECT 1350.260 1159.390 1350.400 1206.475 ;
        RECT 1350.200 1159.070 1350.460 1159.390 ;
        RECT 1352.040 1159.070 1352.300 1159.390 ;
        RECT 1352.100 1111.110 1352.240 1159.070 ;
        RECT 1351.120 1110.790 1351.380 1111.110 ;
        RECT 1352.040 1110.790 1352.300 1111.110 ;
        RECT 1351.180 1077.110 1351.320 1110.790 ;
        RECT 1351.120 1076.790 1351.380 1077.110 ;
        RECT 1351.120 1075.770 1351.380 1076.090 ;
        RECT 1351.180 1028.570 1351.320 1075.770 ;
        RECT 1350.720 1028.430 1351.320 1028.570 ;
        RECT 1347.900 1017.630 1348.160 1017.950 ;
        RECT 1347.440 1010.490 1347.700 1010.810 ;
        RECT 1343.300 1008.110 1343.560 1008.430 ;
        RECT 1340.600 1000.000 1340.900 1000.010 ;
        RECT 1342.740 1000.000 1343.040 1000.010 ;
        RECT 1340.600 999.870 1341.050 1000.000 ;
      LAYER met2 ;
        RECT 1326.150 995.720 1327.150 998.470 ;
      LAYER met2 ;
        RECT 1327.430 996.000 1327.710 999.870 ;
      LAYER met2 ;
        RECT 1327.990 995.720 1329.450 998.470 ;
      LAYER met2 ;
        RECT 1329.730 996.000 1330.010 999.870 ;
      LAYER met2 ;
        RECT 1330.290 995.720 1331.750 998.470 ;
      LAYER met2 ;
        RECT 1332.030 996.000 1332.310 999.870 ;
      LAYER met2 ;
        RECT 1332.590 995.720 1334.050 998.470 ;
      LAYER met2 ;
        RECT 1334.330 996.000 1334.610 999.870 ;
      LAYER met2 ;
        RECT 1334.890 995.720 1335.890 998.470 ;
      LAYER met2 ;
        RECT 1336.170 996.000 1336.450 999.870 ;
      LAYER met2 ;
        RECT 1336.730 995.720 1338.190 998.470 ;
      LAYER met2 ;
        RECT 1338.470 996.000 1338.750 999.870 ;
      LAYER met2 ;
        RECT 1339.030 995.720 1340.490 998.470 ;
      LAYER met2 ;
        RECT 1340.770 996.000 1341.050 999.870 ;
        RECT 1342.610 999.870 1343.040 1000.000 ;
        RECT 1343.360 1000.010 1343.500 1008.110 ;
        RECT 1347.960 1000.010 1348.100 1017.630 ;
        RECT 1350.720 1000.010 1350.860 1028.430 ;
        RECT 1352.040 1017.630 1352.300 1017.950 ;
        RECT 1352.100 1000.010 1352.240 1017.630 ;
        RECT 1352.560 1010.470 1352.700 2051.230 ;
        RECT 1353.020 1012.170 1353.160 2053.950 ;
        RECT 1353.880 2052.930 1354.140 2053.250 ;
        RECT 1353.420 2050.890 1353.680 2051.210 ;
        RECT 1353.480 1014.210 1353.620 2050.890 ;
        RECT 1353.420 1013.890 1353.680 1014.210 ;
        RECT 1352.960 1011.850 1353.220 1012.170 ;
        RECT 1353.940 1011.830 1354.080 2052.930 ;
        RECT 1357.100 1018.310 1357.360 1018.630 ;
        RECT 1355.260 1013.890 1355.520 1014.210 ;
        RECT 1353.880 1011.510 1354.140 1011.830 ;
        RECT 1352.500 1010.150 1352.760 1010.470 ;
        RECT 1355.320 1000.010 1355.460 1013.890 ;
        RECT 1357.160 1000.010 1357.300 1018.310 ;
        RECT 1358.080 1014.210 1358.220 2849.550 ;
        RECT 1358.480 2780.870 1358.740 2781.190 ;
        RECT 1358.020 1013.890 1358.280 1014.210 ;
        RECT 1358.540 1000.010 1358.680 2780.870 ;
        RECT 1365.840 1735.030 1366.100 1735.350 ;
        RECT 1365.900 1000.010 1366.040 1735.030 ;
        RECT 1372.800 1008.770 1372.940 2913.130 ;
        RECT 1379.700 1010.810 1379.840 2914.830 ;
        RECT 1407.240 2914.490 1407.500 2914.810 ;
        RECT 1393.440 2608.150 1393.700 2608.470 ;
        RECT 1392.980 2594.550 1393.240 2594.870 ;
        RECT 1386.540 2485.410 1386.800 2485.730 ;
        RECT 1385.620 1024.430 1385.880 1024.750 ;
        RECT 1376.880 1010.490 1377.140 1010.810 ;
        RECT 1379.640 1010.490 1379.900 1010.810 ;
        RECT 1374.580 1009.810 1374.840 1010.130 ;
        RECT 1368.140 1008.450 1368.400 1008.770 ;
        RECT 1372.740 1008.450 1373.000 1008.770 ;
        RECT 1368.200 1000.010 1368.340 1008.450 ;
        RECT 1374.640 1000.010 1374.780 1009.810 ;
        RECT 1376.940 1000.010 1377.080 1010.490 ;
        RECT 1383.320 1008.450 1383.580 1008.770 ;
        RECT 1383.380 1000.010 1383.520 1008.450 ;
        RECT 1385.680 1000.010 1385.820 1024.430 ;
        RECT 1386.600 1008.770 1386.740 2485.410 ;
        RECT 1386.540 1008.450 1386.800 1008.770 ;
        RECT 1393.040 1000.690 1393.180 2594.550 ;
        RECT 1391.660 1000.550 1393.180 1000.690 ;
        RECT 1391.660 1000.010 1391.800 1000.550 ;
        RECT 1393.500 1000.010 1393.640 2608.150 ;
        RECT 1397.120 2485.070 1397.380 2485.390 ;
        RECT 1397.180 1010.130 1397.320 2485.070 ;
        RECT 1400.340 1017.970 1400.600 1018.290 ;
        RECT 1397.120 1009.810 1397.380 1010.130 ;
        RECT 1400.400 1000.010 1400.540 1017.970 ;
        RECT 1407.300 1010.130 1407.440 2914.490 ;
        RECT 1413.680 2580.610 1413.940 2580.930 ;
        RECT 1411.380 1012.190 1411.640 1012.510 ;
        RECT 1409.080 1010.490 1409.340 1010.810 ;
        RECT 1402.640 1009.810 1402.900 1010.130 ;
        RECT 1407.240 1009.810 1407.500 1010.130 ;
        RECT 1402.700 1000.010 1402.840 1009.810 ;
        RECT 1409.140 1000.010 1409.280 1010.490 ;
        RECT 1411.440 1000.010 1411.580 1012.190 ;
        RECT 1413.740 1010.810 1413.880 2580.610 ;
        RECT 1414.200 1012.510 1414.340 2916.870 ;
        RECT 1479.920 2915.510 1480.180 2915.830 ;
        RECT 1461.520 2914.150 1461.780 2914.470 ;
        RECT 1455.540 2900.890 1455.800 2901.210 ;
        RECT 1434.380 2691.110 1434.640 2691.430 ;
        RECT 1421.040 2488.470 1421.300 2488.790 ;
        RECT 1420.580 2487.790 1420.840 2488.110 ;
        RECT 1414.140 1012.190 1414.400 1012.510 ;
        RECT 1413.680 1010.490 1413.940 1010.810 ;
        RECT 1415.980 1010.490 1416.240 1010.810 ;
        RECT 1416.040 1000.010 1416.180 1010.490 ;
        RECT 1417.820 1007.430 1418.080 1007.750 ;
        RECT 1417.880 1000.010 1418.020 1007.430 ;
        RECT 1420.640 1000.690 1420.780 2487.790 ;
        RECT 1421.100 1007.750 1421.240 2488.470 ;
        RECT 1427.940 2486.090 1428.200 2486.410 ;
        RECT 1428.000 1011.570 1428.140 2486.090 ;
        RECT 1426.620 1011.430 1428.140 1011.570 ;
        RECT 1421.040 1007.430 1421.300 1007.750 ;
        RECT 1420.180 1000.550 1420.780 1000.690 ;
        RECT 1420.180 1000.010 1420.320 1000.550 ;
        RECT 1426.620 1000.010 1426.760 1011.430 ;
        RECT 1427.940 1010.830 1428.200 1011.150 ;
        RECT 1428.000 1000.010 1428.140 1010.830 ;
        RECT 1434.440 1000.690 1434.580 2691.110 ;
        RECT 1455.080 2488.130 1455.340 2488.450 ;
        RECT 1448.640 2486.770 1448.900 2487.090 ;
        RECT 1441.740 2484.730 1442.000 2485.050 ;
        RECT 1434.840 1018.650 1435.100 1018.970 ;
        RECT 1433.060 1000.550 1434.580 1000.690 ;
        RECT 1433.060 1000.010 1433.200 1000.550 ;
        RECT 1434.900 1000.010 1435.040 1018.650 ;
        RECT 1441.280 1011.850 1441.540 1012.170 ;
        RECT 1437.600 1007.430 1437.860 1007.750 ;
        RECT 1437.660 1000.010 1437.800 1007.430 ;
        RECT 1441.340 1000.010 1441.480 1011.850 ;
        RECT 1441.800 1007.750 1441.940 2484.730 ;
        RECT 1444.040 1011.170 1444.300 1011.490 ;
        RECT 1441.740 1007.430 1442.000 1007.750 ;
        RECT 1444.100 1000.010 1444.240 1011.170 ;
        RECT 1448.700 1007.750 1448.840 2486.770 ;
        RECT 1454.620 2486.430 1454.880 2486.750 ;
        RECT 1450.480 1007.770 1450.740 1008.090 ;
        RECT 1446.340 1007.430 1446.600 1007.750 ;
        RECT 1448.640 1007.430 1448.900 1007.750 ;
        RECT 1446.400 1000.010 1446.540 1007.430 ;
        RECT 1450.540 1000.010 1450.680 1007.770 ;
        RECT 1452.780 1007.430 1453.040 1007.750 ;
        RECT 1452.840 1000.010 1452.980 1007.430 ;
        RECT 1454.680 1000.010 1454.820 2486.430 ;
        RECT 1455.140 1008.090 1455.280 2488.130 ;
        RECT 1455.080 1007.770 1455.340 1008.090 ;
        RECT 1455.600 1007.750 1455.740 2900.890 ;
        RECT 1461.060 1007.770 1461.320 1008.090 ;
        RECT 1455.540 1007.430 1455.800 1007.750 ;
        RECT 1459.220 1007.430 1459.480 1007.750 ;
        RECT 1459.280 1000.010 1459.420 1007.430 ;
        RECT 1461.120 1000.010 1461.260 1007.770 ;
        RECT 1343.360 1000.000 1345.040 1000.010 ;
        RECT 1347.340 1000.000 1348.100 1000.010 ;
        RECT 1349.180 1000.000 1350.860 1000.010 ;
        RECT 1351.480 1000.000 1352.240 1000.010 ;
        RECT 1353.780 1000.000 1355.460 1000.010 ;
        RECT 1356.080 1000.000 1357.300 1000.010 ;
        RECT 1357.920 1000.000 1358.680 1000.010 ;
        RECT 1364.360 1000.000 1366.040 1000.010 ;
        RECT 1366.660 1000.000 1368.340 1000.010 ;
        RECT 1373.100 1000.000 1374.780 1000.010 ;
        RECT 1375.400 1000.000 1377.080 1000.010 ;
        RECT 1381.840 1000.000 1383.520 1000.010 ;
        RECT 1384.140 1000.000 1385.820 1000.010 ;
        RECT 1390.580 1000.000 1391.800 1000.010 ;
        RECT 1392.880 1000.000 1393.640 1000.010 ;
        RECT 1399.320 1000.000 1400.540 1000.010 ;
        RECT 1401.620 1000.000 1402.840 1000.010 ;
        RECT 1408.060 1000.000 1409.280 1000.010 ;
        RECT 1409.900 1000.000 1411.580 1000.010 ;
        RECT 1414.500 1000.000 1416.180 1000.010 ;
        RECT 1416.800 1000.000 1418.020 1000.010 ;
        RECT 1418.640 1000.000 1420.320 1000.010 ;
        RECT 1425.080 1000.000 1426.760 1000.010 ;
        RECT 1427.380 1000.000 1428.140 1000.010 ;
        RECT 1431.980 1000.000 1433.200 1000.010 ;
        RECT 1433.820 1000.000 1435.040 1000.010 ;
        RECT 1436.120 1000.000 1437.800 1000.010 ;
        RECT 1440.260 1000.000 1441.480 1000.010 ;
        RECT 1442.560 1000.000 1444.240 1000.010 ;
        RECT 1444.860 1000.000 1446.540 1000.010 ;
        RECT 1449.000 1000.000 1450.680 1000.010 ;
        RECT 1451.300 1000.000 1452.980 1000.010 ;
        RECT 1453.600 1000.000 1454.820 1000.010 ;
        RECT 1457.740 1000.000 1459.420 1000.010 ;
        RECT 1460.040 1000.000 1461.260 1000.010 ;
        RECT 1343.360 999.870 1345.190 1000.000 ;
      LAYER met2 ;
        RECT 1341.330 995.720 1342.330 998.470 ;
      LAYER met2 ;
        RECT 1342.610 996.000 1342.890 999.870 ;
      LAYER met2 ;
        RECT 1343.170 995.720 1344.630 998.470 ;
      LAYER met2 ;
        RECT 1344.910 996.000 1345.190 999.870 ;
        RECT 1347.210 999.870 1348.100 1000.000 ;
        RECT 1349.050 999.870 1350.860 1000.000 ;
        RECT 1351.350 999.870 1352.240 1000.000 ;
        RECT 1353.650 999.870 1355.460 1000.000 ;
        RECT 1355.950 999.870 1357.300 1000.000 ;
        RECT 1357.790 999.870 1358.680 1000.000 ;
      LAYER met2 ;
        RECT 1345.470 995.720 1346.930 998.470 ;
      LAYER met2 ;
        RECT 1347.210 996.000 1347.490 999.870 ;
      LAYER met2 ;
        RECT 1347.770 995.720 1348.770 998.470 ;
      LAYER met2 ;
        RECT 1349.050 996.000 1349.330 999.870 ;
      LAYER met2 ;
        RECT 1349.610 995.720 1351.070 998.470 ;
      LAYER met2 ;
        RECT 1351.350 996.000 1351.630 999.870 ;
      LAYER met2 ;
        RECT 1351.910 995.720 1353.370 998.470 ;
      LAYER met2 ;
        RECT 1353.650 996.000 1353.930 999.870 ;
      LAYER met2 ;
        RECT 1354.210 995.720 1355.670 998.470 ;
      LAYER met2 ;
        RECT 1355.950 996.000 1356.230 999.870 ;
      LAYER met2 ;
        RECT 1356.510 995.720 1357.510 998.470 ;
      LAYER met2 ;
        RECT 1357.790 996.000 1358.070 999.870 ;
      LAYER met2 ;
        RECT 1358.350 995.720 1359.810 998.470 ;
      LAYER met2 ;
        RECT 1360.090 996.000 1360.370 1000.000 ;
      LAYER met2 ;
        RECT 1360.650 995.720 1362.110 998.470 ;
      LAYER met2 ;
        RECT 1362.390 996.000 1362.670 1000.000 ;
        RECT 1364.230 999.870 1366.040 1000.000 ;
        RECT 1366.530 999.870 1368.340 1000.000 ;
      LAYER met2 ;
        RECT 1362.950 995.720 1363.950 998.470 ;
      LAYER met2 ;
        RECT 1364.230 996.000 1364.510 999.870 ;
      LAYER met2 ;
        RECT 1364.790 995.720 1366.250 998.470 ;
      LAYER met2 ;
        RECT 1366.530 996.000 1366.810 999.870 ;
      LAYER met2 ;
        RECT 1367.090 995.720 1368.550 998.470 ;
      LAYER met2 ;
        RECT 1368.830 996.000 1369.110 1000.000 ;
      LAYER met2 ;
        RECT 1369.390 995.720 1370.850 998.470 ;
      LAYER met2 ;
        RECT 1371.130 996.000 1371.410 1000.000 ;
        RECT 1372.970 999.870 1374.780 1000.000 ;
        RECT 1375.270 999.870 1377.080 1000.000 ;
      LAYER met2 ;
        RECT 1371.690 995.720 1372.690 998.470 ;
      LAYER met2 ;
        RECT 1372.970 996.000 1373.250 999.870 ;
      LAYER met2 ;
        RECT 1373.530 995.720 1374.990 998.470 ;
      LAYER met2 ;
        RECT 1375.270 996.000 1375.550 999.870 ;
      LAYER met2 ;
        RECT 1375.830 995.720 1377.290 998.470 ;
      LAYER met2 ;
        RECT 1377.570 996.000 1377.850 1000.000 ;
      LAYER met2 ;
        RECT 1378.130 995.720 1379.130 998.470 ;
      LAYER met2 ;
        RECT 1379.410 996.000 1379.690 1000.000 ;
        RECT 1381.710 999.870 1383.520 1000.000 ;
        RECT 1384.010 999.870 1385.820 1000.000 ;
      LAYER met2 ;
        RECT 1379.970 995.720 1381.430 998.470 ;
      LAYER met2 ;
        RECT 1381.710 996.000 1381.990 999.870 ;
      LAYER met2 ;
        RECT 1382.270 995.720 1383.730 998.470 ;
      LAYER met2 ;
        RECT 1384.010 996.000 1384.290 999.870 ;
      LAYER met2 ;
        RECT 1384.570 995.720 1386.030 998.470 ;
      LAYER met2 ;
        RECT 1386.310 996.000 1386.590 1000.000 ;
      LAYER met2 ;
        RECT 1386.870 995.720 1387.870 998.470 ;
      LAYER met2 ;
        RECT 1388.150 996.000 1388.430 1000.000 ;
        RECT 1390.450 999.870 1391.800 1000.000 ;
        RECT 1392.750 999.870 1393.640 1000.000 ;
      LAYER met2 ;
        RECT 1388.710 995.720 1390.170 998.470 ;
      LAYER met2 ;
        RECT 1390.450 996.000 1390.730 999.870 ;
      LAYER met2 ;
        RECT 1391.010 995.720 1392.470 998.470 ;
      LAYER met2 ;
        RECT 1392.750 996.000 1393.030 999.870 ;
      LAYER met2 ;
        RECT 1393.310 995.720 1394.310 998.470 ;
      LAYER met2 ;
        RECT 1394.590 996.000 1394.870 1000.000 ;
      LAYER met2 ;
        RECT 1395.150 995.720 1396.610 998.470 ;
      LAYER met2 ;
        RECT 1396.890 996.000 1397.170 1000.000 ;
        RECT 1399.190 999.870 1400.540 1000.000 ;
        RECT 1401.490 999.870 1402.840 1000.000 ;
      LAYER met2 ;
        RECT 1397.450 995.720 1398.910 998.470 ;
      LAYER met2 ;
        RECT 1399.190 996.000 1399.470 999.870 ;
      LAYER met2 ;
        RECT 1399.750 995.720 1401.210 998.470 ;
      LAYER met2 ;
        RECT 1401.490 996.000 1401.770 999.870 ;
      LAYER met2 ;
        RECT 1402.050 995.720 1403.050 998.470 ;
      LAYER met2 ;
        RECT 1403.330 996.000 1403.610 1000.000 ;
      LAYER met2 ;
        RECT 1403.890 995.720 1405.350 998.470 ;
      LAYER met2 ;
        RECT 1405.630 996.000 1405.910 1000.000 ;
        RECT 1407.930 999.870 1409.280 1000.000 ;
        RECT 1409.770 999.870 1411.580 1000.000 ;
      LAYER met2 ;
        RECT 1406.190 995.720 1407.650 998.470 ;
      LAYER met2 ;
        RECT 1407.930 996.000 1408.210 999.870 ;
      LAYER met2 ;
        RECT 1408.490 995.720 1409.490 998.470 ;
      LAYER met2 ;
        RECT 1409.770 996.000 1410.050 999.870 ;
      LAYER met2 ;
        RECT 1410.330 995.720 1411.790 998.470 ;
      LAYER met2 ;
        RECT 1412.070 996.000 1412.350 1000.000 ;
        RECT 1414.370 999.870 1416.180 1000.000 ;
        RECT 1416.670 999.870 1418.020 1000.000 ;
        RECT 1418.510 999.870 1420.320 1000.000 ;
      LAYER met2 ;
        RECT 1412.630 995.720 1414.090 998.470 ;
      LAYER met2 ;
        RECT 1414.370 996.000 1414.650 999.870 ;
      LAYER met2 ;
        RECT 1414.930 995.720 1416.390 998.470 ;
      LAYER met2 ;
        RECT 1416.670 996.000 1416.950 999.870 ;
      LAYER met2 ;
        RECT 1417.230 995.720 1418.230 998.470 ;
      LAYER met2 ;
        RECT 1418.510 996.000 1418.790 999.870 ;
      LAYER met2 ;
        RECT 1419.070 995.720 1420.530 998.470 ;
      LAYER met2 ;
        RECT 1420.810 996.000 1421.090 1000.000 ;
      LAYER met2 ;
        RECT 1421.370 995.720 1422.830 998.470 ;
      LAYER met2 ;
        RECT 1423.110 996.000 1423.390 1000.000 ;
        RECT 1424.950 999.870 1426.760 1000.000 ;
        RECT 1427.250 999.870 1428.140 1000.000 ;
      LAYER met2 ;
        RECT 1423.670 995.720 1424.670 998.470 ;
      LAYER met2 ;
        RECT 1424.950 996.000 1425.230 999.870 ;
      LAYER met2 ;
        RECT 1425.510 995.720 1426.970 998.470 ;
      LAYER met2 ;
        RECT 1427.250 996.000 1427.530 999.870 ;
      LAYER met2 ;
        RECT 1427.810 995.720 1429.270 998.470 ;
      LAYER met2 ;
        RECT 1429.550 996.000 1429.830 1000.000 ;
        RECT 1431.850 999.870 1433.200 1000.000 ;
        RECT 1433.690 999.870 1435.040 1000.000 ;
        RECT 1435.990 999.870 1437.800 1000.000 ;
      LAYER met2 ;
        RECT 1430.110 995.720 1431.570 998.470 ;
      LAYER met2 ;
        RECT 1431.850 996.000 1432.130 999.870 ;
      LAYER met2 ;
        RECT 1432.410 995.720 1433.410 998.470 ;
      LAYER met2 ;
        RECT 1433.690 996.000 1433.970 999.870 ;
      LAYER met2 ;
        RECT 1434.250 995.720 1435.710 998.470 ;
      LAYER met2 ;
        RECT 1435.990 996.000 1436.270 999.870 ;
      LAYER met2 ;
        RECT 1436.550 995.720 1438.010 998.470 ;
      LAYER met2 ;
        RECT 1438.290 996.000 1438.570 1000.000 ;
        RECT 1440.130 999.870 1441.480 1000.000 ;
        RECT 1442.430 999.870 1444.240 1000.000 ;
        RECT 1444.730 999.870 1446.540 1000.000 ;
      LAYER met2 ;
        RECT 1438.850 995.720 1439.850 998.470 ;
      LAYER met2 ;
        RECT 1440.130 996.000 1440.410 999.870 ;
      LAYER met2 ;
        RECT 1440.690 995.720 1442.150 998.470 ;
      LAYER met2 ;
        RECT 1442.430 996.000 1442.710 999.870 ;
      LAYER met2 ;
        RECT 1442.990 995.720 1444.450 998.470 ;
      LAYER met2 ;
        RECT 1444.730 996.000 1445.010 999.870 ;
      LAYER met2 ;
        RECT 1445.290 995.720 1446.750 998.470 ;
      LAYER met2 ;
        RECT 1447.030 996.000 1447.310 1000.000 ;
        RECT 1448.870 999.870 1450.680 1000.000 ;
        RECT 1451.170 999.870 1452.980 1000.000 ;
        RECT 1453.470 999.870 1454.820 1000.000 ;
      LAYER met2 ;
        RECT 1447.590 995.720 1448.590 998.470 ;
      LAYER met2 ;
        RECT 1448.870 996.000 1449.150 999.870 ;
      LAYER met2 ;
        RECT 1449.430 995.720 1450.890 998.470 ;
      LAYER met2 ;
        RECT 1451.170 996.000 1451.450 999.870 ;
      LAYER met2 ;
        RECT 1451.730 995.720 1453.190 998.470 ;
      LAYER met2 ;
        RECT 1453.470 996.000 1453.750 999.870 ;
      LAYER met2 ;
        RECT 1454.030 995.720 1455.030 998.470 ;
      LAYER met2 ;
        RECT 1455.310 996.000 1455.590 1000.000 ;
        RECT 1457.610 999.870 1459.420 1000.000 ;
        RECT 1459.910 999.870 1461.260 1000.000 ;
        RECT 1461.580 1000.010 1461.720 2914.150 ;
        RECT 1476.240 2829.150 1476.500 2829.470 ;
        RECT 1468.880 2546.270 1469.140 2546.590 ;
        RECT 1462.440 1019.330 1462.700 1019.650 ;
        RECT 1461.980 1018.990 1462.240 1019.310 ;
        RECT 1462.040 1007.750 1462.180 1018.990 ;
        RECT 1462.500 1008.090 1462.640 1019.330 ;
        RECT 1468.940 1012.510 1469.080 2546.270 ;
        RECT 1472.100 1024.770 1472.360 1025.090 ;
        RECT 1469.340 1020.690 1469.600 1021.010 ;
        RECT 1467.500 1012.190 1467.760 1012.510 ;
        RECT 1468.880 1012.190 1469.140 1012.510 ;
        RECT 1462.440 1007.770 1462.700 1008.090 ;
        RECT 1461.980 1007.430 1462.240 1007.750 ;
        RECT 1467.560 1000.010 1467.700 1012.190 ;
        RECT 1469.400 1000.010 1469.540 1020.690 ;
        RECT 1472.160 1000.010 1472.300 1024.770 ;
        RECT 1476.300 1000.010 1476.440 2829.150 ;
        RECT 1478.540 1016.950 1478.800 1017.270 ;
        RECT 1478.600 1000.010 1478.740 1016.950 ;
        RECT 1479.980 1011.490 1480.120 2915.510 ;
        RECT 1495.560 2915.170 1495.820 2915.490 ;
        RECT 1494.640 2913.810 1494.900 2914.130 ;
        RECT 1493.720 2912.790 1493.980 2913.110 ;
        RECT 1490.030 2850.035 1490.310 2850.405 ;
        RECT 1490.100 2849.870 1490.240 2850.035 ;
        RECT 1490.040 2849.550 1490.300 2849.870 ;
        RECT 1490.030 2830.315 1490.310 2830.685 ;
        RECT 1490.100 2829.470 1490.240 2830.315 ;
        RECT 1490.040 2829.150 1490.300 2829.470 ;
        RECT 1490.030 2801.755 1490.310 2802.125 ;
        RECT 1485.430 2784.075 1485.710 2784.445 ;
        RECT 1485.500 2781.190 1485.640 2784.075 ;
        RECT 1485.440 2780.870 1485.700 2781.190 ;
        RECT 1489.570 2767.755 1489.850 2768.125 ;
        RECT 1487.270 2739.195 1487.550 2739.565 ;
        RECT 1486.810 2720.155 1487.090 2720.525 ;
        RECT 1482.670 2656.915 1482.950 2657.285 ;
        RECT 1482.740 1012.510 1482.880 2656.915 ;
        RECT 1484.510 2548.795 1484.790 2549.165 ;
        RECT 1484.580 2546.590 1484.720 2548.795 ;
        RECT 1484.520 2546.270 1484.780 2546.590 ;
        RECT 1486.880 1460.970 1487.020 2720.155 ;
        RECT 1487.340 1461.310 1487.480 2739.195 ;
        RECT 1489.110 2691.595 1489.390 2691.965 ;
        RECT 1489.180 2691.430 1489.320 2691.595 ;
        RECT 1489.120 2691.110 1489.380 2691.430 ;
        RECT 1489.110 2673.915 1489.390 2674.285 ;
        RECT 1488.190 2629.035 1488.470 2629.405 ;
        RECT 1488.260 2607.530 1488.400 2629.035 ;
        RECT 1488.650 2609.995 1488.930 2610.365 ;
        RECT 1488.720 2608.470 1488.860 2609.995 ;
        RECT 1488.660 2608.150 1488.920 2608.470 ;
        RECT 1488.260 2607.390 1488.860 2607.530 ;
        RECT 1488.190 2595.035 1488.470 2595.405 ;
        RECT 1488.260 2594.870 1488.400 2595.035 ;
        RECT 1488.200 2594.550 1488.460 2594.870 ;
        RECT 1488.190 2580.755 1488.470 2581.125 ;
        RECT 1488.200 2580.610 1488.460 2580.755 ;
        RECT 1488.190 2567.155 1488.470 2567.525 ;
        RECT 1487.730 2518.875 1488.010 2519.245 ;
        RECT 1487.280 1460.990 1487.540 1461.310 ;
        RECT 1486.820 1460.650 1487.080 1460.970 ;
        RECT 1487.800 1013.530 1487.940 2518.875 ;
        RECT 1487.740 1013.210 1488.000 1013.530 ;
        RECT 1480.380 1012.190 1480.640 1012.510 ;
        RECT 1482.680 1012.190 1482.940 1012.510 ;
        RECT 1479.920 1011.170 1480.180 1011.490 ;
        RECT 1480.440 1000.010 1480.580 1012.190 ;
        RECT 1484.980 1011.170 1485.240 1011.490 ;
        RECT 1485.040 1000.010 1485.180 1011.170 ;
        RECT 1487.280 1009.470 1487.540 1009.790 ;
        RECT 1487.340 1000.010 1487.480 1009.470 ;
        RECT 1488.260 1008.090 1488.400 2567.155 ;
        RECT 1488.720 1013.870 1488.860 2607.390 ;
        RECT 1488.660 1013.550 1488.920 1013.870 ;
        RECT 1489.180 1008.770 1489.320 2673.915 ;
        RECT 1489.640 1055.690 1489.780 2767.755 ;
        RECT 1489.580 1055.370 1489.840 1055.690 ;
        RECT 1490.100 1016.590 1490.240 2801.755 ;
        RECT 1490.040 1016.270 1490.300 1016.590 ;
        RECT 1489.580 1012.530 1489.840 1012.850 ;
        RECT 1489.120 1008.450 1489.380 1008.770 ;
        RECT 1488.200 1007.770 1488.460 1008.090 ;
        RECT 1489.640 1000.010 1489.780 1012.530 ;
        RECT 1493.260 1009.810 1493.520 1010.130 ;
        RECT 1493.320 1000.010 1493.460 1009.810 ;
        RECT 1493.780 1009.790 1493.920 2912.790 ;
        RECT 1494.700 2494.230 1494.840 2913.810 ;
        RECT 1495.100 2912.110 1495.360 2912.430 ;
        RECT 1495.160 2494.570 1495.300 2912.110 ;
        RECT 1495.620 2495.250 1495.760 2915.170 ;
        RECT 1496.940 2912.450 1497.200 2912.770 ;
        RECT 1496.480 2898.170 1496.740 2898.490 ;
        RECT 1496.010 2753.475 1496.290 2753.845 ;
        RECT 1495.560 2494.930 1495.820 2495.250 ;
        RECT 1495.100 2494.250 1495.360 2494.570 ;
        RECT 1494.640 2493.910 1494.900 2494.230 ;
        RECT 1495.560 1458.950 1495.820 1459.270 ;
        RECT 1495.100 1019.670 1495.360 1019.990 ;
        RECT 1493.720 1009.470 1493.980 1009.790 ;
        RECT 1495.160 1000.010 1495.300 1019.670 ;
        RECT 1461.580 1000.000 1462.340 1000.010 ;
        RECT 1466.480 1000.000 1467.700 1000.010 ;
        RECT 1468.780 1000.000 1469.540 1000.010 ;
        RECT 1470.620 1000.000 1472.300 1000.010 ;
        RECT 1475.220 1000.000 1476.440 1000.010 ;
        RECT 1477.520 1000.000 1478.740 1000.010 ;
        RECT 1479.360 1000.000 1480.580 1000.010 ;
        RECT 1483.960 1000.000 1485.180 1000.010 ;
        RECT 1485.800 1000.000 1487.480 1000.010 ;
        RECT 1488.100 1000.000 1489.780 1000.010 ;
        RECT 1492.700 1000.000 1493.460 1000.010 ;
        RECT 1494.540 1000.000 1495.300 1000.010 ;
        RECT 1461.580 999.870 1462.490 1000.000 ;
      LAYER met2 ;
        RECT 1455.870 995.720 1457.330 998.470 ;
      LAYER met2 ;
        RECT 1457.610 996.000 1457.890 999.870 ;
      LAYER met2 ;
        RECT 1458.170 995.720 1459.630 998.470 ;
      LAYER met2 ;
        RECT 1459.910 996.000 1460.190 999.870 ;
      LAYER met2 ;
        RECT 1460.470 995.720 1461.930 998.470 ;
      LAYER met2 ;
        RECT 1462.210 996.000 1462.490 999.870 ;
      LAYER met2 ;
        RECT 1462.770 995.720 1463.770 998.470 ;
      LAYER met2 ;
        RECT 1464.050 996.000 1464.330 1000.000 ;
        RECT 1466.350 999.870 1467.700 1000.000 ;
        RECT 1468.650 999.870 1469.540 1000.000 ;
        RECT 1470.490 999.870 1472.300 1000.000 ;
      LAYER met2 ;
        RECT 1464.610 995.720 1466.070 998.470 ;
      LAYER met2 ;
        RECT 1466.350 996.000 1466.630 999.870 ;
      LAYER met2 ;
        RECT 1466.910 995.720 1468.370 998.470 ;
      LAYER met2 ;
        RECT 1468.650 996.000 1468.930 999.870 ;
      LAYER met2 ;
        RECT 1469.210 995.720 1470.210 998.470 ;
      LAYER met2 ;
        RECT 1470.490 996.000 1470.770 999.870 ;
      LAYER met2 ;
        RECT 1471.050 995.720 1472.510 998.470 ;
      LAYER met2 ;
        RECT 1472.790 996.000 1473.070 1000.000 ;
        RECT 1475.090 999.870 1476.440 1000.000 ;
        RECT 1477.390 999.870 1478.740 1000.000 ;
        RECT 1479.230 999.870 1480.580 1000.000 ;
      LAYER met2 ;
        RECT 1473.350 995.720 1474.810 998.470 ;
      LAYER met2 ;
        RECT 1475.090 996.000 1475.370 999.870 ;
      LAYER met2 ;
        RECT 1475.650 995.720 1477.110 998.470 ;
      LAYER met2 ;
        RECT 1477.390 996.000 1477.670 999.870 ;
      LAYER met2 ;
        RECT 1477.950 995.720 1478.950 998.470 ;
      LAYER met2 ;
        RECT 1479.230 996.000 1479.510 999.870 ;
      LAYER met2 ;
        RECT 1479.790 995.720 1481.250 998.470 ;
      LAYER met2 ;
        RECT 1481.530 996.000 1481.810 1000.000 ;
        RECT 1483.830 999.870 1485.180 1000.000 ;
        RECT 1485.670 999.870 1487.480 1000.000 ;
        RECT 1487.970 999.870 1489.780 1000.000 ;
      LAYER met2 ;
        RECT 1482.090 995.720 1483.550 998.470 ;
      LAYER met2 ;
        RECT 1483.830 996.000 1484.110 999.870 ;
      LAYER met2 ;
        RECT 1484.390 995.720 1485.390 998.470 ;
      LAYER met2 ;
        RECT 1485.670 996.000 1485.950 999.870 ;
      LAYER met2 ;
        RECT 1486.230 995.720 1487.690 998.470 ;
      LAYER met2 ;
        RECT 1487.970 996.000 1488.250 999.870 ;
      LAYER met2 ;
        RECT 1488.530 995.720 1489.990 998.470 ;
      LAYER met2 ;
        RECT 1490.270 996.000 1490.550 1000.000 ;
        RECT 1492.570 999.870 1493.460 1000.000 ;
        RECT 1494.410 999.870 1495.300 1000.000 ;
        RECT 1495.620 1000.010 1495.760 1458.950 ;
        RECT 1496.080 1008.430 1496.220 2753.475 ;
        RECT 1496.540 1009.450 1496.680 2898.170 ;
        RECT 1497.000 1013.190 1497.140 2912.450 ;
        RECT 1497.400 2896.470 1497.660 2896.790 ;
        RECT 1496.940 1012.870 1497.200 1013.190 ;
        RECT 1496.480 1009.130 1496.740 1009.450 ;
        RECT 1497.460 1009.110 1497.600 2896.470 ;
        RECT 1501.600 2491.510 1501.740 2917.210 ;
        RECT 1502.000 2913.470 1502.260 2913.790 ;
        RECT 1502.060 2494.910 1502.200 2913.470 ;
        RECT 1502.460 2911.770 1502.720 2912.090 ;
        RECT 1502.000 2494.590 1502.260 2494.910 ;
        RECT 1501.540 2491.190 1501.800 2491.510 ;
        RECT 1502.000 1012.190 1502.260 1012.510 ;
        RECT 1497.400 1008.790 1497.660 1009.110 ;
        RECT 1496.020 1008.110 1496.280 1008.430 ;
        RECT 1502.060 1000.010 1502.200 1012.190 ;
        RECT 1502.520 1009.790 1502.660 2911.770 ;
        RECT 1535.180 2900.055 1535.320 2917.550 ;
        RECT 1546.160 2917.210 1546.420 2917.530 ;
        RECT 1546.220 2900.055 1546.360 2917.210 ;
        RECT 1567.320 2916.870 1567.580 2917.190 ;
        RECT 1567.380 2900.055 1567.520 2916.870 ;
        RECT 1641.840 2915.510 1642.100 2915.830 ;
        RECT 1598.600 2914.830 1598.860 2915.150 ;
        RECT 1598.660 2900.055 1598.800 2914.830 ;
        RECT 1630.800 2914.490 1631.060 2914.810 ;
        RECT 1609.640 2912.110 1609.900 2912.430 ;
        RECT 1609.700 2900.055 1609.840 2912.110 ;
        RECT 1630.860 2900.055 1631.000 2914.490 ;
        RECT 1641.900 2900.055 1642.040 2915.510 ;
        RECT 1705.320 2915.170 1705.580 2915.490 ;
        RECT 1694.280 2914.150 1694.540 2914.470 ;
        RECT 1663.000 2912.450 1663.260 2912.770 ;
        RECT 1663.060 2900.055 1663.200 2912.450 ;
        RECT 1694.340 2900.055 1694.480 2914.150 ;
        RECT 1705.380 2900.055 1705.520 2915.170 ;
        RECT 1768.800 2913.810 1769.060 2914.130 ;
        RECT 1789.960 2913.810 1790.220 2914.130 ;
        RECT 1895.300 2913.810 1895.560 2914.130 ;
        RECT 1758.680 2900.890 1758.940 2901.210 ;
        RECT 1758.740 2900.055 1758.880 2900.890 ;
        RECT 1768.860 2900.055 1769.000 2913.810 ;
        RECT 1779.840 2911.770 1780.100 2912.090 ;
        RECT 1779.900 2900.055 1780.040 2911.770 ;
        RECT 1790.020 2900.055 1790.160 2913.810 ;
        RECT 1812.040 2913.470 1812.300 2913.790 ;
        RECT 1801.000 2912.790 1801.260 2913.110 ;
        RECT 1801.060 2900.055 1801.200 2912.790 ;
        RECT 1812.100 2900.055 1812.240 2913.470 ;
        RECT 1843.320 2913.130 1843.580 2913.450 ;
        RECT 1833.200 2912.790 1833.460 2913.110 ;
        RECT 1833.260 2900.055 1833.400 2912.790 ;
        RECT 1843.380 2900.055 1843.520 2913.130 ;
        RECT 1887.480 2912.790 1887.740 2913.110 ;
        RECT 1854.360 2912.450 1854.620 2912.770 ;
        RECT 1886.560 2912.450 1886.820 2912.770 ;
        RECT 1854.420 2900.055 1854.560 2912.450 ;
        RECT 1864.480 2911.770 1864.740 2912.090 ;
        RECT 1864.540 2900.055 1864.680 2911.770 ;
        RECT 1502.850 2896.530 1503.130 2900.055 ;
        RECT 1524.930 2898.570 1525.210 2900.055 ;
        RECT 1524.140 2898.490 1525.210 2898.570 ;
        RECT 1524.080 2898.430 1525.210 2898.490 ;
        RECT 1524.080 2898.170 1524.340 2898.430 ;
        RECT 1503.380 2896.530 1503.640 2896.790 ;
        RECT 1502.850 2896.470 1503.640 2896.530 ;
        RECT 1502.850 2896.390 1503.580 2896.470 ;
        RECT 1502.850 2896.055 1503.130 2896.390 ;
        RECT 1524.930 2896.055 1525.210 2898.430 ;
        RECT 1535.050 2896.055 1535.330 2900.055 ;
        RECT 1546.090 2896.055 1546.370 2900.055 ;
        RECT 1567.250 2896.055 1567.530 2900.055 ;
        RECT 1598.530 2896.055 1598.810 2900.055 ;
        RECT 1609.570 2896.055 1609.850 2900.055 ;
        RECT 1630.730 2896.055 1631.010 2900.055 ;
        RECT 1641.770 2896.055 1642.050 2900.055 ;
        RECT 1662.930 2896.055 1663.210 2900.055 ;
        RECT 1694.210 2896.055 1694.490 2900.055 ;
        RECT 1705.250 2896.055 1705.530 2900.055 ;
        RECT 1758.610 2896.055 1758.890 2900.055 ;
        RECT 1768.730 2896.055 1769.010 2900.055 ;
        RECT 1779.770 2896.055 1780.050 2900.055 ;
        RECT 1789.890 2896.055 1790.170 2900.055 ;
        RECT 1800.930 2896.055 1801.210 2900.055 ;
        RECT 1811.970 2896.055 1812.250 2900.055 ;
        RECT 1833.130 2896.055 1833.410 2900.055 ;
        RECT 1843.250 2896.055 1843.530 2900.055 ;
        RECT 1854.290 2896.055 1854.570 2900.055 ;
        RECT 1864.410 2896.055 1864.690 2900.055 ;
        RECT 1875.450 2896.530 1875.730 2900.055 ;
        RECT 1876.900 2896.530 1877.160 2896.790 ;
        RECT 1875.450 2896.470 1877.160 2896.530 ;
        RECT 1885.570 2896.530 1885.850 2900.055 ;
        RECT 1875.450 2896.390 1877.100 2896.470 ;
        RECT 1885.570 2896.390 1886.300 2896.530 ;
        RECT 1875.450 2896.055 1875.730 2896.390 ;
        RECT 1885.570 2896.055 1885.850 2896.390 ;
      LAYER met2 ;
        RECT 1503.410 2895.775 1513.610 2896.055 ;
        RECT 1514.450 2895.775 1524.650 2896.055 ;
        RECT 1525.490 2895.775 1534.770 2896.055 ;
        RECT 1535.610 2895.775 1545.810 2896.055 ;
        RECT 1546.650 2895.775 1555.930 2896.055 ;
        RECT 1556.770 2895.775 1566.970 2896.055 ;
        RECT 1567.810 2895.775 1577.090 2896.055 ;
        RECT 1577.930 2895.775 1588.130 2896.055 ;
        RECT 1588.970 2895.775 1598.250 2896.055 ;
        RECT 1599.090 2895.775 1609.290 2896.055 ;
        RECT 1610.130 2895.775 1620.330 2896.055 ;
        RECT 1621.170 2895.775 1630.450 2896.055 ;
        RECT 1631.290 2895.775 1641.490 2896.055 ;
        RECT 1642.330 2895.775 1651.610 2896.055 ;
        RECT 1652.450 2895.775 1662.650 2896.055 ;
        RECT 1663.490 2895.775 1672.770 2896.055 ;
        RECT 1673.610 2895.775 1683.810 2896.055 ;
        RECT 1684.650 2895.775 1693.930 2896.055 ;
        RECT 1694.770 2895.775 1704.970 2896.055 ;
        RECT 1705.810 2895.775 1716.010 2896.055 ;
        RECT 1716.850 2895.775 1726.130 2896.055 ;
        RECT 1726.970 2895.775 1737.170 2896.055 ;
        RECT 1738.010 2895.775 1747.290 2896.055 ;
        RECT 1748.130 2895.775 1758.330 2896.055 ;
        RECT 1759.170 2895.775 1768.450 2896.055 ;
        RECT 1769.290 2895.775 1779.490 2896.055 ;
        RECT 1780.330 2895.775 1789.610 2896.055 ;
        RECT 1790.450 2895.775 1800.650 2896.055 ;
        RECT 1801.490 2895.775 1811.690 2896.055 ;
        RECT 1812.530 2895.775 1821.810 2896.055 ;
        RECT 1822.650 2895.775 1832.850 2896.055 ;
        RECT 1833.690 2895.775 1842.970 2896.055 ;
        RECT 1843.810 2895.775 1854.010 2896.055 ;
        RECT 1854.850 2895.775 1864.130 2896.055 ;
        RECT 1864.970 2895.775 1875.170 2896.055 ;
        RECT 1876.010 2895.775 1885.290 2896.055 ;
        RECT 1502.860 2504.280 1885.840 2895.775 ;
        RECT 1503.410 2504.000 1512.690 2504.280 ;
        RECT 1513.530 2504.000 1523.730 2504.280 ;
        RECT 1524.570 2504.000 1533.850 2504.280 ;
        RECT 1534.690 2504.000 1544.890 2504.280 ;
        RECT 1545.730 2504.000 1555.010 2504.280 ;
        RECT 1555.850 2504.000 1566.050 2504.280 ;
        RECT 1566.890 2504.000 1576.170 2504.280 ;
        RECT 1577.010 2504.000 1587.210 2504.280 ;
        RECT 1588.050 2504.000 1598.250 2504.280 ;
        RECT 1599.090 2504.000 1608.370 2504.280 ;
        RECT 1609.210 2504.000 1619.410 2504.280 ;
        RECT 1620.250 2504.000 1629.530 2504.280 ;
        RECT 1630.370 2504.000 1640.570 2504.280 ;
        RECT 1641.410 2504.000 1650.690 2504.280 ;
        RECT 1651.530 2504.000 1661.730 2504.280 ;
        RECT 1662.570 2504.000 1671.850 2504.280 ;
        RECT 1672.690 2504.000 1682.890 2504.280 ;
        RECT 1683.730 2504.000 1693.930 2504.280 ;
        RECT 1694.770 2504.000 1704.050 2504.280 ;
        RECT 1704.890 2504.000 1715.090 2504.280 ;
        RECT 1715.930 2504.000 1725.210 2504.280 ;
        RECT 1726.050 2504.000 1736.250 2504.280 ;
        RECT 1737.090 2504.000 1746.370 2504.280 ;
        RECT 1747.210 2504.000 1757.410 2504.280 ;
        RECT 1758.250 2504.000 1767.530 2504.280 ;
        RECT 1768.370 2504.000 1778.570 2504.280 ;
        RECT 1779.410 2504.000 1789.610 2504.280 ;
        RECT 1790.450 2504.000 1799.730 2504.280 ;
        RECT 1800.570 2504.000 1810.770 2504.280 ;
        RECT 1811.610 2504.000 1820.890 2504.280 ;
        RECT 1821.730 2504.000 1831.930 2504.280 ;
        RECT 1832.770 2504.000 1842.050 2504.280 ;
        RECT 1842.890 2504.000 1853.090 2504.280 ;
        RECT 1853.930 2504.000 1863.210 2504.280 ;
        RECT 1864.050 2504.000 1874.250 2504.280 ;
        RECT 1875.090 2504.000 1885.290 2504.280 ;
      LAYER met2 ;
        RECT 1524.010 2500.770 1524.290 2504.000 ;
        RECT 1524.010 2500.630 1524.740 2500.770 ;
        RECT 1524.010 2500.000 1524.290 2500.630 ;
        RECT 1514.880 2494.250 1515.140 2494.570 ;
        RECT 1504.300 2491.190 1504.560 2491.510 ;
        RECT 1503.840 1020.010 1504.100 1020.330 ;
        RECT 1502.460 1009.470 1502.720 1009.790 ;
        RECT 1503.900 1000.010 1504.040 1020.010 ;
        RECT 1504.360 1010.470 1504.500 2491.190 ;
        RECT 1514.940 2463.485 1515.080 2494.250 ;
        RECT 1514.870 2463.115 1515.150 2463.485 ;
        RECT 1519.020 1460.990 1519.280 1461.310 ;
        RECT 1512.120 1016.610 1512.380 1016.930 ;
        RECT 1509.360 1013.210 1509.620 1013.530 ;
        RECT 1506.600 1011.510 1506.860 1011.830 ;
        RECT 1504.300 1010.150 1504.560 1010.470 ;
        RECT 1506.660 1000.010 1506.800 1011.510 ;
        RECT 1507.980 1010.150 1508.240 1010.470 ;
        RECT 1495.620 1000.000 1496.840 1000.010 ;
        RECT 1500.980 1000.000 1502.200 1000.010 ;
        RECT 1503.280 1000.000 1504.040 1000.010 ;
        RECT 1505.580 1000.000 1506.800 1000.010 ;
        RECT 1508.040 1000.010 1508.180 1010.150 ;
        RECT 1508.900 1009.810 1509.160 1010.130 ;
        RECT 1508.960 1009.450 1509.100 1009.810 ;
        RECT 1509.420 1009.450 1509.560 1013.210 ;
        RECT 1511.660 1012.870 1511.920 1013.190 ;
        RECT 1508.900 1009.130 1509.160 1009.450 ;
        RECT 1509.360 1009.130 1509.620 1009.450 ;
        RECT 1511.720 1007.750 1511.860 1012.870 ;
        RECT 1511.660 1007.430 1511.920 1007.750 ;
        RECT 1512.180 1000.010 1512.320 1016.610 ;
        RECT 1513.040 1013.890 1513.300 1014.210 ;
        RECT 1512.580 1013.210 1512.840 1013.530 ;
        RECT 1512.640 1010.470 1512.780 1013.210 ;
        RECT 1512.580 1010.150 1512.840 1010.470 ;
        RECT 1508.040 1000.000 1509.720 1000.010 ;
        RECT 1512.020 1000.000 1512.320 1000.010 ;
        RECT 1495.620 999.870 1496.990 1000.000 ;
      LAYER met2 ;
        RECT 1490.830 995.720 1492.290 998.470 ;
      LAYER met2 ;
        RECT 1492.570 996.000 1492.850 999.870 ;
      LAYER met2 ;
        RECT 1493.130 995.720 1494.130 998.470 ;
      LAYER met2 ;
        RECT 1494.410 996.000 1494.690 999.870 ;
      LAYER met2 ;
        RECT 1494.970 995.720 1496.430 998.470 ;
      LAYER met2 ;
        RECT 1496.710 996.000 1496.990 999.870 ;
      LAYER met2 ;
        RECT 1497.270 995.720 1498.730 998.470 ;
      LAYER met2 ;
        RECT 1499.010 996.000 1499.290 1000.000 ;
        RECT 1500.850 999.870 1502.200 1000.000 ;
        RECT 1503.150 999.870 1504.040 1000.000 ;
        RECT 1505.450 999.870 1506.800 1000.000 ;
      LAYER met2 ;
        RECT 1499.570 995.720 1500.570 998.470 ;
      LAYER met2 ;
        RECT 1500.850 996.000 1501.130 999.870 ;
      LAYER met2 ;
        RECT 1501.410 995.720 1502.870 998.470 ;
      LAYER met2 ;
        RECT 1503.150 996.000 1503.430 999.870 ;
      LAYER met2 ;
        RECT 1503.710 995.720 1505.170 998.470 ;
      LAYER met2 ;
        RECT 1505.450 996.000 1505.730 999.870 ;
      LAYER met2 ;
        RECT 1506.010 995.720 1507.010 998.470 ;
      LAYER met2 ;
        RECT 1507.290 996.000 1507.570 1000.000 ;
        RECT 1508.040 999.870 1509.870 1000.000 ;
      LAYER met2 ;
        RECT 1507.850 995.720 1509.310 998.470 ;
      LAYER met2 ;
        RECT 1509.590 996.000 1509.870 999.870 ;
        RECT 1511.890 999.870 1512.320 1000.000 ;
        RECT 1513.100 1000.010 1513.240 1013.890 ;
        RECT 1519.080 1012.850 1519.220 1460.990 ;
        RECT 1519.480 1055.370 1519.740 1055.690 ;
        RECT 1519.020 1012.530 1519.280 1012.850 ;
        RECT 1518.100 1007.770 1518.360 1008.090 ;
        RECT 1518.160 1000.010 1518.300 1007.770 ;
        RECT 1519.540 1000.010 1519.680 1055.370 ;
        RECT 1524.600 1013.190 1524.740 2500.630 ;
        RECT 1534.130 2500.000 1534.410 2504.000 ;
        RECT 1545.170 2500.000 1545.450 2504.000 ;
        RECT 1555.290 2500.090 1555.570 2504.000 ;
        RECT 1553.120 2500.000 1555.570 2500.090 ;
        RECT 1576.450 2500.000 1576.730 2504.000 ;
        RECT 1587.490 2500.000 1587.770 2504.000 ;
        RECT 1608.650 2500.000 1608.930 2504.000 ;
        RECT 1619.690 2500.000 1619.970 2504.000 ;
        RECT 1629.810 2500.090 1630.090 2504.000 ;
        RECT 1640.850 2500.090 1641.130 2504.000 ;
        RECT 1662.010 2500.090 1662.290 2504.000 ;
        RECT 1628.560 2500.000 1630.090 2500.090 ;
        RECT 1635.460 2500.000 1641.130 2500.090 ;
        RECT 1656.160 2500.000 1662.290 2500.090 ;
        RECT 1683.170 2500.000 1683.450 2504.000 ;
        RECT 1704.330 2500.000 1704.610 2504.000 ;
        RECT 1715.370 2500.000 1715.650 2504.000 ;
        RECT 1725.490 2500.000 1725.770 2504.000 ;
        RECT 1746.650 2500.000 1746.930 2504.000 ;
        RECT 1757.690 2500.000 1757.970 2504.000 ;
        RECT 1767.810 2500.090 1768.090 2504.000 ;
        RECT 1766.560 2500.000 1768.090 2500.090 ;
        RECT 1778.850 2500.000 1779.130 2504.000 ;
        RECT 1789.890 2500.000 1790.170 2504.000 ;
        RECT 1811.050 2500.000 1811.330 2504.000 ;
        RECT 1832.210 2500.000 1832.490 2504.000 ;
        RECT 1842.330 2500.000 1842.610 2504.000 ;
        RECT 1853.370 2500.090 1853.650 2504.000 ;
        RECT 1849.360 2500.000 1853.650 2500.090 ;
        RECT 1874.530 2500.000 1874.810 2504.000 ;
        RECT 1885.570 2500.000 1885.850 2504.000 ;
        RECT 1528.220 2485.750 1528.480 2486.070 ;
        RECT 1526.380 1460.650 1526.640 1460.970 ;
        RECT 1524.540 1012.870 1524.800 1013.190 ;
        RECT 1521.320 1012.530 1521.580 1012.850 ;
        RECT 1521.380 1000.010 1521.520 1012.530 ;
        RECT 1526.440 1000.010 1526.580 1460.650 ;
        RECT 1528.280 1013.870 1528.420 2485.750 ;
        RECT 1534.260 2485.390 1534.400 2500.000 ;
        RECT 1544.320 2494.250 1544.580 2494.570 ;
        RECT 1534.200 2485.070 1534.460 2485.390 ;
        RECT 1535.120 2484.390 1535.380 2484.710 ;
        RECT 1532.350 2463.115 1532.630 2463.485 ;
        RECT 1532.420 2429.290 1532.560 2463.115 ;
        RECT 1532.360 2428.970 1532.620 2429.290 ;
        RECT 1532.820 2428.290 1533.080 2428.610 ;
        RECT 1532.880 2381.090 1533.020 2428.290 ;
        RECT 1532.880 2380.950 1533.480 2381.090 ;
        RECT 1533.340 2367.070 1533.480 2380.950 ;
        RECT 1531.900 2366.810 1532.160 2367.070 ;
        RECT 1531.900 2366.750 1532.560 2366.810 ;
        RECT 1533.280 2366.750 1533.540 2367.070 ;
        RECT 1531.960 2366.670 1532.560 2366.750 ;
        RECT 1532.420 2359.930 1532.560 2366.670 ;
        RECT 1532.360 2359.610 1532.620 2359.930 ;
        RECT 1533.280 2359.610 1533.540 2359.930 ;
        RECT 1533.340 2318.790 1533.480 2359.610 ;
        RECT 1533.280 2318.470 1533.540 2318.790 ;
        RECT 1532.820 2318.130 1533.080 2318.450 ;
        RECT 1532.880 2311.730 1533.020 2318.130 ;
        RECT 1532.880 2311.590 1533.480 2311.730 ;
        RECT 1533.340 2270.365 1533.480 2311.590 ;
        RECT 1532.350 2269.995 1532.630 2270.365 ;
        RECT 1533.270 2269.995 1533.550 2270.365 ;
        RECT 1532.420 2263.030 1532.560 2269.995 ;
        RECT 1531.440 2262.710 1531.700 2263.030 ;
        RECT 1532.360 2262.710 1532.620 2263.030 ;
        RECT 1531.500 2215.090 1531.640 2262.710 ;
        RECT 1531.440 2214.770 1531.700 2215.090 ;
        RECT 1532.820 2214.770 1533.080 2215.090 ;
        RECT 1532.880 2187.890 1533.020 2214.770 ;
        RECT 1532.820 2187.570 1533.080 2187.890 ;
        RECT 1532.360 2186.890 1532.620 2187.210 ;
        RECT 1532.420 2173.270 1532.560 2186.890 ;
        RECT 1531.900 2172.950 1532.160 2173.270 ;
        RECT 1532.360 2172.950 1532.620 2173.270 ;
        RECT 1531.960 2166.470 1532.100 2172.950 ;
        RECT 1531.440 2166.150 1531.700 2166.470 ;
        RECT 1531.900 2166.150 1532.160 2166.470 ;
        RECT 1531.500 2124.990 1531.640 2166.150 ;
        RECT 1531.440 2124.670 1531.700 2124.990 ;
        RECT 1532.820 2124.670 1533.080 2124.990 ;
        RECT 1532.880 2111.390 1533.020 2124.670 ;
        RECT 1532.820 2111.070 1533.080 2111.390 ;
        RECT 1533.740 2111.070 1534.000 2111.390 ;
        RECT 1533.800 2063.450 1533.940 2111.070 ;
        RECT 1532.360 2063.130 1532.620 2063.450 ;
        RECT 1533.740 2063.130 1534.000 2063.450 ;
        RECT 1532.420 2062.965 1532.560 2063.130 ;
        RECT 1532.350 2062.595 1532.630 2062.965 ;
        RECT 1532.810 2027.915 1533.090 2028.285 ;
        RECT 1532.880 1980.830 1533.020 2027.915 ;
        RECT 1532.820 1980.510 1533.080 1980.830 ;
        RECT 1532.360 1979.830 1532.620 1980.150 ;
        RECT 1532.420 1932.210 1532.560 1979.830 ;
        RECT 1532.360 1931.890 1532.620 1932.210 ;
        RECT 1532.360 1931.210 1532.620 1931.530 ;
        RECT 1532.420 1883.930 1532.560 1931.210 ;
        RECT 1531.900 1883.610 1532.160 1883.930 ;
        RECT 1532.360 1883.610 1532.620 1883.930 ;
        RECT 1531.960 1835.650 1532.100 1883.610 ;
        RECT 1531.900 1835.330 1532.160 1835.650 ;
        RECT 1532.820 1835.330 1533.080 1835.650 ;
        RECT 1532.880 1786.690 1533.020 1835.330 ;
        RECT 1532.820 1786.370 1533.080 1786.690 ;
        RECT 1534.200 1786.370 1534.460 1786.690 ;
        RECT 1534.260 1739.430 1534.400 1786.370 ;
        RECT 1533.280 1739.170 1533.540 1739.430 ;
        RECT 1532.880 1739.110 1533.540 1739.170 ;
        RECT 1534.200 1739.110 1534.460 1739.430 ;
        RECT 1532.880 1739.030 1533.480 1739.110 ;
        RECT 1532.880 1738.750 1533.020 1739.030 ;
        RECT 1532.820 1738.430 1533.080 1738.750 ;
        RECT 1533.740 1738.430 1534.000 1738.750 ;
        RECT 1533.800 1690.810 1533.940 1738.430 ;
        RECT 1532.820 1690.490 1533.080 1690.810 ;
        RECT 1533.740 1690.490 1534.000 1690.810 ;
        RECT 1532.880 1690.325 1533.020 1690.490 ;
        RECT 1531.430 1689.955 1531.710 1690.325 ;
        RECT 1532.810 1689.955 1533.090 1690.325 ;
        RECT 1531.500 1683.670 1531.640 1689.955 ;
        RECT 1531.440 1683.350 1531.700 1683.670 ;
        RECT 1532.360 1683.350 1532.620 1683.670 ;
        RECT 1532.420 1641.930 1532.560 1683.350 ;
        RECT 1532.420 1641.790 1533.020 1641.930 ;
        RECT 1532.880 1635.390 1533.020 1641.790 ;
        RECT 1532.820 1635.070 1533.080 1635.390 ;
        RECT 1533.740 1635.070 1534.000 1635.390 ;
        RECT 1533.800 1587.110 1533.940 1635.070 ;
        RECT 1533.740 1586.790 1534.000 1587.110 ;
        RECT 1534.200 1586.790 1534.460 1587.110 ;
        RECT 1534.260 1545.970 1534.400 1586.790 ;
        RECT 1534.200 1545.650 1534.460 1545.970 ;
        RECT 1534.200 1544.970 1534.460 1545.290 ;
        RECT 1534.260 1497.690 1534.400 1544.970 ;
        RECT 1532.820 1497.370 1533.080 1497.690 ;
        RECT 1534.200 1497.370 1534.460 1497.690 ;
        RECT 1532.880 1497.205 1533.020 1497.370 ;
        RECT 1532.810 1496.835 1533.090 1497.205 ;
        RECT 1534.190 1496.835 1534.470 1497.205 ;
        RECT 1534.260 1449.605 1534.400 1496.835 ;
        RECT 1534.190 1449.235 1534.470 1449.605 ;
        RECT 1533.270 1448.555 1533.550 1448.925 ;
        RECT 1533.340 1393.730 1533.480 1448.555 ;
        RECT 1532.880 1393.590 1533.480 1393.730 ;
        RECT 1532.880 1387.045 1533.020 1393.590 ;
        RECT 1532.810 1386.675 1533.090 1387.045 ;
        RECT 1533.730 1386.675 1534.010 1387.045 ;
        RECT 1533.800 1338.910 1533.940 1386.675 ;
        RECT 1532.820 1338.590 1533.080 1338.910 ;
        RECT 1533.740 1338.590 1534.000 1338.910 ;
        RECT 1532.880 1249.005 1533.020 1338.590 ;
        RECT 1531.430 1248.635 1531.710 1249.005 ;
        RECT 1532.810 1248.635 1533.090 1249.005 ;
        RECT 1531.500 1206.730 1531.640 1248.635 ;
        RECT 1531.500 1206.590 1533.020 1206.730 ;
        RECT 1532.880 1111.110 1533.020 1206.590 ;
        RECT 1530.980 1110.790 1531.240 1111.110 ;
        RECT 1532.820 1110.790 1533.080 1111.110 ;
        RECT 1531.040 1076.090 1531.180 1110.790 ;
        RECT 1530.980 1075.770 1531.240 1076.090 ;
        RECT 1532.820 1075.770 1533.080 1076.090 ;
        RECT 1530.520 1020.350 1530.780 1020.670 ;
        RECT 1528.220 1013.550 1528.480 1013.870 ;
        RECT 1530.580 1000.010 1530.720 1020.350 ;
        RECT 1530.980 1013.550 1531.240 1013.870 ;
        RECT 1531.040 1009.450 1531.180 1013.550 ;
        RECT 1530.980 1009.130 1531.240 1009.450 ;
        RECT 1531.440 1009.130 1531.700 1009.450 ;
        RECT 1531.500 1000.010 1531.640 1009.130 ;
        RECT 1532.880 1001.290 1533.020 1075.770 ;
        RECT 1534.660 1009.810 1534.920 1010.130 ;
        RECT 1534.720 1008.770 1534.860 1009.810 ;
        RECT 1535.180 1009.450 1535.320 2484.390 ;
        RECT 1544.380 2415.010 1544.520 2494.250 ;
        RECT 1545.300 2484.370 1545.440 2500.000 ;
        RECT 1553.120 2499.950 1555.490 2500.000 ;
        RECT 1552.600 2494.930 1552.860 2495.250 ;
        RECT 1545.240 2484.050 1545.500 2484.370 ;
        RECT 1548.920 2484.050 1549.180 2484.370 ;
        RECT 1544.320 2414.690 1544.580 2415.010 ;
        RECT 1545.240 2414.690 1545.500 2415.010 ;
        RECT 1545.300 2380.670 1545.440 2414.690 ;
        RECT 1545.240 2380.350 1545.500 2380.670 ;
        RECT 1544.780 2380.010 1545.040 2380.330 ;
        RECT 1544.840 2366.810 1544.980 2380.010 ;
        RECT 1544.840 2366.670 1545.440 2366.810 ;
        RECT 1545.300 2332.390 1545.440 2366.670 ;
        RECT 1544.320 2332.070 1544.580 2332.390 ;
        RECT 1545.240 2332.070 1545.500 2332.390 ;
        RECT 1544.380 2318.450 1544.520 2332.070 ;
        RECT 1543.860 2318.130 1544.120 2318.450 ;
        RECT 1544.320 2318.130 1544.580 2318.450 ;
        RECT 1543.920 2283.770 1544.060 2318.130 ;
        RECT 1543.860 2283.450 1544.120 2283.770 ;
        RECT 1544.780 2283.450 1545.040 2283.770 ;
        RECT 1544.840 2270.250 1544.980 2283.450 ;
        RECT 1544.840 2270.110 1545.440 2270.250 ;
        RECT 1545.300 2269.830 1545.440 2270.110 ;
        RECT 1543.860 2269.510 1544.120 2269.830 ;
        RECT 1545.240 2269.510 1545.500 2269.830 ;
        RECT 1543.920 2245.090 1544.060 2269.510 ;
        RECT 1543.920 2244.950 1544.520 2245.090 ;
        RECT 1544.380 2004.630 1544.520 2244.950 ;
        RECT 1543.400 2004.310 1543.660 2004.630 ;
        RECT 1544.320 2004.310 1544.580 2004.630 ;
        RECT 1543.460 1980.490 1543.600 2004.310 ;
        RECT 1543.400 1980.170 1543.660 1980.490 ;
        RECT 1543.860 1980.170 1544.120 1980.490 ;
        RECT 1543.920 1956.350 1544.060 1980.170 ;
        RECT 1543.860 1956.030 1544.120 1956.350 ;
        RECT 1544.780 1956.030 1545.040 1956.350 ;
        RECT 1544.840 1932.290 1544.980 1956.030 ;
        RECT 1544.840 1932.150 1545.440 1932.290 ;
        RECT 1545.300 1931.870 1545.440 1932.150 ;
        RECT 1545.240 1931.550 1545.500 1931.870 ;
        RECT 1544.320 1931.210 1544.580 1931.530 ;
        RECT 1544.380 1897.530 1544.520 1931.210 ;
        RECT 1544.320 1897.210 1544.580 1897.530 ;
        RECT 1545.240 1897.210 1545.500 1897.530 ;
        RECT 1545.300 1859.790 1545.440 1897.210 ;
        RECT 1544.320 1859.470 1544.580 1859.790 ;
        RECT 1545.240 1859.470 1545.500 1859.790 ;
        RECT 1544.380 1822.050 1544.520 1859.470 ;
        RECT 1544.320 1821.730 1544.580 1822.050 ;
        RECT 1545.240 1821.730 1545.500 1822.050 ;
        RECT 1545.300 1773.170 1545.440 1821.730 ;
        RECT 1544.380 1773.030 1545.440 1773.170 ;
        RECT 1544.380 1725.490 1544.520 1773.030 ;
        RECT 1544.320 1725.170 1544.580 1725.490 ;
        RECT 1545.240 1725.170 1545.500 1725.490 ;
        RECT 1545.300 1642.530 1545.440 1725.170 ;
        RECT 1544.320 1642.210 1544.580 1642.530 ;
        RECT 1545.240 1642.210 1545.500 1642.530 ;
        RECT 1544.380 1641.930 1544.520 1642.210 ;
        RECT 1544.380 1641.790 1544.980 1641.930 ;
        RECT 1544.840 1593.910 1544.980 1641.790 ;
        RECT 1543.860 1593.590 1544.120 1593.910 ;
        RECT 1544.780 1593.590 1545.040 1593.910 ;
        RECT 1543.920 1587.110 1544.060 1593.590 ;
        RECT 1543.860 1586.790 1544.120 1587.110 ;
        RECT 1545.240 1586.790 1545.500 1587.110 ;
        RECT 1545.300 1449.410 1545.440 1586.790 ;
        RECT 1544.320 1449.090 1544.580 1449.410 ;
        RECT 1545.240 1449.090 1545.500 1449.410 ;
        RECT 1544.380 1435.470 1544.520 1449.090 ;
        RECT 1544.320 1435.150 1544.580 1435.470 ;
        RECT 1545.240 1435.150 1545.500 1435.470 ;
        RECT 1545.300 1414.130 1545.440 1435.150 ;
        RECT 1544.840 1413.990 1545.440 1414.130 ;
        RECT 1544.840 1400.790 1544.980 1413.990 ;
        RECT 1543.400 1400.470 1543.660 1400.790 ;
        RECT 1544.780 1400.470 1545.040 1400.790 ;
        RECT 1543.460 1352.850 1543.600 1400.470 ;
        RECT 1543.400 1352.530 1543.660 1352.850 ;
        RECT 1544.320 1352.530 1544.580 1352.850 ;
        RECT 1544.380 1345.565 1544.520 1352.530 ;
        RECT 1543.390 1345.195 1543.670 1345.565 ;
        RECT 1544.310 1345.195 1544.590 1345.565 ;
        RECT 1543.460 1297.430 1543.600 1345.195 ;
        RECT 1543.400 1297.110 1543.660 1297.430 ;
        RECT 1545.240 1297.110 1545.500 1297.430 ;
        RECT 1545.300 1270.230 1545.440 1297.110 ;
        RECT 1545.240 1269.910 1545.500 1270.230 ;
        RECT 1544.320 1269.230 1544.580 1269.550 ;
        RECT 1544.380 1221.270 1544.520 1269.230 ;
        RECT 1544.320 1220.950 1544.580 1221.270 ;
        RECT 1544.320 1220.270 1544.580 1220.590 ;
        RECT 1544.380 1159.390 1544.520 1220.270 ;
        RECT 1543.860 1159.070 1544.120 1159.390 ;
        RECT 1544.320 1159.070 1544.580 1159.390 ;
        RECT 1543.920 1124.450 1544.060 1159.070 ;
        RECT 1543.920 1124.310 1544.520 1124.450 ;
        RECT 1544.380 1076.850 1544.520 1124.310 ;
        RECT 1544.380 1076.710 1544.980 1076.850 ;
        RECT 1544.840 1028.570 1544.980 1076.710 ;
        RECT 1544.840 1028.430 1545.440 1028.570 ;
        RECT 1538.340 1013.890 1538.600 1014.210 ;
        RECT 1535.120 1009.130 1535.380 1009.450 ;
        RECT 1534.660 1008.450 1534.920 1008.770 ;
        RECT 1532.820 1000.970 1533.080 1001.290 ;
        RECT 1535.810 1000.970 1536.070 1001.290 ;
        RECT 1513.100 1000.000 1514.320 1000.010 ;
        RECT 1518.160 1000.000 1518.460 1000.010 ;
        RECT 1519.540 1000.000 1520.760 1000.010 ;
        RECT 1521.380 1000.000 1522.600 1000.010 ;
        RECT 1526.440 1000.000 1527.200 1000.010 ;
        RECT 1529.500 1000.000 1530.720 1000.010 ;
        RECT 1531.340 1000.000 1531.640 1000.010 ;
        RECT 1535.870 1000.000 1536.010 1000.970 ;
        RECT 1538.400 1000.010 1538.540 1013.890 ;
        RECT 1542.940 1012.870 1543.200 1013.190 ;
        RECT 1541.560 1012.530 1541.820 1012.850 ;
        RECT 1541.620 1000.010 1541.760 1012.530 ;
        RECT 1537.780 1000.000 1538.540 1000.010 ;
        RECT 1540.080 1000.000 1541.760 1000.010 ;
        RECT 1543.000 1000.010 1543.140 1012.870 ;
        RECT 1545.300 1012.850 1545.440 1028.430 ;
        RECT 1545.240 1012.530 1545.500 1012.850 ;
        RECT 1548.980 1009.110 1549.120 2484.050 ;
        RECT 1550.300 1013.890 1550.560 1014.210 ;
        RECT 1548.920 1008.790 1549.180 1009.110 ;
        RECT 1545.700 1007.430 1545.960 1007.750 ;
        RECT 1545.760 1000.010 1545.900 1007.430 ;
        RECT 1550.360 1000.010 1550.500 1013.890 ;
        RECT 1552.660 1008.770 1552.800 2494.930 ;
        RECT 1553.120 1735.350 1553.260 2499.950 ;
        RECT 1559.500 2494.590 1559.760 2494.910 ;
        RECT 1559.560 2319.325 1559.700 2494.590 ;
        RECT 1573.760 2493.910 1574.020 2494.230 ;
        RECT 1572.380 2485.070 1572.640 2485.390 ;
        RECT 1559.490 2318.955 1559.770 2319.325 ;
        RECT 1559.040 2318.130 1559.300 2318.450 ;
        RECT 1559.490 2318.275 1559.770 2318.645 ;
        RECT 1559.500 2318.130 1559.760 2318.275 ;
        RECT 1559.100 2270.510 1559.240 2318.130 ;
        RECT 1559.040 2270.190 1559.300 2270.510 ;
        RECT 1559.500 2270.190 1559.760 2270.510 ;
        RECT 1559.560 2263.030 1559.700 2270.190 ;
        RECT 1559.500 2262.710 1559.760 2263.030 ;
        RECT 1560.420 2262.710 1560.680 2263.030 ;
        RECT 1560.480 2215.090 1560.620 2262.710 ;
        RECT 1559.500 2214.770 1559.760 2215.090 ;
        RECT 1560.420 2214.770 1560.680 2215.090 ;
        RECT 1559.560 2166.470 1559.700 2214.770 ;
        RECT 1559.500 2166.150 1559.760 2166.470 ;
        RECT 1560.420 2166.150 1560.680 2166.470 ;
        RECT 1560.480 2118.530 1560.620 2166.150 ;
        RECT 1559.500 2118.210 1559.760 2118.530 ;
        RECT 1560.420 2118.210 1560.680 2118.530 ;
        RECT 1559.560 2069.910 1559.700 2118.210 ;
        RECT 1559.500 2069.590 1559.760 2069.910 ;
        RECT 1560.420 2069.590 1560.680 2069.910 ;
        RECT 1560.480 2021.970 1560.620 2069.590 ;
        RECT 1559.500 2021.650 1559.760 2021.970 ;
        RECT 1560.420 2021.650 1560.680 2021.970 ;
        RECT 1559.560 1973.350 1559.700 2021.650 ;
        RECT 1559.500 1973.030 1559.760 1973.350 ;
        RECT 1560.420 1973.030 1560.680 1973.350 ;
        RECT 1560.480 1925.410 1560.620 1973.030 ;
        RECT 1559.500 1925.090 1559.760 1925.410 ;
        RECT 1560.420 1925.090 1560.680 1925.410 ;
        RECT 1559.560 1876.790 1559.700 1925.090 ;
        RECT 1558.580 1876.470 1558.840 1876.790 ;
        RECT 1559.500 1876.470 1559.760 1876.790 ;
        RECT 1558.640 1828.850 1558.780 1876.470 ;
        RECT 1558.580 1828.530 1558.840 1828.850 ;
        RECT 1559.960 1828.530 1560.220 1828.850 ;
        RECT 1560.020 1787.450 1560.160 1828.530 ;
        RECT 1559.560 1787.310 1560.160 1787.450 ;
        RECT 1559.560 1780.230 1559.700 1787.310 ;
        RECT 1559.500 1779.910 1559.760 1780.230 ;
        RECT 1560.420 1779.910 1560.680 1780.230 ;
        RECT 1553.060 1735.030 1553.320 1735.350 ;
        RECT 1560.480 1732.290 1560.620 1779.910 ;
        RECT 1559.500 1731.970 1559.760 1732.290 ;
        RECT 1560.420 1731.970 1560.680 1732.290 ;
        RECT 1559.560 1714.690 1559.700 1731.970 ;
        RECT 1559.100 1714.550 1559.700 1714.690 ;
        RECT 1559.100 1701.010 1559.240 1714.550 ;
        RECT 1559.040 1700.690 1559.300 1701.010 ;
        RECT 1560.420 1700.690 1560.680 1701.010 ;
        RECT 1560.480 1656.210 1560.620 1700.690 ;
        RECT 1559.560 1656.070 1560.620 1656.210 ;
        RECT 1559.560 1593.910 1559.700 1656.070 ;
        RECT 1559.500 1593.590 1559.760 1593.910 ;
        RECT 1560.420 1593.590 1560.680 1593.910 ;
        RECT 1560.480 1545.970 1560.620 1593.590 ;
        RECT 1559.500 1545.650 1559.760 1545.970 ;
        RECT 1560.420 1545.650 1560.680 1545.970 ;
        RECT 1559.560 1497.350 1559.700 1545.650 ;
        RECT 1559.500 1497.030 1559.760 1497.350 ;
        RECT 1560.420 1497.030 1560.680 1497.350 ;
        RECT 1560.480 1449.410 1560.620 1497.030 ;
        RECT 1559.500 1449.090 1559.760 1449.410 ;
        RECT 1560.420 1449.090 1560.680 1449.410 ;
        RECT 1559.560 1400.790 1559.700 1449.090 ;
        RECT 1559.500 1400.470 1559.760 1400.790 ;
        RECT 1560.420 1400.470 1560.680 1400.790 ;
        RECT 1560.480 1352.850 1560.620 1400.470 ;
        RECT 1559.500 1352.530 1559.760 1352.850 ;
        RECT 1560.420 1352.530 1560.680 1352.850 ;
        RECT 1553.060 1013.210 1553.320 1013.530 ;
        RECT 1552.600 1008.450 1552.860 1008.770 ;
        RECT 1553.120 1000.010 1553.260 1013.210 ;
        RECT 1554.440 1008.450 1554.700 1008.770 ;
        RECT 1543.000 1000.000 1544.680 1000.010 ;
        RECT 1545.760 1000.000 1546.520 1000.010 ;
        RECT 1548.820 1000.000 1550.500 1000.010 ;
        RECT 1552.960 1000.000 1553.260 1000.010 ;
        RECT 1513.100 999.870 1514.470 1000.000 ;
      LAYER met2 ;
        RECT 1510.150 995.720 1511.610 998.470 ;
      LAYER met2 ;
        RECT 1511.890 996.000 1512.170 999.870 ;
      LAYER met2 ;
        RECT 1512.450 995.720 1513.910 998.470 ;
      LAYER met2 ;
        RECT 1514.190 996.000 1514.470 999.870 ;
      LAYER met2 ;
        RECT 1514.750 995.720 1515.750 998.470 ;
      LAYER met2 ;
        RECT 1516.030 996.000 1516.310 1000.000 ;
        RECT 1518.160 999.870 1518.610 1000.000 ;
        RECT 1519.540 999.870 1520.910 1000.000 ;
        RECT 1521.380 999.870 1522.750 1000.000 ;
      LAYER met2 ;
        RECT 1516.590 995.720 1518.050 998.470 ;
      LAYER met2 ;
        RECT 1518.330 996.000 1518.610 999.870 ;
      LAYER met2 ;
        RECT 1518.890 995.720 1520.350 998.470 ;
      LAYER met2 ;
        RECT 1520.630 996.000 1520.910 999.870 ;
      LAYER met2 ;
        RECT 1521.190 995.720 1522.190 998.470 ;
      LAYER met2 ;
        RECT 1522.470 996.000 1522.750 999.870 ;
      LAYER met2 ;
        RECT 1523.030 995.720 1524.490 998.470 ;
      LAYER met2 ;
        RECT 1524.770 996.000 1525.050 1000.000 ;
        RECT 1526.440 999.870 1527.350 1000.000 ;
      LAYER met2 ;
        RECT 1525.330 995.720 1526.790 998.470 ;
      LAYER met2 ;
        RECT 1527.070 996.000 1527.350 999.870 ;
        RECT 1529.370 999.870 1530.720 1000.000 ;
        RECT 1531.210 999.870 1531.640 1000.000 ;
      LAYER met2 ;
        RECT 1527.630 995.720 1529.090 998.470 ;
      LAYER met2 ;
        RECT 1529.370 996.000 1529.650 999.870 ;
      LAYER met2 ;
        RECT 1529.930 995.720 1530.930 998.470 ;
      LAYER met2 ;
        RECT 1531.210 996.000 1531.490 999.870 ;
      LAYER met2 ;
        RECT 1531.770 995.720 1533.230 998.470 ;
      LAYER met2 ;
        RECT 1533.510 996.000 1533.790 1000.000 ;
      LAYER met2 ;
        RECT 1534.070 995.720 1535.530 998.470 ;
      LAYER met2 ;
        RECT 1535.810 996.000 1536.090 1000.000 ;
        RECT 1537.650 999.870 1538.540 1000.000 ;
        RECT 1539.950 999.870 1541.760 1000.000 ;
      LAYER met2 ;
        RECT 1536.370 995.720 1537.370 998.470 ;
      LAYER met2 ;
        RECT 1537.650 996.000 1537.930 999.870 ;
      LAYER met2 ;
        RECT 1538.210 995.720 1539.670 998.470 ;
      LAYER met2 ;
        RECT 1539.950 996.000 1540.230 999.870 ;
      LAYER met2 ;
        RECT 1540.510 995.720 1541.970 998.470 ;
      LAYER met2 ;
        RECT 1542.250 996.000 1542.530 1000.000 ;
        RECT 1543.000 999.870 1544.830 1000.000 ;
        RECT 1545.760 999.870 1546.670 1000.000 ;
      LAYER met2 ;
        RECT 1542.810 995.720 1544.270 998.470 ;
      LAYER met2 ;
        RECT 1544.550 996.000 1544.830 999.870 ;
      LAYER met2 ;
        RECT 1545.110 995.720 1546.110 998.470 ;
      LAYER met2 ;
        RECT 1546.390 996.000 1546.670 999.870 ;
        RECT 1548.690 999.870 1550.500 1000.000 ;
      LAYER met2 ;
        RECT 1546.950 995.720 1548.410 998.470 ;
      LAYER met2 ;
        RECT 1548.690 996.000 1548.970 999.870 ;
      LAYER met2 ;
        RECT 1549.250 995.720 1550.710 998.470 ;
      LAYER met2 ;
        RECT 1550.990 996.000 1551.270 1000.000 ;
        RECT 1552.830 999.870 1553.260 1000.000 ;
        RECT 1554.500 1000.010 1554.640 1008.450 ;
        RECT 1555.820 1008.110 1556.080 1008.430 ;
        RECT 1555.880 1000.010 1556.020 1008.110 ;
        RECT 1559.560 1001.290 1559.700 1352.530 ;
        RECT 1571.920 1021.030 1572.180 1021.350 ;
        RECT 1565.480 1017.290 1565.740 1017.610 ;
        RECT 1559.500 1000.970 1559.760 1001.290 ;
        RECT 1561.570 1000.970 1561.830 1001.290 ;
        RECT 1554.500 1000.000 1555.260 1000.010 ;
        RECT 1555.880 1000.000 1557.560 1000.010 ;
        RECT 1561.630 1000.000 1561.770 1000.970 ;
        RECT 1565.540 1000.010 1565.680 1017.290 ;
        RECT 1566.400 1009.130 1566.660 1009.450 ;
        RECT 1566.460 1000.010 1566.600 1009.130 ;
        RECT 1571.980 1000.010 1572.120 1021.030 ;
        RECT 1564.000 1000.000 1565.680 1000.010 ;
        RECT 1566.300 1000.000 1566.600 1000.010 ;
        RECT 1570.440 1000.000 1572.120 1000.010 ;
        RECT 1554.500 999.870 1555.410 1000.000 ;
        RECT 1555.880 999.870 1557.710 1000.000 ;
      LAYER met2 ;
        RECT 1551.550 995.720 1552.550 998.470 ;
      LAYER met2 ;
        RECT 1552.830 996.000 1553.110 999.870 ;
      LAYER met2 ;
        RECT 1553.390 995.720 1554.850 998.470 ;
      LAYER met2 ;
        RECT 1555.130 996.000 1555.410 999.870 ;
      LAYER met2 ;
        RECT 1555.690 995.720 1557.150 998.470 ;
      LAYER met2 ;
        RECT 1557.430 996.000 1557.710 999.870 ;
      LAYER met2 ;
        RECT 1557.990 995.720 1559.450 998.470 ;
      LAYER met2 ;
        RECT 1559.730 996.000 1560.010 1000.000 ;
      LAYER met2 ;
        RECT 1560.290 995.720 1561.290 998.470 ;
      LAYER met2 ;
        RECT 1561.570 996.000 1561.850 1000.000 ;
        RECT 1563.870 999.870 1565.680 1000.000 ;
        RECT 1566.170 999.870 1566.600 1000.000 ;
      LAYER met2 ;
        RECT 1562.130 995.720 1563.590 998.470 ;
      LAYER met2 ;
        RECT 1563.870 996.000 1564.150 999.870 ;
      LAYER met2 ;
        RECT 1564.430 995.720 1565.890 998.470 ;
      LAYER met2 ;
        RECT 1566.170 996.000 1566.450 999.870 ;
      LAYER met2 ;
        RECT 1566.730 995.720 1567.730 998.470 ;
      LAYER met2 ;
        RECT 1568.010 996.000 1568.290 1000.000 ;
        RECT 1570.310 999.870 1572.120 1000.000 ;
        RECT 1572.440 1000.010 1572.580 2485.070 ;
        RECT 1573.820 2319.325 1573.960 2493.910 ;
        RECT 1576.580 2484.710 1576.720 2500.000 ;
        RECT 1586.640 2494.590 1586.900 2494.910 ;
        RECT 1576.520 2484.390 1576.780 2484.710 ;
        RECT 1573.750 2318.955 1574.030 2319.325 ;
        RECT 1573.750 2318.275 1574.030 2318.645 ;
        RECT 1573.820 1883.590 1573.960 2318.275 ;
        RECT 1573.760 1883.270 1574.020 1883.590 ;
        RECT 1574.680 1883.270 1574.940 1883.590 ;
        RECT 1574.740 1835.845 1574.880 1883.270 ;
        RECT 1573.750 1835.475 1574.030 1835.845 ;
        RECT 1574.670 1835.475 1574.950 1835.845 ;
        RECT 1573.820 1787.030 1573.960 1835.475 ;
        RECT 1573.760 1786.710 1574.020 1787.030 ;
        RECT 1574.680 1786.710 1574.940 1787.030 ;
        RECT 1574.740 1739.285 1574.880 1786.710 ;
        RECT 1573.750 1738.915 1574.030 1739.285 ;
        RECT 1574.670 1738.915 1574.950 1739.285 ;
        RECT 1573.820 1691.150 1573.960 1738.915 ;
        RECT 1573.760 1690.830 1574.020 1691.150 ;
        RECT 1574.220 1690.490 1574.480 1690.810 ;
        RECT 1574.280 1683.670 1574.420 1690.490 ;
        RECT 1572.840 1683.350 1573.100 1683.670 ;
        RECT 1574.220 1683.350 1574.480 1683.670 ;
        RECT 1572.900 1635.730 1573.040 1683.350 ;
        RECT 1572.840 1635.410 1573.100 1635.730 ;
        RECT 1573.760 1635.410 1574.020 1635.730 ;
        RECT 1573.820 1593.650 1573.960 1635.410 ;
        RECT 1573.820 1593.510 1574.420 1593.650 ;
        RECT 1574.280 1545.970 1574.420 1593.510 ;
        RECT 1573.760 1545.650 1574.020 1545.970 ;
        RECT 1574.220 1545.650 1574.480 1545.970 ;
        RECT 1573.820 1497.090 1573.960 1545.650 ;
        RECT 1573.820 1496.950 1574.420 1497.090 ;
        RECT 1574.280 1449.410 1574.420 1496.950 ;
        RECT 1573.760 1449.090 1574.020 1449.410 ;
        RECT 1574.220 1449.090 1574.480 1449.410 ;
        RECT 1573.820 1400.530 1573.960 1449.090 ;
        RECT 1573.820 1400.390 1574.420 1400.530 ;
        RECT 1574.280 1352.850 1574.420 1400.390 ;
        RECT 1573.760 1352.530 1574.020 1352.850 ;
        RECT 1574.220 1352.530 1574.480 1352.850 ;
        RECT 1573.820 1014.405 1573.960 1352.530 ;
        RECT 1573.750 1014.035 1574.030 1014.405 ;
        RECT 1575.590 1014.035 1575.870 1014.405 ;
        RECT 1573.300 1009.810 1573.560 1010.130 ;
        RECT 1573.360 1000.010 1573.500 1009.810 ;
        RECT 1575.660 1000.010 1575.800 1014.035 ;
        RECT 1586.700 1010.470 1586.840 2494.590 ;
        RECT 1587.620 2485.730 1587.760 2500.000 ;
        RECT 1600.440 2494.930 1600.700 2495.250 ;
        RECT 1593.540 2489.150 1593.800 2489.470 ;
        RECT 1587.560 2485.410 1587.820 2485.730 ;
        RECT 1593.600 1010.470 1593.740 2489.150 ;
        RECT 1600.500 1010.470 1600.640 2494.930 ;
        RECT 1608.780 2485.050 1608.920 2500.000 ;
        RECT 1608.720 2484.730 1608.980 2485.050 ;
        RECT 1619.820 2484.370 1619.960 2500.000 ;
        RECT 1628.560 2499.950 1630.010 2500.000 ;
        RECT 1635.460 2499.950 1641.050 2500.000 ;
        RECT 1656.160 2499.950 1662.210 2500.000 ;
        RECT 1621.140 2495.270 1621.400 2495.590 ;
        RECT 1611.020 2484.050 1611.280 2484.370 ;
        RECT 1619.760 2484.050 1620.020 2484.370 ;
        RECT 1611.080 1012.170 1611.220 2484.050 ;
        RECT 1614.240 1459.290 1614.500 1459.610 ;
        RECT 1611.020 1011.850 1611.280 1012.170 ;
        RECT 1582.500 1010.150 1582.760 1010.470 ;
        RECT 1586.640 1010.150 1586.900 1010.470 ;
        RECT 1591.240 1010.150 1591.500 1010.470 ;
        RECT 1593.540 1010.150 1593.800 1010.470 ;
        RECT 1599.060 1010.150 1599.320 1010.470 ;
        RECT 1600.440 1010.150 1600.700 1010.470 ;
        RECT 1582.560 1000.010 1582.700 1010.150 ;
        RECT 1582.960 1009.470 1583.220 1009.790 ;
        RECT 1572.440 1000.000 1572.740 1000.010 ;
        RECT 1573.360 1000.000 1575.040 1000.010 ;
        RECT 1575.660 1000.000 1576.880 1000.010 ;
        RECT 1581.480 1000.000 1582.700 1000.010 ;
        RECT 1572.440 999.870 1572.890 1000.000 ;
        RECT 1573.360 999.870 1575.190 1000.000 ;
        RECT 1575.660 999.870 1577.030 1000.000 ;
      LAYER met2 ;
        RECT 1568.570 995.720 1570.030 998.470 ;
      LAYER met2 ;
        RECT 1570.310 996.000 1570.590 999.870 ;
      LAYER met2 ;
        RECT 1570.870 995.720 1572.330 998.470 ;
      LAYER met2 ;
        RECT 1572.610 996.000 1572.890 999.870 ;
      LAYER met2 ;
        RECT 1573.170 995.720 1574.630 998.470 ;
      LAYER met2 ;
        RECT 1574.910 996.000 1575.190 999.870 ;
      LAYER met2 ;
        RECT 1575.470 995.720 1576.470 998.470 ;
      LAYER met2 ;
        RECT 1576.750 996.000 1577.030 999.870 ;
      LAYER met2 ;
        RECT 1577.310 995.720 1578.770 998.470 ;
      LAYER met2 ;
        RECT 1579.050 996.000 1579.330 1000.000 ;
        RECT 1581.350 999.870 1582.700 1000.000 ;
        RECT 1583.020 1000.010 1583.160 1009.470 ;
        RECT 1591.300 1000.010 1591.440 1010.150 ;
        RECT 1593.080 1009.810 1593.340 1010.130 ;
        RECT 1593.140 1000.010 1593.280 1009.810 ;
        RECT 1599.120 1000.010 1599.260 1010.150 ;
        RECT 1600.900 1009.470 1601.160 1009.790 ;
        RECT 1600.960 1000.010 1601.100 1009.470 ;
        RECT 1605.960 1008.790 1606.220 1009.110 ;
        RECT 1583.020 1000.000 1583.320 1000.010 ;
        RECT 1590.220 1000.000 1591.440 1000.010 ;
        RECT 1592.060 1000.000 1593.280 1000.010 ;
        RECT 1598.500 1000.000 1599.260 1000.010 ;
        RECT 1600.800 1000.000 1601.100 1000.010 ;
        RECT 1606.020 1000.010 1606.160 1008.790 ;
        RECT 1614.300 1007.750 1614.440 1459.290 ;
        RECT 1611.020 1007.430 1611.280 1007.750 ;
        RECT 1614.240 1007.430 1614.500 1007.750 ;
        RECT 1617.460 1007.430 1617.720 1007.750 ;
        RECT 1611.080 1000.010 1611.220 1007.430 ;
        RECT 1617.520 1000.010 1617.660 1007.430 ;
        RECT 1621.200 1000.690 1621.340 2495.270 ;
        RECT 1622.980 1016.270 1623.240 1016.590 ;
        RECT 1619.820 1000.550 1621.340 1000.690 ;
        RECT 1619.820 1000.010 1619.960 1000.550 ;
        RECT 1606.020 1000.000 1607.240 1000.010 ;
        RECT 1609.540 1000.000 1611.220 1000.010 ;
        RECT 1615.980 1000.000 1617.660 1000.010 ;
        RECT 1618.280 1000.000 1619.960 1000.010 ;
        RECT 1623.040 1000.010 1623.180 1016.270 ;
        RECT 1625.280 1012.870 1625.540 1013.190 ;
        RECT 1625.340 1000.010 1625.480 1012.870 ;
        RECT 1628.560 1012.850 1628.700 2499.950 ;
        RECT 1628.500 1012.530 1628.760 1012.850 ;
        RECT 1635.460 1007.750 1635.600 2499.950 ;
        RECT 1645.520 2488.810 1645.780 2489.130 ;
        RECT 1645.580 1010.130 1645.720 2488.810 ;
        RECT 1656.160 1016.930 1656.300 2499.950 ;
        RECT 1683.300 2489.810 1683.440 2500.000 ;
        RECT 1679.560 2489.490 1679.820 2489.810 ;
        RECT 1683.240 2489.490 1683.500 2489.810 ;
        RECT 1679.620 2484.370 1679.760 2489.490 ;
        RECT 1673.120 2484.050 1673.380 2484.370 ;
        RECT 1679.560 2484.050 1679.820 2484.370 ;
        RECT 1680.020 2484.050 1680.280 2484.370 ;
        RECT 1662.540 1814.590 1662.800 1814.910 ;
        RECT 1656.100 1016.610 1656.360 1016.930 ;
        RECT 1660.700 1010.150 1660.960 1010.470 ;
        RECT 1645.520 1009.810 1645.780 1010.130 ;
        RECT 1635.400 1007.430 1635.660 1007.750 ;
        RECT 1660.760 1000.010 1660.900 1010.150 ;
        RECT 1662.600 1000.010 1662.740 1814.590 ;
        RECT 1669.440 1735.030 1669.700 1735.350 ;
        RECT 1669.500 1012.170 1669.640 1735.030 ;
        RECT 1673.180 1013.530 1673.320 2484.050 ;
        RECT 1673.120 1013.210 1673.380 1013.530 ;
        RECT 1665.300 1011.850 1665.560 1012.170 ;
        RECT 1669.440 1011.850 1669.700 1012.170 ;
        RECT 1669.900 1011.850 1670.160 1012.170 ;
        RECT 1665.360 1000.010 1665.500 1011.850 ;
        RECT 1669.960 1010.470 1670.100 1011.850 ;
        RECT 1680.080 1010.810 1680.220 2484.050 ;
        RECT 1703.940 1735.710 1704.200 1736.030 ;
        RECT 1680.020 1010.490 1680.280 1010.810 ;
        RECT 1669.900 1010.150 1670.160 1010.470 ;
        RECT 1704.000 1000.010 1704.140 1735.710 ;
        RECT 1704.460 1021.010 1704.600 2500.000 ;
        RECT 1715.500 2484.370 1715.640 2500.000 ;
        RECT 1725.620 2486.410 1725.760 2500.000 ;
        RECT 1725.560 2486.090 1725.820 2486.410 ;
        RECT 1746.780 2485.390 1746.920 2500.000 ;
        RECT 1757.820 2486.750 1757.960 2500.000 ;
        RECT 1766.560 2499.950 1768.010 2500.000 ;
        RECT 1757.760 2486.430 1758.020 2486.750 ;
        RECT 1746.720 2485.070 1746.980 2485.390 ;
        RECT 1715.440 2484.050 1715.700 2484.370 ;
        RECT 1724.640 1928.490 1724.900 1928.810 ;
        RECT 1717.280 1925.770 1717.540 1926.090 ;
        RECT 1704.400 1020.690 1704.660 1021.010 ;
        RECT 1716.820 1020.690 1717.080 1021.010 ;
        RECT 1708.540 1013.210 1708.800 1013.530 ;
        RECT 1708.600 1000.010 1708.740 1013.210 ;
        RECT 1712.680 1009.810 1712.940 1010.130 ;
        RECT 1712.740 1000.010 1712.880 1009.810 ;
        RECT 1716.880 1000.010 1717.020 1020.690 ;
        RECT 1717.340 1010.130 1717.480 1925.770 ;
        RECT 1724.180 1012.870 1724.440 1013.190 ;
        RECT 1721.420 1012.530 1721.680 1012.850 ;
        RECT 1717.280 1009.810 1717.540 1010.130 ;
        RECT 1721.480 1000.010 1721.620 1012.530 ;
        RECT 1623.040 1000.000 1624.720 1000.010 ;
        RECT 1625.340 1000.000 1627.020 1000.010 ;
        RECT 1659.220 1000.000 1660.900 1000.010 ;
        RECT 1661.520 1000.000 1662.740 1000.010 ;
        RECT 1663.820 1000.000 1665.500 1000.010 ;
        RECT 1702.920 1000.000 1704.140 1000.010 ;
        RECT 1707.060 1000.000 1708.740 1000.010 ;
        RECT 1711.200 1000.000 1712.880 1000.010 ;
        RECT 1715.800 1000.000 1717.020 1000.010 ;
        RECT 1719.940 1000.000 1721.620 1000.010 ;
        RECT 1724.240 1000.010 1724.380 1012.870 ;
        RECT 1724.700 1012.850 1724.840 1928.490 ;
        RECT 1745.340 1927.470 1745.600 1927.790 ;
        RECT 1738.440 1926.110 1738.700 1926.430 ;
        RECT 1731.540 1849.270 1731.800 1849.590 ;
        RECT 1731.600 1062.830 1731.740 1849.270 ;
        RECT 1730.620 1062.510 1730.880 1062.830 ;
        RECT 1731.540 1062.510 1731.800 1062.830 ;
        RECT 1724.640 1012.530 1724.900 1012.850 ;
        RECT 1730.680 1000.690 1730.820 1062.510 ;
        RECT 1737.980 1010.490 1738.240 1010.810 ;
        RECT 1734.300 1009.810 1734.560 1010.130 ;
        RECT 1730.220 1000.550 1730.820 1000.690 ;
        RECT 1730.220 1000.010 1730.360 1000.550 ;
        RECT 1734.360 1000.010 1734.500 1009.810 ;
        RECT 1738.040 1000.010 1738.180 1010.490 ;
        RECT 1738.500 1010.130 1738.640 1926.110 ;
        RECT 1745.400 1012.850 1745.540 1927.470 ;
        RECT 1759.140 1926.450 1759.400 1926.770 ;
        RECT 1752.240 1883.610 1752.500 1883.930 ;
        RECT 1751.780 1736.730 1752.040 1737.050 ;
        RECT 1751.320 1013.045 1751.580 1013.190 ;
        RECT 1743.040 1012.530 1743.300 1012.850 ;
        RECT 1745.340 1012.530 1745.600 1012.850 ;
        RECT 1747.640 1012.530 1747.900 1012.850 ;
        RECT 1751.310 1012.675 1751.590 1013.045 ;
        RECT 1751.840 1012.850 1751.980 1736.730 ;
        RECT 1751.780 1012.530 1752.040 1012.850 ;
        RECT 1738.440 1009.810 1738.700 1010.130 ;
        RECT 1743.100 1000.010 1743.240 1012.530 ;
        RECT 1747.700 1000.010 1747.840 1012.530 ;
        RECT 1752.300 1000.690 1752.440 1883.610 ;
        RECT 1753.160 1013.045 1753.420 1013.190 ;
        RECT 1753.150 1012.675 1753.430 1013.045 ;
        RECT 1755.920 1010.150 1756.180 1010.470 ;
        RECT 1751.840 1000.550 1752.440 1000.690 ;
        RECT 1751.840 1000.010 1751.980 1000.550 ;
        RECT 1755.980 1000.010 1756.120 1010.150 ;
        RECT 1759.200 1000.010 1759.340 1926.450 ;
        RECT 1766.040 1766.310 1766.300 1766.630 ;
        RECT 1766.100 1076.170 1766.240 1766.310 ;
        RECT 1765.180 1076.030 1766.240 1076.170 ;
        RECT 1765.180 1028.570 1765.320 1076.030 ;
        RECT 1764.720 1028.430 1765.320 1028.570 ;
        RECT 1762.820 1013.890 1763.080 1014.210 ;
        RECT 1762.880 1013.530 1763.020 1013.890 ;
        RECT 1762.820 1013.210 1763.080 1013.530 ;
        RECT 1764.720 1000.010 1764.860 1028.430 ;
        RECT 1766.560 1017.270 1766.700 2499.950 ;
        RECT 1778.980 2489.470 1779.120 2500.000 ;
        RECT 1778.920 2489.150 1779.180 2489.470 ;
        RECT 1790.020 2489.130 1790.160 2500.000 ;
        RECT 1789.960 2488.810 1790.220 2489.130 ;
        RECT 1811.180 2486.070 1811.320 2500.000 ;
        RECT 1832.340 2487.090 1832.480 2500.000 ;
        RECT 1842.460 2488.790 1842.600 2500.000 ;
        RECT 1849.360 2499.950 1853.570 2500.000 ;
        RECT 1842.400 2488.470 1842.660 2488.790 ;
        RECT 1832.280 2486.770 1832.540 2487.090 ;
        RECT 1811.120 2485.750 1811.380 2486.070 ;
        RECT 1828.140 1927.810 1828.400 1928.130 ;
        RECT 1779.840 1927.130 1780.100 1927.450 ;
        RECT 1772.940 1925.430 1773.200 1925.750 ;
        RECT 1772.480 1736.390 1772.740 1736.710 ;
        RECT 1766.500 1016.950 1766.760 1017.270 ;
        RECT 1772.540 1008.770 1772.680 1736.390 ;
        RECT 1769.260 1008.450 1769.520 1008.770 ;
        RECT 1772.480 1008.450 1772.740 1008.770 ;
        RECT 1769.320 1000.010 1769.460 1008.450 ;
        RECT 1773.000 1000.010 1773.140 1925.430 ;
        RECT 1779.900 1014.210 1780.040 1927.130 ;
        RECT 1786.740 1926.790 1787.000 1927.110 ;
        RECT 1786.800 1703.130 1786.940 1926.790 ;
        RECT 1827.680 1925.090 1827.940 1925.410 ;
        RECT 1821.240 1870.010 1821.500 1870.330 ;
        RECT 1820.780 1738.430 1821.040 1738.750 ;
        RECT 1800.540 1738.090 1800.800 1738.410 ;
        RECT 1793.640 1737.410 1793.900 1737.730 ;
        RECT 1786.340 1702.990 1786.940 1703.130 ;
        RECT 1786.340 1701.090 1786.480 1702.990 ;
        RECT 1786.340 1700.950 1786.940 1701.090 ;
        RECT 1777.540 1013.890 1777.800 1014.210 ;
        RECT 1779.840 1013.890 1780.100 1014.210 ;
        RECT 1777.600 1000.010 1777.740 1013.890 ;
        RECT 1786.280 1009.810 1786.540 1010.130 ;
        RECT 1782.140 1008.450 1782.400 1008.770 ;
        RECT 1782.200 1000.010 1782.340 1008.450 ;
        RECT 1786.340 1000.010 1786.480 1009.810 ;
        RECT 1786.800 1008.770 1786.940 1700.950 ;
        RECT 1790.420 1014.230 1790.680 1014.550 ;
        RECT 1790.480 1013.530 1790.620 1014.230 ;
        RECT 1793.700 1013.530 1793.840 1737.410 ;
        RECT 1800.080 1735.370 1800.340 1735.690 ;
        RECT 1790.420 1013.210 1790.680 1013.530 ;
        RECT 1790.880 1013.210 1791.140 1013.530 ;
        RECT 1793.640 1013.210 1793.900 1013.530 ;
        RECT 1794.100 1013.210 1794.360 1013.530 ;
        RECT 1786.740 1008.450 1787.000 1008.770 ;
        RECT 1790.940 1000.010 1791.080 1013.210 ;
        RECT 1794.160 1010.810 1794.300 1013.210 ;
        RECT 1794.100 1010.490 1794.360 1010.810 ;
        RECT 1795.020 1010.490 1795.280 1010.810 ;
        RECT 1795.080 1000.010 1795.220 1010.490 ;
        RECT 1800.140 1000.690 1800.280 1735.370 ;
        RECT 1800.600 1010.810 1800.740 1738.090 ;
        RECT 1814.340 1737.750 1814.600 1738.070 ;
        RECT 1807.440 1737.070 1807.700 1737.390 ;
        RECT 1806.980 1736.050 1807.240 1736.370 ;
        RECT 1800.540 1010.490 1800.800 1010.810 ;
        RECT 1807.040 1007.750 1807.180 1736.050 ;
        RECT 1803.760 1007.430 1804.020 1007.750 ;
        RECT 1806.980 1007.430 1807.240 1007.750 ;
        RECT 1799.220 1000.550 1800.280 1000.690 ;
        RECT 1799.220 1000.010 1799.360 1000.550 ;
        RECT 1803.820 1000.010 1803.960 1007.430 ;
        RECT 1807.500 1000.010 1807.640 1737.070 ;
        RECT 1814.400 1000.690 1814.540 1737.750 ;
        RECT 1815.490 1000.970 1815.750 1001.290 ;
        RECT 1812.560 1000.550 1814.540 1000.690 ;
        RECT 1812.560 1000.010 1812.700 1000.550 ;
        RECT 1724.240 1000.000 1724.540 1000.010 ;
        RECT 1728.680 1000.000 1730.360 1000.010 ;
        RECT 1733.280 1000.000 1734.500 1000.010 ;
        RECT 1737.420 1000.000 1738.180 1000.010 ;
        RECT 1741.560 1000.000 1743.240 1000.010 ;
        RECT 1746.160 1000.000 1747.840 1000.010 ;
        RECT 1750.300 1000.000 1751.980 1000.010 ;
        RECT 1754.900 1000.000 1756.120 1000.010 ;
        RECT 1759.040 1000.000 1759.340 1000.010 ;
        RECT 1763.640 1000.000 1764.860 1000.010 ;
        RECT 1767.780 1000.000 1769.460 1000.010 ;
        RECT 1771.920 1000.000 1773.140 1000.010 ;
        RECT 1776.520 1000.000 1777.740 1000.010 ;
        RECT 1780.660 1000.000 1782.340 1000.010 ;
        RECT 1785.260 1000.000 1786.480 1000.010 ;
        RECT 1789.400 1000.000 1791.080 1000.010 ;
        RECT 1794.000 1000.000 1795.220 1000.010 ;
        RECT 1798.140 1000.000 1799.360 1000.010 ;
        RECT 1802.280 1000.000 1803.960 1000.010 ;
        RECT 1806.880 1000.000 1807.640 1000.010 ;
        RECT 1811.020 1000.000 1812.700 1000.010 ;
        RECT 1815.550 1000.000 1815.690 1000.970 ;
        RECT 1820.840 1000.010 1820.980 1738.430 ;
        RECT 1821.300 1001.290 1821.440 1870.010 ;
        RECT 1823.540 1010.490 1823.800 1010.810 ;
        RECT 1821.240 1000.970 1821.500 1001.290 ;
        RECT 1823.600 1000.010 1823.740 1010.490 ;
        RECT 1827.740 1000.010 1827.880 1925.090 ;
        RECT 1828.200 1010.810 1828.340 1927.810 ;
        RECT 1849.360 1018.630 1849.500 2499.950 ;
        RECT 1869.540 2493.910 1869.800 2494.230 ;
        RECT 1849.300 1018.310 1849.560 1018.630 ;
        RECT 1869.600 1010.810 1869.740 2493.910 ;
        RECT 1874.660 2488.110 1874.800 2500.000 ;
        RECT 1885.700 2488.450 1885.840 2500.000 ;
        RECT 1885.640 2488.130 1885.900 2488.450 ;
        RECT 1874.600 2487.790 1874.860 2488.110 ;
        RECT 1870.000 1014.570 1870.260 1014.890 ;
        RECT 1870.060 1014.210 1870.200 1014.570 ;
        RECT 1870.000 1013.890 1870.260 1014.210 ;
        RECT 1886.160 1013.870 1886.300 2896.390 ;
        RECT 1886.620 1014.890 1886.760 2912.450 ;
        RECT 1887.540 2494.910 1887.680 2912.790 ;
        RECT 1894.840 2911.770 1895.100 2912.090 ;
        RECT 1887.940 2896.470 1888.200 2896.790 ;
        RECT 1888.000 2495.250 1888.140 2896.470 ;
        RECT 1890.690 2848.335 1890.970 2848.705 ;
        RECT 1887.940 2494.930 1888.200 2495.250 ;
        RECT 1887.480 2494.590 1887.740 2494.910 ;
        RECT 1890.760 1017.610 1890.900 2848.335 ;
        RECT 1891.150 2832.015 1891.430 2832.385 ;
        RECT 1890.700 1017.290 1890.960 1017.610 ;
        RECT 1886.560 1014.570 1886.820 1014.890 ;
        RECT 1886.100 1013.550 1886.360 1013.870 ;
        RECT 1872.820 1012.170 1874.340 1012.250 ;
        RECT 1875.520 1012.190 1875.780 1012.510 ;
        RECT 1872.760 1012.110 1874.400 1012.170 ;
        RECT 1872.760 1011.850 1873.020 1012.110 ;
        RECT 1874.140 1011.850 1874.400 1012.110 ;
        RECT 1873.220 1011.510 1873.480 1011.830 ;
        RECT 1828.140 1010.490 1828.400 1010.810 ;
        RECT 1867.700 1010.490 1867.960 1010.810 ;
        RECT 1869.540 1010.490 1869.800 1010.810 ;
        RECT 1831.820 1009.470 1832.080 1009.790 ;
        RECT 1831.880 1000.010 1832.020 1009.470 ;
        RECT 1867.760 1000.010 1867.900 1010.490 ;
        RECT 1873.280 1009.450 1873.420 1011.510 ;
        RECT 1873.220 1009.130 1873.480 1009.450 ;
        RECT 1875.580 1000.010 1875.720 1012.190 ;
        RECT 1891.220 1011.150 1891.360 2832.015 ;
        RECT 1891.610 2817.055 1891.890 2817.425 ;
        RECT 1891.680 1025.090 1891.820 2817.055 ;
        RECT 1892.070 2797.675 1892.350 2798.045 ;
        RECT 1891.620 1024.770 1891.880 1025.090 ;
        RECT 1892.140 1024.750 1892.280 2797.675 ;
        RECT 1892.530 2782.715 1892.810 2783.085 ;
        RECT 1892.080 1024.430 1892.340 1024.750 ;
        RECT 1892.600 1011.830 1892.740 2782.715 ;
        RECT 1893.920 2780.870 1894.180 2781.190 ;
        RECT 1893.450 2753.475 1893.730 2753.845 ;
        RECT 1892.990 2718.795 1893.270 2719.165 ;
        RECT 1893.060 1018.970 1893.200 2718.795 ;
        RECT 1893.520 1459.610 1893.660 2753.475 ;
        RECT 1893.460 1459.290 1893.720 1459.610 ;
        RECT 1893.000 1018.650 1893.260 1018.970 ;
        RECT 1893.980 1012.510 1894.120 2780.870 ;
        RECT 1894.370 2735.115 1894.650 2735.485 ;
        RECT 1894.440 1459.270 1894.580 2735.115 ;
        RECT 1894.900 2494.570 1895.040 2911.770 ;
        RECT 1895.360 2495.590 1895.500 2913.810 ;
        RECT 2094.020 2781.210 2094.280 2781.530 ;
        RECT 2556.320 2781.210 2556.580 2781.530 ;
        RECT 1897.590 2767.075 1897.870 2767.445 ;
        RECT 1895.300 2495.270 1895.560 2495.590 ;
        RECT 1894.840 2494.250 1895.100 2494.570 ;
        RECT 1894.380 1458.950 1894.640 1459.270 ;
        RECT 1897.660 1020.330 1897.800 2767.075 ;
        RECT 1898.050 2687.515 1898.330 2687.885 ;
        RECT 1897.600 1020.010 1897.860 1020.330 ;
        RECT 1898.120 1019.310 1898.260 2687.515 ;
        RECT 1898.510 2672.555 1898.790 2672.925 ;
        RECT 1898.580 1019.650 1898.720 2672.555 ;
        RECT 1898.970 2656.915 1899.250 2657.285 ;
        RECT 1898.520 1019.330 1898.780 1019.650 ;
        RECT 1898.060 1018.990 1898.320 1019.310 ;
        RECT 1899.040 1018.290 1899.180 2656.915 ;
        RECT 1899.430 2624.955 1899.710 2625.325 ;
        RECT 1898.980 1017.970 1899.240 1018.290 ;
        RECT 1899.500 1017.950 1899.640 2624.955 ;
        RECT 1899.890 2608.635 1900.170 2609.005 ;
        RECT 1899.440 1017.630 1899.700 1017.950 ;
        RECT 1893.920 1012.190 1894.180 1012.510 ;
        RECT 1892.540 1011.510 1892.800 1011.830 ;
        RECT 1899.960 1011.490 1900.100 2608.635 ;
        RECT 1900.350 2577.355 1900.630 2577.725 ;
        RECT 1899.900 1011.170 1900.160 1011.490 ;
        RECT 1891.160 1010.830 1891.420 1011.150 ;
        RECT 1879.660 1010.490 1879.920 1010.810 ;
        RECT 1879.720 1000.010 1879.860 1010.490 ;
        RECT 1900.420 1009.450 1900.560 2577.355 ;
        RECT 1900.810 2562.395 1901.090 2562.765 ;
        RECT 1900.880 1021.350 1901.020 2562.395 ;
        RECT 1901.270 2547.435 1901.550 2547.805 ;
        RECT 1900.820 1021.030 1901.080 1021.350 ;
        RECT 1901.340 1019.990 1901.480 2547.435 ;
        RECT 1903.570 2514.795 1903.850 2515.165 ;
        RECT 1903.640 1020.670 1903.780 2514.795 ;
        RECT 2076.540 1946.510 2076.800 1946.830 ;
        RECT 2044.340 1928.490 2044.600 1928.810 ;
        RECT 1964.300 1927.810 1964.560 1928.130 ;
        RECT 1929.340 1927.470 1929.600 1927.790 ;
        RECT 1929.400 1917.095 1929.540 1927.470 ;
        RECT 1952.340 1925.090 1952.600 1925.410 ;
        RECT 1952.400 1917.095 1952.540 1925.090 ;
        RECT 1964.360 1917.095 1964.500 1927.810 ;
        RECT 1998.340 1927.130 1998.600 1927.450 ;
        RECT 1987.300 1926.110 1987.560 1926.430 ;
        RECT 1975.340 1925.770 1975.600 1926.090 ;
        RECT 1975.400 1917.095 1975.540 1925.770 ;
        RECT 1987.360 1917.095 1987.500 1926.110 ;
        RECT 1998.400 1917.095 1998.540 1927.130 ;
        RECT 2033.300 1926.790 2033.560 1927.110 ;
        RECT 2010.300 1926.450 2010.560 1926.770 ;
        RECT 2010.360 1917.095 2010.500 1926.450 ;
        RECT 2033.360 1917.095 2033.500 1926.790 ;
        RECT 2044.400 1917.095 2044.540 1928.490 ;
        RECT 2067.340 1925.430 2067.600 1925.750 ;
        RECT 2067.400 1917.095 2067.540 1925.430 ;
        RECT 1929.290 1913.095 1929.570 1917.095 ;
        RECT 1952.290 1913.095 1952.570 1917.095 ;
        RECT 1964.250 1913.095 1964.530 1917.095 ;
        RECT 1975.290 1913.095 1975.570 1917.095 ;
        RECT 1987.250 1913.095 1987.530 1917.095 ;
        RECT 1998.290 1913.095 1998.570 1917.095 ;
        RECT 2010.250 1913.095 2010.530 1917.095 ;
        RECT 2033.250 1913.095 2033.530 1917.095 ;
        RECT 2044.290 1913.095 2044.570 1917.095 ;
        RECT 2067.290 1913.095 2067.570 1917.095 ;
      LAYER met2 ;
        RECT 1922.860 1912.815 1929.010 1913.095 ;
        RECT 1929.850 1912.815 1940.970 1913.095 ;
        RECT 1941.810 1912.815 1952.010 1913.095 ;
        RECT 1952.850 1912.815 1963.970 1913.095 ;
        RECT 1964.810 1912.815 1975.010 1913.095 ;
        RECT 1975.850 1912.815 1986.970 1913.095 ;
        RECT 1987.810 1912.815 1998.010 1913.095 ;
        RECT 1998.850 1912.815 2009.970 1913.095 ;
        RECT 2010.810 1912.815 2021.010 1913.095 ;
        RECT 2021.850 1912.815 2032.970 1913.095 ;
        RECT 2033.810 1912.815 2044.010 1913.095 ;
        RECT 2044.850 1912.815 2055.970 1913.095 ;
        RECT 2056.810 1912.815 2067.010 1913.095 ;
        RECT 2067.850 1912.815 2072.160 1913.095 ;
      LAYER met2 ;
        RECT 1904.490 1885.795 1904.770 1886.165 ;
        RECT 1904.560 1883.930 1904.700 1885.795 ;
        RECT 1904.500 1883.610 1904.760 1883.930 ;
        RECT 1904.490 1870.155 1904.770 1870.525 ;
        RECT 1904.500 1870.010 1904.760 1870.155 ;
        RECT 1904.490 1851.795 1904.770 1852.165 ;
        RECT 1904.560 1849.590 1904.700 1851.795 ;
        RECT 1904.500 1849.270 1904.760 1849.590 ;
        RECT 1904.490 1817.795 1904.770 1818.165 ;
        RECT 1904.560 1814.910 1904.700 1817.795 ;
        RECT 1904.500 1814.590 1904.760 1814.910 ;
        RECT 1904.490 1767.475 1904.770 1767.845 ;
        RECT 1904.560 1766.630 1904.700 1767.475 ;
        RECT 1904.500 1766.310 1904.760 1766.630 ;
      LAYER met2 ;
        RECT 1922.860 1754.280 2072.160 1912.815 ;
        RECT 1923.410 1754.000 1933.610 1754.280 ;
        RECT 1934.450 1754.000 1944.650 1754.280 ;
        RECT 1945.490 1754.000 1956.610 1754.280 ;
        RECT 1957.450 1754.000 1967.650 1754.280 ;
        RECT 1968.490 1754.000 1979.610 1754.280 ;
        RECT 1980.450 1754.000 1990.650 1754.280 ;
        RECT 1991.490 1754.000 2002.610 1754.280 ;
        RECT 2003.450 1754.000 2013.650 1754.280 ;
        RECT 2014.490 1754.000 2025.610 1754.280 ;
        RECT 2026.450 1754.000 2036.650 1754.280 ;
        RECT 2037.490 1754.000 2048.610 1754.280 ;
        RECT 2049.450 1754.000 2059.650 1754.280 ;
        RECT 2060.490 1754.000 2071.610 1754.280 ;
      LAYER met2 ;
        RECT 1933.890 1750.000 1934.170 1754.000 ;
        RECT 1944.930 1750.000 1945.210 1754.000 ;
        RECT 1956.890 1750.000 1957.170 1754.000 ;
        RECT 1967.930 1750.000 1968.210 1754.000 ;
        RECT 1979.890 1750.000 1980.170 1754.000 ;
        RECT 1990.930 1750.000 1991.210 1754.000 ;
        RECT 2002.890 1750.000 2003.170 1754.000 ;
        RECT 2013.930 1750.000 2014.210 1754.000 ;
        RECT 2036.930 1750.000 2037.210 1754.000 ;
        RECT 2059.930 1750.000 2060.210 1754.000 ;
        RECT 2071.890 1750.000 2072.170 1754.000 ;
        RECT 1934.000 1738.750 1934.140 1750.000 ;
        RECT 1933.940 1738.430 1934.200 1738.750 ;
        RECT 1945.040 1736.030 1945.180 1750.000 ;
        RECT 1957.000 1738.410 1957.140 1750.000 ;
        RECT 1956.940 1738.090 1957.200 1738.410 ;
        RECT 1968.040 1737.730 1968.180 1750.000 ;
        RECT 1967.980 1737.410 1968.240 1737.730 ;
        RECT 1980.000 1737.050 1980.140 1750.000 ;
        RECT 1991.040 1738.070 1991.180 1750.000 ;
        RECT 1990.980 1737.750 1991.240 1738.070 ;
        RECT 1979.940 1736.730 1980.200 1737.050 ;
        RECT 2003.000 1736.710 2003.140 1750.000 ;
        RECT 2014.040 1737.390 2014.180 1750.000 ;
        RECT 2013.980 1737.070 2014.240 1737.390 ;
        RECT 2002.940 1736.390 2003.200 1736.710 ;
        RECT 2037.040 1736.370 2037.180 1750.000 ;
        RECT 2036.980 1736.050 2037.240 1736.370 ;
        RECT 1944.980 1735.710 1945.240 1736.030 ;
        RECT 2060.040 1735.350 2060.180 1750.000 ;
        RECT 2072.000 1735.690 2072.140 1750.000 ;
        RECT 2071.940 1735.370 2072.200 1735.690 ;
        RECT 2059.980 1735.030 2060.240 1735.350 ;
        RECT 2000.640 1687.770 2000.900 1688.090 ;
        RECT 1903.580 1020.350 1903.840 1020.670 ;
        RECT 1901.280 1019.670 1901.540 1019.990 ;
        RECT 2000.700 1013.870 2000.840 1687.770 ;
        RECT 2048.940 1687.430 2049.200 1687.750 ;
        RECT 2042.040 1687.090 2042.300 1687.410 ;
        RECT 1998.340 1013.550 1998.600 1013.870 ;
        RECT 2000.640 1013.550 2000.900 1013.870 ;
        RECT 1900.360 1009.130 1900.620 1009.450 ;
        RECT 1998.400 1000.010 1998.540 1013.550 ;
        RECT 2000.640 1012.190 2000.900 1012.510 ;
        RECT 2000.700 1000.010 2000.840 1012.190 ;
        RECT 2041.580 1010.830 2041.840 1011.150 ;
        RECT 2037.900 1009.130 2038.160 1009.450 ;
        RECT 2037.960 1000.010 2038.100 1009.130 ;
        RECT 2041.640 1000.010 2041.780 1010.830 ;
        RECT 2042.100 1009.450 2042.240 1687.090 ;
        RECT 2049.000 1012.170 2049.140 1687.430 ;
        RECT 2069.640 1686.750 2069.900 1687.070 ;
        RECT 2061.820 1013.890 2062.080 1014.210 ;
        RECT 2057.220 1013.550 2057.480 1013.870 ;
        RECT 2046.640 1011.850 2046.900 1012.170 ;
        RECT 2048.940 1011.850 2049.200 1012.170 ;
        RECT 2042.040 1009.130 2042.300 1009.450 ;
        RECT 2046.700 1000.010 2046.840 1011.850 ;
        RECT 2053.080 1011.170 2053.340 1011.490 ;
        RECT 2053.140 1000.010 2053.280 1011.170 ;
        RECT 2057.280 1000.010 2057.420 1013.550 ;
        RECT 2061.880 1000.010 2062.020 1013.890 ;
        RECT 2069.180 1011.510 2069.440 1011.830 ;
        RECT 2065.960 1009.130 2066.220 1009.450 ;
        RECT 2066.020 1000.010 2066.160 1009.130 ;
        RECT 2069.240 1000.010 2069.380 1011.510 ;
        RECT 2069.700 1009.450 2069.840 1686.750 ;
        RECT 2076.600 1076.170 2076.740 1946.510 ;
        RECT 2082.980 1946.170 2083.240 1946.490 ;
        RECT 2075.220 1076.030 2076.740 1076.170 ;
        RECT 2075.220 1028.570 2075.360 1076.030 ;
        RECT 2074.760 1028.430 2075.360 1028.570 ;
        RECT 2069.640 1009.130 2069.900 1009.450 ;
        RECT 2074.760 1000.010 2074.900 1028.430 ;
        RECT 2079.300 1009.130 2079.560 1009.450 ;
        RECT 2079.360 1000.010 2079.500 1009.130 ;
        RECT 2083.040 1000.010 2083.180 1946.170 ;
        RECT 2083.440 1945.830 2083.700 1946.150 ;
        RECT 2083.500 1009.450 2083.640 1945.830 ;
        RECT 2087.110 1884.435 2087.390 1884.805 ;
        RECT 2084.350 1850.435 2084.630 1850.805 ;
        RECT 2084.420 1021.010 2084.560 1850.435 ;
        RECT 2084.810 1835.475 2085.090 1835.845 ;
        RECT 2084.360 1020.690 2084.620 1021.010 ;
        RECT 2084.880 1010.130 2085.020 1835.475 ;
        RECT 2085.270 1816.435 2085.550 1816.805 ;
        RECT 2085.340 1012.850 2085.480 1816.435 ;
        RECT 2085.730 1800.795 2086.010 1801.165 ;
        RECT 2085.800 1013.190 2085.940 1800.795 ;
        RECT 2086.190 1782.435 2086.470 1782.805 ;
        RECT 2086.260 1013.530 2086.400 1782.435 ;
        RECT 2086.650 1766.795 2086.930 1767.165 ;
        RECT 2086.200 1013.210 2086.460 1013.530 ;
        RECT 2085.740 1012.870 2086.000 1013.190 ;
        RECT 2085.280 1012.530 2085.540 1012.850 ;
        RECT 2086.720 1010.470 2086.860 1766.795 ;
        RECT 2087.180 1012.170 2087.320 1884.435 ;
        RECT 2087.120 1011.850 2087.380 1012.170 ;
        RECT 2086.660 1010.150 2086.920 1010.470 ;
        RECT 2084.820 1009.810 2085.080 1010.130 ;
        RECT 2083.440 1009.130 2083.700 1009.450 ;
        RECT 2094.080 1009.110 2094.220 2781.210 ;
        RECT 2422.000 2780.870 2422.260 2781.190 ;
        RECT 2422.060 2773.820 2422.200 2780.870 ;
        RECT 2556.380 2773.820 2556.520 2781.210 ;
        RECT 2422.060 2773.380 2422.380 2773.820 ;
        RECT 2556.380 2773.380 2556.700 2773.820 ;
        RECT 2422.100 2769.820 2422.380 2773.380 ;
        RECT 2556.420 2769.820 2556.700 2773.380 ;
      LAYER met2 ;
        RECT 2400.030 2769.540 2421.820 2769.820 ;
        RECT 2422.660 2769.540 2556.140 2769.820 ;
        RECT 2400.030 2604.280 2556.690 2769.540 ;
        RECT 2400.580 2604.000 2534.060 2604.280 ;
        RECT 2534.900 2604.000 2556.690 2604.280 ;
      LAYER met2 ;
        RECT 2400.020 2600.730 2400.300 2604.000 ;
        RECT 2394.460 2600.590 2400.300 2600.730 ;
        RECT 2534.340 2600.660 2534.620 2604.000 ;
        RECT 2394.460 2494.230 2394.600 2600.590 ;
        RECT 2400.020 2600.000 2400.300 2600.590 ;
        RECT 2534.300 2600.000 2534.620 2600.660 ;
        RECT 2534.300 2587.730 2534.440 2600.000 ;
        RECT 2528.720 2587.410 2528.980 2587.730 ;
        RECT 2534.240 2587.410 2534.500 2587.730 ;
        RECT 2394.400 2493.910 2394.660 2494.230 ;
        RECT 2294.120 1946.850 2294.380 1947.170 ;
        RECT 2380.140 1946.850 2380.400 1947.170 ;
        RECT 2287.210 1876.955 2287.490 1877.325 ;
        RECT 2287.280 1014.210 2287.420 1876.955 ;
        RECT 2287.670 1789.915 2287.950 1790.285 ;
        RECT 2287.220 1013.890 2287.480 1014.210 ;
        RECT 2287.740 1013.870 2287.880 1789.915 ;
        RECT 2287.680 1013.550 2287.940 1013.870 ;
        RECT 2294.180 1012.510 2294.320 1946.850 ;
        RECT 2321.260 1946.510 2321.520 1946.830 ;
        RECT 2321.320 1939.270 2321.460 1946.510 ;
        RECT 2380.200 1939.270 2380.340 1946.850 ;
        RECT 2438.100 1946.170 2438.360 1946.490 ;
        RECT 2438.160 1939.270 2438.300 1946.170 ;
        RECT 2496.980 1945.830 2497.240 1946.150 ;
        RECT 2497.040 1939.270 2497.180 1945.830 ;
        RECT 2321.250 1935.270 2321.530 1939.270 ;
        RECT 2380.130 1935.270 2380.410 1939.270 ;
        RECT 2438.090 1935.270 2438.370 1939.270 ;
        RECT 2496.970 1935.270 2497.250 1939.270 ;
      LAYER met2 ;
        RECT 2302.860 1934.990 2320.970 1935.270 ;
        RECT 2321.810 1934.990 2379.850 1935.270 ;
        RECT 2380.690 1934.990 2437.810 1935.270 ;
        RECT 2438.650 1934.990 2496.690 1935.270 ;
        RECT 2497.530 1934.990 2519.320 1935.270 ;
        RECT 2302.860 1704.280 2519.320 1934.990 ;
        RECT 2303.410 1704.000 2360.530 1704.280 ;
        RECT 2361.370 1704.000 2419.410 1704.280 ;
        RECT 2420.250 1704.000 2477.370 1704.280 ;
        RECT 2478.210 1704.000 2519.320 1704.280 ;
      LAYER met2 ;
        RECT 2302.850 1700.000 2303.130 1704.000 ;
        RECT 2360.810 1700.000 2361.090 1704.000 ;
        RECT 2419.690 1700.000 2419.970 1704.000 ;
        RECT 2477.650 1700.000 2477.930 1704.000 ;
        RECT 2302.920 1688.090 2303.060 1700.000 ;
        RECT 2302.860 1687.770 2303.120 1688.090 ;
        RECT 2360.880 1687.750 2361.020 1700.000 ;
        RECT 2360.820 1687.430 2361.080 1687.750 ;
        RECT 2419.760 1687.410 2419.900 1700.000 ;
        RECT 2419.700 1687.090 2419.960 1687.410 ;
        RECT 2477.720 1687.070 2477.860 1700.000 ;
        RECT 2477.660 1686.750 2477.920 1687.070 ;
        RECT 2294.120 1012.190 2294.380 1012.510 ;
        RECT 2528.780 1010.810 2528.920 2587.410 ;
        RECT 2539.290 1891.915 2539.570 1892.285 ;
        RECT 2539.360 1011.150 2539.500 1891.915 ;
        RECT 2539.750 1804.875 2540.030 1805.245 ;
        RECT 2539.820 1011.490 2539.960 1804.875 ;
        RECT 2540.210 1719.195 2540.490 1719.565 ;
        RECT 2540.280 1011.830 2540.420 1719.195 ;
        RECT 2540.220 1011.510 2540.480 1011.830 ;
        RECT 2539.760 1011.170 2540.020 1011.490 ;
        RECT 2539.300 1010.830 2539.560 1011.150 ;
        RECT 2528.720 1010.490 2528.980 1010.810 ;
        RECT 2094.020 1008.790 2094.280 1009.110 ;
        RECT 1819.760 1000.000 1820.980 1000.010 ;
        RECT 1822.060 1000.000 1823.740 1000.010 ;
        RECT 1826.200 1000.000 1827.880 1000.010 ;
        RECT 1830.800 1000.000 1832.020 1000.010 ;
        RECT 1867.600 1000.000 1867.900 1000.010 ;
        RECT 1874.040 1000.000 1875.720 1000.010 ;
        RECT 1878.180 1000.000 1879.860 1000.010 ;
        RECT 1997.780 1000.000 1998.540 1000.010 ;
        RECT 1999.620 1000.000 2000.840 1000.010 ;
        RECT 2036.420 1000.000 2038.100 1000.010 ;
        RECT 2041.020 1000.000 2041.780 1000.010 ;
        RECT 2045.160 1000.000 2046.840 1000.010 ;
        RECT 2051.600 1000.000 2053.280 1000.010 ;
        RECT 2056.200 1000.000 2057.420 1000.010 ;
        RECT 2060.340 1000.000 2062.020 1000.010 ;
        RECT 2064.940 1000.000 2066.160 1000.010 ;
        RECT 2069.080 1000.000 2069.380 1000.010 ;
        RECT 2073.220 1000.000 2074.900 1000.010 ;
        RECT 2077.820 1000.000 2079.500 1000.010 ;
        RECT 2081.960 1000.000 2083.180 1000.010 ;
        RECT 1583.020 999.870 1583.470 1000.000 ;
      LAYER met2 ;
        RECT 1579.610 995.720 1581.070 998.470 ;
      LAYER met2 ;
        RECT 1581.350 996.000 1581.630 999.870 ;
      LAYER met2 ;
        RECT 1581.910 995.720 1582.910 998.470 ;
      LAYER met2 ;
        RECT 1583.190 996.000 1583.470 999.870 ;
      LAYER met2 ;
        RECT 1583.750 995.720 1585.210 998.470 ;
      LAYER met2 ;
        RECT 1585.490 996.000 1585.770 1000.000 ;
      LAYER met2 ;
        RECT 1586.050 995.720 1587.510 998.470 ;
      LAYER met2 ;
        RECT 1587.790 996.000 1588.070 1000.000 ;
        RECT 1590.090 999.870 1591.440 1000.000 ;
        RECT 1591.930 999.870 1593.280 1000.000 ;
      LAYER met2 ;
        RECT 1588.350 995.720 1589.810 998.470 ;
      LAYER met2 ;
        RECT 1590.090 996.000 1590.370 999.870 ;
      LAYER met2 ;
        RECT 1590.650 995.720 1591.650 998.470 ;
      LAYER met2 ;
        RECT 1591.930 996.000 1592.210 999.870 ;
      LAYER met2 ;
        RECT 1592.490 995.720 1593.950 998.470 ;
      LAYER met2 ;
        RECT 1594.230 996.000 1594.510 1000.000 ;
      LAYER met2 ;
        RECT 1594.790 995.720 1596.250 998.470 ;
      LAYER met2 ;
        RECT 1596.530 996.000 1596.810 1000.000 ;
        RECT 1598.370 999.870 1599.260 1000.000 ;
        RECT 1600.670 999.870 1601.100 1000.000 ;
      LAYER met2 ;
        RECT 1597.090 995.720 1598.090 998.470 ;
      LAYER met2 ;
        RECT 1598.370 996.000 1598.650 999.870 ;
      LAYER met2 ;
        RECT 1598.930 995.720 1600.390 998.470 ;
      LAYER met2 ;
        RECT 1600.670 996.000 1600.950 999.870 ;
      LAYER met2 ;
        RECT 1601.230 995.720 1602.690 998.470 ;
      LAYER met2 ;
        RECT 1602.970 996.000 1603.250 1000.000 ;
      LAYER met2 ;
        RECT 1603.530 995.720 1604.990 998.470 ;
      LAYER met2 ;
        RECT 1605.270 996.000 1605.550 1000.000 ;
        RECT 1606.020 999.870 1607.390 1000.000 ;
      LAYER met2 ;
        RECT 1605.830 995.720 1606.830 998.470 ;
      LAYER met2 ;
        RECT 1607.110 996.000 1607.390 999.870 ;
        RECT 1609.410 999.870 1611.220 1000.000 ;
      LAYER met2 ;
        RECT 1607.670 995.720 1609.130 998.470 ;
      LAYER met2 ;
        RECT 1609.410 996.000 1609.690 999.870 ;
      LAYER met2 ;
        RECT 1609.970 995.720 1611.430 998.470 ;
      LAYER met2 ;
        RECT 1611.710 996.000 1611.990 1000.000 ;
      LAYER met2 ;
        RECT 1612.270 995.720 1613.270 998.470 ;
      LAYER met2 ;
        RECT 1613.550 996.000 1613.830 1000.000 ;
        RECT 1615.850 999.870 1617.660 1000.000 ;
        RECT 1618.150 999.870 1619.960 1000.000 ;
      LAYER met2 ;
        RECT 1614.110 995.720 1615.570 998.470 ;
      LAYER met2 ;
        RECT 1615.850 996.000 1616.130 999.870 ;
      LAYER met2 ;
        RECT 1616.410 995.720 1617.870 998.470 ;
      LAYER met2 ;
        RECT 1618.150 996.000 1618.430 999.870 ;
      LAYER met2 ;
        RECT 1618.710 995.720 1620.170 998.470 ;
      LAYER met2 ;
        RECT 1620.450 996.000 1620.730 1000.000 ;
      LAYER met2 ;
        RECT 1621.010 995.720 1622.010 998.470 ;
      LAYER met2 ;
        RECT 1622.290 996.000 1622.570 1000.000 ;
        RECT 1623.040 999.870 1624.870 1000.000 ;
        RECT 1625.340 999.870 1627.170 1000.000 ;
      LAYER met2 ;
        RECT 1622.850 995.720 1624.310 998.470 ;
      LAYER met2 ;
        RECT 1624.590 996.000 1624.870 999.870 ;
      LAYER met2 ;
        RECT 1625.150 995.720 1626.610 998.470 ;
      LAYER met2 ;
        RECT 1626.890 996.000 1627.170 999.870 ;
      LAYER met2 ;
        RECT 1627.450 995.720 1628.450 998.470 ;
      LAYER met2 ;
        RECT 1628.730 996.000 1629.010 1000.000 ;
      LAYER met2 ;
        RECT 1629.290 995.720 1630.750 998.470 ;
      LAYER met2 ;
        RECT 1631.030 996.000 1631.310 1000.000 ;
      LAYER met2 ;
        RECT 1631.590 995.720 1633.050 998.470 ;
      LAYER met2 ;
        RECT 1633.330 996.000 1633.610 1000.000 ;
      LAYER met2 ;
        RECT 1633.890 995.720 1635.350 998.470 ;
      LAYER met2 ;
        RECT 1635.630 996.000 1635.910 1000.000 ;
      LAYER met2 ;
        RECT 1636.190 995.720 1637.190 998.470 ;
      LAYER met2 ;
        RECT 1637.470 996.000 1637.750 1000.000 ;
      LAYER met2 ;
        RECT 1638.030 995.720 1639.490 998.470 ;
      LAYER met2 ;
        RECT 1639.770 996.000 1640.050 1000.000 ;
      LAYER met2 ;
        RECT 1640.330 995.720 1641.790 998.470 ;
      LAYER met2 ;
        RECT 1642.070 996.000 1642.350 1000.000 ;
      LAYER met2 ;
        RECT 1642.630 995.720 1643.630 998.470 ;
      LAYER met2 ;
        RECT 1643.910 996.000 1644.190 1000.000 ;
      LAYER met2 ;
        RECT 1644.470 995.720 1645.930 998.470 ;
      LAYER met2 ;
        RECT 1646.210 996.000 1646.490 1000.000 ;
      LAYER met2 ;
        RECT 1646.770 995.720 1648.230 998.470 ;
      LAYER met2 ;
        RECT 1648.510 996.000 1648.790 1000.000 ;
      LAYER met2 ;
        RECT 1649.070 995.720 1650.530 998.470 ;
      LAYER met2 ;
        RECT 1650.810 996.000 1651.090 1000.000 ;
      LAYER met2 ;
        RECT 1651.370 995.720 1652.370 998.470 ;
      LAYER met2 ;
        RECT 1652.650 996.000 1652.930 1000.000 ;
      LAYER met2 ;
        RECT 1653.210 995.720 1654.670 998.470 ;
      LAYER met2 ;
        RECT 1654.950 996.000 1655.230 1000.000 ;
      LAYER met2 ;
        RECT 1655.510 995.720 1656.970 998.470 ;
      LAYER met2 ;
        RECT 1657.250 996.000 1657.530 1000.000 ;
        RECT 1659.090 999.870 1660.900 1000.000 ;
        RECT 1661.390 999.870 1662.740 1000.000 ;
        RECT 1663.690 999.870 1665.500 1000.000 ;
      LAYER met2 ;
        RECT 1657.810 995.720 1658.810 998.470 ;
      LAYER met2 ;
        RECT 1659.090 996.000 1659.370 999.870 ;
      LAYER met2 ;
        RECT 1659.650 995.720 1661.110 998.470 ;
      LAYER met2 ;
        RECT 1661.390 996.000 1661.670 999.870 ;
      LAYER met2 ;
        RECT 1661.950 995.720 1663.410 998.470 ;
      LAYER met2 ;
        RECT 1663.690 996.000 1663.970 999.870 ;
      LAYER met2 ;
        RECT 1664.250 995.720 1665.710 998.470 ;
      LAYER met2 ;
        RECT 1665.990 996.000 1666.270 1000.000 ;
      LAYER met2 ;
        RECT 1666.550 995.720 1667.550 998.470 ;
      LAYER met2 ;
        RECT 1667.830 996.000 1668.110 1000.000 ;
      LAYER met2 ;
        RECT 1668.390 995.720 1669.850 998.470 ;
      LAYER met2 ;
        RECT 1670.130 996.000 1670.410 1000.000 ;
      LAYER met2 ;
        RECT 1670.690 995.720 1672.150 998.470 ;
      LAYER met2 ;
        RECT 1672.430 996.000 1672.710 1000.000 ;
      LAYER met2 ;
        RECT 1672.990 995.720 1673.990 998.470 ;
      LAYER met2 ;
        RECT 1674.270 996.000 1674.550 1000.000 ;
      LAYER met2 ;
        RECT 1674.830 995.720 1676.290 998.470 ;
      LAYER met2 ;
        RECT 1676.570 996.000 1676.850 1000.000 ;
      LAYER met2 ;
        RECT 1677.130 995.720 1678.590 998.470 ;
      LAYER met2 ;
        RECT 1678.870 996.000 1679.150 1000.000 ;
      LAYER met2 ;
        RECT 1679.430 995.720 1680.430 998.470 ;
      LAYER met2 ;
        RECT 1680.710 996.000 1680.990 1000.000 ;
      LAYER met2 ;
        RECT 1681.270 995.720 1682.730 998.470 ;
      LAYER met2 ;
        RECT 1683.010 996.000 1683.290 1000.000 ;
      LAYER met2 ;
        RECT 1683.570 995.720 1685.030 998.470 ;
      LAYER met2 ;
        RECT 1685.310 996.000 1685.590 1000.000 ;
      LAYER met2 ;
        RECT 1685.870 995.720 1687.330 998.470 ;
      LAYER met2 ;
        RECT 1687.610 996.000 1687.890 1000.000 ;
      LAYER met2 ;
        RECT 1688.170 995.720 1689.170 998.470 ;
      LAYER met2 ;
        RECT 1689.450 996.000 1689.730 1000.000 ;
      LAYER met2 ;
        RECT 1690.010 995.720 1691.470 998.470 ;
      LAYER met2 ;
        RECT 1691.750 996.000 1692.030 1000.000 ;
      LAYER met2 ;
        RECT 1692.310 995.720 1693.770 998.470 ;
      LAYER met2 ;
        RECT 1694.050 996.000 1694.330 1000.000 ;
      LAYER met2 ;
        RECT 1694.610 995.720 1695.610 998.470 ;
      LAYER met2 ;
        RECT 1695.890 996.000 1696.170 1000.000 ;
      LAYER met2 ;
        RECT 1696.450 995.720 1697.910 998.470 ;
      LAYER met2 ;
        RECT 1698.190 996.000 1698.470 1000.000 ;
      LAYER met2 ;
        RECT 1698.750 995.720 1700.210 998.470 ;
      LAYER met2 ;
        RECT 1700.490 996.000 1700.770 1000.000 ;
        RECT 1702.790 999.870 1704.140 1000.000 ;
      LAYER met2 ;
        RECT 1701.050 995.720 1702.510 998.470 ;
      LAYER met2 ;
        RECT 1702.790 996.000 1703.070 999.870 ;
      LAYER met2 ;
        RECT 1703.350 995.720 1704.350 998.470 ;
      LAYER met2 ;
        RECT 1704.630 996.000 1704.910 1000.000 ;
        RECT 1706.930 999.870 1708.740 1000.000 ;
      LAYER met2 ;
        RECT 1705.190 995.720 1706.650 998.470 ;
      LAYER met2 ;
        RECT 1706.930 996.000 1707.210 999.870 ;
      LAYER met2 ;
        RECT 1707.490 995.720 1708.950 998.470 ;
      LAYER met2 ;
        RECT 1709.230 996.000 1709.510 1000.000 ;
        RECT 1711.070 999.870 1712.880 1000.000 ;
      LAYER met2 ;
        RECT 1709.790 995.720 1710.790 998.470 ;
      LAYER met2 ;
        RECT 1711.070 996.000 1711.350 999.870 ;
      LAYER met2 ;
        RECT 1711.630 995.720 1713.090 998.470 ;
      LAYER met2 ;
        RECT 1713.370 996.000 1713.650 1000.000 ;
        RECT 1715.670 999.870 1717.020 1000.000 ;
      LAYER met2 ;
        RECT 1713.930 995.720 1715.390 998.470 ;
      LAYER met2 ;
        RECT 1715.670 996.000 1715.950 999.870 ;
      LAYER met2 ;
        RECT 1716.230 995.720 1717.690 998.470 ;
      LAYER met2 ;
        RECT 1717.970 996.000 1718.250 1000.000 ;
        RECT 1719.810 999.870 1721.620 1000.000 ;
      LAYER met2 ;
        RECT 1718.530 995.720 1719.530 998.470 ;
      LAYER met2 ;
        RECT 1719.810 996.000 1720.090 999.870 ;
      LAYER met2 ;
        RECT 1720.370 995.720 1721.830 998.470 ;
      LAYER met2 ;
        RECT 1722.110 996.000 1722.390 1000.000 ;
        RECT 1724.240 999.870 1724.690 1000.000 ;
      LAYER met2 ;
        RECT 1722.670 995.720 1724.130 998.470 ;
      LAYER met2 ;
        RECT 1724.410 996.000 1724.690 999.870 ;
      LAYER met2 ;
        RECT 1724.970 995.720 1725.970 998.470 ;
      LAYER met2 ;
        RECT 1726.250 996.000 1726.530 1000.000 ;
        RECT 1728.550 999.870 1730.360 1000.000 ;
      LAYER met2 ;
        RECT 1726.810 995.720 1728.270 998.470 ;
      LAYER met2 ;
        RECT 1728.550 996.000 1728.830 999.870 ;
      LAYER met2 ;
        RECT 1729.110 995.720 1730.570 998.470 ;
      LAYER met2 ;
        RECT 1730.850 996.000 1731.130 1000.000 ;
        RECT 1733.150 999.870 1734.500 1000.000 ;
      LAYER met2 ;
        RECT 1731.410 995.720 1732.870 998.470 ;
      LAYER met2 ;
        RECT 1733.150 996.000 1733.430 999.870 ;
      LAYER met2 ;
        RECT 1733.710 995.720 1734.710 998.470 ;
      LAYER met2 ;
        RECT 1734.990 996.000 1735.270 1000.000 ;
        RECT 1737.290 999.870 1738.180 1000.000 ;
      LAYER met2 ;
        RECT 1735.550 995.720 1737.010 998.470 ;
      LAYER met2 ;
        RECT 1737.290 996.000 1737.570 999.870 ;
      LAYER met2 ;
        RECT 1737.850 995.720 1739.310 998.470 ;
      LAYER met2 ;
        RECT 1739.590 996.000 1739.870 1000.000 ;
        RECT 1741.430 999.870 1743.240 1000.000 ;
      LAYER met2 ;
        RECT 1740.150 995.720 1741.150 998.470 ;
      LAYER met2 ;
        RECT 1741.430 996.000 1741.710 999.870 ;
      LAYER met2 ;
        RECT 1741.990 995.720 1743.450 998.470 ;
      LAYER met2 ;
        RECT 1743.730 996.000 1744.010 1000.000 ;
        RECT 1746.030 999.870 1747.840 1000.000 ;
      LAYER met2 ;
        RECT 1744.290 995.720 1745.750 998.470 ;
      LAYER met2 ;
        RECT 1746.030 996.000 1746.310 999.870 ;
      LAYER met2 ;
        RECT 1746.590 995.720 1748.050 998.470 ;
      LAYER met2 ;
        RECT 1748.330 996.000 1748.610 1000.000 ;
        RECT 1750.170 999.870 1751.980 1000.000 ;
      LAYER met2 ;
        RECT 1748.890 995.720 1749.890 998.470 ;
      LAYER met2 ;
        RECT 1750.170 996.000 1750.450 999.870 ;
      LAYER met2 ;
        RECT 1750.730 995.720 1752.190 998.470 ;
      LAYER met2 ;
        RECT 1752.470 996.000 1752.750 1000.000 ;
        RECT 1754.770 999.870 1756.120 1000.000 ;
      LAYER met2 ;
        RECT 1753.030 995.720 1754.490 998.470 ;
      LAYER met2 ;
        RECT 1754.770 996.000 1755.050 999.870 ;
      LAYER met2 ;
        RECT 1755.330 995.720 1756.330 998.470 ;
      LAYER met2 ;
        RECT 1756.610 996.000 1756.890 1000.000 ;
        RECT 1758.910 999.870 1759.340 1000.000 ;
      LAYER met2 ;
        RECT 1757.170 995.720 1758.630 998.470 ;
      LAYER met2 ;
        RECT 1758.910 996.000 1759.190 999.870 ;
      LAYER met2 ;
        RECT 1759.470 995.720 1760.930 998.470 ;
      LAYER met2 ;
        RECT 1761.210 996.000 1761.490 1000.000 ;
        RECT 1763.510 999.870 1764.860 1000.000 ;
      LAYER met2 ;
        RECT 1761.770 995.720 1763.230 998.470 ;
      LAYER met2 ;
        RECT 1763.510 996.000 1763.790 999.870 ;
      LAYER met2 ;
        RECT 1764.070 995.720 1765.070 998.470 ;
      LAYER met2 ;
        RECT 1765.350 996.000 1765.630 1000.000 ;
        RECT 1767.650 999.870 1769.460 1000.000 ;
      LAYER met2 ;
        RECT 1765.910 995.720 1767.370 998.470 ;
      LAYER met2 ;
        RECT 1767.650 996.000 1767.930 999.870 ;
      LAYER met2 ;
        RECT 1768.210 995.720 1769.670 998.470 ;
      LAYER met2 ;
        RECT 1769.950 996.000 1770.230 1000.000 ;
        RECT 1771.790 999.870 1773.140 1000.000 ;
      LAYER met2 ;
        RECT 1770.510 995.720 1771.510 998.470 ;
      LAYER met2 ;
        RECT 1771.790 996.000 1772.070 999.870 ;
      LAYER met2 ;
        RECT 1772.350 995.720 1773.810 998.470 ;
      LAYER met2 ;
        RECT 1774.090 996.000 1774.370 1000.000 ;
        RECT 1776.390 999.870 1777.740 1000.000 ;
      LAYER met2 ;
        RECT 1774.650 995.720 1776.110 998.470 ;
      LAYER met2 ;
        RECT 1776.390 996.000 1776.670 999.870 ;
      LAYER met2 ;
        RECT 1776.950 995.720 1778.410 998.470 ;
      LAYER met2 ;
        RECT 1778.690 996.000 1778.970 1000.000 ;
        RECT 1780.530 999.870 1782.340 1000.000 ;
      LAYER met2 ;
        RECT 1779.250 995.720 1780.250 998.470 ;
      LAYER met2 ;
        RECT 1780.530 996.000 1780.810 999.870 ;
      LAYER met2 ;
        RECT 1781.090 995.720 1782.550 998.470 ;
      LAYER met2 ;
        RECT 1782.830 996.000 1783.110 1000.000 ;
        RECT 1785.130 999.870 1786.480 1000.000 ;
      LAYER met2 ;
        RECT 1783.390 995.720 1784.850 998.470 ;
      LAYER met2 ;
        RECT 1785.130 996.000 1785.410 999.870 ;
      LAYER met2 ;
        RECT 1785.690 995.720 1786.690 998.470 ;
      LAYER met2 ;
        RECT 1786.970 996.000 1787.250 1000.000 ;
        RECT 1789.270 999.870 1791.080 1000.000 ;
      LAYER met2 ;
        RECT 1787.530 995.720 1788.990 998.470 ;
      LAYER met2 ;
        RECT 1789.270 996.000 1789.550 999.870 ;
      LAYER met2 ;
        RECT 1789.830 995.720 1791.290 998.470 ;
      LAYER met2 ;
        RECT 1791.570 996.000 1791.850 1000.000 ;
        RECT 1793.870 999.870 1795.220 1000.000 ;
      LAYER met2 ;
        RECT 1792.130 995.720 1793.590 998.470 ;
      LAYER met2 ;
        RECT 1793.870 996.000 1794.150 999.870 ;
      LAYER met2 ;
        RECT 1794.430 995.720 1795.430 998.470 ;
      LAYER met2 ;
        RECT 1795.710 996.000 1795.990 1000.000 ;
        RECT 1798.010 999.870 1799.360 1000.000 ;
      LAYER met2 ;
        RECT 1796.270 995.720 1797.730 998.470 ;
      LAYER met2 ;
        RECT 1798.010 996.000 1798.290 999.870 ;
      LAYER met2 ;
        RECT 1798.570 995.720 1800.030 998.470 ;
      LAYER met2 ;
        RECT 1800.310 996.000 1800.590 1000.000 ;
        RECT 1802.150 999.870 1803.960 1000.000 ;
      LAYER met2 ;
        RECT 1800.870 995.720 1801.870 998.470 ;
      LAYER met2 ;
        RECT 1802.150 996.000 1802.430 999.870 ;
      LAYER met2 ;
        RECT 1802.710 995.720 1804.170 998.470 ;
      LAYER met2 ;
        RECT 1804.450 996.000 1804.730 1000.000 ;
        RECT 1806.750 999.870 1807.640 1000.000 ;
      LAYER met2 ;
        RECT 1805.010 995.720 1806.470 998.470 ;
      LAYER met2 ;
        RECT 1806.750 996.000 1807.030 999.870 ;
      LAYER met2 ;
        RECT 1807.310 995.720 1808.770 998.470 ;
      LAYER met2 ;
        RECT 1809.050 996.000 1809.330 1000.000 ;
        RECT 1810.890 999.870 1812.700 1000.000 ;
      LAYER met2 ;
        RECT 1809.610 995.720 1810.610 998.470 ;
      LAYER met2 ;
        RECT 1810.890 996.000 1811.170 999.870 ;
      LAYER met2 ;
        RECT 1811.450 995.720 1812.910 998.470 ;
      LAYER met2 ;
        RECT 1813.190 996.000 1813.470 1000.000 ;
      LAYER met2 ;
        RECT 1813.750 995.720 1815.210 998.470 ;
      LAYER met2 ;
        RECT 1815.490 996.000 1815.770 1000.000 ;
      LAYER met2 ;
        RECT 1816.050 995.720 1817.050 998.470 ;
      LAYER met2 ;
        RECT 1817.330 996.000 1817.610 1000.000 ;
        RECT 1819.630 999.870 1820.980 1000.000 ;
        RECT 1821.930 999.870 1823.740 1000.000 ;
      LAYER met2 ;
        RECT 1817.890 995.720 1819.350 998.470 ;
      LAYER met2 ;
        RECT 1819.630 996.000 1819.910 999.870 ;
      LAYER met2 ;
        RECT 1820.190 995.720 1821.650 998.470 ;
      LAYER met2 ;
        RECT 1821.930 996.000 1822.210 999.870 ;
      LAYER met2 ;
        RECT 1822.490 995.720 1823.950 998.470 ;
      LAYER met2 ;
        RECT 1824.230 996.000 1824.510 1000.000 ;
        RECT 1826.070 999.870 1827.880 1000.000 ;
      LAYER met2 ;
        RECT 1824.790 995.720 1825.790 998.470 ;
      LAYER met2 ;
        RECT 1826.070 996.000 1826.350 999.870 ;
      LAYER met2 ;
        RECT 1826.630 995.720 1828.090 998.470 ;
      LAYER met2 ;
        RECT 1828.370 996.000 1828.650 1000.000 ;
        RECT 1830.670 999.870 1832.020 1000.000 ;
      LAYER met2 ;
        RECT 1828.930 995.720 1830.390 998.470 ;
      LAYER met2 ;
        RECT 1830.670 996.000 1830.950 999.870 ;
      LAYER met2 ;
        RECT 1831.230 995.720 1832.230 998.470 ;
      LAYER met2 ;
        RECT 1832.510 996.000 1832.790 1000.000 ;
      LAYER met2 ;
        RECT 1833.070 995.720 1834.530 998.470 ;
      LAYER met2 ;
        RECT 1834.810 996.000 1835.090 1000.000 ;
      LAYER met2 ;
        RECT 1835.370 995.720 1836.830 998.470 ;
      LAYER met2 ;
        RECT 1837.110 996.000 1837.390 1000.000 ;
      LAYER met2 ;
        RECT 1837.670 995.720 1838.670 998.470 ;
      LAYER met2 ;
        RECT 1838.950 996.000 1839.230 1000.000 ;
      LAYER met2 ;
        RECT 1839.510 995.720 1840.970 998.470 ;
      LAYER met2 ;
        RECT 1841.250 996.000 1841.530 1000.000 ;
      LAYER met2 ;
        RECT 1841.810 995.720 1843.270 998.470 ;
      LAYER met2 ;
        RECT 1843.550 996.000 1843.830 1000.000 ;
      LAYER met2 ;
        RECT 1844.110 995.720 1845.570 998.470 ;
      LAYER met2 ;
        RECT 1845.850 996.000 1846.130 1000.000 ;
      LAYER met2 ;
        RECT 1846.410 995.720 1847.410 998.470 ;
      LAYER met2 ;
        RECT 1847.690 996.000 1847.970 1000.000 ;
      LAYER met2 ;
        RECT 1848.250 995.720 1849.710 998.470 ;
      LAYER met2 ;
        RECT 1849.990 996.000 1850.270 1000.000 ;
      LAYER met2 ;
        RECT 1850.550 995.720 1852.010 998.470 ;
      LAYER met2 ;
        RECT 1852.290 996.000 1852.570 1000.000 ;
      LAYER met2 ;
        RECT 1852.850 995.720 1853.850 998.470 ;
      LAYER met2 ;
        RECT 1854.130 996.000 1854.410 1000.000 ;
      LAYER met2 ;
        RECT 1854.690 995.720 1856.150 998.470 ;
      LAYER met2 ;
        RECT 1856.430 996.000 1856.710 1000.000 ;
      LAYER met2 ;
        RECT 1856.990 995.720 1858.450 998.470 ;
      LAYER met2 ;
        RECT 1858.730 996.000 1859.010 1000.000 ;
      LAYER met2 ;
        RECT 1859.290 995.720 1860.750 998.470 ;
      LAYER met2 ;
        RECT 1861.030 996.000 1861.310 1000.000 ;
      LAYER met2 ;
        RECT 1861.590 995.720 1862.590 998.470 ;
      LAYER met2 ;
        RECT 1862.870 996.000 1863.150 1000.000 ;
      LAYER met2 ;
        RECT 1863.430 995.720 1864.890 998.470 ;
      LAYER met2 ;
        RECT 1865.170 996.000 1865.450 1000.000 ;
        RECT 1867.470 999.870 1867.900 1000.000 ;
      LAYER met2 ;
        RECT 1865.730 995.720 1867.190 998.470 ;
      LAYER met2 ;
        RECT 1867.470 996.000 1867.750 999.870 ;
      LAYER met2 ;
        RECT 1868.030 995.720 1869.030 998.470 ;
      LAYER met2 ;
        RECT 1869.310 996.000 1869.590 1000.000 ;
      LAYER met2 ;
        RECT 1869.870 995.720 1871.330 998.470 ;
      LAYER met2 ;
        RECT 1871.610 996.000 1871.890 1000.000 ;
        RECT 1873.910 999.870 1875.720 1000.000 ;
      LAYER met2 ;
        RECT 1872.170 995.720 1873.630 998.470 ;
      LAYER met2 ;
        RECT 1873.910 996.000 1874.190 999.870 ;
      LAYER met2 ;
        RECT 1874.470 995.720 1875.930 998.470 ;
      LAYER met2 ;
        RECT 1876.210 996.000 1876.490 1000.000 ;
        RECT 1878.050 999.870 1879.860 1000.000 ;
      LAYER met2 ;
        RECT 1876.770 995.720 1877.770 998.470 ;
      LAYER met2 ;
        RECT 1878.050 996.000 1878.330 999.870 ;
      LAYER met2 ;
        RECT 1878.610 995.720 1880.070 998.470 ;
      LAYER met2 ;
        RECT 1880.350 996.000 1880.630 1000.000 ;
      LAYER met2 ;
        RECT 1880.910 995.720 1882.370 998.470 ;
      LAYER met2 ;
        RECT 1882.650 996.000 1882.930 1000.000 ;
      LAYER met2 ;
        RECT 1883.210 995.720 1884.210 998.470 ;
      LAYER met2 ;
        RECT 1884.490 996.000 1884.770 1000.000 ;
      LAYER met2 ;
        RECT 1885.050 995.720 1886.510 998.470 ;
      LAYER met2 ;
        RECT 1886.790 996.000 1887.070 1000.000 ;
      LAYER met2 ;
        RECT 1887.350 995.720 1888.810 998.470 ;
      LAYER met2 ;
        RECT 1889.090 996.000 1889.370 1000.000 ;
      LAYER met2 ;
        RECT 1889.650 995.720 1891.110 998.470 ;
      LAYER met2 ;
        RECT 1891.390 996.000 1891.670 1000.000 ;
      LAYER met2 ;
        RECT 1891.950 995.720 1892.950 998.470 ;
      LAYER met2 ;
        RECT 1893.230 996.000 1893.510 1000.000 ;
      LAYER met2 ;
        RECT 1893.790 995.720 1895.250 998.470 ;
      LAYER met2 ;
        RECT 1895.530 996.000 1895.810 1000.000 ;
      LAYER met2 ;
        RECT 1896.090 995.720 1897.550 998.470 ;
      LAYER met2 ;
        RECT 1897.830 996.000 1898.110 1000.000 ;
      LAYER met2 ;
        RECT 1898.390 995.720 1899.390 998.470 ;
      LAYER met2 ;
        RECT 1899.670 996.000 1899.950 1000.000 ;
      LAYER met2 ;
        RECT 1900.230 995.720 1901.690 998.470 ;
      LAYER met2 ;
        RECT 1901.970 996.000 1902.250 1000.000 ;
      LAYER met2 ;
        RECT 1902.530 995.720 1903.990 998.470 ;
      LAYER met2 ;
        RECT 1904.270 996.000 1904.550 1000.000 ;
      LAYER met2 ;
        RECT 1904.830 995.720 1906.290 998.470 ;
      LAYER met2 ;
        RECT 1906.570 996.000 1906.850 1000.000 ;
      LAYER met2 ;
        RECT 1907.130 995.720 1908.130 998.470 ;
      LAYER met2 ;
        RECT 1908.410 996.000 1908.690 1000.000 ;
      LAYER met2 ;
        RECT 1908.970 995.720 1910.430 998.470 ;
      LAYER met2 ;
        RECT 1910.710 996.000 1910.990 1000.000 ;
      LAYER met2 ;
        RECT 1911.270 995.720 1912.730 998.470 ;
      LAYER met2 ;
        RECT 1913.010 996.000 1913.290 1000.000 ;
      LAYER met2 ;
        RECT 1913.570 995.720 1914.570 998.470 ;
      LAYER met2 ;
        RECT 1914.850 996.000 1915.130 1000.000 ;
      LAYER met2 ;
        RECT 1915.410 995.720 1916.870 998.470 ;
      LAYER met2 ;
        RECT 1917.150 996.000 1917.430 1000.000 ;
      LAYER met2 ;
        RECT 1917.710 995.720 1919.170 998.470 ;
      LAYER met2 ;
        RECT 1919.450 996.000 1919.730 1000.000 ;
      LAYER met2 ;
        RECT 1920.010 995.720 1921.470 998.470 ;
      LAYER met2 ;
        RECT 1921.750 996.000 1922.030 1000.000 ;
      LAYER met2 ;
        RECT 1922.310 995.720 1923.310 998.470 ;
      LAYER met2 ;
        RECT 1923.590 996.000 1923.870 1000.000 ;
      LAYER met2 ;
        RECT 1924.150 995.720 1925.610 998.470 ;
      LAYER met2 ;
        RECT 1925.890 996.000 1926.170 1000.000 ;
      LAYER met2 ;
        RECT 1926.450 995.720 1927.910 998.470 ;
      LAYER met2 ;
        RECT 1928.190 996.000 1928.470 1000.000 ;
      LAYER met2 ;
        RECT 1928.750 995.720 1929.750 998.470 ;
      LAYER met2 ;
        RECT 1930.030 996.000 1930.310 1000.000 ;
      LAYER met2 ;
        RECT 1930.590 995.720 1932.050 998.470 ;
      LAYER met2 ;
        RECT 1932.330 996.000 1932.610 1000.000 ;
      LAYER met2 ;
        RECT 1932.890 995.720 1934.350 998.470 ;
      LAYER met2 ;
        RECT 1934.630 996.000 1934.910 1000.000 ;
      LAYER met2 ;
        RECT 1935.190 995.720 1936.650 998.470 ;
      LAYER met2 ;
        RECT 1936.930 996.000 1937.210 1000.000 ;
      LAYER met2 ;
        RECT 1937.490 995.720 1938.490 998.470 ;
      LAYER met2 ;
        RECT 1938.770 996.000 1939.050 1000.000 ;
      LAYER met2 ;
        RECT 1939.330 995.720 1940.790 998.470 ;
      LAYER met2 ;
        RECT 1941.070 996.000 1941.350 1000.000 ;
      LAYER met2 ;
        RECT 1941.630 995.720 1943.090 998.470 ;
      LAYER met2 ;
        RECT 1943.370 996.000 1943.650 1000.000 ;
      LAYER met2 ;
        RECT 1943.930 995.720 1944.930 998.470 ;
      LAYER met2 ;
        RECT 1945.210 996.000 1945.490 1000.000 ;
      LAYER met2 ;
        RECT 1945.770 995.720 1947.230 998.470 ;
      LAYER met2 ;
        RECT 1947.510 996.000 1947.790 1000.000 ;
      LAYER met2 ;
        RECT 1948.070 995.720 1949.530 998.470 ;
      LAYER met2 ;
        RECT 1949.810 996.000 1950.090 1000.000 ;
      LAYER met2 ;
        RECT 1950.370 995.720 1951.830 998.470 ;
      LAYER met2 ;
        RECT 1952.110 996.000 1952.390 1000.000 ;
      LAYER met2 ;
        RECT 1952.670 995.720 1953.670 998.470 ;
      LAYER met2 ;
        RECT 1953.950 996.000 1954.230 1000.000 ;
      LAYER met2 ;
        RECT 1954.510 995.720 1955.970 998.470 ;
      LAYER met2 ;
        RECT 1956.250 996.000 1956.530 1000.000 ;
      LAYER met2 ;
        RECT 1956.810 995.720 1958.270 998.470 ;
      LAYER met2 ;
        RECT 1958.550 996.000 1958.830 1000.000 ;
      LAYER met2 ;
        RECT 1959.110 995.720 1960.110 998.470 ;
      LAYER met2 ;
        RECT 1960.390 996.000 1960.670 1000.000 ;
      LAYER met2 ;
        RECT 1960.950 995.720 1962.410 998.470 ;
      LAYER met2 ;
        RECT 1962.690 996.000 1962.970 1000.000 ;
      LAYER met2 ;
        RECT 1963.250 995.720 1964.710 998.470 ;
      LAYER met2 ;
        RECT 1964.990 996.000 1965.270 1000.000 ;
      LAYER met2 ;
        RECT 1965.550 995.720 1967.010 998.470 ;
      LAYER met2 ;
        RECT 1967.290 996.000 1967.570 1000.000 ;
      LAYER met2 ;
        RECT 1967.850 995.720 1968.850 998.470 ;
      LAYER met2 ;
        RECT 1969.130 996.000 1969.410 1000.000 ;
      LAYER met2 ;
        RECT 1969.690 995.720 1971.150 998.470 ;
      LAYER met2 ;
        RECT 1971.430 996.000 1971.710 1000.000 ;
      LAYER met2 ;
        RECT 1971.990 995.720 1973.450 998.470 ;
      LAYER met2 ;
        RECT 1973.730 996.000 1974.010 1000.000 ;
      LAYER met2 ;
        RECT 1974.290 995.720 1975.290 998.470 ;
      LAYER met2 ;
        RECT 1975.570 996.000 1975.850 1000.000 ;
      LAYER met2 ;
        RECT 1976.130 995.720 1977.590 998.470 ;
      LAYER met2 ;
        RECT 1977.870 996.000 1978.150 1000.000 ;
      LAYER met2 ;
        RECT 1978.430 995.720 1979.890 998.470 ;
      LAYER met2 ;
        RECT 1980.170 996.000 1980.450 1000.000 ;
      LAYER met2 ;
        RECT 1980.730 995.720 1982.190 998.470 ;
      LAYER met2 ;
        RECT 1982.470 996.000 1982.750 1000.000 ;
      LAYER met2 ;
        RECT 1983.030 995.720 1984.030 998.470 ;
      LAYER met2 ;
        RECT 1984.310 996.000 1984.590 1000.000 ;
      LAYER met2 ;
        RECT 1984.870 995.720 1986.330 998.470 ;
      LAYER met2 ;
        RECT 1986.610 996.000 1986.890 1000.000 ;
      LAYER met2 ;
        RECT 1987.170 995.720 1988.630 998.470 ;
      LAYER met2 ;
        RECT 1988.910 996.000 1989.190 1000.000 ;
      LAYER met2 ;
        RECT 1989.470 995.720 1990.470 998.470 ;
      LAYER met2 ;
        RECT 1990.750 996.000 1991.030 1000.000 ;
      LAYER met2 ;
        RECT 1991.310 995.720 1992.770 998.470 ;
      LAYER met2 ;
        RECT 1993.050 996.000 1993.330 1000.000 ;
      LAYER met2 ;
        RECT 1993.610 995.720 1995.070 998.470 ;
      LAYER met2 ;
        RECT 1995.350 996.000 1995.630 1000.000 ;
        RECT 1997.650 999.870 1998.540 1000.000 ;
        RECT 1999.490 999.870 2000.840 1000.000 ;
      LAYER met2 ;
        RECT 1995.910 995.720 1997.370 998.470 ;
      LAYER met2 ;
        RECT 1997.650 996.000 1997.930 999.870 ;
      LAYER met2 ;
        RECT 1998.210 995.720 1999.210 998.470 ;
      LAYER met2 ;
        RECT 1999.490 996.000 1999.770 999.870 ;
      LAYER met2 ;
        RECT 2000.050 995.720 2001.510 998.470 ;
      LAYER met2 ;
        RECT 2001.790 996.000 2002.070 1000.000 ;
      LAYER met2 ;
        RECT 2002.350 995.720 2003.810 998.470 ;
      LAYER met2 ;
        RECT 2004.090 996.000 2004.370 1000.000 ;
      LAYER met2 ;
        RECT 2004.650 995.720 2005.650 998.470 ;
      LAYER met2 ;
        RECT 2005.930 996.000 2006.210 1000.000 ;
      LAYER met2 ;
        RECT 2006.490 995.720 2007.950 998.470 ;
      LAYER met2 ;
        RECT 2008.230 996.000 2008.510 1000.000 ;
      LAYER met2 ;
        RECT 2008.790 995.720 2010.250 998.470 ;
      LAYER met2 ;
        RECT 2010.530 996.000 2010.810 1000.000 ;
      LAYER met2 ;
        RECT 2011.090 995.720 2012.090 998.470 ;
      LAYER met2 ;
        RECT 2012.370 996.000 2012.650 1000.000 ;
      LAYER met2 ;
        RECT 2012.930 995.720 2014.390 998.470 ;
      LAYER met2 ;
        RECT 2014.670 996.000 2014.950 1000.000 ;
      LAYER met2 ;
        RECT 2015.230 995.720 2016.690 998.470 ;
      LAYER met2 ;
        RECT 2016.970 996.000 2017.250 1000.000 ;
      LAYER met2 ;
        RECT 2017.530 995.720 2018.990 998.470 ;
      LAYER met2 ;
        RECT 2019.270 996.000 2019.550 1000.000 ;
      LAYER met2 ;
        RECT 2019.830 995.720 2020.830 998.470 ;
      LAYER met2 ;
        RECT 2021.110 996.000 2021.390 1000.000 ;
      LAYER met2 ;
        RECT 2021.670 995.720 2023.130 998.470 ;
      LAYER met2 ;
        RECT 2023.410 996.000 2023.690 1000.000 ;
      LAYER met2 ;
        RECT 2023.970 995.720 2025.430 998.470 ;
      LAYER met2 ;
        RECT 2025.710 996.000 2025.990 1000.000 ;
      LAYER met2 ;
        RECT 2026.270 995.720 2027.270 998.470 ;
      LAYER met2 ;
        RECT 2027.550 996.000 2027.830 1000.000 ;
      LAYER met2 ;
        RECT 2028.110 995.720 2029.570 998.470 ;
      LAYER met2 ;
        RECT 2029.850 996.000 2030.130 1000.000 ;
      LAYER met2 ;
        RECT 2030.410 995.720 2031.870 998.470 ;
      LAYER met2 ;
        RECT 2032.150 996.000 2032.430 1000.000 ;
      LAYER met2 ;
        RECT 2032.710 995.720 2034.170 998.470 ;
      LAYER met2 ;
        RECT 2034.450 996.000 2034.730 1000.000 ;
        RECT 2036.290 999.870 2038.100 1000.000 ;
      LAYER met2 ;
        RECT 2035.010 995.720 2036.010 998.470 ;
      LAYER met2 ;
        RECT 2036.290 996.000 2036.570 999.870 ;
      LAYER met2 ;
        RECT 2036.850 995.720 2038.310 998.470 ;
      LAYER met2 ;
        RECT 2038.590 996.000 2038.870 1000.000 ;
        RECT 2040.890 999.870 2041.780 1000.000 ;
      LAYER met2 ;
        RECT 2039.150 995.720 2040.610 998.470 ;
      LAYER met2 ;
        RECT 2040.890 996.000 2041.170 999.870 ;
      LAYER met2 ;
        RECT 2041.450 995.720 2042.450 998.470 ;
      LAYER met2 ;
        RECT 2042.730 996.000 2043.010 1000.000 ;
        RECT 2045.030 999.870 2046.840 1000.000 ;
      LAYER met2 ;
        RECT 2043.290 995.720 2044.750 998.470 ;
      LAYER met2 ;
        RECT 2045.030 996.000 2045.310 999.870 ;
      LAYER met2 ;
        RECT 2045.590 995.720 2047.050 998.470 ;
      LAYER met2 ;
        RECT 2047.330 996.000 2047.610 1000.000 ;
      LAYER met2 ;
        RECT 2047.890 995.720 2049.350 998.470 ;
      LAYER met2 ;
        RECT 2049.630 996.000 2049.910 1000.000 ;
        RECT 2051.470 999.870 2053.280 1000.000 ;
      LAYER met2 ;
        RECT 2050.190 995.720 2051.190 998.470 ;
      LAYER met2 ;
        RECT 2051.470 996.000 2051.750 999.870 ;
      LAYER met2 ;
        RECT 2052.030 995.720 2053.490 998.470 ;
      LAYER met2 ;
        RECT 2053.770 996.000 2054.050 1000.000 ;
        RECT 2056.070 999.870 2057.420 1000.000 ;
      LAYER met2 ;
        RECT 2054.330 995.720 2055.790 998.470 ;
      LAYER met2 ;
        RECT 2056.070 996.000 2056.350 999.870 ;
      LAYER met2 ;
        RECT 2056.630 995.720 2057.630 998.470 ;
      LAYER met2 ;
        RECT 2057.910 996.000 2058.190 1000.000 ;
        RECT 2060.210 999.870 2062.020 1000.000 ;
      LAYER met2 ;
        RECT 2058.470 995.720 2059.930 998.470 ;
      LAYER met2 ;
        RECT 2060.210 996.000 2060.490 999.870 ;
      LAYER met2 ;
        RECT 2060.770 995.720 2062.230 998.470 ;
      LAYER met2 ;
        RECT 2062.510 996.000 2062.790 1000.000 ;
        RECT 2064.810 999.870 2066.160 1000.000 ;
      LAYER met2 ;
        RECT 2063.070 995.720 2064.530 998.470 ;
      LAYER met2 ;
        RECT 2064.810 996.000 2065.090 999.870 ;
      LAYER met2 ;
        RECT 2065.370 995.720 2066.370 998.470 ;
      LAYER met2 ;
        RECT 2066.650 996.000 2066.930 1000.000 ;
        RECT 2068.950 999.870 2069.380 1000.000 ;
      LAYER met2 ;
        RECT 2067.210 995.720 2068.670 998.470 ;
      LAYER met2 ;
        RECT 2068.950 996.000 2069.230 999.870 ;
      LAYER met2 ;
        RECT 2069.510 995.720 2070.970 998.470 ;
      LAYER met2 ;
        RECT 2071.250 996.000 2071.530 1000.000 ;
        RECT 2073.090 999.870 2074.900 1000.000 ;
      LAYER met2 ;
        RECT 2071.810 995.720 2072.810 998.470 ;
      LAYER met2 ;
        RECT 2073.090 996.000 2073.370 999.870 ;
      LAYER met2 ;
        RECT 2073.650 995.720 2075.110 998.470 ;
      LAYER met2 ;
        RECT 2075.390 996.000 2075.670 1000.000 ;
        RECT 2077.690 999.870 2079.500 1000.000 ;
      LAYER met2 ;
        RECT 2075.950 995.720 2077.410 998.470 ;
      LAYER met2 ;
        RECT 2077.690 996.000 2077.970 999.870 ;
      LAYER met2 ;
        RECT 2078.250 995.720 2079.710 998.470 ;
      LAYER met2 ;
        RECT 2079.990 996.000 2080.270 1000.000 ;
        RECT 2081.830 999.870 2083.180 1000.000 ;
      LAYER met2 ;
        RECT 2080.550 995.720 2081.550 998.470 ;
      LAYER met2 ;
        RECT 2081.830 996.000 2082.110 999.870 ;
      LAYER met2 ;
        RECT 2082.390 995.720 2083.850 998.470 ;
      LAYER met2 ;
        RECT 2084.130 996.000 2084.410 1000.000 ;
      LAYER met2 ;
        RECT 2084.690 995.720 2086.150 998.470 ;
      LAYER met2 ;
        RECT 2086.430 996.000 2086.710 1000.000 ;
      LAYER met2 ;
        RECT 2086.990 995.720 2087.990 998.470 ;
      LAYER met2 ;
        RECT 2088.270 996.000 2088.550 1000.000 ;
      LAYER met2 ;
        RECT 2088.830 995.720 2090.290 998.470 ;
      LAYER met2 ;
        RECT 2090.570 996.000 2090.850 1000.000 ;
      LAYER met2 ;
        RECT 2091.130 995.720 2092.590 998.470 ;
      LAYER met2 ;
        RECT 2092.870 996.000 2093.150 1000.000 ;
      LAYER met2 ;
        RECT 2093.430 995.720 2094.890 998.470 ;
      LAYER met2 ;
        RECT 2095.170 996.000 2095.450 1000.000 ;
      LAYER met2 ;
        RECT 2095.730 995.720 2096.730 998.470 ;
      LAYER met2 ;
        RECT 2097.010 996.000 2097.290 1000.000 ;
      LAYER met2 ;
        RECT 2097.570 995.720 2099.030 998.470 ;
      LAYER met2 ;
        RECT 2099.310 996.000 2099.590 1000.000 ;
      LAYER met2 ;
        RECT 2099.870 995.720 2101.330 998.470 ;
      LAYER met2 ;
        RECT 2101.610 996.000 2101.890 1000.000 ;
      LAYER met2 ;
        RECT 2102.170 995.720 2103.170 998.470 ;
      LAYER met2 ;
        RECT 2103.450 996.000 2103.730 1000.000 ;
      LAYER met2 ;
        RECT 2104.010 995.720 2105.470 998.470 ;
      LAYER met2 ;
        RECT 2105.750 996.000 2106.030 1000.000 ;
      LAYER met2 ;
        RECT 2106.310 995.720 2107.770 998.470 ;
      LAYER met2 ;
        RECT 2108.050 996.000 2108.330 1000.000 ;
      LAYER met2 ;
        RECT 2108.610 995.720 2110.070 998.470 ;
      LAYER met2 ;
        RECT 2110.350 996.000 2110.630 1000.000 ;
      LAYER met2 ;
        RECT 2110.910 995.720 2111.910 998.470 ;
      LAYER met2 ;
        RECT 2112.190 996.000 2112.470 1000.000 ;
      LAYER met2 ;
        RECT 2112.750 995.720 2114.210 998.470 ;
      LAYER met2 ;
        RECT 2114.490 996.000 2114.770 1000.000 ;
      LAYER met2 ;
        RECT 2115.050 995.720 2116.510 998.470 ;
      LAYER met2 ;
        RECT 2116.790 996.000 2117.070 1000.000 ;
      LAYER met2 ;
        RECT 2117.350 995.720 2118.350 998.470 ;
      LAYER met2 ;
        RECT 2118.630 996.000 2118.910 1000.000 ;
      LAYER met2 ;
        RECT 2119.190 995.720 2120.650 998.470 ;
      LAYER met2 ;
        RECT 2120.930 996.000 2121.210 1000.000 ;
      LAYER met2 ;
        RECT 2121.490 995.720 2122.950 998.470 ;
      LAYER met2 ;
        RECT 2123.230 996.000 2123.510 1000.000 ;
      LAYER met2 ;
        RECT 2123.790 995.720 2125.250 998.470 ;
      LAYER met2 ;
        RECT 2125.530 996.000 2125.810 1000.000 ;
      LAYER met2 ;
        RECT 2126.090 995.720 2127.090 998.470 ;
      LAYER met2 ;
        RECT 2127.370 996.000 2127.650 1000.000 ;
      LAYER met2 ;
        RECT 2127.930 995.720 2129.390 998.470 ;
      LAYER met2 ;
        RECT 2129.670 996.000 2129.950 1000.000 ;
      LAYER met2 ;
        RECT 2130.230 995.720 2131.690 998.470 ;
      LAYER met2 ;
        RECT 2131.970 996.000 2132.250 1000.000 ;
      LAYER met2 ;
        RECT 2132.530 995.720 2133.530 998.470 ;
      LAYER met2 ;
        RECT 2133.810 996.000 2134.090 1000.000 ;
      LAYER met2 ;
        RECT 2134.370 995.720 2135.830 998.470 ;
      LAYER met2 ;
        RECT 2136.110 996.000 2136.390 1000.000 ;
      LAYER met2 ;
        RECT 2136.670 995.720 2138.130 998.470 ;
      LAYER met2 ;
        RECT 2138.410 996.000 2138.690 1000.000 ;
      LAYER met2 ;
        RECT 2138.970 995.720 2140.430 998.470 ;
      LAYER met2 ;
        RECT 2140.710 996.000 2140.990 1000.000 ;
      LAYER met2 ;
        RECT 2141.270 995.720 2142.270 998.470 ;
      LAYER met2 ;
        RECT 2142.550 996.000 2142.830 1000.000 ;
      LAYER met2 ;
        RECT 2143.110 995.720 2144.570 998.470 ;
      LAYER met2 ;
        RECT 2144.850 996.000 2145.130 1000.000 ;
      LAYER met2 ;
        RECT 2145.410 995.720 2146.870 998.470 ;
      LAYER met2 ;
        RECT 2147.150 996.000 2147.430 1000.000 ;
      LAYER met2 ;
        RECT 2147.710 995.720 2148.710 998.470 ;
      LAYER met2 ;
        RECT 2148.990 996.000 2149.270 1000.000 ;
      LAYER met2 ;
        RECT 2149.550 995.720 2151.010 998.470 ;
      LAYER met2 ;
        RECT 2151.290 996.000 2151.570 1000.000 ;
      LAYER met2 ;
        RECT 2151.850 995.720 2153.310 998.470 ;
      LAYER met2 ;
        RECT 2153.590 996.000 2153.870 1000.000 ;
      LAYER met2 ;
        RECT 2154.150 995.720 2155.610 998.470 ;
      LAYER met2 ;
        RECT 2155.890 996.000 2156.170 1000.000 ;
      LAYER met2 ;
        RECT 2156.450 995.720 2157.450 998.470 ;
      LAYER met2 ;
        RECT 2157.730 996.000 2158.010 1000.000 ;
      LAYER met2 ;
        RECT 2158.290 995.720 2159.750 998.470 ;
      LAYER met2 ;
        RECT 2160.030 996.000 2160.310 1000.000 ;
      LAYER met2 ;
        RECT 2160.590 995.720 2162.050 998.470 ;
      LAYER met2 ;
        RECT 2162.330 996.000 2162.610 1000.000 ;
      LAYER met2 ;
        RECT 2162.890 995.720 2163.890 998.470 ;
      LAYER met2 ;
        RECT 2164.170 996.000 2164.450 1000.000 ;
        RECT 2166.470 996.000 2166.750 1000.000 ;
        RECT 2168.770 996.000 2169.050 1000.000 ;
      LAYER met2 ;
        RECT 670.100 604.280 2164.380 995.720 ;
        RECT 670.100 602.195 671.190 604.280 ;
        RECT 672.030 602.195 673.950 604.280 ;
        RECT 674.790 602.195 677.170 604.280 ;
        RECT 678.010 602.195 679.930 604.280 ;
        RECT 680.770 602.195 683.150 604.280 ;
        RECT 683.990 602.195 686.370 604.280 ;
        RECT 687.210 602.195 689.130 604.280 ;
        RECT 689.970 602.195 692.350 604.280 ;
        RECT 693.190 602.195 695.570 604.280 ;
        RECT 696.410 602.195 698.330 604.280 ;
        RECT 699.170 602.195 701.550 604.280 ;
        RECT 702.390 602.195 704.770 604.280 ;
        RECT 705.610 602.195 707.530 604.280 ;
        RECT 708.370 602.195 710.750 604.280 ;
        RECT 711.590 602.195 713.510 604.280 ;
        RECT 714.350 602.195 716.730 604.280 ;
        RECT 717.570 602.195 719.950 604.280 ;
        RECT 720.790 602.195 722.710 604.280 ;
        RECT 723.550 602.195 725.930 604.280 ;
        RECT 726.770 602.195 729.150 604.280 ;
        RECT 729.990 602.195 731.910 604.280 ;
        RECT 732.750 602.195 735.130 604.280 ;
        RECT 735.970 602.195 738.350 604.280 ;
        RECT 739.190 602.195 741.110 604.280 ;
        RECT 741.950 602.195 744.330 604.280 ;
        RECT 745.170 602.195 747.550 604.280 ;
        RECT 748.390 602.195 750.310 604.280 ;
        RECT 751.150 602.195 753.530 604.280 ;
        RECT 754.370 602.195 756.290 604.280 ;
        RECT 757.130 602.195 759.510 604.280 ;
        RECT 760.350 602.195 762.730 604.280 ;
        RECT 763.570 602.195 765.490 604.280 ;
        RECT 766.330 602.195 768.710 604.280 ;
        RECT 769.550 602.195 771.930 604.280 ;
        RECT 772.770 602.195 774.690 604.280 ;
        RECT 775.530 602.195 777.910 604.280 ;
        RECT 778.750 602.195 781.130 604.280 ;
        RECT 781.970 602.195 783.890 604.280 ;
        RECT 784.730 602.195 787.110 604.280 ;
        RECT 787.950 602.195 790.330 604.280 ;
        RECT 791.170 602.195 793.090 604.280 ;
        RECT 793.930 602.195 796.310 604.280 ;
        RECT 797.150 602.195 799.070 604.280 ;
        RECT 799.910 602.195 802.290 604.280 ;
        RECT 803.130 602.195 805.510 604.280 ;
        RECT 806.350 602.195 808.270 604.280 ;
        RECT 809.110 602.195 811.490 604.280 ;
        RECT 812.330 602.195 814.710 604.280 ;
        RECT 815.550 602.195 817.470 604.280 ;
        RECT 818.310 602.195 820.690 604.280 ;
        RECT 821.530 602.195 823.910 604.280 ;
        RECT 824.750 602.195 826.670 604.280 ;
        RECT 827.510 602.195 829.890 604.280 ;
        RECT 830.730 602.195 833.110 604.280 ;
        RECT 833.950 602.195 835.870 604.280 ;
        RECT 836.710 602.195 839.090 604.280 ;
        RECT 839.930 602.195 841.850 604.280 ;
        RECT 842.690 602.195 845.070 604.280 ;
        RECT 845.910 602.195 848.290 604.280 ;
        RECT 849.130 602.195 851.050 604.280 ;
        RECT 851.890 602.195 854.270 604.280 ;
        RECT 855.110 602.195 857.490 604.280 ;
        RECT 858.330 602.195 860.250 604.280 ;
        RECT 861.090 602.195 863.470 604.280 ;
        RECT 864.310 602.195 866.690 604.280 ;
        RECT 867.530 602.195 869.450 604.280 ;
        RECT 870.290 602.195 872.670 604.280 ;
        RECT 873.510 602.195 875.430 604.280 ;
        RECT 876.270 602.195 878.650 604.280 ;
        RECT 879.490 602.195 881.870 604.280 ;
        RECT 882.710 602.195 884.630 604.280 ;
        RECT 885.470 602.195 887.850 604.280 ;
        RECT 888.690 602.195 891.070 604.280 ;
        RECT 891.910 602.195 893.830 604.280 ;
        RECT 894.670 602.195 897.050 604.280 ;
        RECT 897.890 602.195 900.270 604.280 ;
        RECT 901.110 602.195 903.030 604.280 ;
        RECT 903.870 602.195 906.250 604.280 ;
        RECT 907.090 602.195 909.470 604.280 ;
        RECT 910.310 602.195 912.230 604.280 ;
        RECT 913.070 602.195 915.450 604.280 ;
        RECT 916.290 602.195 918.210 604.280 ;
        RECT 919.050 602.195 921.430 604.280 ;
        RECT 922.270 602.195 924.650 604.280 ;
        RECT 925.490 602.195 927.410 604.280 ;
        RECT 928.250 602.195 930.630 604.280 ;
        RECT 931.470 602.195 933.850 604.280 ;
        RECT 934.690 602.195 936.610 604.280 ;
        RECT 937.450 602.195 939.830 604.280 ;
        RECT 940.670 602.195 943.050 604.280 ;
        RECT 943.890 602.195 945.810 604.280 ;
        RECT 946.650 602.195 949.030 604.280 ;
        RECT 949.870 602.195 952.250 604.280 ;
        RECT 953.090 602.195 955.010 604.280 ;
        RECT 955.850 602.195 958.230 604.280 ;
        RECT 959.070 602.195 960.990 604.280 ;
        RECT 961.830 602.195 964.210 604.280 ;
        RECT 965.050 602.195 967.430 604.280 ;
        RECT 968.270 602.195 970.190 604.280 ;
        RECT 971.030 602.195 973.410 604.280 ;
        RECT 974.250 602.195 976.630 604.280 ;
        RECT 977.470 602.195 979.390 604.280 ;
        RECT 980.230 602.195 982.610 604.280 ;
        RECT 983.450 602.195 985.830 604.280 ;
        RECT 986.670 602.195 988.590 604.280 ;
        RECT 989.430 602.195 991.810 604.280 ;
        RECT 992.650 602.195 995.030 604.280 ;
        RECT 995.870 602.195 997.790 604.280 ;
        RECT 998.630 602.195 1001.010 604.280 ;
        RECT 1001.850 602.195 1003.770 604.280 ;
        RECT 1004.610 602.195 1006.990 604.280 ;
        RECT 1007.830 602.195 1010.210 604.280 ;
        RECT 1011.050 602.195 1012.970 604.280 ;
        RECT 1013.810 602.195 1016.190 604.280 ;
        RECT 1017.030 602.195 1019.410 604.280 ;
        RECT 1020.250 602.195 1022.170 604.280 ;
        RECT 1023.010 602.195 1025.390 604.280 ;
        RECT 1026.230 602.195 1028.610 604.280 ;
        RECT 1029.450 602.195 1031.370 604.280 ;
        RECT 1032.210 602.195 1034.590 604.280 ;
        RECT 1035.430 602.195 1037.350 604.280 ;
        RECT 1038.190 602.195 1040.570 604.280 ;
        RECT 1041.410 602.195 1043.790 604.280 ;
        RECT 1044.630 602.195 1046.550 604.280 ;
        RECT 1047.390 602.195 1049.770 604.280 ;
        RECT 1050.610 602.195 1052.990 604.280 ;
        RECT 1053.830 602.195 1055.750 604.280 ;
        RECT 1056.590 602.195 1058.970 604.280 ;
        RECT 1059.810 602.195 1062.190 604.280 ;
        RECT 1063.030 602.195 1064.950 604.280 ;
        RECT 1065.790 602.195 1068.170 604.280 ;
        RECT 1069.010 602.195 1071.390 604.280 ;
        RECT 1072.230 602.195 1074.150 604.280 ;
        RECT 1074.990 602.195 1077.370 604.280 ;
        RECT 1078.210 602.195 1080.130 604.280 ;
        RECT 1080.970 602.195 1083.350 604.280 ;
        RECT 1084.190 602.195 1086.570 604.280 ;
        RECT 1087.410 602.195 1089.330 604.280 ;
        RECT 1090.170 602.195 1092.550 604.280 ;
        RECT 1093.390 602.195 1095.770 604.280 ;
        RECT 1096.610 602.195 1098.530 604.280 ;
        RECT 1099.370 602.195 1101.750 604.280 ;
        RECT 1102.590 602.195 1104.970 604.280 ;
        RECT 1105.810 602.195 1107.730 604.280 ;
        RECT 1108.570 602.195 1110.950 604.280 ;
        RECT 1111.790 602.195 1114.170 604.280 ;
        RECT 1115.010 602.195 1116.930 604.280 ;
        RECT 1117.770 602.195 1120.150 604.280 ;
        RECT 1120.990 602.195 1122.910 604.280 ;
        RECT 1123.750 602.195 1126.130 604.280 ;
        RECT 1126.970 602.195 1129.350 604.280 ;
        RECT 1130.190 602.195 1132.110 604.280 ;
        RECT 1132.950 602.195 1135.330 604.280 ;
        RECT 1136.170 602.195 1138.550 604.280 ;
        RECT 1139.390 602.195 1141.310 604.280 ;
        RECT 1142.150 602.195 1144.530 604.280 ;
        RECT 1145.370 602.195 1147.750 604.280 ;
        RECT 1148.590 602.195 1150.510 604.280 ;
        RECT 1151.350 602.195 1153.730 604.280 ;
        RECT 1154.570 602.195 1156.950 604.280 ;
        RECT 1157.790 602.195 1159.710 604.280 ;
        RECT 1160.550 602.195 1162.930 604.280 ;
        RECT 1163.770 602.195 1165.690 604.280 ;
        RECT 1166.530 602.195 1168.910 604.280 ;
        RECT 1169.750 602.195 1172.130 604.280 ;
        RECT 1172.970 602.195 1174.890 604.280 ;
        RECT 1175.730 602.195 1178.110 604.280 ;
        RECT 1178.950 602.195 1181.330 604.280 ;
        RECT 1182.170 602.195 1184.090 604.280 ;
        RECT 1184.930 602.195 1187.310 604.280 ;
        RECT 1188.150 602.195 1190.530 604.280 ;
        RECT 1191.370 602.195 1193.290 604.280 ;
        RECT 1194.130 602.195 1196.510 604.280 ;
        RECT 1197.350 602.195 1199.270 604.280 ;
        RECT 1200.110 602.195 1202.490 604.280 ;
        RECT 1203.330 602.195 1205.710 604.280 ;
        RECT 1206.550 602.195 1208.470 604.280 ;
        RECT 1209.310 602.195 1211.690 604.280 ;
        RECT 1212.530 602.195 1214.910 604.280 ;
        RECT 1215.750 602.195 1217.670 604.280 ;
        RECT 1218.510 602.195 1220.890 604.280 ;
        RECT 1221.730 602.195 1224.110 604.280 ;
        RECT 1224.950 602.195 1226.870 604.280 ;
        RECT 1227.710 602.195 1230.090 604.280 ;
        RECT 1230.930 602.195 1233.310 604.280 ;
        RECT 1234.150 602.195 1236.070 604.280 ;
        RECT 1236.910 602.195 1239.290 604.280 ;
        RECT 1240.130 602.195 1242.050 604.280 ;
        RECT 1242.890 602.195 1245.270 604.280 ;
        RECT 1246.110 602.195 1248.490 604.280 ;
        RECT 1249.330 602.195 1251.250 604.280 ;
        RECT 1252.090 602.195 1254.470 604.280 ;
        RECT 1255.310 602.195 1257.690 604.280 ;
        RECT 1258.530 602.195 1260.450 604.280 ;
        RECT 1261.290 602.195 1263.670 604.280 ;
        RECT 1264.510 602.195 1266.890 604.280 ;
        RECT 1267.730 602.195 1269.650 604.280 ;
        RECT 1270.490 602.195 1272.870 604.280 ;
        RECT 1273.710 602.195 1276.090 604.280 ;
        RECT 1276.930 602.195 1278.850 604.280 ;
        RECT 1279.690 602.195 1282.070 604.280 ;
        RECT 1282.910 602.195 1284.830 604.280 ;
        RECT 1285.670 602.195 1288.050 604.280 ;
        RECT 1288.890 602.195 1291.270 604.280 ;
        RECT 1292.110 602.195 1294.030 604.280 ;
        RECT 1294.870 602.195 1297.250 604.280 ;
        RECT 1298.090 602.195 1300.470 604.280 ;
        RECT 1301.310 602.195 1303.230 604.280 ;
        RECT 1304.070 602.195 1306.450 604.280 ;
        RECT 1307.290 602.195 1309.670 604.280 ;
        RECT 1310.510 602.195 1312.430 604.280 ;
        RECT 1313.270 602.195 1315.650 604.280 ;
        RECT 1316.490 602.195 1318.870 604.280 ;
        RECT 1319.710 602.195 1321.630 604.280 ;
        RECT 1322.470 602.195 1324.850 604.280 ;
        RECT 1325.690 602.195 1327.610 604.280 ;
        RECT 1328.450 602.195 1330.830 604.280 ;
        RECT 1331.670 602.195 1334.050 604.280 ;
        RECT 1334.890 602.195 1336.810 604.280 ;
        RECT 1337.650 602.195 1340.030 604.280 ;
        RECT 1340.870 602.195 1343.250 604.280 ;
        RECT 1344.090 602.195 1346.010 604.280 ;
        RECT 1346.850 602.195 1349.230 604.280 ;
        RECT 1350.070 602.195 1352.450 604.280 ;
        RECT 1353.290 602.195 1355.210 604.280 ;
        RECT 1356.050 602.195 1358.430 604.280 ;
        RECT 1359.270 602.195 1361.190 604.280 ;
        RECT 1362.030 602.195 1364.410 604.280 ;
        RECT 1365.250 602.195 1367.630 604.280 ;
        RECT 1368.470 602.195 1370.390 604.280 ;
        RECT 1371.230 602.195 1373.610 604.280 ;
        RECT 1374.450 602.195 1376.830 604.280 ;
        RECT 1377.670 602.195 1379.590 604.280 ;
        RECT 1380.430 602.195 1382.810 604.280 ;
        RECT 1383.650 602.195 1386.030 604.280 ;
        RECT 1386.870 602.195 1388.790 604.280 ;
        RECT 1389.630 602.195 1392.010 604.280 ;
        RECT 1392.850 602.195 1395.230 604.280 ;
        RECT 1396.070 602.195 1397.990 604.280 ;
        RECT 1398.830 602.195 1401.210 604.280 ;
        RECT 1402.050 602.195 1403.970 604.280 ;
        RECT 1404.810 602.195 1407.190 604.280 ;
        RECT 1408.030 602.195 1410.410 604.280 ;
        RECT 1411.250 602.195 1413.170 604.280 ;
        RECT 1414.010 602.195 1416.390 604.280 ;
        RECT 1417.230 602.195 1419.610 604.280 ;
        RECT 1420.450 602.195 1422.370 604.280 ;
        RECT 1423.210 602.195 1425.590 604.280 ;
        RECT 1426.430 602.195 1428.810 604.280 ;
        RECT 1429.650 602.195 1431.570 604.280 ;
        RECT 1432.410 602.195 1434.790 604.280 ;
        RECT 1435.630 602.195 1438.010 604.280 ;
        RECT 1438.850 602.195 1440.770 604.280 ;
        RECT 1441.610 602.195 1443.990 604.280 ;
        RECT 1444.830 602.195 1446.750 604.280 ;
        RECT 1447.590 602.195 1449.970 604.280 ;
        RECT 1450.810 602.195 1453.190 604.280 ;
        RECT 1454.030 602.195 1455.950 604.280 ;
        RECT 1456.790 602.195 1459.170 604.280 ;
        RECT 1460.010 602.195 1462.390 604.280 ;
        RECT 1463.230 602.195 1465.150 604.280 ;
        RECT 1465.990 602.195 1468.370 604.280 ;
        RECT 1469.210 602.195 1471.590 604.280 ;
        RECT 1472.430 602.195 1474.350 604.280 ;
        RECT 1475.190 602.195 1477.570 604.280 ;
        RECT 1478.410 602.195 1480.790 604.280 ;
        RECT 1481.630 602.195 1483.550 604.280 ;
        RECT 1484.390 602.195 1486.770 604.280 ;
        RECT 1487.610 602.195 1489.530 604.280 ;
        RECT 1490.370 602.195 1492.750 604.280 ;
        RECT 1493.590 602.195 1495.970 604.280 ;
        RECT 1496.810 602.195 1498.730 604.280 ;
        RECT 1499.570 602.195 1501.950 604.280 ;
        RECT 1502.790 602.195 1505.170 604.280 ;
        RECT 1506.010 602.195 1507.930 604.280 ;
        RECT 1508.770 602.195 1511.150 604.280 ;
        RECT 1511.990 602.195 1514.370 604.280 ;
        RECT 1515.210 602.195 1517.130 604.280 ;
        RECT 1517.970 602.195 1520.350 604.280 ;
        RECT 1521.190 602.195 1523.110 604.280 ;
        RECT 1523.950 602.195 1526.330 604.280 ;
        RECT 1527.170 602.195 1529.550 604.280 ;
        RECT 1530.390 602.195 1532.310 604.280 ;
        RECT 1533.150 602.195 1535.530 604.280 ;
        RECT 1536.370 602.195 1538.750 604.280 ;
        RECT 1539.590 602.195 1541.510 604.280 ;
        RECT 1542.350 602.195 1544.730 604.280 ;
        RECT 1545.570 602.195 1547.950 604.280 ;
        RECT 1548.790 602.195 1550.710 604.280 ;
        RECT 1551.550 602.195 1553.930 604.280 ;
        RECT 1554.770 602.195 1557.150 604.280 ;
        RECT 1557.990 602.195 1559.910 604.280 ;
        RECT 1560.750 602.195 1563.130 604.280 ;
        RECT 1563.970 602.195 1565.890 604.280 ;
        RECT 1566.730 602.195 1569.110 604.280 ;
        RECT 1569.950 602.195 1572.330 604.280 ;
        RECT 1573.170 602.195 1575.090 604.280 ;
        RECT 1575.930 602.195 1578.310 604.280 ;
        RECT 1579.150 602.195 1581.530 604.280 ;
        RECT 1582.370 602.195 1584.290 604.280 ;
        RECT 1585.130 602.195 1587.510 604.280 ;
        RECT 1588.350 602.195 1590.730 604.280 ;
        RECT 1591.570 602.195 1593.490 604.280 ;
        RECT 1594.330 602.195 1596.710 604.280 ;
        RECT 1597.550 602.195 1599.930 604.280 ;
        RECT 1600.770 602.195 1602.690 604.280 ;
        RECT 1603.530 602.195 1605.910 604.280 ;
        RECT 1606.750 602.195 1608.670 604.280 ;
        RECT 1609.510 602.195 1611.890 604.280 ;
        RECT 1612.730 602.195 1615.110 604.280 ;
        RECT 1615.950 602.195 1617.870 604.280 ;
        RECT 1618.710 602.195 1621.090 604.280 ;
        RECT 1621.930 602.195 1624.310 604.280 ;
        RECT 1625.150 602.195 1627.070 604.280 ;
        RECT 1627.910 602.195 1630.290 604.280 ;
        RECT 1631.130 602.195 1633.510 604.280 ;
        RECT 1634.350 602.195 1636.270 604.280 ;
        RECT 1637.110 602.195 1639.490 604.280 ;
        RECT 1640.330 602.195 1642.710 604.280 ;
        RECT 1643.550 602.195 1645.470 604.280 ;
        RECT 1646.310 602.195 1648.690 604.280 ;
        RECT 1649.530 602.195 1651.450 604.280 ;
        RECT 1652.290 602.195 1654.670 604.280 ;
        RECT 1655.510 602.195 1657.890 604.280 ;
        RECT 1658.730 602.195 1660.650 604.280 ;
        RECT 1661.490 602.195 1663.870 604.280 ;
        RECT 1664.710 602.195 1667.090 604.280 ;
        RECT 1667.930 602.195 1669.850 604.280 ;
        RECT 1670.690 602.195 1673.070 604.280 ;
        RECT 1673.910 602.195 1676.290 604.280 ;
        RECT 1677.130 602.195 1679.050 604.280 ;
        RECT 1679.890 602.195 1682.270 604.280 ;
        RECT 1683.110 602.195 1685.030 604.280 ;
        RECT 1685.870 602.195 1688.250 604.280 ;
        RECT 1689.090 602.195 1691.470 604.280 ;
        RECT 1692.310 602.195 1694.230 604.280 ;
        RECT 1695.070 602.195 1697.450 604.280 ;
        RECT 1698.290 602.195 1700.670 604.280 ;
        RECT 1701.510 602.195 1703.430 604.280 ;
        RECT 1704.270 602.195 1706.650 604.280 ;
        RECT 1707.490 602.195 1709.870 604.280 ;
        RECT 1710.710 602.195 1712.630 604.280 ;
        RECT 1713.470 602.195 1715.850 604.280 ;
        RECT 1716.690 602.195 1719.070 604.280 ;
        RECT 1719.910 602.195 1721.830 604.280 ;
        RECT 1722.670 602.195 1725.050 604.280 ;
        RECT 1725.890 602.195 1727.810 604.280 ;
        RECT 1728.650 602.195 1731.030 604.280 ;
        RECT 1731.870 602.195 1734.250 604.280 ;
        RECT 1735.090 602.195 1737.010 604.280 ;
        RECT 1737.850 602.195 1740.230 604.280 ;
        RECT 1741.070 602.195 1743.450 604.280 ;
        RECT 1744.290 602.195 1746.210 604.280 ;
        RECT 1747.050 602.195 1749.430 604.280 ;
        RECT 1750.270 602.195 1752.650 604.280 ;
        RECT 1753.490 602.195 1755.410 604.280 ;
        RECT 1756.250 602.195 1758.630 604.280 ;
        RECT 1759.470 602.195 1761.850 604.280 ;
        RECT 1762.690 602.195 1764.610 604.280 ;
        RECT 1765.450 602.195 1767.830 604.280 ;
        RECT 1768.670 602.195 1770.590 604.280 ;
        RECT 1771.430 602.195 1773.810 604.280 ;
        RECT 1774.650 602.195 1777.030 604.280 ;
        RECT 1777.870 602.195 1779.790 604.280 ;
        RECT 1780.630 602.195 1783.010 604.280 ;
        RECT 1783.850 602.195 1786.230 604.280 ;
        RECT 1787.070 602.195 1788.990 604.280 ;
        RECT 1789.830 602.195 1792.210 604.280 ;
        RECT 1793.050 602.195 1795.430 604.280 ;
        RECT 1796.270 602.195 1798.190 604.280 ;
        RECT 1799.030 602.195 1801.410 604.280 ;
        RECT 1802.250 602.195 1804.630 604.280 ;
        RECT 1805.470 602.195 1807.390 604.280 ;
        RECT 1808.230 602.195 1810.610 604.280 ;
        RECT 1811.450 602.195 1813.370 604.280 ;
        RECT 1814.210 602.195 1816.590 604.280 ;
        RECT 1817.430 602.195 1819.810 604.280 ;
        RECT 1820.650 602.195 1822.570 604.280 ;
        RECT 1823.410 602.195 1825.790 604.280 ;
        RECT 1826.630 602.195 1829.010 604.280 ;
        RECT 1829.850 602.195 1831.770 604.280 ;
        RECT 1832.610 602.195 1834.990 604.280 ;
        RECT 1835.830 602.195 1838.210 604.280 ;
        RECT 1839.050 602.195 1840.970 604.280 ;
        RECT 1841.810 602.195 1844.190 604.280 ;
        RECT 1845.030 602.195 1846.950 604.280 ;
        RECT 1847.790 602.195 1850.170 604.280 ;
        RECT 1851.010 602.195 1853.390 604.280 ;
        RECT 1854.230 602.195 1856.150 604.280 ;
        RECT 1856.990 602.195 1859.370 604.280 ;
        RECT 1860.210 602.195 1862.590 604.280 ;
        RECT 1863.430 602.195 1865.350 604.280 ;
        RECT 1866.190 602.195 1868.570 604.280 ;
        RECT 1869.410 602.195 1871.790 604.280 ;
        RECT 1872.630 602.195 1874.550 604.280 ;
        RECT 1875.390 602.195 1877.770 604.280 ;
        RECT 1878.610 602.195 1880.990 604.280 ;
        RECT 1881.830 602.195 1883.750 604.280 ;
        RECT 1884.590 602.195 1886.970 604.280 ;
        RECT 1887.810 602.195 1889.730 604.280 ;
        RECT 1890.570 602.195 1892.950 604.280 ;
        RECT 1893.790 602.195 1896.170 604.280 ;
        RECT 1897.010 602.195 1898.930 604.280 ;
        RECT 1899.770 602.195 1902.150 604.280 ;
        RECT 1902.990 602.195 1905.370 604.280 ;
        RECT 1906.210 602.195 1908.130 604.280 ;
        RECT 1908.970 602.195 1911.350 604.280 ;
        RECT 1912.190 602.195 1914.570 604.280 ;
        RECT 1915.410 602.195 1917.330 604.280 ;
        RECT 1918.170 602.195 1920.550 604.280 ;
        RECT 1921.390 602.195 1923.770 604.280 ;
        RECT 1924.610 602.195 1926.530 604.280 ;
        RECT 1927.370 602.195 1929.750 604.280 ;
        RECT 1930.590 602.195 1932.510 604.280 ;
        RECT 1933.350 602.195 1935.730 604.280 ;
        RECT 1936.570 602.195 1938.950 604.280 ;
        RECT 1939.790 602.195 1941.710 604.280 ;
        RECT 1942.550 602.195 1944.930 604.280 ;
        RECT 1945.770 602.195 1948.150 604.280 ;
        RECT 1948.990 602.195 1950.910 604.280 ;
        RECT 1951.750 602.195 1954.130 604.280 ;
        RECT 1954.970 602.195 1957.350 604.280 ;
        RECT 1958.190 602.195 1960.110 604.280 ;
        RECT 1960.950 602.195 1963.330 604.280 ;
        RECT 1964.170 602.195 1966.550 604.280 ;
        RECT 1967.390 602.195 1969.310 604.280 ;
        RECT 1970.150 602.195 1972.530 604.280 ;
        RECT 1973.370 602.195 1975.290 604.280 ;
        RECT 1976.130 602.195 1978.510 604.280 ;
        RECT 1979.350 602.195 1981.730 604.280 ;
        RECT 1982.570 602.195 1984.490 604.280 ;
        RECT 1985.330 602.195 1987.710 604.280 ;
        RECT 1988.550 602.195 1990.930 604.280 ;
        RECT 1991.770 602.195 1993.690 604.280 ;
        RECT 1994.530 602.195 1996.910 604.280 ;
        RECT 1997.750 602.195 2000.130 604.280 ;
        RECT 2000.970 602.195 2002.890 604.280 ;
        RECT 2003.730 602.195 2006.110 604.280 ;
        RECT 2006.950 602.195 2008.870 604.280 ;
        RECT 2009.710 602.195 2012.090 604.280 ;
        RECT 2012.930 602.195 2015.310 604.280 ;
        RECT 2016.150 602.195 2018.070 604.280 ;
        RECT 2018.910 602.195 2021.290 604.280 ;
        RECT 2022.130 602.195 2024.510 604.280 ;
        RECT 2025.350 602.195 2027.270 604.280 ;
        RECT 2028.110 602.195 2030.490 604.280 ;
        RECT 2031.330 602.195 2033.710 604.280 ;
        RECT 2034.550 602.195 2036.470 604.280 ;
        RECT 2037.310 602.195 2039.690 604.280 ;
        RECT 2040.530 602.195 2042.910 604.280 ;
        RECT 2043.750 602.195 2045.670 604.280 ;
        RECT 2046.510 602.195 2048.890 604.280 ;
        RECT 2049.730 602.195 2051.650 604.280 ;
        RECT 2052.490 602.195 2054.870 604.280 ;
        RECT 2055.710 602.195 2058.090 604.280 ;
        RECT 2058.930 602.195 2060.850 604.280 ;
        RECT 2061.690 602.195 2064.070 604.280 ;
        RECT 2064.910 602.195 2067.290 604.280 ;
        RECT 2068.130 602.195 2070.050 604.280 ;
        RECT 2070.890 602.195 2073.270 604.280 ;
        RECT 2074.110 602.195 2076.490 604.280 ;
        RECT 2077.330 602.195 2079.250 604.280 ;
        RECT 2080.090 602.195 2082.470 604.280 ;
        RECT 2083.310 602.195 2085.690 604.280 ;
        RECT 2086.530 602.195 2088.450 604.280 ;
        RECT 2089.290 602.195 2091.670 604.280 ;
        RECT 2092.510 602.195 2094.430 604.280 ;
        RECT 2095.270 602.195 2097.650 604.280 ;
        RECT 2098.490 602.195 2100.870 604.280 ;
        RECT 2101.710 602.195 2103.630 604.280 ;
        RECT 2104.470 602.195 2106.850 604.280 ;
        RECT 2107.690 602.195 2110.070 604.280 ;
        RECT 2110.910 602.195 2112.830 604.280 ;
        RECT 2113.670 602.195 2116.050 604.280 ;
        RECT 2116.890 602.195 2119.270 604.280 ;
        RECT 2120.110 602.195 2122.030 604.280 ;
        RECT 2122.870 602.195 2125.250 604.280 ;
        RECT 2126.090 602.195 2128.470 604.280 ;
        RECT 2129.310 602.195 2131.230 604.280 ;
        RECT 2132.070 602.195 2134.450 604.280 ;
        RECT 2135.290 602.195 2137.210 604.280 ;
        RECT 2138.050 602.195 2140.430 604.280 ;
        RECT 2141.270 602.195 2143.650 604.280 ;
        RECT 2144.490 602.195 2146.410 604.280 ;
        RECT 2147.250 602.195 2149.630 604.280 ;
        RECT 2150.470 602.195 2152.850 604.280 ;
        RECT 2153.690 602.195 2155.610 604.280 ;
        RECT 2156.450 602.195 2158.830 604.280 ;
        RECT 2159.670 602.195 2162.050 604.280 ;
        RECT 2162.890 602.195 2164.380 604.280 ;
      LAYER met2 ;
        RECT 2168.310 600.000 2168.590 604.000 ;
      LAYER via2 ;
        RECT 1351.110 2842.600 1351.390 2842.880 ;
        RECT 1352.950 2842.600 1353.230 2842.880 ;
        RECT 420.530 2729.040 420.810 2729.320 ;
        RECT 420.070 2707.280 420.350 2707.560 ;
        RECT 588.890 2686.880 589.170 2687.160 ;
        RECT 588.890 2666.480 589.170 2666.760 ;
        RECT 978.970 1014.080 979.250 1014.360 ;
        RECT 978.510 1012.040 978.790 1012.320 ;
        RECT 979.430 1011.360 979.710 1011.640 ;
        RECT 985.410 1012.720 985.690 1013.000 ;
        RECT 993.230 2783.440 993.510 2783.720 ;
        RECT 992.770 2739.240 993.050 2739.520 ;
        RECT 992.310 2718.840 992.590 2719.120 ;
        RECT 987.250 2646.080 987.530 2646.360 ;
        RECT 991.850 2622.960 992.130 2623.240 ;
        RECT 991.390 1955.880 991.670 1956.160 ;
        RECT 990.930 1935.480 991.210 1935.760 ;
        RECT 990.470 1893.320 990.750 1893.600 ;
        RECT 990.010 1871.560 990.290 1871.840 ;
        RECT 989.550 1851.160 989.830 1851.440 ;
        RECT 989.090 1809.000 989.370 1809.280 ;
        RECT 988.630 1787.240 988.910 1787.520 ;
        RECT 988.170 1766.840 988.450 1767.120 ;
        RECT 987.710 1745.080 987.990 1745.360 ;
        RECT 986.330 1010.680 986.610 1010.960 ;
        RECT 985.870 1010.000 986.150 1010.280 ;
        RECT 993.690 2760.320 993.970 2760.600 ;
        RECT 994.150 2692.320 994.430 2692.600 ;
        RECT 994.610 2670.560 994.890 2670.840 ;
        RECT 994.150 1013.400 994.430 1013.680 ;
        RECT 993.230 1009.320 993.510 1009.600 ;
        RECT 995.070 2018.440 995.350 2018.720 ;
        RECT 995.530 1998.040 995.810 1998.320 ;
        RECT 995.990 1976.280 996.270 1976.560 ;
        RECT 996.450 1913.720 996.730 1914.000 ;
        RECT 996.910 1829.400 997.190 1829.680 ;
        RECT 997.370 1724.680 997.650 1724.960 ;
        RECT 1110.990 2780.720 1111.270 2781.000 ;
        RECT 1097.190 2644.720 1097.470 2645.000 ;
        RECT 1097.650 2622.280 1097.930 2622.560 ;
        RECT 1111.450 2760.320 1111.730 2760.600 ;
        RECT 1111.910 2734.480 1112.190 2734.760 ;
        RECT 1112.370 2712.720 1112.650 2713.000 ;
        RECT 1112.830 2691.640 1113.110 2691.920 ;
        RECT 1113.290 2666.480 1113.570 2666.760 ;
        RECT 1350.190 2601.200 1350.470 2601.480 ;
        RECT 1351.110 2601.200 1351.390 2601.480 ;
        RECT 1351.570 2559.720 1351.850 2560.000 ;
        RECT 1350.190 2559.040 1350.470 2559.320 ;
        RECT 1351.110 2463.160 1351.390 2463.440 ;
        RECT 1352.030 2463.160 1352.310 2463.440 ;
        RECT 1350.190 2270.040 1350.470 2270.320 ;
        RECT 1351.110 2270.040 1351.390 2270.320 ;
        RECT 1350.190 2173.480 1350.470 2173.760 ;
        RECT 1351.110 2173.480 1351.390 2173.760 ;
        RECT 1065.910 1009.320 1066.190 1009.600 ;
        RECT 1087.530 1010.000 1087.810 1010.280 ;
        RECT 1100.870 1014.080 1101.150 1014.360 ;
        RECT 1124.790 1013.400 1125.070 1013.680 ;
        RECT 1117.890 1012.040 1118.170 1012.320 ;
        RECT 1128.930 1012.720 1129.210 1013.000 ;
        RECT 1141.810 1011.360 1142.090 1011.640 ;
        RECT 1166.190 1010.680 1166.470 1010.960 ;
        RECT 1334.090 1998.040 1334.370 1998.320 ;
        RECT 1334.550 1787.240 1334.830 1787.520 ;
        RECT 1336.850 1745.080 1337.130 1745.360 ;
        RECT 1337.310 1724.680 1337.590 1724.960 ;
        RECT 1338.690 2018.440 1338.970 2018.720 ;
        RECT 1339.150 1976.280 1339.430 1976.560 ;
        RECT 1339.610 1955.880 1339.890 1956.160 ;
        RECT 1340.070 1934.120 1340.350 1934.400 ;
        RECT 1340.530 1913.720 1340.810 1914.000 ;
        RECT 1340.990 1891.960 1341.270 1892.240 ;
        RECT 1341.450 1871.560 1341.730 1871.840 ;
        RECT 1341.910 1849.800 1342.190 1850.080 ;
        RECT 1342.370 1829.400 1342.650 1829.680 ;
        RECT 1342.830 1807.640 1343.110 1807.920 ;
        RECT 1343.290 1766.840 1343.570 1767.120 ;
        RECT 1352.030 1883.800 1352.310 1884.080 ;
        RECT 1350.190 1882.440 1350.470 1882.720 ;
        RECT 1351.110 1607.720 1351.390 1608.000 ;
        RECT 1351.570 1607.040 1351.850 1607.320 ;
        RECT 1350.650 1255.480 1350.930 1255.760 ;
        RECT 1351.570 1255.480 1351.850 1255.760 ;
        RECT 1351.570 1207.200 1351.850 1207.480 ;
        RECT 1350.190 1206.520 1350.470 1206.800 ;
        RECT 1490.030 2850.080 1490.310 2850.360 ;
        RECT 1490.030 2830.360 1490.310 2830.640 ;
        RECT 1490.030 2801.800 1490.310 2802.080 ;
        RECT 1485.430 2784.120 1485.710 2784.400 ;
        RECT 1489.570 2767.800 1489.850 2768.080 ;
        RECT 1487.270 2739.240 1487.550 2739.520 ;
        RECT 1486.810 2720.200 1487.090 2720.480 ;
        RECT 1482.670 2656.960 1482.950 2657.240 ;
        RECT 1484.510 2548.840 1484.790 2549.120 ;
        RECT 1489.110 2691.640 1489.390 2691.920 ;
        RECT 1489.110 2673.960 1489.390 2674.240 ;
        RECT 1488.190 2629.080 1488.470 2629.360 ;
        RECT 1488.650 2610.040 1488.930 2610.320 ;
        RECT 1488.190 2595.080 1488.470 2595.360 ;
        RECT 1488.190 2580.800 1488.470 2581.080 ;
        RECT 1488.190 2567.200 1488.470 2567.480 ;
        RECT 1487.730 2518.920 1488.010 2519.200 ;
        RECT 1496.010 2753.520 1496.290 2753.800 ;
        RECT 1514.870 2463.160 1515.150 2463.440 ;
        RECT 1532.350 2463.160 1532.630 2463.440 ;
        RECT 1532.350 2270.040 1532.630 2270.320 ;
        RECT 1533.270 2270.040 1533.550 2270.320 ;
        RECT 1532.350 2062.640 1532.630 2062.920 ;
        RECT 1532.810 2027.960 1533.090 2028.240 ;
        RECT 1531.430 1690.000 1531.710 1690.280 ;
        RECT 1532.810 1690.000 1533.090 1690.280 ;
        RECT 1532.810 1496.880 1533.090 1497.160 ;
        RECT 1534.190 1496.880 1534.470 1497.160 ;
        RECT 1534.190 1449.280 1534.470 1449.560 ;
        RECT 1533.270 1448.600 1533.550 1448.880 ;
        RECT 1532.810 1386.720 1533.090 1387.000 ;
        RECT 1533.730 1386.720 1534.010 1387.000 ;
        RECT 1531.430 1248.680 1531.710 1248.960 ;
        RECT 1532.810 1248.680 1533.090 1248.960 ;
        RECT 1543.390 1345.240 1543.670 1345.520 ;
        RECT 1544.310 1345.240 1544.590 1345.520 ;
        RECT 1559.490 2319.000 1559.770 2319.280 ;
        RECT 1559.490 2318.320 1559.770 2318.600 ;
        RECT 1573.750 2319.000 1574.030 2319.280 ;
        RECT 1573.750 2318.320 1574.030 2318.600 ;
        RECT 1573.750 1835.520 1574.030 1835.800 ;
        RECT 1574.670 1835.520 1574.950 1835.800 ;
        RECT 1573.750 1738.960 1574.030 1739.240 ;
        RECT 1574.670 1738.960 1574.950 1739.240 ;
        RECT 1573.750 1014.080 1574.030 1014.360 ;
        RECT 1575.590 1014.080 1575.870 1014.360 ;
        RECT 1751.310 1012.720 1751.590 1013.000 ;
        RECT 1753.150 1012.720 1753.430 1013.000 ;
        RECT 1890.690 2848.380 1890.970 2848.660 ;
        RECT 1891.150 2832.060 1891.430 2832.340 ;
        RECT 1891.610 2817.100 1891.890 2817.380 ;
        RECT 1892.070 2797.720 1892.350 2798.000 ;
        RECT 1892.530 2782.760 1892.810 2783.040 ;
        RECT 1893.450 2753.520 1893.730 2753.800 ;
        RECT 1892.990 2718.840 1893.270 2719.120 ;
        RECT 1894.370 2735.160 1894.650 2735.440 ;
        RECT 1897.590 2767.120 1897.870 2767.400 ;
        RECT 1898.050 2687.560 1898.330 2687.840 ;
        RECT 1898.510 2672.600 1898.790 2672.880 ;
        RECT 1898.970 2656.960 1899.250 2657.240 ;
        RECT 1899.430 2625.000 1899.710 2625.280 ;
        RECT 1899.890 2608.680 1900.170 2608.960 ;
        RECT 1900.350 2577.400 1900.630 2577.680 ;
        RECT 1900.810 2562.440 1901.090 2562.720 ;
        RECT 1901.270 2547.480 1901.550 2547.760 ;
        RECT 1903.570 2514.840 1903.850 2515.120 ;
        RECT 1904.490 1885.840 1904.770 1886.120 ;
        RECT 1904.490 1870.200 1904.770 1870.480 ;
        RECT 1904.490 1851.840 1904.770 1852.120 ;
        RECT 1904.490 1817.840 1904.770 1818.120 ;
        RECT 1904.490 1767.520 1904.770 1767.800 ;
        RECT 2087.110 1884.480 2087.390 1884.760 ;
        RECT 2084.350 1850.480 2084.630 1850.760 ;
        RECT 2084.810 1835.520 2085.090 1835.800 ;
        RECT 2085.270 1816.480 2085.550 1816.760 ;
        RECT 2085.730 1800.840 2086.010 1801.120 ;
        RECT 2086.190 1782.480 2086.470 1782.760 ;
        RECT 2086.650 1766.840 2086.930 1767.120 ;
        RECT 2287.210 1877.000 2287.490 1877.280 ;
        RECT 2287.670 1789.960 2287.950 1790.240 ;
        RECT 2539.290 1891.960 2539.570 1892.240 ;
        RECT 2539.750 1804.920 2540.030 1805.200 ;
        RECT 2540.210 1719.240 2540.490 1719.520 ;
      LAYER met3 ;
        RECT 1504.000 2881.840 1885.335 2889.125 ;
        RECT 1504.400 2880.480 1885.335 2881.840 ;
        RECT 1504.400 2880.440 1884.935 2880.480 ;
        RECT 1504.000 2879.080 1884.935 2880.440 ;
        RECT 1504.000 2865.520 1885.335 2879.080 ;
        RECT 1504.400 2864.160 1885.335 2865.520 ;
        RECT 1504.400 2864.120 1884.935 2864.160 ;
        RECT 1504.000 2862.760 1884.935 2864.120 ;
        RECT 1504.000 2850.560 1885.335 2862.760 ;
      LAYER met3 ;
        RECT 1490.005 2850.370 1490.335 2850.385 ;
        RECT 1490.005 2850.160 1500.210 2850.370 ;
        RECT 1490.005 2850.070 1504.000 2850.160 ;
        RECT 1490.005 2850.055 1490.335 2850.070 ;
        RECT 1499.910 2849.880 1504.000 2850.070 ;
        RECT 1500.000 2849.560 1504.000 2849.880 ;
      LAYER met3 ;
        RECT 1504.400 2849.200 1885.335 2850.560 ;
        RECT 1504.400 2849.160 1884.935 2849.200 ;
        RECT 1504.000 2847.800 1884.935 2849.160 ;
      LAYER met3 ;
        RECT 1885.335 2848.670 1889.335 2848.800 ;
        RECT 1890.665 2848.670 1890.995 2848.685 ;
        RECT 1885.335 2848.370 1890.995 2848.670 ;
        RECT 1885.335 2848.200 1889.335 2848.370 ;
        RECT 1890.665 2848.355 1890.995 2848.370 ;
        RECT 1351.085 2842.890 1351.415 2842.905 ;
        RECT 1352.925 2842.890 1353.255 2842.905 ;
        RECT 1351.085 2842.590 1353.255 2842.890 ;
        RECT 1351.085 2842.575 1351.415 2842.590 ;
        RECT 1352.925 2842.575 1353.255 2842.590 ;
      LAYER met3 ;
        RECT 1504.000 2834.240 1885.335 2847.800 ;
      LAYER met3 ;
        RECT 1500.000 2833.560 1504.000 2833.840 ;
        RECT 1499.910 2833.240 1504.000 2833.560 ;
        RECT 1490.005 2830.650 1490.335 2830.665 ;
        RECT 1499.910 2830.650 1500.210 2833.240 ;
      LAYER met3 ;
        RECT 1504.400 2832.880 1885.335 2834.240 ;
        RECT 1504.400 2832.840 1884.935 2832.880 ;
      LAYER met3 ;
        RECT 1490.005 2830.350 1500.210 2830.650 ;
      LAYER met3 ;
        RECT 1504.000 2831.480 1884.935 2832.840 ;
      LAYER met3 ;
        RECT 1885.335 2832.350 1889.335 2832.480 ;
        RECT 1891.125 2832.350 1891.455 2832.365 ;
        RECT 1885.335 2832.050 1891.455 2832.350 ;
        RECT 1885.335 2831.880 1889.335 2832.050 ;
        RECT 1891.125 2832.035 1891.455 2832.050 ;
        RECT 1490.005 2830.335 1490.335 2830.350 ;
      LAYER met3 ;
        RECT 1504.000 2819.280 1885.335 2831.480 ;
        RECT 1504.400 2817.920 1885.335 2819.280 ;
        RECT 1504.400 2817.880 1884.935 2817.920 ;
        RECT 1504.000 2816.520 1884.935 2817.880 ;
      LAYER met3 ;
        RECT 1885.335 2817.390 1889.335 2817.520 ;
        RECT 1891.585 2817.390 1891.915 2817.405 ;
        RECT 1885.335 2817.090 1891.915 2817.390 ;
        RECT 1885.335 2816.920 1889.335 2817.090 ;
        RECT 1891.585 2817.075 1891.915 2817.090 ;
      LAYER met3 ;
        RECT 1504.000 2802.960 1885.335 2816.520 ;
      LAYER met3 ;
        RECT 1500.000 2802.280 1504.000 2802.560 ;
        RECT 1490.005 2802.090 1490.335 2802.105 ;
        RECT 1499.910 2802.090 1504.000 2802.280 ;
        RECT 1490.005 2801.960 1504.000 2802.090 ;
        RECT 1490.005 2801.790 1500.210 2801.960 ;
        RECT 1490.005 2801.775 1490.335 2801.790 ;
      LAYER met3 ;
        RECT 1504.400 2801.600 1885.335 2802.960 ;
        RECT 1504.400 2801.560 1884.935 2801.600 ;
        RECT 1504.000 2800.200 1884.935 2801.560 ;
      LAYER met3 ;
        RECT 1885.335 2800.920 1889.335 2801.200 ;
        RECT 1885.335 2800.600 1889.370 2800.920 ;
      LAYER met3 ;
        RECT 1504.000 2788.000 1885.335 2800.200 ;
      LAYER met3 ;
        RECT 1889.070 2798.010 1889.370 2800.600 ;
        RECT 1892.045 2798.010 1892.375 2798.025 ;
        RECT 1889.070 2797.710 1892.375 2798.010 ;
        RECT 1892.045 2797.695 1892.375 2797.710 ;
      LAYER met3 ;
        RECT 1004.000 2787.360 1096.000 2787.845 ;
      LAYER met3 ;
        RECT 1000.000 2786.360 1004.000 2786.960 ;
        RECT 993.205 2783.730 993.535 2783.745 ;
        RECT 1000.350 2783.730 1000.650 2786.360 ;
      LAYER met3 ;
        RECT 1004.400 2785.960 1096.000 2787.360 ;
      LAYER met3 ;
        RECT 1500.000 2787.320 1504.000 2787.600 ;
        RECT 993.205 2783.430 1000.650 2783.730 ;
      LAYER met3 ;
        RECT 1004.000 2784.640 1096.000 2785.960 ;
      LAYER met3 ;
        RECT 1499.910 2787.000 1504.000 2787.320 ;
        RECT 993.205 2783.415 993.535 2783.430 ;
      LAYER met3 ;
        RECT 1004.000 2783.240 1095.600 2784.640 ;
      LAYER met3 ;
        RECT 1485.405 2784.410 1485.735 2784.425 ;
        RECT 1499.910 2784.410 1500.210 2787.000 ;
      LAYER met3 ;
        RECT 1504.400 2786.640 1885.335 2788.000 ;
        RECT 1504.400 2786.600 1884.935 2786.640 ;
      LAYER met3 ;
        RECT 1096.000 2783.920 1100.000 2784.240 ;
        RECT 1485.405 2784.110 1500.210 2784.410 ;
      LAYER met3 ;
        RECT 1504.000 2785.240 1884.935 2786.600 ;
      LAYER met3 ;
        RECT 1885.335 2785.960 1889.335 2786.240 ;
        RECT 1885.335 2785.640 1889.370 2785.960 ;
        RECT 1485.405 2784.095 1485.735 2784.110 ;
        RECT 1096.000 2783.640 1100.010 2783.920 ;
      LAYER met3 ;
        RECT 1004.000 2764.240 1096.000 2783.240 ;
      LAYER met3 ;
        RECT 1099.710 2781.010 1100.010 2783.640 ;
        RECT 1110.965 2781.010 1111.295 2781.025 ;
        RECT 1099.710 2780.710 1111.295 2781.010 ;
        RECT 1110.965 2780.695 1111.295 2780.710 ;
      LAYER met3 ;
        RECT 1504.000 2771.680 1885.335 2785.240 ;
      LAYER met3 ;
        RECT 1889.070 2783.050 1889.370 2785.640 ;
        RECT 1892.505 2783.050 1892.835 2783.065 ;
        RECT 1889.070 2782.750 1892.835 2783.050 ;
        RECT 1892.505 2782.735 1892.835 2782.750 ;
        RECT 1500.000 2771.000 1504.000 2771.280 ;
        RECT 1499.910 2770.680 1504.000 2771.000 ;
        RECT 1489.545 2768.090 1489.875 2768.105 ;
        RECT 1499.910 2768.090 1500.210 2770.680 ;
      LAYER met3 ;
        RECT 1504.400 2770.320 1885.335 2771.680 ;
        RECT 1504.400 2770.280 1884.935 2770.320 ;
      LAYER met3 ;
        RECT 1489.545 2767.790 1500.210 2768.090 ;
      LAYER met3 ;
        RECT 1504.000 2768.920 1884.935 2770.280 ;
      LAYER met3 ;
        RECT 1885.335 2769.640 1889.335 2769.920 ;
        RECT 1885.335 2769.320 1889.370 2769.640 ;
        RECT 1489.545 2767.775 1489.875 2767.790 ;
        RECT 1000.000 2763.240 1004.000 2763.840 ;
        RECT 993.665 2760.610 993.995 2760.625 ;
        RECT 1000.350 2760.610 1000.650 2763.240 ;
      LAYER met3 ;
        RECT 1004.400 2762.840 1096.000 2764.240 ;
      LAYER met3 ;
        RECT 993.665 2760.310 1000.650 2760.610 ;
      LAYER met3 ;
        RECT 1004.000 2761.520 1096.000 2762.840 ;
      LAYER met3 ;
        RECT 993.665 2760.295 993.995 2760.310 ;
      LAYER met3 ;
        RECT 1004.000 2760.120 1095.600 2761.520 ;
      LAYER met3 ;
        RECT 1096.000 2760.800 1100.000 2761.120 ;
        RECT 1096.000 2760.610 1100.010 2760.800 ;
        RECT 1111.425 2760.610 1111.755 2760.625 ;
        RECT 1096.000 2760.520 1111.755 2760.610 ;
        RECT 1099.710 2760.310 1111.755 2760.520 ;
        RECT 1111.425 2760.295 1111.755 2760.310 ;
      LAYER met3 ;
        RECT 434.400 2751.960 574.800 2752.825 ;
        RECT 434.000 2734.320 574.800 2751.960 ;
        RECT 1004.000 2741.120 1096.000 2760.120 ;
        RECT 1504.000 2755.360 1885.335 2768.920 ;
      LAYER met3 ;
        RECT 1889.070 2767.410 1889.370 2769.320 ;
        RECT 1897.565 2767.410 1897.895 2767.425 ;
        RECT 1889.070 2767.110 1897.895 2767.410 ;
        RECT 1897.565 2767.095 1897.895 2767.110 ;
        RECT 1500.000 2754.680 1504.000 2754.960 ;
        RECT 1499.910 2754.360 1504.000 2754.680 ;
        RECT 1495.985 2753.810 1496.315 2753.825 ;
        RECT 1499.910 2753.810 1500.210 2754.360 ;
      LAYER met3 ;
        RECT 1504.400 2754.000 1885.335 2755.360 ;
        RECT 1504.400 2753.960 1884.935 2754.000 ;
      LAYER met3 ;
        RECT 1495.985 2753.510 1500.210 2753.810 ;
        RECT 1495.985 2753.495 1496.315 2753.510 ;
        RECT 1000.000 2740.120 1004.000 2740.720 ;
        RECT 992.745 2739.530 993.075 2739.545 ;
        RECT 1000.350 2739.530 1000.650 2740.120 ;
      LAYER met3 ;
        RECT 1004.400 2739.720 1096.000 2741.120 ;
        RECT 1504.000 2752.600 1884.935 2753.960 ;
      LAYER met3 ;
        RECT 1893.425 2753.810 1893.755 2753.825 ;
        RECT 1889.070 2753.600 1893.755 2753.810 ;
        RECT 1885.335 2753.510 1893.755 2753.600 ;
        RECT 1885.335 2753.320 1889.370 2753.510 ;
        RECT 1893.425 2753.495 1893.755 2753.510 ;
        RECT 1885.335 2753.000 1889.335 2753.320 ;
      LAYER met3 ;
        RECT 1504.000 2740.400 1885.335 2752.600 ;
      LAYER met3 ;
        RECT 1500.000 2739.720 1504.000 2740.000 ;
        RECT 992.745 2739.230 1000.650 2739.530 ;
        RECT 992.745 2739.215 993.075 2739.230 ;
      LAYER met3 ;
        RECT 1004.000 2738.400 1096.000 2739.720 ;
      LAYER met3 ;
        RECT 1487.245 2739.530 1487.575 2739.545 ;
        RECT 1499.910 2739.530 1504.000 2739.720 ;
        RECT 1487.245 2739.400 1504.000 2739.530 ;
        RECT 1487.245 2739.230 1500.210 2739.400 ;
        RECT 1487.245 2739.215 1487.575 2739.230 ;
      LAYER met3 ;
        RECT 1504.400 2739.040 1885.335 2740.400 ;
        RECT 1504.400 2739.000 1884.935 2739.040 ;
        RECT 1004.000 2737.000 1095.600 2738.400 ;
      LAYER met3 ;
        RECT 1096.000 2737.680 1100.000 2738.000 ;
        RECT 1096.000 2737.400 1100.010 2737.680 ;
      LAYER met3 ;
        RECT 434.000 2732.960 574.400 2734.320 ;
        RECT 434.400 2732.920 574.400 2732.960 ;
      LAYER met3 ;
        RECT 430.000 2732.240 434.000 2732.560 ;
        RECT 429.950 2731.960 434.000 2732.240 ;
        RECT 420.505 2729.330 420.835 2729.345 ;
        RECT 429.950 2729.330 430.250 2731.960 ;
      LAYER met3 ;
        RECT 434.400 2731.560 574.800 2732.920 ;
      LAYER met3 ;
        RECT 420.505 2729.030 430.250 2729.330 ;
        RECT 420.505 2729.015 420.835 2729.030 ;
      LAYER met3 ;
        RECT 434.000 2712.560 574.800 2731.560 ;
        RECT 1004.000 2719.360 1096.000 2737.000 ;
      LAYER met3 ;
        RECT 1099.710 2734.770 1100.010 2737.400 ;
      LAYER met3 ;
        RECT 1504.000 2737.640 1884.935 2739.000 ;
      LAYER met3 ;
        RECT 1885.335 2738.360 1889.335 2738.640 ;
        RECT 1885.335 2738.040 1889.370 2738.360 ;
        RECT 1111.885 2734.770 1112.215 2734.785 ;
        RECT 1099.710 2734.470 1112.215 2734.770 ;
        RECT 1111.885 2734.455 1112.215 2734.470 ;
      LAYER met3 ;
        RECT 1504.000 2724.080 1885.335 2737.640 ;
      LAYER met3 ;
        RECT 1889.070 2735.450 1889.370 2738.040 ;
        RECT 1894.345 2735.450 1894.675 2735.465 ;
        RECT 1889.070 2735.150 1894.675 2735.450 ;
        RECT 1894.345 2735.135 1894.675 2735.150 ;
        RECT 1500.000 2723.400 1504.000 2723.680 ;
        RECT 1499.910 2723.080 1504.000 2723.400 ;
        RECT 1486.785 2720.490 1487.115 2720.505 ;
        RECT 1499.910 2720.490 1500.210 2723.080 ;
      LAYER met3 ;
        RECT 1504.400 2722.720 1885.335 2724.080 ;
        RECT 1504.400 2722.680 1884.935 2722.720 ;
      LAYER met3 ;
        RECT 1486.785 2720.190 1500.210 2720.490 ;
      LAYER met3 ;
        RECT 1504.000 2721.320 1884.935 2722.680 ;
      LAYER met3 ;
        RECT 1885.335 2722.040 1889.335 2722.320 ;
        RECT 1885.335 2721.720 1889.370 2722.040 ;
        RECT 1486.785 2720.175 1487.115 2720.190 ;
        RECT 992.285 2719.130 992.615 2719.145 ;
        RECT 992.285 2718.960 1000.650 2719.130 ;
        RECT 992.285 2718.830 1004.000 2718.960 ;
        RECT 992.285 2718.815 992.615 2718.830 ;
        RECT 1000.000 2718.360 1004.000 2718.830 ;
      LAYER met3 ;
        RECT 1004.400 2717.960 1096.000 2719.360 ;
        RECT 1004.000 2716.640 1096.000 2717.960 ;
        RECT 1004.000 2715.240 1095.600 2716.640 ;
      LAYER met3 ;
        RECT 1096.000 2715.920 1100.000 2716.240 ;
        RECT 1096.000 2715.640 1100.010 2715.920 ;
      LAYER met3 ;
        RECT 434.000 2711.200 574.400 2712.560 ;
        RECT 434.400 2711.160 574.400 2711.200 ;
      LAYER met3 ;
        RECT 430.000 2710.480 434.000 2710.800 ;
        RECT 429.950 2710.200 434.000 2710.480 ;
        RECT 420.045 2707.570 420.375 2707.585 ;
        RECT 429.950 2707.570 430.250 2710.200 ;
      LAYER met3 ;
        RECT 434.400 2709.800 574.800 2711.160 ;
      LAYER met3 ;
        RECT 420.045 2707.270 430.250 2707.570 ;
        RECT 420.045 2707.255 420.375 2707.270 ;
      LAYER met3 ;
        RECT 434.000 2690.800 574.800 2709.800 ;
        RECT 1004.000 2696.240 1096.000 2715.240 ;
      LAYER met3 ;
        RECT 1099.710 2713.010 1100.010 2715.640 ;
        RECT 1112.345 2713.010 1112.675 2713.025 ;
        RECT 1099.710 2712.710 1112.675 2713.010 ;
        RECT 1112.345 2712.695 1112.675 2712.710 ;
      LAYER met3 ;
        RECT 1504.000 2709.120 1885.335 2721.320 ;
      LAYER met3 ;
        RECT 1889.070 2719.130 1889.370 2721.720 ;
        RECT 1892.965 2719.130 1893.295 2719.145 ;
        RECT 1889.070 2718.830 1893.295 2719.130 ;
        RECT 1892.965 2718.815 1893.295 2718.830 ;
      LAYER met3 ;
        RECT 1504.400 2707.760 1885.335 2709.120 ;
        RECT 1504.400 2707.720 1884.935 2707.760 ;
      LAYER met3 ;
        RECT 1000.000 2695.240 1004.000 2695.840 ;
        RECT 994.125 2692.610 994.455 2692.625 ;
        RECT 1000.350 2692.610 1000.650 2695.240 ;
      LAYER met3 ;
        RECT 1004.400 2694.840 1096.000 2696.240 ;
      LAYER met3 ;
        RECT 994.125 2692.310 1000.650 2692.610 ;
      LAYER met3 ;
        RECT 1004.000 2693.520 1096.000 2694.840 ;
        RECT 1504.000 2706.360 1884.935 2707.720 ;
      LAYER met3 ;
        RECT 994.125 2692.295 994.455 2692.310 ;
      LAYER met3 ;
        RECT 1004.000 2692.120 1095.600 2693.520 ;
      LAYER met3 ;
        RECT 1096.000 2692.800 1100.000 2693.120 ;
      LAYER met3 ;
        RECT 1504.000 2692.800 1885.335 2706.360 ;
      LAYER met3 ;
        RECT 1096.000 2692.520 1100.010 2692.800 ;
      LAYER met3 ;
        RECT 434.000 2689.440 574.400 2690.800 ;
      LAYER met3 ;
        RECT 574.800 2689.800 578.800 2690.400 ;
      LAYER met3 ;
        RECT 434.400 2689.400 574.400 2689.440 ;
        RECT 434.400 2688.040 574.800 2689.400 ;
        RECT 434.000 2670.400 574.800 2688.040 ;
      LAYER met3 ;
        RECT 578.070 2687.170 578.370 2689.800 ;
        RECT 588.865 2687.170 589.195 2687.185 ;
        RECT 578.070 2686.870 589.195 2687.170 ;
        RECT 588.865 2686.855 589.195 2686.870 ;
      LAYER met3 ;
        RECT 1004.000 2673.120 1096.000 2692.120 ;
      LAYER met3 ;
        RECT 1099.710 2691.930 1100.010 2692.520 ;
        RECT 1500.000 2692.120 1504.000 2692.400 ;
        RECT 1112.805 2691.930 1113.135 2691.945 ;
        RECT 1099.710 2691.630 1113.135 2691.930 ;
        RECT 1112.805 2691.615 1113.135 2691.630 ;
        RECT 1489.085 2691.930 1489.415 2691.945 ;
        RECT 1499.910 2691.930 1504.000 2692.120 ;
        RECT 1489.085 2691.800 1504.000 2691.930 ;
        RECT 1489.085 2691.630 1500.210 2691.800 ;
        RECT 1489.085 2691.615 1489.415 2691.630 ;
      LAYER met3 ;
        RECT 1504.400 2691.440 1885.335 2692.800 ;
        RECT 1504.400 2691.400 1884.935 2691.440 ;
        RECT 1504.000 2690.040 1884.935 2691.400 ;
      LAYER met3 ;
        RECT 1885.335 2690.760 1889.335 2691.040 ;
        RECT 1885.335 2690.440 1889.370 2690.760 ;
      LAYER met3 ;
        RECT 1504.000 2677.840 1885.335 2690.040 ;
      LAYER met3 ;
        RECT 1889.070 2687.850 1889.370 2690.440 ;
        RECT 1898.025 2687.850 1898.355 2687.865 ;
        RECT 1889.070 2687.550 1898.355 2687.850 ;
        RECT 1898.025 2687.535 1898.355 2687.550 ;
        RECT 1500.000 2677.160 1504.000 2677.440 ;
        RECT 1499.910 2676.840 1504.000 2677.160 ;
        RECT 1489.085 2674.250 1489.415 2674.265 ;
        RECT 1499.910 2674.250 1500.210 2676.840 ;
      LAYER met3 ;
        RECT 1504.400 2676.480 1885.335 2677.840 ;
        RECT 1504.400 2676.440 1884.935 2676.480 ;
      LAYER met3 ;
        RECT 1489.085 2673.950 1500.210 2674.250 ;
      LAYER met3 ;
        RECT 1504.000 2675.080 1884.935 2676.440 ;
      LAYER met3 ;
        RECT 1885.335 2675.800 1889.335 2676.080 ;
        RECT 1885.335 2675.480 1889.370 2675.800 ;
        RECT 1489.085 2673.935 1489.415 2673.950 ;
        RECT 1000.000 2672.120 1004.000 2672.720 ;
        RECT 994.585 2670.850 994.915 2670.865 ;
        RECT 1000.350 2670.850 1000.650 2672.120 ;
      LAYER met3 ;
        RECT 1004.400 2671.720 1096.000 2673.120 ;
      LAYER met3 ;
        RECT 994.585 2670.550 1000.650 2670.850 ;
        RECT 994.585 2670.535 994.915 2670.550 ;
      LAYER met3 ;
        RECT 1004.000 2670.400 1096.000 2671.720 ;
        RECT 434.000 2669.040 574.400 2670.400 ;
      LAYER met3 ;
        RECT 574.800 2669.400 578.800 2670.000 ;
      LAYER met3 ;
        RECT 434.400 2669.000 574.400 2669.040 ;
        RECT 434.400 2667.640 574.800 2669.000 ;
        RECT 434.000 2648.640 574.800 2667.640 ;
      LAYER met3 ;
        RECT 578.070 2666.770 578.370 2669.400 ;
      LAYER met3 ;
        RECT 1004.000 2669.000 1095.600 2670.400 ;
      LAYER met3 ;
        RECT 1096.000 2669.680 1100.000 2670.000 ;
        RECT 1096.000 2669.400 1100.010 2669.680 ;
        RECT 588.865 2666.770 589.195 2666.785 ;
        RECT 578.070 2666.470 589.195 2666.770 ;
        RECT 588.865 2666.455 589.195 2666.470 ;
      LAYER met3 ;
        RECT 1004.000 2650.000 1096.000 2669.000 ;
      LAYER met3 ;
        RECT 1099.710 2666.770 1100.010 2669.400 ;
        RECT 1113.265 2666.770 1113.595 2666.785 ;
        RECT 1099.710 2666.470 1113.595 2666.770 ;
        RECT 1113.265 2666.455 1113.595 2666.470 ;
      LAYER met3 ;
        RECT 1504.000 2661.520 1885.335 2675.080 ;
      LAYER met3 ;
        RECT 1889.070 2672.890 1889.370 2675.480 ;
        RECT 1898.485 2672.890 1898.815 2672.905 ;
        RECT 1889.070 2672.590 1898.815 2672.890 ;
        RECT 1898.485 2672.575 1898.815 2672.590 ;
        RECT 1500.000 2660.840 1504.000 2661.120 ;
        RECT 1499.910 2660.520 1504.000 2660.840 ;
        RECT 1482.645 2657.250 1482.975 2657.265 ;
        RECT 1499.910 2657.250 1500.210 2660.520 ;
      LAYER met3 ;
        RECT 1504.400 2660.160 1885.335 2661.520 ;
        RECT 1504.400 2660.120 1884.935 2660.160 ;
      LAYER met3 ;
        RECT 1482.645 2656.950 1500.210 2657.250 ;
      LAYER met3 ;
        RECT 1504.000 2658.760 1884.935 2660.120 ;
      LAYER met3 ;
        RECT 1885.335 2659.480 1889.335 2659.760 ;
        RECT 1885.335 2659.160 1889.370 2659.480 ;
        RECT 1482.645 2656.935 1482.975 2656.950 ;
        RECT 1000.000 2649.000 1004.000 2649.600 ;
      LAYER met3 ;
        RECT 434.000 2647.280 574.400 2648.640 ;
        RECT 434.400 2647.240 574.400 2647.280 ;
        RECT 434.400 2645.880 574.800 2647.240 ;
      LAYER met3 ;
        RECT 987.225 2646.370 987.555 2646.385 ;
        RECT 1000.350 2646.370 1000.650 2649.000 ;
      LAYER met3 ;
        RECT 1004.400 2648.600 1096.000 2650.000 ;
      LAYER met3 ;
        RECT 987.225 2646.070 1000.650 2646.370 ;
      LAYER met3 ;
        RECT 1004.000 2647.280 1096.000 2648.600 ;
      LAYER met3 ;
        RECT 987.225 2646.055 987.555 2646.070 ;
      LAYER met3 ;
        RECT 434.000 2626.880 574.800 2645.880 ;
        RECT 1004.000 2645.880 1095.600 2647.280 ;
      LAYER met3 ;
        RECT 1096.000 2646.280 1100.000 2646.880 ;
      LAYER met3 ;
        RECT 1504.000 2646.560 1885.335 2658.760 ;
      LAYER met3 ;
        RECT 1889.070 2657.250 1889.370 2659.160 ;
        RECT 1898.945 2657.250 1899.275 2657.265 ;
        RECT 1889.070 2656.950 1899.275 2657.250 ;
        RECT 1898.945 2656.935 1899.275 2656.950 ;
      LAYER met3 ;
        RECT 1004.000 2626.880 1096.000 2645.880 ;
      LAYER met3 ;
        RECT 1096.950 2645.025 1097.250 2646.280 ;
      LAYER met3 ;
        RECT 1504.400 2645.200 1885.335 2646.560 ;
        RECT 1504.400 2645.160 1884.935 2645.200 ;
      LAYER met3 ;
        RECT 1096.950 2644.710 1097.495 2645.025 ;
        RECT 1097.165 2644.695 1097.495 2644.710 ;
      LAYER met3 ;
        RECT 1504.000 2643.800 1884.935 2645.160 ;
        RECT 1504.000 2630.240 1885.335 2643.800 ;
      LAYER met3 ;
        RECT 1500.000 2629.560 1504.000 2629.840 ;
        RECT 1488.165 2629.370 1488.495 2629.385 ;
        RECT 1499.910 2629.370 1504.000 2629.560 ;
        RECT 1488.165 2629.240 1504.000 2629.370 ;
        RECT 1488.165 2629.070 1500.210 2629.240 ;
        RECT 1488.165 2629.055 1488.495 2629.070 ;
      LAYER met3 ;
        RECT 1504.400 2628.880 1885.335 2630.240 ;
        RECT 1504.400 2628.840 1884.935 2628.880 ;
        RECT 434.000 2625.520 574.400 2626.880 ;
      LAYER met3 ;
        RECT 1000.000 2625.880 1004.000 2626.480 ;
      LAYER met3 ;
        RECT 434.400 2625.480 574.400 2625.520 ;
        RECT 434.400 2624.120 574.800 2625.480 ;
        RECT 434.000 2606.480 574.800 2624.120 ;
      LAYER met3 ;
        RECT 991.825 2623.250 992.155 2623.265 ;
        RECT 1000.350 2623.250 1000.650 2625.880 ;
      LAYER met3 ;
        RECT 1004.400 2625.480 1096.000 2626.880 ;
      LAYER met3 ;
        RECT 991.825 2622.950 1000.650 2623.250 ;
      LAYER met3 ;
        RECT 1004.000 2624.160 1096.000 2625.480 ;
        RECT 1504.000 2627.480 1884.935 2628.840 ;
      LAYER met3 ;
        RECT 1885.335 2628.200 1889.335 2628.480 ;
        RECT 1885.335 2627.880 1889.370 2628.200 ;
        RECT 991.825 2622.935 992.155 2622.950 ;
      LAYER met3 ;
        RECT 1004.000 2622.760 1095.600 2624.160 ;
      LAYER met3 ;
        RECT 1096.000 2623.160 1100.000 2623.760 ;
      LAYER met3 ;
        RECT 1004.000 2610.715 1096.000 2622.760 ;
      LAYER met3 ;
        RECT 1097.870 2622.585 1098.170 2623.160 ;
        RECT 1097.625 2622.270 1098.170 2622.585 ;
        RECT 1097.625 2622.255 1097.955 2622.270 ;
      LAYER met3 ;
        RECT 1504.000 2613.920 1885.335 2627.480 ;
      LAYER met3 ;
        RECT 1889.070 2625.290 1889.370 2627.880 ;
        RECT 1899.405 2625.290 1899.735 2625.305 ;
        RECT 1889.070 2624.990 1899.735 2625.290 ;
        RECT 1899.405 2624.975 1899.735 2624.990 ;
        RECT 1500.000 2613.240 1504.000 2613.520 ;
        RECT 1499.910 2612.920 1504.000 2613.240 ;
        RECT 1488.625 2610.330 1488.955 2610.345 ;
        RECT 1499.910 2610.330 1500.210 2612.920 ;
      LAYER met3 ;
        RECT 1504.400 2612.560 1885.335 2613.920 ;
        RECT 1504.400 2612.520 1884.935 2612.560 ;
      LAYER met3 ;
        RECT 1488.625 2610.030 1500.210 2610.330 ;
      LAYER met3 ;
        RECT 1504.000 2611.160 1884.935 2612.520 ;
      LAYER met3 ;
        RECT 1885.335 2611.880 1889.335 2612.160 ;
        RECT 1885.335 2611.560 1889.370 2611.880 ;
        RECT 1488.625 2610.015 1488.955 2610.030 ;
      LAYER met3 ;
        RECT 434.000 2605.080 574.400 2606.480 ;
        RECT 434.000 2604.255 574.800 2605.080 ;
      LAYER met3 ;
        RECT 1350.165 2601.490 1350.495 2601.505 ;
        RECT 1351.085 2601.490 1351.415 2601.505 ;
        RECT 1350.165 2601.190 1351.415 2601.490 ;
        RECT 1350.165 2601.175 1350.495 2601.190 ;
        RECT 1351.085 2601.175 1351.415 2601.190 ;
      LAYER met3 ;
        RECT 1504.000 2598.960 1885.335 2611.160 ;
      LAYER met3 ;
        RECT 1889.070 2608.970 1889.370 2611.560 ;
      LAYER met3 ;
        RECT 2427.190 2610.715 2529.990 2760.645 ;
      LAYER met3 ;
        RECT 1899.865 2608.970 1900.195 2608.985 ;
        RECT 1889.070 2608.670 1900.195 2608.970 ;
        RECT 1899.865 2608.655 1900.195 2608.670 ;
        RECT 1500.000 2598.280 1504.000 2598.560 ;
        RECT 1499.910 2597.960 1504.000 2598.280 ;
        RECT 1488.165 2595.370 1488.495 2595.385 ;
        RECT 1499.910 2595.370 1500.210 2597.960 ;
      LAYER met3 ;
        RECT 1504.400 2597.600 1885.335 2598.960 ;
        RECT 1504.400 2597.560 1884.935 2597.600 ;
      LAYER met3 ;
        RECT 1488.165 2595.070 1500.210 2595.370 ;
      LAYER met3 ;
        RECT 1504.000 2596.200 1884.935 2597.560 ;
      LAYER met3 ;
        RECT 1488.165 2595.055 1488.495 2595.070 ;
      LAYER met3 ;
        RECT 1504.000 2582.640 1885.335 2596.200 ;
      LAYER met3 ;
        RECT 1500.000 2581.960 1504.000 2582.240 ;
        RECT 1499.910 2581.640 1504.000 2581.960 ;
        RECT 1488.165 2581.090 1488.495 2581.105 ;
        RECT 1499.910 2581.090 1500.210 2581.640 ;
      LAYER met3 ;
        RECT 1504.400 2581.280 1885.335 2582.640 ;
        RECT 1504.400 2581.240 1884.935 2581.280 ;
      LAYER met3 ;
        RECT 1488.165 2580.790 1500.210 2581.090 ;
        RECT 1488.165 2580.775 1488.495 2580.790 ;
      LAYER met3 ;
        RECT 1504.000 2579.880 1884.935 2581.240 ;
      LAYER met3 ;
        RECT 1885.335 2580.600 1889.335 2580.880 ;
        RECT 1885.335 2580.280 1889.370 2580.600 ;
      LAYER met3 ;
        RECT 1504.000 2567.680 1885.335 2579.880 ;
      LAYER met3 ;
        RECT 1889.070 2577.690 1889.370 2580.280 ;
        RECT 1900.325 2577.690 1900.655 2577.705 ;
        RECT 1889.070 2577.390 1900.655 2577.690 ;
        RECT 1900.325 2577.375 1900.655 2577.390 ;
        RECT 1488.165 2567.490 1488.495 2567.505 ;
        RECT 1488.165 2567.280 1500.210 2567.490 ;
        RECT 1488.165 2567.190 1504.000 2567.280 ;
        RECT 1488.165 2567.175 1488.495 2567.190 ;
        RECT 1499.910 2567.000 1504.000 2567.190 ;
        RECT 1500.000 2566.680 1504.000 2567.000 ;
      LAYER met3 ;
        RECT 1504.400 2566.320 1885.335 2567.680 ;
        RECT 1504.400 2566.280 1884.935 2566.320 ;
        RECT 1504.000 2564.920 1884.935 2566.280 ;
      LAYER met3 ;
        RECT 1885.335 2565.640 1889.335 2565.920 ;
        RECT 1885.335 2565.320 1889.370 2565.640 ;
        RECT 1351.545 2560.010 1351.875 2560.025 ;
        RECT 1351.545 2559.695 1352.090 2560.010 ;
        RECT 1350.165 2559.330 1350.495 2559.345 ;
        RECT 1351.790 2559.330 1352.090 2559.695 ;
        RECT 1350.165 2559.030 1352.090 2559.330 ;
        RECT 1350.165 2559.015 1350.495 2559.030 ;
      LAYER met3 ;
        RECT 1504.000 2551.360 1885.335 2564.920 ;
      LAYER met3 ;
        RECT 1889.070 2562.730 1889.370 2565.320 ;
        RECT 1900.785 2562.730 1901.115 2562.745 ;
        RECT 1889.070 2562.430 1901.115 2562.730 ;
        RECT 1900.785 2562.415 1901.115 2562.430 ;
        RECT 1500.000 2550.680 1504.000 2550.960 ;
        RECT 1499.910 2550.360 1504.000 2550.680 ;
        RECT 1484.485 2549.130 1484.815 2549.145 ;
        RECT 1499.910 2549.130 1500.210 2550.360 ;
      LAYER met3 ;
        RECT 1504.400 2550.000 1885.335 2551.360 ;
        RECT 1504.400 2549.960 1884.935 2550.000 ;
      LAYER met3 ;
        RECT 1484.485 2548.830 1500.210 2549.130 ;
        RECT 1484.485 2548.815 1484.815 2548.830 ;
      LAYER met3 ;
        RECT 1504.000 2548.600 1884.935 2549.960 ;
      LAYER met3 ;
        RECT 1885.335 2549.320 1889.335 2549.600 ;
        RECT 1885.335 2549.000 1889.370 2549.320 ;
      LAYER met3 ;
        RECT 1504.000 2536.400 1885.335 2548.600 ;
      LAYER met3 ;
        RECT 1889.070 2547.770 1889.370 2549.000 ;
        RECT 1901.245 2547.770 1901.575 2547.785 ;
        RECT 1889.070 2547.470 1901.575 2547.770 ;
        RECT 1901.245 2547.455 1901.575 2547.470 ;
      LAYER met3 ;
        RECT 1504.400 2535.040 1885.335 2536.400 ;
        RECT 1504.400 2535.000 1884.935 2535.040 ;
        RECT 1504.000 2533.640 1884.935 2535.000 ;
        RECT 1504.000 2520.080 1885.335 2533.640 ;
      LAYER met3 ;
        RECT 1500.000 2519.400 1504.000 2519.680 ;
        RECT 1487.705 2519.210 1488.035 2519.225 ;
        RECT 1499.910 2519.210 1504.000 2519.400 ;
        RECT 1487.705 2519.080 1504.000 2519.210 ;
        RECT 1487.705 2518.910 1500.210 2519.080 ;
        RECT 1487.705 2518.895 1488.035 2518.910 ;
      LAYER met3 ;
        RECT 1504.400 2518.720 1885.335 2520.080 ;
        RECT 1504.400 2518.680 1884.935 2518.720 ;
        RECT 1504.000 2517.320 1884.935 2518.680 ;
      LAYER met3 ;
        RECT 1885.335 2518.040 1889.335 2518.320 ;
        RECT 1885.335 2517.720 1889.370 2518.040 ;
      LAYER met3 ;
        RECT 1504.000 2510.715 1885.335 2517.320 ;
      LAYER met3 ;
        RECT 1889.070 2515.130 1889.370 2517.720 ;
        RECT 1903.545 2515.130 1903.875 2515.145 ;
        RECT 1889.070 2514.830 1903.875 2515.130 ;
        RECT 1903.545 2514.815 1903.875 2514.830 ;
        RECT 1351.085 2463.450 1351.415 2463.465 ;
        RECT 1352.005 2463.450 1352.335 2463.465 ;
        RECT 1351.085 2463.150 1352.335 2463.450 ;
        RECT 1351.085 2463.135 1351.415 2463.150 ;
        RECT 1352.005 2463.135 1352.335 2463.150 ;
        RECT 1514.845 2463.450 1515.175 2463.465 ;
        RECT 1532.325 2463.450 1532.655 2463.465 ;
        RECT 1514.845 2463.150 1532.655 2463.450 ;
        RECT 1514.845 2463.135 1515.175 2463.150 ;
        RECT 1532.325 2463.135 1532.655 2463.150 ;
        RECT 1559.465 2319.290 1559.795 2319.305 ;
        RECT 1558.790 2318.990 1559.795 2319.290 ;
        RECT 1558.790 2318.610 1559.090 2318.990 ;
        RECT 1559.465 2318.975 1559.795 2318.990 ;
        RECT 1573.725 2319.290 1574.055 2319.305 ;
        RECT 1573.725 2318.990 1574.730 2319.290 ;
        RECT 1573.725 2318.975 1574.055 2318.990 ;
        RECT 1559.465 2318.610 1559.795 2318.625 ;
        RECT 1558.790 2318.310 1559.795 2318.610 ;
        RECT 1559.465 2318.295 1559.795 2318.310 ;
        RECT 1573.725 2318.610 1574.055 2318.625 ;
        RECT 1574.430 2318.610 1574.730 2318.990 ;
        RECT 1573.725 2318.310 1574.730 2318.610 ;
        RECT 1573.725 2318.295 1574.055 2318.310 ;
        RECT 1350.165 2270.330 1350.495 2270.345 ;
        RECT 1351.085 2270.330 1351.415 2270.345 ;
        RECT 1350.165 2270.030 1351.415 2270.330 ;
        RECT 1350.165 2270.015 1350.495 2270.030 ;
        RECT 1351.085 2270.015 1351.415 2270.030 ;
        RECT 1532.325 2270.330 1532.655 2270.345 ;
        RECT 1533.245 2270.330 1533.575 2270.345 ;
        RECT 1532.325 2270.030 1533.575 2270.330 ;
        RECT 1532.325 2270.015 1532.655 2270.030 ;
        RECT 1533.245 2270.015 1533.575 2270.030 ;
        RECT 1350.165 2173.770 1350.495 2173.785 ;
        RECT 1351.085 2173.770 1351.415 2173.785 ;
        RECT 1350.165 2173.470 1351.415 2173.770 ;
        RECT 1350.165 2173.455 1350.495 2173.470 ;
        RECT 1351.085 2173.455 1351.415 2173.470 ;
        RECT 1532.325 2062.940 1532.655 2062.945 ;
        RECT 1532.070 2062.930 1532.655 2062.940 ;
        RECT 1532.070 2062.630 1532.880 2062.930 ;
        RECT 1532.070 2062.620 1532.655 2062.630 ;
        RECT 1532.325 2062.615 1532.655 2062.620 ;
      LAYER met3 ;
        RECT 1004.000 2019.280 1329.390 2032.005 ;
      LAYER met3 ;
        RECT 1532.070 2028.250 1532.450 2028.260 ;
        RECT 1532.785 2028.250 1533.115 2028.265 ;
        RECT 1532.070 2027.950 1533.115 2028.250 ;
        RECT 1532.070 2027.940 1532.450 2027.950 ;
        RECT 1532.785 2027.935 1533.115 2027.950 ;
        RECT 995.045 2018.730 995.375 2018.745 ;
        RECT 1000.000 2018.730 1004.000 2018.880 ;
        RECT 995.045 2018.430 1004.000 2018.730 ;
        RECT 995.045 2018.415 995.375 2018.430 ;
        RECT 1000.000 2018.280 1004.000 2018.430 ;
      LAYER met3 ;
        RECT 1004.400 2017.880 1328.990 2019.280 ;
      LAYER met3 ;
        RECT 1329.390 2018.730 1333.390 2018.880 ;
        RECT 1338.665 2018.730 1338.995 2018.745 ;
        RECT 1329.390 2018.430 1338.995 2018.730 ;
        RECT 1329.390 2018.280 1333.390 2018.430 ;
        RECT 1338.665 2018.415 1338.995 2018.430 ;
      LAYER met3 ;
        RECT 1004.000 1998.880 1329.390 2017.880 ;
      LAYER met3 ;
        RECT 995.505 1998.330 995.835 1998.345 ;
        RECT 1000.000 1998.330 1004.000 1998.480 ;
        RECT 995.505 1998.030 1004.000 1998.330 ;
        RECT 995.505 1998.015 995.835 1998.030 ;
        RECT 1000.000 1997.880 1004.000 1998.030 ;
      LAYER met3 ;
        RECT 1004.400 1997.480 1328.990 1998.880 ;
      LAYER met3 ;
        RECT 1329.390 1998.330 1333.390 1998.480 ;
        RECT 1334.065 1998.330 1334.395 1998.345 ;
        RECT 1329.390 1998.030 1334.395 1998.330 ;
        RECT 1329.390 1997.880 1333.390 1998.030 ;
        RECT 1334.065 1998.015 1334.395 1998.030 ;
      LAYER met3 ;
        RECT 1004.000 1977.120 1329.390 1997.480 ;
      LAYER met3 ;
        RECT 995.965 1976.570 996.295 1976.585 ;
        RECT 1000.000 1976.570 1004.000 1976.720 ;
        RECT 995.965 1976.270 1004.000 1976.570 ;
        RECT 995.965 1976.255 996.295 1976.270 ;
        RECT 1000.000 1976.120 1004.000 1976.270 ;
      LAYER met3 ;
        RECT 1004.400 1975.720 1328.990 1977.120 ;
      LAYER met3 ;
        RECT 1329.390 1976.570 1333.390 1976.720 ;
        RECT 1339.125 1976.570 1339.455 1976.585 ;
        RECT 1329.390 1976.270 1339.455 1976.570 ;
        RECT 1329.390 1976.120 1333.390 1976.270 ;
        RECT 1339.125 1976.255 1339.455 1976.270 ;
      LAYER met3 ;
        RECT 364.000 1963.520 627.030 1969.445 ;
        RECT 364.400 1962.120 627.030 1963.520 ;
        RECT 364.000 1940.400 627.030 1962.120 ;
        RECT 1004.000 1956.720 1329.390 1975.720 ;
      LAYER met3 ;
        RECT 991.365 1956.170 991.695 1956.185 ;
        RECT 1000.000 1956.170 1004.000 1956.320 ;
        RECT 991.365 1955.870 1004.000 1956.170 ;
        RECT 991.365 1955.855 991.695 1955.870 ;
        RECT 1000.000 1955.720 1004.000 1955.870 ;
      LAYER met3 ;
        RECT 1004.400 1955.320 1328.990 1956.720 ;
      LAYER met3 ;
        RECT 1329.390 1956.170 1333.390 1956.320 ;
        RECT 1339.585 1956.170 1339.915 1956.185 ;
        RECT 1329.390 1955.870 1339.915 1956.170 ;
        RECT 1329.390 1955.720 1333.390 1955.870 ;
        RECT 1339.585 1955.855 1339.915 1955.870 ;
      LAYER met3 ;
        RECT 364.000 1939.000 626.630 1940.400 ;
        RECT 364.000 1926.800 627.030 1939.000 ;
        RECT 1004.000 1936.320 1329.390 1955.320 ;
      LAYER met3 ;
        RECT 990.905 1935.770 991.235 1935.785 ;
        RECT 1000.000 1935.770 1004.000 1935.920 ;
        RECT 990.905 1935.470 1004.000 1935.770 ;
        RECT 990.905 1935.455 991.235 1935.470 ;
        RECT 1000.000 1935.320 1004.000 1935.470 ;
      LAYER met3 ;
        RECT 1004.400 1934.960 1329.390 1936.320 ;
        RECT 1004.400 1934.920 1328.990 1934.960 ;
        RECT 364.400 1925.400 627.030 1926.800 ;
        RECT 364.000 1903.680 627.030 1925.400 ;
        RECT 1004.000 1933.560 1328.990 1934.920 ;
      LAYER met3 ;
        RECT 1329.390 1934.410 1333.390 1934.560 ;
        RECT 1340.045 1934.410 1340.375 1934.425 ;
        RECT 1329.390 1934.110 1340.375 1934.410 ;
        RECT 1329.390 1933.960 1333.390 1934.110 ;
        RECT 1340.045 1934.095 1340.375 1934.110 ;
      LAYER met3 ;
        RECT 1004.000 1914.560 1329.390 1933.560 ;
      LAYER met3 ;
        RECT 996.425 1914.010 996.755 1914.025 ;
        RECT 1000.000 1914.010 1004.000 1914.160 ;
        RECT 996.425 1913.710 1004.000 1914.010 ;
        RECT 996.425 1913.695 996.755 1913.710 ;
        RECT 1000.000 1913.560 1004.000 1913.710 ;
      LAYER met3 ;
        RECT 1004.400 1913.160 1328.990 1914.560 ;
      LAYER met3 ;
        RECT 1329.390 1914.010 1333.390 1914.160 ;
        RECT 1340.505 1914.010 1340.835 1914.025 ;
        RECT 1329.390 1913.710 1340.835 1914.010 ;
        RECT 1329.390 1913.560 1333.390 1913.710 ;
        RECT 1340.505 1913.695 1340.835 1913.710 ;
      LAYER met3 ;
        RECT 364.000 1902.280 626.630 1903.680 ;
        RECT 364.000 1890.080 627.030 1902.280 ;
        RECT 1004.000 1894.160 1329.390 1913.160 ;
        RECT 1924.400 1906.040 2072.375 1906.905 ;
      LAYER met3 ;
        RECT 990.445 1893.610 990.775 1893.625 ;
        RECT 1000.000 1893.610 1004.000 1893.760 ;
        RECT 990.445 1893.310 1004.000 1893.610 ;
        RECT 990.445 1893.295 990.775 1893.310 ;
        RECT 1000.000 1893.160 1004.000 1893.310 ;
      LAYER met3 ;
        RECT 1004.400 1892.800 1329.390 1894.160 ;
        RECT 1924.000 1904.720 2072.375 1906.040 ;
        RECT 1924.000 1903.320 2071.975 1904.720 ;
        RECT 1004.400 1892.760 1328.990 1892.800 ;
        RECT 364.400 1888.680 627.030 1890.080 ;
        RECT 364.000 1866.960 627.030 1888.680 ;
        RECT 1004.000 1891.400 1328.990 1892.760 ;
      LAYER met3 ;
        RECT 1329.390 1892.250 1333.390 1892.400 ;
        RECT 1340.965 1892.250 1341.295 1892.265 ;
        RECT 1329.390 1891.950 1341.295 1892.250 ;
        RECT 1329.390 1891.800 1333.390 1891.950 ;
        RECT 1340.965 1891.935 1341.295 1891.950 ;
      LAYER met3 ;
        RECT 1004.000 1872.400 1329.390 1891.400 ;
        RECT 1924.000 1889.760 2072.375 1903.320 ;
      LAYER met3 ;
        RECT 1920.000 1888.760 1924.000 1889.360 ;
        RECT 1904.465 1886.130 1904.795 1886.145 ;
        RECT 1920.350 1886.130 1920.650 1888.760 ;
      LAYER met3 ;
        RECT 1924.400 1888.400 2072.375 1889.760 ;
        RECT 2304.000 1892.800 2524.550 1925.925 ;
        RECT 2304.000 1891.400 2524.150 1892.800 ;
      LAYER met3 ;
        RECT 2524.550 1892.250 2528.550 1892.400 ;
        RECT 2539.265 1892.250 2539.595 1892.265 ;
        RECT 2524.550 1891.950 2539.595 1892.250 ;
        RECT 2524.550 1891.800 2528.550 1891.950 ;
        RECT 2539.265 1891.935 2539.595 1891.950 ;
      LAYER met3 ;
        RECT 1924.400 1888.360 2071.975 1888.400 ;
      LAYER met3 ;
        RECT 1904.465 1885.830 1920.650 1886.130 ;
      LAYER met3 ;
        RECT 1924.000 1887.000 2071.975 1888.360 ;
      LAYER met3 ;
        RECT 2072.375 1887.400 2076.375 1888.000 ;
        RECT 1904.465 1885.815 1904.795 1885.830 ;
        RECT 1352.005 1884.090 1352.335 1884.105 ;
        RECT 1351.790 1883.775 1352.335 1884.090 ;
        RECT 1350.165 1882.730 1350.495 1882.745 ;
        RECT 1351.790 1882.730 1352.090 1883.775 ;
        RECT 1350.165 1882.430 1352.090 1882.730 ;
        RECT 1350.165 1882.415 1350.495 1882.430 ;
      LAYER met3 ;
        RECT 1924.000 1873.440 2072.375 1887.000 ;
      LAYER met3 ;
        RECT 2075.830 1884.770 2076.130 1887.400 ;
        RECT 2087.085 1884.770 2087.415 1884.785 ;
        RECT 2075.830 1884.470 2087.415 1884.770 ;
        RECT 2087.085 1884.455 2087.415 1884.470 ;
      LAYER met3 ;
        RECT 2304.000 1877.840 2524.550 1891.400 ;
      LAYER met3 ;
        RECT 2287.185 1877.290 2287.515 1877.305 ;
        RECT 2300.000 1877.290 2304.000 1877.440 ;
        RECT 2287.185 1876.990 2304.000 1877.290 ;
        RECT 2287.185 1876.975 2287.515 1876.990 ;
        RECT 2300.000 1876.840 2304.000 1876.990 ;
      LAYER met3 ;
        RECT 2304.400 1876.440 2524.550 1877.840 ;
      LAYER met3 ;
        RECT 1920.000 1872.440 1924.000 1873.040 ;
        RECT 989.985 1871.850 990.315 1871.865 ;
        RECT 1000.000 1871.850 1004.000 1872.000 ;
        RECT 989.985 1871.550 1004.000 1871.850 ;
        RECT 989.985 1871.535 990.315 1871.550 ;
        RECT 1000.000 1871.400 1004.000 1871.550 ;
      LAYER met3 ;
        RECT 1004.400 1871.000 1328.990 1872.400 ;
      LAYER met3 ;
        RECT 1329.390 1871.850 1333.390 1872.000 ;
        RECT 1341.425 1871.850 1341.755 1871.865 ;
        RECT 1329.390 1871.550 1341.755 1871.850 ;
        RECT 1329.390 1871.400 1333.390 1871.550 ;
        RECT 1341.425 1871.535 1341.755 1871.550 ;
      LAYER met3 ;
        RECT 364.000 1865.560 626.630 1866.960 ;
        RECT 364.000 1852.000 627.030 1865.560 ;
        RECT 1004.000 1852.000 1329.390 1871.000 ;
      LAYER met3 ;
        RECT 1904.465 1870.490 1904.795 1870.505 ;
        RECT 1920.350 1870.490 1920.650 1872.440 ;
      LAYER met3 ;
        RECT 1924.400 1872.040 2072.375 1873.440 ;
      LAYER met3 ;
        RECT 1904.465 1870.190 1920.650 1870.490 ;
      LAYER met3 ;
        RECT 1924.000 1870.720 2072.375 1872.040 ;
      LAYER met3 ;
        RECT 1904.465 1870.175 1904.795 1870.190 ;
      LAYER met3 ;
        RECT 1924.000 1869.320 2071.975 1870.720 ;
        RECT 1924.000 1855.760 2072.375 1869.320 ;
      LAYER met3 ;
        RECT 1920.000 1854.760 1924.000 1855.360 ;
      LAYER met3 ;
        RECT 364.400 1850.600 627.030 1852.000 ;
      LAYER met3 ;
        RECT 989.525 1851.450 989.855 1851.465 ;
        RECT 1000.000 1851.450 1004.000 1851.600 ;
        RECT 989.525 1851.150 1004.000 1851.450 ;
        RECT 989.525 1851.135 989.855 1851.150 ;
        RECT 1000.000 1851.000 1004.000 1851.150 ;
      LAYER met3 ;
        RECT 1004.400 1850.640 1329.390 1852.000 ;
      LAYER met3 ;
        RECT 1904.465 1852.130 1904.795 1852.145 ;
        RECT 1920.350 1852.130 1920.650 1854.760 ;
      LAYER met3 ;
        RECT 1924.400 1854.400 2072.375 1855.760 ;
        RECT 1924.400 1854.360 2071.975 1854.400 ;
      LAYER met3 ;
        RECT 1904.465 1851.830 1920.650 1852.130 ;
      LAYER met3 ;
        RECT 1924.000 1853.000 2071.975 1854.360 ;
      LAYER met3 ;
        RECT 2072.375 1853.400 2076.375 1854.000 ;
        RECT 1904.465 1851.815 1904.795 1851.830 ;
      LAYER met3 ;
        RECT 1004.400 1850.600 1328.990 1850.640 ;
        RECT 364.000 1830.240 627.030 1850.600 ;
        RECT 1004.000 1849.240 1328.990 1850.600 ;
      LAYER met3 ;
        RECT 1329.390 1850.090 1333.390 1850.240 ;
        RECT 1341.885 1850.090 1342.215 1850.105 ;
        RECT 1329.390 1849.790 1342.215 1850.090 ;
        RECT 1329.390 1849.640 1333.390 1849.790 ;
        RECT 1341.885 1849.775 1342.215 1849.790 ;
      LAYER met3 ;
        RECT 1004.000 1830.240 1329.390 1849.240 ;
        RECT 1924.000 1839.440 2072.375 1853.000 ;
      LAYER met3 ;
        RECT 2075.830 1850.770 2076.130 1853.400 ;
        RECT 2084.325 1850.770 2084.655 1850.785 ;
        RECT 2075.830 1850.470 2084.655 1850.770 ;
        RECT 2084.325 1850.455 2084.655 1850.470 ;
      LAYER met3 ;
        RECT 1924.400 1838.040 2072.375 1839.440 ;
        RECT 1924.000 1836.720 2072.375 1838.040 ;
      LAYER met3 ;
        RECT 1573.725 1835.810 1574.055 1835.825 ;
        RECT 1574.645 1835.810 1574.975 1835.825 ;
        RECT 1573.725 1835.510 1574.975 1835.810 ;
        RECT 1573.725 1835.495 1574.055 1835.510 ;
        RECT 1574.645 1835.495 1574.975 1835.510 ;
      LAYER met3 ;
        RECT 1924.000 1835.320 2071.975 1836.720 ;
      LAYER met3 ;
        RECT 2072.375 1835.810 2076.375 1836.320 ;
        RECT 2084.785 1835.810 2085.115 1835.825 ;
        RECT 2072.375 1835.720 2085.115 1835.810 ;
        RECT 2075.830 1835.510 2085.115 1835.720 ;
        RECT 2084.785 1835.495 2085.115 1835.510 ;
      LAYER met3 ;
        RECT 364.000 1828.840 626.630 1830.240 ;
      LAYER met3 ;
        RECT 996.885 1829.690 997.215 1829.705 ;
        RECT 1000.000 1829.690 1004.000 1829.840 ;
        RECT 996.885 1829.390 1004.000 1829.690 ;
        RECT 996.885 1829.375 997.215 1829.390 ;
        RECT 1000.000 1829.240 1004.000 1829.390 ;
      LAYER met3 ;
        RECT 1004.400 1828.840 1328.990 1830.240 ;
      LAYER met3 ;
        RECT 1329.390 1829.690 1333.390 1829.840 ;
        RECT 1342.345 1829.690 1342.675 1829.705 ;
        RECT 1329.390 1829.390 1342.675 1829.690 ;
        RECT 1329.390 1829.240 1333.390 1829.390 ;
        RECT 1342.345 1829.375 1342.675 1829.390 ;
      LAYER met3 ;
        RECT 364.000 1815.280 627.030 1828.840 ;
        RECT 364.400 1813.880 627.030 1815.280 ;
        RECT 364.000 1792.160 627.030 1813.880 ;
        RECT 1004.000 1809.840 1329.390 1828.840 ;
        RECT 1924.000 1821.760 2072.375 1835.320 ;
      LAYER met3 ;
        RECT 1920.000 1820.760 1924.000 1821.360 ;
        RECT 1904.465 1818.130 1904.795 1818.145 ;
        RECT 1920.350 1818.130 1920.650 1820.760 ;
      LAYER met3 ;
        RECT 1924.400 1820.400 2072.375 1821.760 ;
        RECT 1924.400 1820.360 2071.975 1820.400 ;
      LAYER met3 ;
        RECT 1904.465 1817.830 1920.650 1818.130 ;
      LAYER met3 ;
        RECT 1924.000 1819.000 2071.975 1820.360 ;
      LAYER met3 ;
        RECT 2072.375 1819.400 2076.375 1820.000 ;
        RECT 1904.465 1817.815 1904.795 1817.830 ;
        RECT 989.065 1809.290 989.395 1809.305 ;
        RECT 1000.000 1809.290 1004.000 1809.440 ;
        RECT 989.065 1808.990 1004.000 1809.290 ;
        RECT 989.065 1808.975 989.395 1808.990 ;
        RECT 1000.000 1808.840 1004.000 1808.990 ;
      LAYER met3 ;
        RECT 1004.400 1808.480 1329.390 1809.840 ;
        RECT 1004.400 1808.440 1328.990 1808.480 ;
        RECT 1004.000 1807.080 1328.990 1808.440 ;
      LAYER met3 ;
        RECT 1329.390 1807.930 1333.390 1808.080 ;
        RECT 1342.805 1807.930 1343.135 1807.945 ;
        RECT 1329.390 1807.630 1343.135 1807.930 ;
        RECT 1329.390 1807.480 1333.390 1807.630 ;
        RECT 1342.805 1807.615 1343.135 1807.630 ;
      LAYER met3 ;
        RECT 364.000 1790.760 626.630 1792.160 ;
        RECT 364.000 1778.560 627.030 1790.760 ;
        RECT 1004.000 1788.080 1329.390 1807.080 ;
        RECT 1924.000 1805.440 2072.375 1819.000 ;
      LAYER met3 ;
        RECT 2075.830 1816.770 2076.130 1819.400 ;
        RECT 2085.245 1816.770 2085.575 1816.785 ;
        RECT 2075.830 1816.470 2085.575 1816.770 ;
        RECT 2085.245 1816.455 2085.575 1816.470 ;
      LAYER met3 ;
        RECT 1924.400 1804.040 2072.375 1805.440 ;
        RECT 1924.000 1802.720 2072.375 1804.040 ;
        RECT 2304.000 1805.760 2524.550 1876.440 ;
        RECT 2304.000 1804.360 2524.150 1805.760 ;
      LAYER met3 ;
        RECT 2524.550 1805.210 2528.550 1805.360 ;
        RECT 2539.725 1805.210 2540.055 1805.225 ;
        RECT 2524.550 1804.910 2540.055 1805.210 ;
        RECT 2524.550 1804.760 2528.550 1804.910 ;
        RECT 2539.725 1804.895 2540.055 1804.910 ;
      LAYER met3 ;
        RECT 1924.000 1801.320 2071.975 1802.720 ;
      LAYER met3 ;
        RECT 2072.375 1801.720 2076.375 1802.320 ;
        RECT 988.605 1787.530 988.935 1787.545 ;
        RECT 1000.000 1787.530 1004.000 1787.680 ;
        RECT 988.605 1787.230 1004.000 1787.530 ;
        RECT 988.605 1787.215 988.935 1787.230 ;
        RECT 1000.000 1787.080 1004.000 1787.230 ;
      LAYER met3 ;
        RECT 1004.400 1786.680 1328.990 1788.080 ;
        RECT 1924.000 1787.760 2072.375 1801.320 ;
      LAYER met3 ;
        RECT 2075.830 1801.130 2076.130 1801.720 ;
        RECT 2085.705 1801.130 2086.035 1801.145 ;
        RECT 2075.830 1800.830 2086.035 1801.130 ;
        RECT 2085.705 1800.815 2086.035 1800.830 ;
      LAYER met3 ;
        RECT 2304.000 1790.800 2524.550 1804.360 ;
      LAYER met3 ;
        RECT 2287.645 1790.250 2287.975 1790.265 ;
        RECT 2300.000 1790.250 2304.000 1790.400 ;
        RECT 2287.645 1789.950 2304.000 1790.250 ;
        RECT 2287.645 1789.935 2287.975 1789.950 ;
        RECT 2300.000 1789.800 2304.000 1789.950 ;
      LAYER met3 ;
        RECT 2304.400 1789.400 2524.550 1790.800 ;
      LAYER met3 ;
        RECT 1329.390 1787.530 1333.390 1787.680 ;
        RECT 1334.525 1787.530 1334.855 1787.545 ;
        RECT 1329.390 1787.230 1334.855 1787.530 ;
        RECT 1329.390 1787.080 1333.390 1787.230 ;
        RECT 1334.525 1787.215 1334.855 1787.230 ;
      LAYER met3 ;
        RECT 364.400 1777.160 627.030 1778.560 ;
        RECT 364.000 1755.440 627.030 1777.160 ;
        RECT 1004.000 1767.680 1329.390 1786.680 ;
        RECT 1924.400 1786.400 2072.375 1787.760 ;
        RECT 1924.400 1786.360 2071.975 1786.400 ;
        RECT 1924.000 1785.000 2071.975 1786.360 ;
      LAYER met3 ;
        RECT 2072.375 1785.400 2076.375 1786.000 ;
      LAYER met3 ;
        RECT 1924.000 1771.440 2072.375 1785.000 ;
      LAYER met3 ;
        RECT 2075.830 1782.770 2076.130 1785.400 ;
        RECT 2086.165 1782.770 2086.495 1782.785 ;
        RECT 2075.830 1782.470 2086.495 1782.770 ;
        RECT 2086.165 1782.455 2086.495 1782.470 ;
        RECT 1920.000 1770.440 1924.000 1771.040 ;
        RECT 1904.465 1767.810 1904.795 1767.825 ;
        RECT 1920.350 1767.810 1920.650 1770.440 ;
      LAYER met3 ;
        RECT 1924.400 1770.040 2072.375 1771.440 ;
      LAYER met3 ;
        RECT 988.145 1767.130 988.475 1767.145 ;
        RECT 1000.000 1767.130 1004.000 1767.280 ;
        RECT 988.145 1766.830 1004.000 1767.130 ;
        RECT 988.145 1766.815 988.475 1766.830 ;
        RECT 1000.000 1766.680 1004.000 1766.830 ;
      LAYER met3 ;
        RECT 1004.400 1766.280 1328.990 1767.680 ;
      LAYER met3 ;
        RECT 1904.465 1767.510 1920.650 1767.810 ;
      LAYER met3 ;
        RECT 1924.000 1768.720 2072.375 1770.040 ;
      LAYER met3 ;
        RECT 1904.465 1767.495 1904.795 1767.510 ;
      LAYER met3 ;
        RECT 1924.000 1767.320 2071.975 1768.720 ;
      LAYER met3 ;
        RECT 2072.375 1767.720 2076.375 1768.320 ;
        RECT 1329.390 1767.130 1333.390 1767.280 ;
        RECT 1343.265 1767.130 1343.595 1767.145 ;
        RECT 1329.390 1766.830 1343.595 1767.130 ;
        RECT 1329.390 1766.680 1333.390 1766.830 ;
        RECT 1343.265 1766.815 1343.595 1766.830 ;
      LAYER met3 ;
        RECT 364.000 1754.040 626.630 1755.440 ;
        RECT 364.000 1741.840 627.030 1754.040 ;
        RECT 1004.000 1745.920 1329.390 1766.280 ;
        RECT 1924.000 1760.715 2072.375 1767.320 ;
      LAYER met3 ;
        RECT 2075.830 1767.130 2076.130 1767.720 ;
        RECT 2086.625 1767.130 2086.955 1767.145 ;
        RECT 2075.830 1766.830 2086.955 1767.130 ;
        RECT 2086.625 1766.815 2086.955 1766.830 ;
        RECT 987.685 1745.370 988.015 1745.385 ;
        RECT 1000.000 1745.370 1004.000 1745.520 ;
        RECT 987.685 1745.070 1004.000 1745.370 ;
        RECT 987.685 1745.055 988.015 1745.070 ;
        RECT 1000.000 1744.920 1004.000 1745.070 ;
      LAYER met3 ;
        RECT 1004.400 1744.520 1328.990 1745.920 ;
      LAYER met3 ;
        RECT 1329.390 1745.370 1333.390 1745.520 ;
        RECT 1336.825 1745.370 1337.155 1745.385 ;
        RECT 1329.390 1745.070 1337.155 1745.370 ;
        RECT 1329.390 1744.920 1333.390 1745.070 ;
        RECT 1336.825 1745.055 1337.155 1745.070 ;
      LAYER met3 ;
        RECT 364.400 1740.440 627.030 1741.840 ;
        RECT 364.000 1718.720 627.030 1740.440 ;
        RECT 1004.000 1725.520 1329.390 1744.520 ;
      LAYER met3 ;
        RECT 1573.725 1739.250 1574.055 1739.265 ;
        RECT 1574.645 1739.250 1574.975 1739.265 ;
        RECT 1573.725 1738.950 1574.975 1739.250 ;
        RECT 1573.725 1738.935 1574.055 1738.950 ;
        RECT 1574.645 1738.935 1574.975 1738.950 ;
        RECT 997.345 1724.970 997.675 1724.985 ;
        RECT 1000.000 1724.970 1004.000 1725.120 ;
        RECT 997.345 1724.670 1004.000 1724.970 ;
        RECT 997.345 1724.655 997.675 1724.670 ;
        RECT 1000.000 1724.520 1004.000 1724.670 ;
      LAYER met3 ;
        RECT 1004.400 1724.120 1328.990 1725.520 ;
      LAYER met3 ;
        RECT 1329.390 1724.970 1333.390 1725.120 ;
        RECT 1337.285 1724.970 1337.615 1724.985 ;
        RECT 1329.390 1724.670 1337.615 1724.970 ;
        RECT 1329.390 1724.520 1333.390 1724.670 ;
        RECT 1337.285 1724.655 1337.615 1724.670 ;
      LAYER met3 ;
        RECT 364.000 1717.320 626.630 1718.720 ;
        RECT 364.000 1704.255 627.030 1717.320 ;
        RECT 1004.000 1710.715 1329.390 1724.120 ;
        RECT 2304.000 1720.080 2524.550 1789.400 ;
        RECT 2304.000 1718.680 2524.150 1720.080 ;
      LAYER met3 ;
        RECT 2524.550 1719.530 2528.550 1719.680 ;
        RECT 2540.185 1719.530 2540.515 1719.545 ;
        RECT 2524.550 1719.230 2540.515 1719.530 ;
        RECT 2524.550 1719.080 2528.550 1719.230 ;
        RECT 2540.185 1719.215 2540.515 1719.230 ;
      LAYER met3 ;
        RECT 2304.000 1710.715 2524.550 1718.680 ;
      LAYER met3 ;
        RECT 1531.405 1690.290 1531.735 1690.305 ;
        RECT 1532.785 1690.290 1533.115 1690.305 ;
        RECT 1531.405 1689.990 1533.115 1690.290 ;
        RECT 1531.405 1689.975 1531.735 1689.990 ;
        RECT 1532.785 1689.975 1533.115 1689.990 ;
        RECT 1351.085 1608.010 1351.415 1608.025 ;
        RECT 1351.085 1607.710 1352.090 1608.010 ;
        RECT 1351.085 1607.695 1351.415 1607.710 ;
        RECT 1351.790 1607.345 1352.090 1607.710 ;
        RECT 1351.545 1607.030 1352.090 1607.345 ;
        RECT 1351.545 1607.015 1351.875 1607.030 ;
        RECT 1532.785 1497.170 1533.115 1497.185 ;
        RECT 1534.165 1497.170 1534.495 1497.185 ;
        RECT 1532.785 1496.870 1534.495 1497.170 ;
        RECT 1532.785 1496.855 1533.115 1496.870 ;
        RECT 1534.165 1496.855 1534.495 1496.870 ;
        RECT 1534.165 1449.570 1534.495 1449.585 ;
        RECT 1533.950 1449.255 1534.495 1449.570 ;
        RECT 1533.245 1448.890 1533.575 1448.905 ;
        RECT 1533.950 1448.890 1534.250 1449.255 ;
        RECT 1533.245 1448.590 1534.250 1448.890 ;
        RECT 1533.245 1448.575 1533.575 1448.590 ;
        RECT 1532.785 1387.010 1533.115 1387.025 ;
        RECT 1533.705 1387.010 1534.035 1387.025 ;
        RECT 1532.785 1386.710 1534.035 1387.010 ;
        RECT 1532.785 1386.695 1533.115 1386.710 ;
        RECT 1533.705 1386.695 1534.035 1386.710 ;
        RECT 1543.365 1345.530 1543.695 1345.545 ;
        RECT 1544.285 1345.530 1544.615 1345.545 ;
        RECT 1543.365 1345.230 1544.615 1345.530 ;
        RECT 1543.365 1345.215 1543.695 1345.230 ;
        RECT 1544.285 1345.215 1544.615 1345.230 ;
        RECT 1350.625 1255.770 1350.955 1255.785 ;
        RECT 1351.545 1255.770 1351.875 1255.785 ;
        RECT 1350.625 1255.470 1351.875 1255.770 ;
        RECT 1350.625 1255.455 1350.955 1255.470 ;
        RECT 1351.545 1255.455 1351.875 1255.470 ;
        RECT 1531.405 1248.970 1531.735 1248.985 ;
        RECT 1532.785 1248.970 1533.115 1248.985 ;
        RECT 1531.405 1248.670 1533.115 1248.970 ;
        RECT 1531.405 1248.655 1531.735 1248.670 ;
        RECT 1532.785 1248.655 1533.115 1248.670 ;
        RECT 1351.545 1207.490 1351.875 1207.505 ;
        RECT 1351.545 1207.175 1352.090 1207.490 ;
        RECT 1350.165 1206.810 1350.495 1206.825 ;
        RECT 1351.790 1206.810 1352.090 1207.175 ;
        RECT 1350.165 1206.510 1352.090 1206.810 ;
        RECT 1350.165 1206.495 1350.495 1206.510 ;
        RECT 978.945 1014.370 979.275 1014.385 ;
        RECT 1100.845 1014.370 1101.175 1014.385 ;
        RECT 978.945 1014.070 1101.175 1014.370 ;
        RECT 978.945 1014.055 979.275 1014.070 ;
        RECT 1100.845 1014.055 1101.175 1014.070 ;
        RECT 1573.725 1014.370 1574.055 1014.385 ;
        RECT 1575.565 1014.370 1575.895 1014.385 ;
        RECT 1573.725 1014.070 1575.895 1014.370 ;
        RECT 1573.725 1014.055 1574.055 1014.070 ;
        RECT 1575.565 1014.055 1575.895 1014.070 ;
        RECT 994.125 1013.690 994.455 1013.705 ;
        RECT 1124.765 1013.690 1125.095 1013.705 ;
        RECT 994.125 1013.390 1125.095 1013.690 ;
        RECT 994.125 1013.375 994.455 1013.390 ;
        RECT 1124.765 1013.375 1125.095 1013.390 ;
        RECT 985.385 1013.010 985.715 1013.025 ;
        RECT 1128.905 1013.010 1129.235 1013.025 ;
        RECT 985.385 1012.710 1129.235 1013.010 ;
        RECT 985.385 1012.695 985.715 1012.710 ;
        RECT 1128.905 1012.695 1129.235 1012.710 ;
        RECT 1751.285 1013.010 1751.615 1013.025 ;
        RECT 1753.125 1013.010 1753.455 1013.025 ;
        RECT 1751.285 1012.710 1753.455 1013.010 ;
        RECT 1751.285 1012.695 1751.615 1012.710 ;
        RECT 1753.125 1012.695 1753.455 1012.710 ;
        RECT 978.485 1012.330 978.815 1012.345 ;
        RECT 1117.865 1012.330 1118.195 1012.345 ;
        RECT 978.485 1012.030 1118.195 1012.330 ;
        RECT 978.485 1012.015 978.815 1012.030 ;
        RECT 1117.865 1012.015 1118.195 1012.030 ;
        RECT 979.405 1011.650 979.735 1011.665 ;
        RECT 1141.785 1011.650 1142.115 1011.665 ;
        RECT 979.405 1011.350 1142.115 1011.650 ;
        RECT 979.405 1011.335 979.735 1011.350 ;
        RECT 1141.785 1011.335 1142.115 1011.350 ;
        RECT 986.305 1010.970 986.635 1010.985 ;
        RECT 1166.165 1010.970 1166.495 1010.985 ;
        RECT 986.305 1010.670 1166.495 1010.970 ;
        RECT 986.305 1010.655 986.635 1010.670 ;
        RECT 1166.165 1010.655 1166.495 1010.670 ;
        RECT 985.845 1010.290 986.175 1010.305 ;
        RECT 1087.505 1010.290 1087.835 1010.305 ;
        RECT 985.845 1009.990 1087.835 1010.290 ;
        RECT 985.845 1009.975 986.175 1009.990 ;
        RECT 1087.505 1009.975 1087.835 1009.990 ;
        RECT 993.205 1009.610 993.535 1009.625 ;
        RECT 1065.885 1009.610 1066.215 1009.625 ;
        RECT 993.205 1009.310 1066.215 1009.610 ;
        RECT 993.205 1009.295 993.535 1009.310 ;
        RECT 1065.885 1009.295 1066.215 1009.310 ;
        RECT 670.000 996.480 674.000 997.080 ;
        RECT 2166.000 994.440 2170.000 995.040 ;
      LAYER met3 ;
        RECT 674.000 992.720 2166.000 992.865 ;
      LAYER met3 ;
        RECT 670.000 991.720 674.000 992.320 ;
      LAYER met3 ;
        RECT 674.400 991.320 2166.000 992.720 ;
        RECT 674.000 987.280 2166.000 991.320 ;
      LAYER met3 ;
        RECT 670.000 986.280 674.000 986.880 ;
      LAYER met3 ;
        RECT 674.400 985.880 2166.000 987.280 ;
        RECT 674.000 985.240 2166.000 985.880 ;
        RECT 674.000 983.840 2165.600 985.240 ;
      LAYER met3 ;
        RECT 2166.000 984.240 2170.000 984.840 ;
      LAYER met3 ;
        RECT 674.000 982.520 2166.000 983.840 ;
        RECT 674.400 981.120 2166.000 982.520 ;
        RECT 674.000 977.080 2166.000 981.120 ;
        RECT 674.400 975.680 2166.000 977.080 ;
        RECT 674.000 975.040 2166.000 975.680 ;
        RECT 674.000 973.640 2165.600 975.040 ;
        RECT 674.000 972.320 2166.000 973.640 ;
        RECT 674.400 970.920 2166.000 972.320 ;
        RECT 674.000 966.880 2166.000 970.920 ;
        RECT 674.400 965.520 2166.000 966.880 ;
        RECT 674.400 965.480 2165.600 965.520 ;
        RECT 674.000 964.120 2165.600 965.480 ;
        RECT 674.000 962.120 2166.000 964.120 ;
        RECT 674.400 960.720 2166.000 962.120 ;
        RECT 674.000 957.360 2166.000 960.720 ;
        RECT 674.400 955.960 2166.000 957.360 ;
        RECT 674.000 955.320 2166.000 955.960 ;
        RECT 674.000 953.920 2165.600 955.320 ;
        RECT 674.000 951.920 2166.000 953.920 ;
        RECT 674.400 950.520 2166.000 951.920 ;
        RECT 674.000 947.160 2166.000 950.520 ;
        RECT 674.400 945.760 2166.000 947.160 ;
        RECT 674.000 945.120 2166.000 945.760 ;
        RECT 674.000 943.720 2165.600 945.120 ;
        RECT 674.000 941.720 2166.000 943.720 ;
        RECT 674.400 940.320 2166.000 941.720 ;
        RECT 674.000 936.960 2166.000 940.320 ;
        RECT 674.400 935.600 2166.000 936.960 ;
        RECT 674.400 935.560 2165.600 935.600 ;
        RECT 674.000 934.200 2165.600 935.560 ;
        RECT 674.000 931.520 2166.000 934.200 ;
        RECT 674.400 930.120 2166.000 931.520 ;
        RECT 674.000 926.760 2166.000 930.120 ;
        RECT 674.400 925.400 2166.000 926.760 ;
        RECT 674.400 925.360 2165.600 925.400 ;
        RECT 674.000 924.000 2165.600 925.360 ;
        RECT 674.000 921.320 2166.000 924.000 ;
        RECT 674.400 919.920 2166.000 921.320 ;
        RECT 674.000 916.560 2166.000 919.920 ;
        RECT 674.400 915.200 2166.000 916.560 ;
        RECT 674.400 915.160 2165.600 915.200 ;
        RECT 674.000 913.800 2165.600 915.160 ;
        RECT 674.000 911.800 2166.000 913.800 ;
        RECT 674.400 910.400 2166.000 911.800 ;
        RECT 674.000 906.360 2166.000 910.400 ;
        RECT 674.400 905.680 2166.000 906.360 ;
        RECT 674.400 904.960 2165.600 905.680 ;
        RECT 674.000 904.280 2165.600 904.960 ;
        RECT 674.000 901.600 2166.000 904.280 ;
        RECT 674.400 900.200 2166.000 901.600 ;
        RECT 674.000 896.160 2166.000 900.200 ;
        RECT 674.400 895.480 2166.000 896.160 ;
        RECT 674.400 894.760 2165.600 895.480 ;
        RECT 674.000 894.080 2165.600 894.760 ;
        RECT 674.000 891.400 2166.000 894.080 ;
        RECT 674.400 890.000 2166.000 891.400 ;
        RECT 674.000 885.960 2166.000 890.000 ;
        RECT 674.400 885.280 2166.000 885.960 ;
        RECT 674.400 884.560 2165.600 885.280 ;
        RECT 674.000 883.880 2165.600 884.560 ;
        RECT 674.000 881.200 2166.000 883.880 ;
        RECT 674.400 879.800 2166.000 881.200 ;
        RECT 674.000 875.760 2166.000 879.800 ;
        RECT 674.400 875.080 2166.000 875.760 ;
        RECT 674.400 874.360 2165.600 875.080 ;
        RECT 674.000 873.680 2165.600 874.360 ;
        RECT 674.000 871.000 2166.000 873.680 ;
        RECT 674.400 869.600 2166.000 871.000 ;
        RECT 674.000 866.240 2166.000 869.600 ;
        RECT 674.400 865.560 2166.000 866.240 ;
        RECT 674.400 864.840 2165.600 865.560 ;
        RECT 674.000 864.160 2165.600 864.840 ;
        RECT 674.000 860.800 2166.000 864.160 ;
        RECT 674.400 859.400 2166.000 860.800 ;
        RECT 674.000 856.040 2166.000 859.400 ;
        RECT 674.400 855.360 2166.000 856.040 ;
        RECT 674.400 854.640 2165.600 855.360 ;
        RECT 674.000 853.960 2165.600 854.640 ;
        RECT 674.000 850.600 2166.000 853.960 ;
        RECT 674.400 849.200 2166.000 850.600 ;
        RECT 674.000 845.840 2166.000 849.200 ;
        RECT 674.400 845.160 2166.000 845.840 ;
        RECT 674.400 844.440 2165.600 845.160 ;
        RECT 674.000 843.760 2165.600 844.440 ;
        RECT 674.000 840.400 2166.000 843.760 ;
        RECT 674.400 839.000 2166.000 840.400 ;
        RECT 674.000 835.640 2166.000 839.000 ;
        RECT 674.400 834.240 2165.600 835.640 ;
        RECT 674.000 830.200 2166.000 834.240 ;
        RECT 674.400 828.800 2166.000 830.200 ;
        RECT 674.000 825.440 2166.000 828.800 ;
        RECT 674.400 824.040 2165.600 825.440 ;
        RECT 674.000 820.680 2166.000 824.040 ;
        RECT 674.400 819.280 2166.000 820.680 ;
        RECT 674.000 815.240 2166.000 819.280 ;
        RECT 674.400 813.840 2165.600 815.240 ;
        RECT 674.000 810.480 2166.000 813.840 ;
        RECT 674.400 809.080 2166.000 810.480 ;
        RECT 674.000 805.720 2166.000 809.080 ;
        RECT 674.000 805.040 2165.600 805.720 ;
        RECT 674.400 804.320 2165.600 805.040 ;
        RECT 674.400 803.640 2166.000 804.320 ;
        RECT 674.000 800.280 2166.000 803.640 ;
        RECT 674.400 798.880 2166.000 800.280 ;
        RECT 674.000 795.520 2166.000 798.880 ;
        RECT 674.000 794.840 2165.600 795.520 ;
        RECT 674.400 794.120 2165.600 794.840 ;
        RECT 674.400 793.440 2166.000 794.120 ;
        RECT 674.000 790.080 2166.000 793.440 ;
        RECT 674.400 788.680 2166.000 790.080 ;
        RECT 674.000 785.320 2166.000 788.680 ;
        RECT 674.000 784.640 2165.600 785.320 ;
        RECT 674.400 783.920 2165.600 784.640 ;
        RECT 674.400 783.240 2166.000 783.920 ;
        RECT 674.000 779.880 2166.000 783.240 ;
        RECT 674.400 778.480 2166.000 779.880 ;
        RECT 674.000 775.120 2166.000 778.480 ;
        RECT 674.400 773.720 2165.600 775.120 ;
        RECT 674.000 769.680 2166.000 773.720 ;
        RECT 674.400 768.280 2166.000 769.680 ;
        RECT 674.000 765.600 2166.000 768.280 ;
        RECT 674.000 764.920 2165.600 765.600 ;
        RECT 674.400 764.200 2165.600 764.920 ;
        RECT 674.400 763.520 2166.000 764.200 ;
        RECT 674.000 759.480 2166.000 763.520 ;
        RECT 674.400 758.080 2166.000 759.480 ;
        RECT 674.000 755.400 2166.000 758.080 ;
        RECT 674.000 754.720 2165.600 755.400 ;
        RECT 674.400 754.000 2165.600 754.720 ;
        RECT 674.400 753.320 2166.000 754.000 ;
        RECT 674.000 749.280 2166.000 753.320 ;
        RECT 674.400 747.880 2166.000 749.280 ;
        RECT 674.000 745.200 2166.000 747.880 ;
        RECT 674.000 744.520 2165.600 745.200 ;
        RECT 674.400 743.800 2165.600 744.520 ;
        RECT 674.400 743.120 2166.000 743.800 ;
        RECT 674.000 739.080 2166.000 743.120 ;
        RECT 674.400 737.680 2166.000 739.080 ;
        RECT 674.000 735.680 2166.000 737.680 ;
        RECT 674.000 734.320 2165.600 735.680 ;
        RECT 674.400 734.280 2165.600 734.320 ;
        RECT 674.400 732.920 2166.000 734.280 ;
        RECT 674.000 729.560 2166.000 732.920 ;
        RECT 674.400 728.160 2166.000 729.560 ;
        RECT 674.000 725.480 2166.000 728.160 ;
        RECT 674.000 724.120 2165.600 725.480 ;
        RECT 674.400 724.080 2165.600 724.120 ;
        RECT 674.400 722.720 2166.000 724.080 ;
        RECT 674.000 719.360 2166.000 722.720 ;
        RECT 674.400 717.960 2166.000 719.360 ;
        RECT 674.000 715.280 2166.000 717.960 ;
        RECT 674.000 713.920 2165.600 715.280 ;
        RECT 674.400 713.880 2165.600 713.920 ;
        RECT 674.400 712.520 2166.000 713.880 ;
        RECT 674.000 709.160 2166.000 712.520 ;
        RECT 674.400 707.760 2166.000 709.160 ;
        RECT 674.000 705.760 2166.000 707.760 ;
        RECT 674.000 704.360 2165.600 705.760 ;
        RECT 674.000 703.720 2166.000 704.360 ;
        RECT 674.400 702.320 2166.000 703.720 ;
        RECT 674.000 698.960 2166.000 702.320 ;
        RECT 674.400 697.560 2166.000 698.960 ;
        RECT 674.000 695.560 2166.000 697.560 ;
        RECT 674.000 694.160 2165.600 695.560 ;
        RECT 674.000 693.520 2166.000 694.160 ;
        RECT 674.400 692.120 2166.000 693.520 ;
        RECT 674.000 688.760 2166.000 692.120 ;
        RECT 674.400 687.360 2166.000 688.760 ;
        RECT 674.000 685.360 2166.000 687.360 ;
        RECT 674.000 684.000 2165.600 685.360 ;
        RECT 674.400 683.960 2165.600 684.000 ;
        RECT 674.400 682.600 2166.000 683.960 ;
        RECT 674.000 678.560 2166.000 682.600 ;
        RECT 674.400 677.160 2166.000 678.560 ;
        RECT 674.000 675.160 2166.000 677.160 ;
        RECT 674.000 673.800 2165.600 675.160 ;
        RECT 674.400 673.760 2165.600 673.800 ;
        RECT 674.400 672.400 2166.000 673.760 ;
        RECT 674.000 668.360 2166.000 672.400 ;
        RECT 674.400 666.960 2166.000 668.360 ;
        RECT 674.000 665.640 2166.000 666.960 ;
        RECT 674.000 664.240 2165.600 665.640 ;
        RECT 674.000 663.600 2166.000 664.240 ;
        RECT 674.400 662.200 2166.000 663.600 ;
        RECT 674.000 658.160 2166.000 662.200 ;
        RECT 674.400 656.760 2166.000 658.160 ;
        RECT 674.000 655.440 2166.000 656.760 ;
        RECT 674.000 654.040 2165.600 655.440 ;
        RECT 674.000 653.400 2166.000 654.040 ;
        RECT 674.400 652.000 2166.000 653.400 ;
        RECT 674.000 647.960 2166.000 652.000 ;
        RECT 674.400 646.560 2166.000 647.960 ;
        RECT 674.000 645.240 2166.000 646.560 ;
        RECT 674.000 643.840 2165.600 645.240 ;
        RECT 674.000 643.200 2166.000 643.840 ;
        RECT 674.400 641.800 2166.000 643.200 ;
        RECT 674.000 638.440 2166.000 641.800 ;
        RECT 674.400 637.040 2166.000 638.440 ;
        RECT 674.000 635.720 2166.000 637.040 ;
        RECT 674.000 634.320 2165.600 635.720 ;
        RECT 674.000 633.000 2166.000 634.320 ;
        RECT 674.400 631.600 2166.000 633.000 ;
        RECT 674.000 628.240 2166.000 631.600 ;
        RECT 674.400 626.840 2166.000 628.240 ;
        RECT 674.000 625.520 2166.000 626.840 ;
        RECT 674.000 624.120 2165.600 625.520 ;
        RECT 674.000 622.800 2166.000 624.120 ;
        RECT 674.400 621.400 2166.000 622.800 ;
        RECT 674.000 618.040 2166.000 621.400 ;
        RECT 674.400 616.640 2166.000 618.040 ;
        RECT 674.000 615.320 2166.000 616.640 ;
        RECT 674.000 613.920 2165.600 615.320 ;
        RECT 674.000 612.600 2166.000 613.920 ;
        RECT 674.400 611.200 2166.000 612.600 ;
        RECT 674.000 607.840 2166.000 611.200 ;
        RECT 674.400 606.440 2166.000 607.840 ;
        RECT 674.000 605.800 2166.000 606.440 ;
        RECT 674.000 604.400 2165.600 605.800 ;
        RECT 674.000 603.080 2166.000 604.400 ;
        RECT 674.400 602.215 2166.000 603.080 ;
      LAYER via3 ;
        RECT 1532.100 2062.620 1532.420 2062.940 ;
        RECT 1532.100 2027.940 1532.420 2028.260 ;
      LAYER met4 ;
        RECT 459.645 2610.640 480.165 2747.120 ;
        RECT 482.565 2610.640 550.935 2747.120 ;
        RECT 1036.375 2610.640 1080.450 2787.920 ;
        RECT 1600.575 2510.640 1829.840 2889.200 ;
        RECT 2477.790 2610.640 2529.990 2760.720 ;
      LAYER met4 ;
        RECT 1532.095 2062.615 1532.425 2062.945 ;
      LAYER met4 ;
        RECT 534.640 1710.640 613.040 1969.520 ;
        RECT 1174.640 1710.640 1253.040 2032.080 ;
      LAYER met4 ;
        RECT 1532.110 2028.265 1532.410 2062.615 ;
        RECT 1532.095 2027.935 1532.425 2028.265 ;
      LAYER met4 ;
        RECT 1997.170 1760.640 2047.070 1905.280 ;
        RECT 2474.640 1710.640 2476.240 1926.000 ;
        RECT 808.295 610.640 2151.840 990.825 ;
  END
END user_project_wrapper
END LIBRARY

