VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vga_clock
  CLASS BLOCK ;
  FOREIGN vga_clock ;
  ORIGIN 0.000 0.000 ;
  SIZE 228.550 BY 239.270 ;
  PIN adj_hrs
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END adj_hrs
  PIN adj_min
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 224.550 191.800 228.550 192.400 ;
    END
  END adj_min
  PIN adj_sec
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END adj_sec
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END clk
  PIN hsync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 224.550 104.760 228.550 105.360 ;
    END
  END hsync
  PIN reset_n
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 235.270 80.410 239.270 ;
    END
  END reset_n
  PIN rrggbb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END rrggbb[0]
  PIN rrggbb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END rrggbb[1]
  PIN rrggbb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 224.550 19.080 228.550 19.680 ;
    END
  END rrggbb[2]
  PIN rrggbb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.250 235.270 21.530 239.270 ;
    END
  END rrggbb[3]
  PIN rrggbb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.970 235.270 197.250 239.270 ;
    END
  END rrggbb[4]
  PIN rrggbb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.090 235.270 138.370 239.270 ;
    END
  END rrggbb[5]
  PIN vsync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END vsync
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 226.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 226.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 222.640 225.845 ;
      LAYER met1 ;
        RECT 2.830 10.640 222.640 226.000 ;
      LAYER met2 ;
        RECT 2.860 234.990 20.970 235.270 ;
        RECT 21.810 234.990 79.850 235.270 ;
        RECT 80.690 234.990 137.810 235.270 ;
        RECT 138.650 234.990 196.690 235.270 ;
        RECT 197.530 234.990 219.320 235.270 ;
        RECT 2.860 4.280 219.320 234.990 ;
        RECT 3.410 4.000 60.530 4.280 ;
        RECT 61.370 4.000 119.410 4.280 ;
        RECT 120.250 4.000 177.370 4.280 ;
        RECT 178.210 4.000 219.320 4.280 ;
      LAYER met3 ;
        RECT 4.000 192.800 224.550 225.925 ;
        RECT 4.000 191.400 224.150 192.800 ;
        RECT 4.000 177.840 224.550 191.400 ;
        RECT 4.400 176.440 224.550 177.840 ;
        RECT 4.000 105.760 224.550 176.440 ;
        RECT 4.000 104.360 224.150 105.760 ;
        RECT 4.000 90.800 224.550 104.360 ;
        RECT 4.400 89.400 224.550 90.800 ;
        RECT 4.000 20.080 224.550 89.400 ;
        RECT 4.000 18.680 224.150 20.080 ;
        RECT 4.000 10.715 224.550 18.680 ;
      LAYER met4 ;
        RECT 174.640 10.640 176.240 226.000 ;
  END
END vga_clock
END LIBRARY

