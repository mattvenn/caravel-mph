VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2183.690 89.660 2184.010 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2183.690 89.520 2899.310 89.660 ;
        RECT 2183.690 89.460 2184.010 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2183.720 89.460 2183.980 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2183.710 601.955 2183.990 602.325 ;
        RECT 2183.780 89.750 2183.920 601.955 ;
        RECT 2183.720 89.430 2183.980 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2183.710 602.000 2183.990 602.280 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2166.000 604.800 2170.000 605.400 ;
        RECT 2169.670 602.290 2169.970 604.800 ;
        RECT 2183.685 602.290 2184.015 602.305 ;
        RECT 2169.670 601.990 2184.015 602.290 ;
        RECT 2183.685 601.975 2184.015 601.990 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2191.510 2429.200 2191.830 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 2191.510 2429.060 2901.150 2429.200 ;
        RECT 2191.510 2429.000 2191.830 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 2180.470 710.500 2180.790 710.560 ;
        RECT 2191.510 710.500 2191.830 710.560 ;
        RECT 2180.470 710.360 2191.830 710.500 ;
        RECT 2180.470 710.300 2180.790 710.360 ;
        RECT 2191.510 710.300 2191.830 710.360 ;
      LAYER via ;
        RECT 2191.540 2429.000 2191.800 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 2180.500 710.300 2180.760 710.560 ;
        RECT 2191.540 710.300 2191.800 710.560 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 2191.540 2428.970 2191.800 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 2191.600 710.590 2191.740 2428.970 ;
        RECT 2180.500 710.445 2180.760 710.590 ;
        RECT 2180.490 710.075 2180.770 710.445 ;
        RECT 2191.540 710.270 2191.800 710.590 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 2180.490 710.120 2180.770 710.400 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2180.465 710.410 2180.795 710.425 ;
        RECT 2169.670 710.120 2180.795 710.410 ;
        RECT 2166.000 710.110 2180.795 710.120 ;
        RECT 2166.000 709.520 2170.000 710.110 ;
        RECT 2180.465 710.095 2180.795 710.110 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 724.440 2187.230 724.500 ;
        RECT 2901.290 724.440 2901.610 724.500 ;
        RECT 2186.910 724.300 2901.610 724.440 ;
        RECT 2186.910 724.240 2187.230 724.300 ;
        RECT 2901.290 724.240 2901.610 724.300 ;
      LAYER via ;
        RECT 2186.940 724.240 2187.200 724.500 ;
        RECT 2901.320 724.240 2901.580 724.500 ;
      LAYER met2 ;
        RECT 2901.310 2669.155 2901.590 2669.525 ;
        RECT 2901.380 724.530 2901.520 2669.155 ;
        RECT 2186.940 724.210 2187.200 724.530 ;
        RECT 2901.320 724.210 2901.580 724.530 ;
        RECT 2187.000 722.685 2187.140 724.210 ;
        RECT 2186.930 722.315 2187.210 722.685 ;
      LAYER via2 ;
        RECT 2901.310 2669.200 2901.590 2669.480 ;
        RECT 2186.930 722.360 2187.210 722.640 ;
      LAYER met3 ;
        RECT 2901.285 2669.490 2901.615 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2901.285 2669.190 2924.800 2669.490 ;
        RECT 2901.285 2669.175 2901.615 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2186.905 722.650 2187.235 722.665 ;
        RECT 2169.670 722.350 2187.235 722.650 ;
        RECT 2169.670 721.000 2169.970 722.350 ;
        RECT 2186.905 722.335 2187.235 722.350 ;
        RECT 2166.000 720.400 2170.000 721.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2191.050 2898.400 2191.370 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2191.050 2898.260 2901.150 2898.400 ;
        RECT 2191.050 2898.200 2191.370 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2180.470 731.240 2180.790 731.300 ;
        RECT 2191.050 731.240 2191.370 731.300 ;
        RECT 2180.470 731.100 2191.370 731.240 ;
        RECT 2180.470 731.040 2180.790 731.100 ;
        RECT 2191.050 731.040 2191.370 731.100 ;
      LAYER via ;
        RECT 2191.080 2898.200 2191.340 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2180.500 731.040 2180.760 731.300 ;
        RECT 2191.080 731.040 2191.340 731.300 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2191.080 2898.170 2191.340 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2180.490 731.155 2180.770 731.525 ;
        RECT 2191.140 731.330 2191.280 2898.170 ;
        RECT 2180.500 731.010 2180.760 731.155 ;
        RECT 2191.080 731.010 2191.340 731.330 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 2180.490 731.200 2180.770 731.480 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2180.465 731.490 2180.795 731.505 ;
        RECT 2169.670 731.200 2180.795 731.490 ;
        RECT 2166.000 731.190 2180.795 731.200 ;
        RECT 2166.000 730.600 2170.000 731.190 ;
        RECT 2180.465 731.175 2180.795 731.190 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2197.490 3133.000 2197.810 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2197.490 3132.860 2901.150 3133.000 ;
        RECT 2197.490 3132.800 2197.810 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 2180.930 744.500 2181.250 744.560 ;
        RECT 2197.490 744.500 2197.810 744.560 ;
        RECT 2180.930 744.360 2197.810 744.500 ;
        RECT 2180.930 744.300 2181.250 744.360 ;
        RECT 2197.490 744.300 2197.810 744.360 ;
      LAYER via ;
        RECT 2197.520 3132.800 2197.780 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 2180.960 744.300 2181.220 744.560 ;
        RECT 2197.520 744.300 2197.780 744.560 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2197.520 3132.770 2197.780 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 2197.580 744.590 2197.720 3132.770 ;
        RECT 2180.960 744.445 2181.220 744.590 ;
        RECT 2180.950 744.075 2181.230 744.445 ;
        RECT 2197.520 744.270 2197.780 744.590 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 2180.950 744.120 2181.230 744.400 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2180.925 744.410 2181.255 744.425 ;
        RECT 2169.670 744.110 2181.255 744.410 ;
        RECT 2169.670 742.080 2169.970 744.110 ;
        RECT 2180.925 744.095 2181.255 744.110 ;
        RECT 2166.000 741.480 2170.000 742.080 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2204.390 3367.600 2204.710 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2204.390 3367.460 2901.150 3367.600 ;
        RECT 2204.390 3367.400 2204.710 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 2185.070 751.640 2185.390 751.700 ;
        RECT 2204.390 751.640 2204.710 751.700 ;
        RECT 2185.070 751.500 2204.710 751.640 ;
        RECT 2185.070 751.440 2185.390 751.500 ;
        RECT 2204.390 751.440 2204.710 751.500 ;
      LAYER via ;
        RECT 2204.420 3367.400 2204.680 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 2185.100 751.440 2185.360 751.700 ;
        RECT 2204.420 751.440 2204.680 751.700 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2204.420 3367.370 2204.680 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 2204.480 751.730 2204.620 3367.370 ;
        RECT 2185.100 751.410 2185.360 751.730 ;
        RECT 2204.420 751.410 2204.680 751.730 ;
        RECT 2185.160 751.245 2185.300 751.410 ;
        RECT 2185.090 750.875 2185.370 751.245 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 2185.090 750.920 2185.370 751.200 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2166.000 751.680 2170.000 752.280 ;
        RECT 2169.670 751.210 2169.970 751.680 ;
        RECT 2185.065 751.210 2185.395 751.225 ;
        RECT 2169.670 750.910 2185.395 751.210 ;
        RECT 2185.065 750.895 2185.395 750.910 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2211.290 3502.240 2211.610 3502.300 ;
        RECT 2798.250 3502.240 2798.570 3502.300 ;
        RECT 2211.290 3502.100 2798.570 3502.240 ;
        RECT 2211.290 3502.040 2211.610 3502.100 ;
        RECT 2798.250 3502.040 2798.570 3502.100 ;
        RECT 2186.910 759.800 2187.230 759.860 ;
        RECT 2211.290 759.800 2211.610 759.860 ;
        RECT 2186.910 759.660 2211.610 759.800 ;
        RECT 2186.910 759.600 2187.230 759.660 ;
        RECT 2211.290 759.600 2211.610 759.660 ;
      LAYER via ;
        RECT 2211.320 3502.040 2211.580 3502.300 ;
        RECT 2798.280 3502.040 2798.540 3502.300 ;
        RECT 2186.940 759.600 2187.200 759.860 ;
        RECT 2211.320 759.600 2211.580 759.860 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3502.330 2798.480 3517.600 ;
        RECT 2211.320 3502.010 2211.580 3502.330 ;
        RECT 2798.280 3502.010 2798.540 3502.330 ;
        RECT 2186.930 761.075 2187.210 761.445 ;
        RECT 2187.000 759.890 2187.140 761.075 ;
        RECT 2211.380 759.890 2211.520 3502.010 ;
        RECT 2186.940 759.570 2187.200 759.890 ;
        RECT 2211.320 759.570 2211.580 759.890 ;
      LAYER via2 ;
        RECT 2186.930 761.120 2187.210 761.400 ;
      LAYER met3 ;
        RECT 2166.000 762.560 2170.000 763.160 ;
        RECT 2169.670 761.410 2169.970 762.560 ;
        RECT 2186.905 761.410 2187.235 761.425 ;
        RECT 2169.670 761.110 2187.235 761.410 ;
        RECT 2186.905 761.095 2187.235 761.110 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2190.590 3503.260 2190.910 3503.320 ;
        RECT 2473.950 3503.260 2474.270 3503.320 ;
        RECT 2190.590 3503.120 2474.270 3503.260 ;
        RECT 2190.590 3503.060 2190.910 3503.120 ;
        RECT 2473.950 3503.060 2474.270 3503.120 ;
        RECT 2180.470 778.160 2180.790 778.220 ;
        RECT 2190.590 778.160 2190.910 778.220 ;
        RECT 2180.470 778.020 2190.910 778.160 ;
        RECT 2180.470 777.960 2180.790 778.020 ;
        RECT 2190.590 777.960 2190.910 778.020 ;
      LAYER via ;
        RECT 2190.620 3503.060 2190.880 3503.320 ;
        RECT 2473.980 3503.060 2474.240 3503.320 ;
        RECT 2180.500 777.960 2180.760 778.220 ;
        RECT 2190.620 777.960 2190.880 778.220 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3503.350 2474.180 3517.600 ;
        RECT 2190.620 3503.030 2190.880 3503.350 ;
        RECT 2473.980 3503.030 2474.240 3503.350 ;
        RECT 2190.680 778.250 2190.820 3503.030 ;
        RECT 2180.500 777.930 2180.760 778.250 ;
        RECT 2190.620 777.930 2190.880 778.250 ;
        RECT 2180.560 775.725 2180.700 777.930 ;
        RECT 2180.490 775.355 2180.770 775.725 ;
      LAYER via2 ;
        RECT 2180.490 775.400 2180.770 775.680 ;
      LAYER met3 ;
        RECT 2180.465 775.690 2180.795 775.705 ;
        RECT 2169.670 775.390 2180.795 775.690 ;
        RECT 2169.670 773.360 2169.970 775.390 ;
        RECT 2180.465 775.375 2180.795 775.390 ;
        RECT 2166.000 772.760 2170.000 773.360 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2149.190 3498.500 2149.510 3498.560 ;
        RECT 2169.430 3498.500 2169.750 3498.560 ;
        RECT 2149.190 3498.360 2169.750 3498.500 ;
        RECT 2149.190 3498.300 2149.510 3498.360 ;
        RECT 2169.430 3498.300 2169.750 3498.360 ;
      LAYER via ;
        RECT 2149.220 3498.300 2149.480 3498.560 ;
        RECT 2169.460 3498.300 2169.720 3498.560 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3498.590 2149.420 3517.600 ;
        RECT 2149.220 3498.270 2149.480 3498.590 ;
        RECT 2169.460 3498.270 2169.720 3498.590 ;
        RECT 2169.520 786.605 2169.660 3498.270 ;
        RECT 2169.450 786.235 2169.730 786.605 ;
      LAYER via2 ;
        RECT 2169.450 786.280 2169.730 786.560 ;
      LAYER met3 ;
        RECT 2169.425 786.570 2169.755 786.585 ;
        RECT 2169.425 786.255 2169.970 786.570 ;
        RECT 2169.670 784.240 2169.970 786.255 ;
        RECT 2166.000 783.640 2170.000 784.240 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3504.620 1825.210 3504.680 ;
        RECT 2169.890 3504.620 2170.210 3504.680 ;
        RECT 1824.890 3504.480 2170.210 3504.620 ;
        RECT 1824.890 3504.420 1825.210 3504.480 ;
        RECT 2169.890 3504.420 2170.210 3504.480 ;
      LAYER via ;
        RECT 1824.920 3504.420 1825.180 3504.680 ;
        RECT 2169.920 3504.420 2170.180 3504.680 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3504.710 1825.120 3517.600 ;
        RECT 1824.920 3504.390 1825.180 3504.710 ;
        RECT 2169.920 3504.390 2170.180 3504.710 ;
        RECT 2169.980 796.805 2170.120 3504.390 ;
        RECT 2169.910 796.435 2170.190 796.805 ;
      LAYER via2 ;
        RECT 2169.910 796.480 2170.190 796.760 ;
      LAYER met3 ;
        RECT 2169.885 796.770 2170.215 796.785 ;
        RECT 2169.670 796.455 2170.215 796.770 ;
        RECT 2169.670 794.440 2169.970 796.455 ;
        RECT 2166.000 793.840 2170.000 794.440 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3500.880 1500.910 3500.940 ;
        RECT 2180.470 3500.880 2180.790 3500.940 ;
        RECT 1500.590 3500.740 2180.790 3500.880 ;
        RECT 1500.590 3500.680 1500.910 3500.740 ;
        RECT 2180.470 3500.680 2180.790 3500.740 ;
      LAYER via ;
        RECT 1500.620 3500.680 1500.880 3500.940 ;
        RECT 2180.500 3500.680 2180.760 3500.940 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3500.970 1500.820 3517.600 ;
        RECT 1500.620 3500.650 1500.880 3500.970 ;
        RECT 2180.500 3500.650 2180.760 3500.970 ;
        RECT 2180.560 806.325 2180.700 3500.650 ;
        RECT 2180.490 805.955 2180.770 806.325 ;
      LAYER via2 ;
        RECT 2180.490 806.000 2180.770 806.280 ;
      LAYER met3 ;
        RECT 2180.465 806.290 2180.795 806.305 ;
        RECT 2169.670 805.990 2180.795 806.290 ;
        RECT 2169.670 805.320 2169.970 805.990 ;
        RECT 2180.465 805.975 2180.795 805.990 ;
        RECT 2166.000 804.720 2170.000 805.320 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2184.150 324.260 2184.470 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2184.150 324.120 2899.310 324.260 ;
        RECT 2184.150 324.060 2184.470 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2184.180 324.060 2184.440 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2184.170 614.195 2184.450 614.565 ;
        RECT 2184.240 324.350 2184.380 614.195 ;
        RECT 2184.180 324.030 2184.440 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2184.170 614.240 2184.450 614.520 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2166.000 615.000 2170.000 615.600 ;
        RECT 2169.670 614.530 2169.970 615.000 ;
        RECT 2184.145 614.530 2184.475 614.545 ;
        RECT 2169.670 614.230 2184.475 614.530 ;
        RECT 2184.145 614.215 2184.475 614.230 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3504.960 1176.150 3505.020 ;
        RECT 2170.350 3504.960 2170.670 3505.020 ;
        RECT 1175.830 3504.820 2170.670 3504.960 ;
        RECT 1175.830 3504.760 1176.150 3504.820 ;
        RECT 2170.350 3504.760 2170.670 3504.820 ;
      LAYER via ;
        RECT 1175.860 3504.760 1176.120 3505.020 ;
        RECT 2170.380 3504.760 2170.640 3505.020 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3505.050 1176.060 3517.600 ;
        RECT 1175.860 3504.730 1176.120 3505.050 ;
        RECT 2170.380 3504.730 2170.640 3505.050 ;
        RECT 2170.440 817.885 2170.580 3504.730 ;
        RECT 2170.370 817.515 2170.650 817.885 ;
      LAYER via2 ;
        RECT 2170.370 817.560 2170.650 817.840 ;
      LAYER met3 ;
        RECT 2170.345 817.850 2170.675 817.865 ;
        RECT 2169.670 817.550 2170.675 817.850 ;
        RECT 2169.670 815.520 2169.970 817.550 ;
        RECT 2170.345 817.535 2170.675 817.550 ;
        RECT 2166.000 814.920 2170.000 815.520 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3503.940 851.850 3504.000 ;
        RECT 2170.810 3503.940 2171.130 3504.000 ;
        RECT 851.530 3503.800 2171.130 3503.940 ;
        RECT 851.530 3503.740 851.850 3503.800 ;
        RECT 2170.810 3503.740 2171.130 3503.800 ;
      LAYER via ;
        RECT 851.560 3503.740 851.820 3504.000 ;
        RECT 2170.840 3503.740 2171.100 3504.000 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3504.030 851.760 3517.600 ;
        RECT 851.560 3503.710 851.820 3504.030 ;
        RECT 2170.840 3503.710 2171.100 3504.030 ;
        RECT 2170.900 828.085 2171.040 3503.710 ;
        RECT 2170.830 827.715 2171.110 828.085 ;
      LAYER via2 ;
        RECT 2170.830 827.760 2171.110 828.040 ;
      LAYER met3 ;
        RECT 2170.805 828.050 2171.135 828.065 ;
        RECT 2169.670 827.750 2171.135 828.050 ;
        RECT 2169.670 825.720 2169.970 827.750 ;
        RECT 2170.805 827.735 2171.135 827.750 ;
        RECT 2166.000 825.120 2170.000 825.720 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.260 527.550 3503.320 ;
        RECT 2171.730 3503.260 2172.050 3503.320 ;
        RECT 527.230 3503.120 2172.050 3503.260 ;
        RECT 527.230 3503.060 527.550 3503.120 ;
        RECT 2171.730 3503.060 2172.050 3503.120 ;
      LAYER via ;
        RECT 527.260 3503.060 527.520 3503.320 ;
        RECT 2171.760 3503.060 2172.020 3503.320 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.350 527.460 3517.600 ;
        RECT 527.260 3503.030 527.520 3503.350 ;
        RECT 2171.760 3503.030 2172.020 3503.350 ;
        RECT 2171.820 838.965 2171.960 3503.030 ;
        RECT 2171.750 838.595 2172.030 838.965 ;
      LAYER via2 ;
        RECT 2171.750 838.640 2172.030 838.920 ;
      LAYER met3 ;
        RECT 2171.725 838.930 2172.055 838.945 ;
        RECT 2169.670 838.630 2172.055 838.930 ;
        RECT 2169.670 836.600 2169.970 838.630 ;
        RECT 2171.725 838.615 2172.055 838.630 ;
        RECT 2166.000 836.000 2170.000 836.600 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.240 202.790 3502.300 ;
        RECT 2172.190 3502.240 2172.510 3502.300 ;
        RECT 202.470 3502.100 2172.510 3502.240 ;
        RECT 202.470 3502.040 202.790 3502.100 ;
        RECT 2172.190 3502.040 2172.510 3502.100 ;
      LAYER via ;
        RECT 202.500 3502.040 202.760 3502.300 ;
        RECT 2172.220 3502.040 2172.480 3502.300 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.330 202.700 3517.600 ;
        RECT 202.500 3502.010 202.760 3502.330 ;
        RECT 2172.220 3502.010 2172.480 3502.330 ;
        RECT 2172.280 848.485 2172.420 3502.010 ;
        RECT 2172.210 848.115 2172.490 848.485 ;
      LAYER via2 ;
        RECT 2172.210 848.160 2172.490 848.440 ;
      LAYER met3 ;
        RECT 2172.185 848.450 2172.515 848.465 ;
        RECT 2169.670 848.150 2172.515 848.450 ;
        RECT 2169.670 846.800 2169.970 848.150 ;
        RECT 2172.185 848.135 2172.515 848.150 ;
        RECT 2166.000 846.200 2170.000 846.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.930 3408.740 19.250 3408.800 ;
        RECT 2172.650 3408.740 2172.970 3408.800 ;
        RECT 18.930 3408.600 2172.970 3408.740 ;
        RECT 18.930 3408.540 19.250 3408.600 ;
        RECT 2172.650 3408.540 2172.970 3408.600 ;
      LAYER via ;
        RECT 18.960 3408.540 19.220 3408.800 ;
        RECT 2172.680 3408.540 2172.940 3408.800 ;
      LAYER met2 ;
        RECT 18.950 3411.035 19.230 3411.405 ;
        RECT 19.020 3408.830 19.160 3411.035 ;
        RECT 18.960 3408.510 19.220 3408.830 ;
        RECT 2172.680 3408.510 2172.940 3408.830 ;
        RECT 2172.740 860.045 2172.880 3408.510 ;
        RECT 2172.670 859.675 2172.950 860.045 ;
      LAYER via2 ;
        RECT 18.950 3411.080 19.230 3411.360 ;
        RECT 2172.670 859.720 2172.950 860.000 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 18.925 3411.370 19.255 3411.385 ;
        RECT -4.800 3411.070 19.255 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 18.925 3411.055 19.255 3411.070 ;
        RECT 2172.645 860.010 2172.975 860.025 ;
        RECT 2169.670 859.710 2172.975 860.010 ;
        RECT 2169.670 857.680 2169.970 859.710 ;
        RECT 2172.645 859.695 2172.975 859.710 ;
        RECT 2166.000 857.080 2170.000 857.680 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 3119.060 15.570 3119.120 ;
        RECT 2171.270 3119.060 2171.590 3119.120 ;
        RECT 15.250 3118.920 2171.590 3119.060 ;
        RECT 15.250 3118.860 15.570 3118.920 ;
        RECT 2171.270 3118.860 2171.590 3118.920 ;
      LAYER via ;
        RECT 15.280 3118.860 15.540 3119.120 ;
        RECT 2171.300 3118.860 2171.560 3119.120 ;
      LAYER met2 ;
        RECT 15.270 3124.075 15.550 3124.445 ;
        RECT 15.340 3119.150 15.480 3124.075 ;
        RECT 15.280 3118.830 15.540 3119.150 ;
        RECT 2171.300 3118.830 2171.560 3119.150 ;
        RECT 2171.360 869.565 2171.500 3118.830 ;
        RECT 2171.290 869.195 2171.570 869.565 ;
      LAYER via2 ;
        RECT 15.270 3124.120 15.550 3124.400 ;
        RECT 2171.290 869.240 2171.570 869.520 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 15.245 3124.410 15.575 3124.425 ;
        RECT -4.800 3124.110 15.575 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 15.245 3124.095 15.575 3124.110 ;
        RECT 2171.265 869.530 2171.595 869.545 ;
        RECT 2169.670 869.230 2171.595 869.530 ;
        RECT 2169.670 867.880 2169.970 869.230 ;
        RECT 2171.265 869.215 2171.595 869.230 ;
        RECT 2166.000 867.280 2170.000 867.880 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 1005.620 19.710 1005.680 ;
        RECT 2182.770 1005.620 2183.090 1005.680 ;
        RECT 19.390 1005.480 2183.090 1005.620 ;
        RECT 19.390 1005.420 19.710 1005.480 ;
        RECT 2182.770 1005.420 2183.090 1005.480 ;
      LAYER via ;
        RECT 19.420 1005.420 19.680 1005.680 ;
        RECT 2182.800 1005.420 2183.060 1005.680 ;
      LAYER met2 ;
        RECT 19.410 2836.435 19.690 2836.805 ;
        RECT 19.480 1005.710 19.620 2836.435 ;
        RECT 19.420 1005.390 19.680 1005.710 ;
        RECT 2182.800 1005.390 2183.060 1005.710 ;
        RECT 2182.860 881.125 2183.000 1005.390 ;
        RECT 2182.790 880.755 2183.070 881.125 ;
      LAYER via2 ;
        RECT 19.410 2836.480 19.690 2836.760 ;
        RECT 2182.790 880.800 2183.070 881.080 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 19.385 2836.770 19.715 2836.785 ;
        RECT -4.800 2836.470 19.715 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 19.385 2836.455 19.715 2836.470 ;
        RECT 2182.765 881.090 2183.095 881.105 ;
        RECT 2169.670 880.790 2183.095 881.090 ;
        RECT 2169.670 878.760 2169.970 880.790 ;
        RECT 2182.765 880.775 2183.095 880.790 ;
        RECT 2166.000 878.160 2170.000 878.760 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 1005.960 20.630 1006.020 ;
        RECT 2183.230 1005.960 2183.550 1006.020 ;
        RECT 20.310 1005.820 2183.550 1005.960 ;
        RECT 20.310 1005.760 20.630 1005.820 ;
        RECT 2183.230 1005.760 2183.550 1005.820 ;
      LAYER via ;
        RECT 20.340 1005.760 20.600 1006.020 ;
        RECT 2183.260 1005.760 2183.520 1006.020 ;
      LAYER met2 ;
        RECT 20.330 2549.475 20.610 2549.845 ;
        RECT 20.400 1006.050 20.540 2549.475 ;
        RECT 20.340 1005.730 20.600 1006.050 ;
        RECT 2183.260 1005.730 2183.520 1006.050 ;
        RECT 2183.320 889.965 2183.460 1005.730 ;
        RECT 2183.250 889.595 2183.530 889.965 ;
      LAYER via2 ;
        RECT 20.330 2549.520 20.610 2549.800 ;
        RECT 2183.250 889.640 2183.530 889.920 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 20.305 2549.810 20.635 2549.825 ;
        RECT -4.800 2549.510 20.635 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 20.305 2549.495 20.635 2549.510 ;
        RECT 2183.225 889.930 2183.555 889.945 ;
        RECT 2169.670 889.630 2183.555 889.930 ;
        RECT 2169.670 888.960 2169.970 889.630 ;
        RECT 2183.225 889.615 2183.555 889.630 ;
        RECT 2166.000 888.360 2170.000 888.960 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 2256.820 16.490 2256.880 ;
        RECT 1306.470 2256.820 1306.790 2256.880 ;
        RECT 16.170 2256.680 1306.790 2256.820 ;
        RECT 16.170 2256.620 16.490 2256.680 ;
        RECT 1306.470 2256.620 1306.790 2256.680 ;
        RECT 1306.470 2235.400 1306.790 2235.460 ;
        RECT 1329.930 2235.400 1330.250 2235.460 ;
        RECT 1306.470 2235.260 1330.250 2235.400 ;
        RECT 1306.470 2235.200 1306.790 2235.260 ;
        RECT 1329.930 2235.200 1330.250 2235.260 ;
        RECT 1329.930 2221.800 1330.250 2221.860 ;
        RECT 1330.390 2221.800 1330.710 2221.860 ;
        RECT 1329.930 2221.660 1330.710 2221.800 ;
        RECT 1329.930 2221.600 1330.250 2221.660 ;
        RECT 1330.390 2221.600 1330.710 2221.660 ;
        RECT 1330.390 2187.460 1330.710 2187.520 ;
        RECT 1330.020 2187.320 1330.710 2187.460 ;
        RECT 1330.020 2187.180 1330.160 2187.320 ;
        RECT 1330.390 2187.260 1330.710 2187.320 ;
        RECT 1329.930 2186.920 1330.250 2187.180 ;
        RECT 1329.010 2149.380 1329.330 2149.440 ;
        RECT 1330.390 2149.380 1330.710 2149.440 ;
        RECT 1329.010 2149.240 1330.710 2149.380 ;
        RECT 1329.010 2149.180 1329.330 2149.240 ;
        RECT 1330.390 2149.180 1330.710 2149.240 ;
        RECT 1329.010 2125.920 1329.330 2125.980 ;
        RECT 1329.930 2125.920 1330.250 2125.980 ;
        RECT 1329.010 2125.780 1330.250 2125.920 ;
        RECT 1329.010 2125.720 1329.330 2125.780 ;
        RECT 1329.930 2125.720 1330.250 2125.780 ;
        RECT 1329.930 2125.240 1330.250 2125.300 ;
        RECT 1330.850 2125.240 1331.170 2125.300 ;
        RECT 1329.930 2125.100 1331.170 2125.240 ;
        RECT 1329.930 2125.040 1330.250 2125.100 ;
        RECT 1330.850 2125.040 1331.170 2125.100 ;
        RECT 1328.550 2055.880 1328.870 2055.940 ;
        RECT 1329.470 2055.880 1329.790 2055.940 ;
        RECT 1328.550 2055.740 1329.790 2055.880 ;
        RECT 1328.550 2055.680 1328.870 2055.740 ;
        RECT 1329.470 2055.680 1329.790 2055.740 ;
        RECT 1328.550 2041.940 1328.870 2042.000 ;
        RECT 1330.390 2041.940 1330.710 2042.000 ;
        RECT 1328.550 2041.800 1330.710 2041.940 ;
        RECT 1328.550 2041.740 1328.870 2041.800 ;
        RECT 1330.390 2041.740 1330.710 2041.800 ;
        RECT 1330.850 1963.060 1331.170 1963.120 ;
        RECT 2180.930 1963.060 2181.250 1963.120 ;
        RECT 1330.850 1962.920 2181.250 1963.060 ;
        RECT 1330.850 1962.860 1331.170 1962.920 ;
        RECT 2180.930 1962.860 2181.250 1962.920 ;
      LAYER via ;
        RECT 16.200 2256.620 16.460 2256.880 ;
        RECT 1306.500 2256.620 1306.760 2256.880 ;
        RECT 1306.500 2235.200 1306.760 2235.460 ;
        RECT 1329.960 2235.200 1330.220 2235.460 ;
        RECT 1329.960 2221.600 1330.220 2221.860 ;
        RECT 1330.420 2221.600 1330.680 2221.860 ;
        RECT 1330.420 2187.260 1330.680 2187.520 ;
        RECT 1329.960 2186.920 1330.220 2187.180 ;
        RECT 1329.040 2149.180 1329.300 2149.440 ;
        RECT 1330.420 2149.180 1330.680 2149.440 ;
        RECT 1329.040 2125.720 1329.300 2125.980 ;
        RECT 1329.960 2125.720 1330.220 2125.980 ;
        RECT 1329.960 2125.040 1330.220 2125.300 ;
        RECT 1330.880 2125.040 1331.140 2125.300 ;
        RECT 1328.580 2055.680 1328.840 2055.940 ;
        RECT 1329.500 2055.680 1329.760 2055.940 ;
        RECT 1328.580 2041.740 1328.840 2042.000 ;
        RECT 1330.420 2041.740 1330.680 2042.000 ;
        RECT 1330.880 1962.860 1331.140 1963.120 ;
        RECT 2180.960 1962.860 2181.220 1963.120 ;
      LAYER met2 ;
        RECT 16.190 2261.835 16.470 2262.205 ;
        RECT 16.260 2256.910 16.400 2261.835 ;
        RECT 16.200 2256.590 16.460 2256.910 ;
        RECT 1306.500 2256.590 1306.760 2256.910 ;
        RECT 1306.560 2235.490 1306.700 2256.590 ;
        RECT 1306.500 2235.170 1306.760 2235.490 ;
        RECT 1329.960 2235.170 1330.220 2235.490 ;
        RECT 1330.020 2221.890 1330.160 2235.170 ;
        RECT 1329.960 2221.570 1330.220 2221.890 ;
        RECT 1330.420 2221.570 1330.680 2221.890 ;
        RECT 1330.480 2187.550 1330.620 2221.570 ;
        RECT 1330.420 2187.230 1330.680 2187.550 ;
        RECT 1329.960 2186.890 1330.220 2187.210 ;
        RECT 1330.020 2173.690 1330.160 2186.890 ;
        RECT 1330.020 2173.550 1330.620 2173.690 ;
        RECT 1330.480 2149.470 1330.620 2173.550 ;
        RECT 1329.040 2149.150 1329.300 2149.470 ;
        RECT 1330.420 2149.150 1330.680 2149.470 ;
        RECT 1329.100 2126.010 1329.240 2149.150 ;
        RECT 1329.040 2125.690 1329.300 2126.010 ;
        RECT 1329.960 2125.690 1330.220 2126.010 ;
        RECT 1330.020 2125.330 1330.160 2125.690 ;
        RECT 1329.960 2125.010 1330.220 2125.330 ;
        RECT 1330.880 2125.010 1331.140 2125.330 ;
        RECT 1330.940 2077.245 1331.080 2125.010 ;
        RECT 1329.950 2077.130 1330.230 2077.245 ;
        RECT 1329.560 2076.990 1330.230 2077.130 ;
        RECT 1329.560 2055.970 1329.700 2076.990 ;
        RECT 1329.950 2076.875 1330.230 2076.990 ;
        RECT 1330.870 2076.875 1331.150 2077.245 ;
        RECT 1328.580 2055.650 1328.840 2055.970 ;
        RECT 1329.500 2055.650 1329.760 2055.970 ;
        RECT 1328.640 2042.030 1328.780 2055.650 ;
        RECT 1328.580 2041.710 1328.840 2042.030 ;
        RECT 1330.420 2041.710 1330.680 2042.030 ;
        RECT 1330.480 1994.170 1330.620 2041.710 ;
        RECT 1330.480 1994.030 1331.080 1994.170 ;
        RECT 1330.940 1963.150 1331.080 1994.030 ;
        RECT 1330.880 1962.830 1331.140 1963.150 ;
        RECT 2180.960 1962.830 2181.220 1963.150 ;
        RECT 2181.020 901.525 2181.160 1962.830 ;
        RECT 2180.950 901.155 2181.230 901.525 ;
      LAYER via2 ;
        RECT 16.190 2261.880 16.470 2262.160 ;
        RECT 1329.950 2076.920 1330.230 2077.200 ;
        RECT 1330.870 2076.920 1331.150 2077.200 ;
        RECT 2180.950 901.200 2181.230 901.480 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 16.165 2262.170 16.495 2262.185 ;
        RECT -4.800 2261.870 16.495 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 16.165 2261.855 16.495 2261.870 ;
        RECT 1329.925 2077.210 1330.255 2077.225 ;
        RECT 1330.845 2077.210 1331.175 2077.225 ;
        RECT 1329.925 2076.910 1331.175 2077.210 ;
        RECT 1329.925 2076.895 1330.255 2076.910 ;
        RECT 1330.845 2076.895 1331.175 2076.910 ;
        RECT 2180.925 901.490 2181.255 901.505 ;
        RECT 2169.670 901.190 2181.255 901.490 ;
        RECT 2169.670 899.840 2169.970 901.190 ;
        RECT 2180.925 901.175 2181.255 901.190 ;
        RECT 2166.000 899.240 2170.000 899.840 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.870 1052.200 14.190 1052.260 ;
        RECT 15.250 1052.200 15.570 1052.260 ;
        RECT 13.870 1052.060 15.570 1052.200 ;
        RECT 13.870 1052.000 14.190 1052.060 ;
        RECT 15.250 1052.000 15.570 1052.060 ;
        RECT 13.870 1005.280 14.190 1005.340 ;
        RECT 2183.690 1005.280 2184.010 1005.340 ;
        RECT 13.870 1005.140 2184.010 1005.280 ;
        RECT 13.870 1005.080 14.190 1005.140 ;
        RECT 2183.690 1005.080 2184.010 1005.140 ;
      LAYER via ;
        RECT 13.900 1052.000 14.160 1052.260 ;
        RECT 15.280 1052.000 15.540 1052.260 ;
        RECT 13.900 1005.080 14.160 1005.340 ;
        RECT 2183.720 1005.080 2183.980 1005.340 ;
      LAYER met2 ;
        RECT 15.270 1974.875 15.550 1975.245 ;
        RECT 15.340 1052.290 15.480 1974.875 ;
        RECT 13.900 1051.970 14.160 1052.290 ;
        RECT 15.280 1051.970 15.540 1052.290 ;
        RECT 13.960 1005.370 14.100 1051.970 ;
        RECT 13.900 1005.050 14.160 1005.370 ;
        RECT 2183.720 1005.050 2183.980 1005.370 ;
        RECT 2183.780 910.365 2183.920 1005.050 ;
        RECT 2183.710 909.995 2183.990 910.365 ;
      LAYER via2 ;
        RECT 15.270 1974.920 15.550 1975.200 ;
        RECT 2183.710 910.040 2183.990 910.320 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.245 1975.210 15.575 1975.225 ;
        RECT -4.800 1974.910 15.575 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.245 1974.895 15.575 1974.910 ;
        RECT 2183.685 910.330 2184.015 910.345 ;
        RECT 2169.670 910.040 2184.015 910.330 ;
        RECT 2166.000 910.030 2184.015 910.040 ;
        RECT 2166.000 909.440 2170.000 910.030 ;
        RECT 2183.685 910.015 2184.015 910.030 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2184.610 558.860 2184.930 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2184.610 558.720 2899.310 558.860 ;
        RECT 2184.610 558.660 2184.930 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2184.640 558.660 2184.900 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2184.630 622.355 2184.910 622.725 ;
        RECT 2184.700 558.950 2184.840 622.355 ;
        RECT 2184.640 558.630 2184.900 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2184.630 622.400 2184.910 622.680 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2166.000 625.200 2170.000 625.800 ;
        RECT 2169.670 622.690 2169.970 625.200 ;
        RECT 2184.605 622.690 2184.935 622.705 ;
        RECT 2169.670 622.390 2184.935 622.690 ;
        RECT 2184.605 622.375 2184.935 622.390 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 14.790 1683.920 15.110 1683.980 ;
        RECT 2173.570 1683.920 2173.890 1683.980 ;
        RECT 14.790 1683.780 2173.890 1683.920 ;
        RECT 14.790 1683.720 15.110 1683.780 ;
        RECT 2173.570 1683.720 2173.890 1683.780 ;
      LAYER via ;
        RECT 14.820 1683.720 15.080 1683.980 ;
        RECT 2173.600 1683.720 2173.860 1683.980 ;
      LAYER met2 ;
        RECT 14.810 1687.235 15.090 1687.605 ;
        RECT 14.880 1684.010 15.020 1687.235 ;
        RECT 14.820 1683.690 15.080 1684.010 ;
        RECT 2173.600 1683.690 2173.860 1684.010 ;
        RECT 2173.660 923.285 2173.800 1683.690 ;
        RECT 2173.590 922.915 2173.870 923.285 ;
      LAYER via2 ;
        RECT 14.810 1687.280 15.090 1687.560 ;
        RECT 2173.590 922.960 2173.870 923.240 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 14.785 1687.570 15.115 1687.585 ;
        RECT -4.800 1687.270 15.115 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 14.785 1687.255 15.115 1687.270 ;
        RECT 2173.565 923.250 2173.895 923.265 ;
        RECT 2169.670 922.950 2173.895 923.250 ;
        RECT 2169.670 920.920 2169.970 922.950 ;
        RECT 2173.565 922.935 2173.895 922.950 ;
        RECT 2166.000 920.320 2170.000 920.920 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 14.790 1470.060 15.110 1470.120 ;
        RECT 2174.030 1470.060 2174.350 1470.120 ;
        RECT 14.790 1469.920 2174.350 1470.060 ;
        RECT 14.790 1469.860 15.110 1469.920 ;
        RECT 2174.030 1469.860 2174.350 1469.920 ;
      LAYER via ;
        RECT 14.820 1469.860 15.080 1470.120 ;
        RECT 2174.060 1469.860 2174.320 1470.120 ;
      LAYER met2 ;
        RECT 14.810 1471.675 15.090 1472.045 ;
        RECT 14.880 1470.150 15.020 1471.675 ;
        RECT 14.820 1469.830 15.080 1470.150 ;
        RECT 2174.060 1469.830 2174.320 1470.150 ;
        RECT 2174.120 931.445 2174.260 1469.830 ;
        RECT 2174.050 931.075 2174.330 931.445 ;
      LAYER via2 ;
        RECT 14.810 1471.720 15.090 1472.000 ;
        RECT 2174.050 931.120 2174.330 931.400 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 14.785 1472.010 15.115 1472.025 ;
        RECT -4.800 1471.710 15.115 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 14.785 1471.695 15.115 1471.710 ;
        RECT 2174.025 931.410 2174.355 931.425 ;
        RECT 2169.670 931.120 2174.355 931.410 ;
        RECT 2166.000 931.110 2174.355 931.120 ;
        RECT 2166.000 930.520 2170.000 931.110 ;
        RECT 2174.025 931.095 2174.355 931.110 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 14.330 1256.200 14.650 1256.260 ;
        RECT 2174.490 1256.200 2174.810 1256.260 ;
        RECT 14.330 1256.060 2174.810 1256.200 ;
        RECT 14.330 1256.000 14.650 1256.060 ;
        RECT 2174.490 1256.000 2174.810 1256.060 ;
      LAYER via ;
        RECT 14.360 1256.000 14.620 1256.260 ;
        RECT 2174.520 1256.000 2174.780 1256.260 ;
      LAYER met2 ;
        RECT 14.350 1256.115 14.630 1256.485 ;
        RECT 14.360 1255.970 14.620 1256.115 ;
        RECT 2174.520 1255.970 2174.780 1256.290 ;
        RECT 2174.580 944.365 2174.720 1255.970 ;
        RECT 2174.510 943.995 2174.790 944.365 ;
      LAYER via2 ;
        RECT 14.350 1256.160 14.630 1256.440 ;
        RECT 2174.510 944.040 2174.790 944.320 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 14.325 1256.450 14.655 1256.465 ;
        RECT -4.800 1256.150 14.655 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 14.325 1256.135 14.655 1256.150 ;
        RECT 2174.485 944.330 2174.815 944.345 ;
        RECT 2169.670 944.030 2174.815 944.330 ;
        RECT 2169.670 942.000 2169.970 944.030 ;
        RECT 2174.485 944.015 2174.815 944.030 ;
        RECT 2166.000 941.400 2170.000 942.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 1035.200 15.570 1035.260 ;
        RECT 2174.950 1035.200 2175.270 1035.260 ;
        RECT 15.250 1035.060 2175.270 1035.200 ;
        RECT 15.250 1035.000 15.570 1035.060 ;
        RECT 2174.950 1035.000 2175.270 1035.060 ;
      LAYER via ;
        RECT 15.280 1035.000 15.540 1035.260 ;
        RECT 2174.980 1035.000 2175.240 1035.260 ;
      LAYER met2 ;
        RECT 15.270 1040.555 15.550 1040.925 ;
        RECT 15.340 1035.290 15.480 1040.555 ;
        RECT 15.280 1034.970 15.540 1035.290 ;
        RECT 2174.980 1034.970 2175.240 1035.290 ;
        RECT 2175.040 951.165 2175.180 1034.970 ;
        RECT 2174.970 950.795 2175.250 951.165 ;
      LAYER via2 ;
        RECT 15.270 1040.600 15.550 1040.880 ;
        RECT 2174.970 950.840 2175.250 951.120 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 15.245 1040.890 15.575 1040.905 ;
        RECT -4.800 1040.590 15.575 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 15.245 1040.575 15.575 1040.590 ;
        RECT 2166.000 951.600 2170.000 952.200 ;
        RECT 2169.670 951.130 2169.970 951.600 ;
        RECT 2174.945 951.130 2175.275 951.145 ;
        RECT 2169.670 950.830 2175.275 951.130 ;
        RECT 2174.945 950.815 2175.275 950.830 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.870 999.160 14.190 999.220 ;
        RECT 2181.390 999.160 2181.710 999.220 ;
        RECT 13.870 999.020 2181.710 999.160 ;
        RECT 13.870 998.960 14.190 999.020 ;
        RECT 2181.390 998.960 2181.710 999.020 ;
      LAYER via ;
        RECT 13.900 998.960 14.160 999.220 ;
        RECT 2181.420 998.960 2181.680 999.220 ;
      LAYER met2 ;
        RECT 13.900 998.930 14.160 999.250 ;
        RECT 2181.420 998.930 2181.680 999.250 ;
        RECT 13.960 825.365 14.100 998.930 ;
        RECT 2181.480 965.445 2181.620 998.930 ;
        RECT 2181.410 965.075 2181.690 965.445 ;
        RECT 13.890 824.995 14.170 825.365 ;
      LAYER via2 ;
        RECT 2181.410 965.120 2181.690 965.400 ;
        RECT 13.890 825.040 14.170 825.320 ;
      LAYER met3 ;
        RECT 2181.385 965.410 2181.715 965.425 ;
        RECT 2169.670 965.110 2181.715 965.410 ;
        RECT 2169.670 963.080 2169.970 965.110 ;
        RECT 2181.385 965.095 2181.715 965.110 ;
        RECT 2166.000 962.480 2170.000 963.080 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 13.865 825.330 14.195 825.345 ;
        RECT -4.800 825.030 14.195 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 13.865 825.015 14.195 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 603.060 16.490 603.120 ;
        RECT 2182.310 603.060 2182.630 603.120 ;
        RECT 16.170 602.920 2182.630 603.060 ;
        RECT 16.170 602.860 16.490 602.920 ;
        RECT 2182.310 602.860 2182.630 602.920 ;
      LAYER via ;
        RECT 16.200 602.860 16.460 603.120 ;
        RECT 2182.340 602.860 2182.600 603.120 ;
      LAYER met2 ;
        RECT 2182.330 969.835 2182.610 970.205 ;
        RECT 16.190 610.115 16.470 610.485 ;
        RECT 16.260 603.150 16.400 610.115 ;
        RECT 2182.400 603.150 2182.540 969.835 ;
        RECT 16.200 602.830 16.460 603.150 ;
        RECT 2182.340 602.830 2182.600 603.150 ;
      LAYER via2 ;
        RECT 2182.330 969.880 2182.610 970.160 ;
        RECT 16.190 610.160 16.470 610.440 ;
      LAYER met3 ;
        RECT 2166.000 972.680 2170.000 973.280 ;
        RECT 2169.670 970.170 2169.970 972.680 ;
        RECT 2182.305 970.170 2182.635 970.185 ;
        RECT 2169.670 969.870 2182.635 970.170 ;
        RECT 2182.305 969.855 2182.635 969.870 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 16.165 610.450 16.495 610.465 ;
        RECT -4.800 610.150 16.495 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 16.165 610.135 16.495 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 400.080 16.030 400.140 ;
        RECT 2181.850 400.080 2182.170 400.140 ;
        RECT 15.710 399.940 2182.170 400.080 ;
        RECT 15.710 399.880 16.030 399.940 ;
        RECT 2181.850 399.880 2182.170 399.940 ;
      LAYER via ;
        RECT 15.740 399.880 16.000 400.140 ;
        RECT 2181.880 399.880 2182.140 400.140 ;
      LAYER met2 ;
        RECT 2181.870 980.715 2182.150 981.085 ;
        RECT 2181.940 400.170 2182.080 980.715 ;
        RECT 15.740 399.850 16.000 400.170 ;
        RECT 2181.880 399.850 2182.140 400.170 ;
        RECT 15.800 394.925 15.940 399.850 ;
        RECT 15.730 394.555 16.010 394.925 ;
      LAYER via2 ;
        RECT 2181.870 980.760 2182.150 981.040 ;
        RECT 15.730 394.600 16.010 394.880 ;
      LAYER met3 ;
        RECT 2166.000 983.560 2170.000 984.160 ;
        RECT 2169.670 981.050 2169.970 983.560 ;
        RECT 2181.845 981.050 2182.175 981.065 ;
        RECT 2169.670 980.750 2182.175 981.050 ;
        RECT 2181.845 980.735 2182.175 980.750 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 15.705 394.890 16.035 394.905 ;
        RECT -4.800 394.590 16.035 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 15.705 394.575 16.035 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2181.390 964.820 2181.710 964.880 ;
        RECT 2184.150 964.820 2184.470 964.880 ;
        RECT 2181.390 964.680 2184.470 964.820 ;
        RECT 2181.390 964.620 2181.710 964.680 ;
        RECT 2184.150 964.620 2184.470 964.680 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 2181.390 179.420 2181.710 179.480 ;
        RECT 17.090 179.280 2181.710 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 2181.390 179.220 2181.710 179.280 ;
      LAYER via ;
        RECT 2181.420 964.620 2181.680 964.880 ;
        RECT 2184.180 964.620 2184.440 964.880 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 2181.420 179.220 2181.680 179.480 ;
      LAYER met2 ;
        RECT 2184.170 994.315 2184.450 994.685 ;
        RECT 2184.240 964.910 2184.380 994.315 ;
        RECT 2181.420 964.590 2181.680 964.910 ;
        RECT 2184.180 964.590 2184.440 964.910 ;
        RECT 2181.480 179.510 2181.620 964.590 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 2181.420 179.190 2181.680 179.510 ;
      LAYER via2 ;
        RECT 2184.170 994.360 2184.450 994.640 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 2184.145 994.650 2184.475 994.665 ;
        RECT 2169.670 994.360 2184.475 994.650 ;
        RECT 2166.000 994.350 2184.475 994.360 ;
        RECT 2166.000 993.760 2170.000 994.350 ;
        RECT 2184.145 994.335 2184.475 994.350 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.470 641.480 2180.790 641.540 ;
        RECT 2903.130 641.480 2903.450 641.540 ;
        RECT 2180.470 641.340 2903.450 641.480 ;
        RECT 2180.470 641.280 2180.790 641.340 ;
        RECT 2903.130 641.280 2903.450 641.340 ;
      LAYER via ;
        RECT 2180.500 641.280 2180.760 641.540 ;
        RECT 2903.160 641.280 2903.420 641.540 ;
      LAYER met2 ;
        RECT 2903.150 791.675 2903.430 792.045 ;
        RECT 2903.220 641.570 2903.360 791.675 ;
        RECT 2180.500 641.250 2180.760 641.570 ;
        RECT 2903.160 641.250 2903.420 641.570 ;
        RECT 2180.560 639.045 2180.700 641.250 ;
        RECT 2180.490 638.675 2180.770 639.045 ;
      LAYER via2 ;
        RECT 2903.150 791.720 2903.430 792.000 ;
        RECT 2180.490 638.720 2180.770 639.000 ;
      LAYER met3 ;
        RECT 2903.125 792.010 2903.455 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2903.125 791.710 2924.800 792.010 ;
        RECT 2903.125 791.695 2903.455 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2180.465 639.010 2180.795 639.025 ;
        RECT 2169.670 638.710 2180.795 639.010 ;
        RECT 2169.670 636.680 2169.970 638.710 ;
        RECT 2180.465 638.695 2180.795 638.710 ;
        RECT 2166.000 636.080 2170.000 636.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 648.620 2187.230 648.680 ;
        RECT 2900.370 648.620 2900.690 648.680 ;
        RECT 2186.910 648.480 2900.690 648.620 ;
        RECT 2186.910 648.420 2187.230 648.480 ;
        RECT 2900.370 648.420 2900.690 648.480 ;
      LAYER via ;
        RECT 2186.940 648.420 2187.200 648.680 ;
        RECT 2900.400 648.420 2900.660 648.680 ;
      LAYER met2 ;
        RECT 2900.390 1026.275 2900.670 1026.645 ;
        RECT 2900.460 648.710 2900.600 1026.275 ;
        RECT 2186.940 648.390 2187.200 648.710 ;
        RECT 2900.400 648.390 2900.660 648.710 ;
        RECT 2187.000 647.885 2187.140 648.390 ;
        RECT 2186.930 647.515 2187.210 647.885 ;
      LAYER via2 ;
        RECT 2900.390 1026.320 2900.670 1026.600 ;
        RECT 2186.930 647.560 2187.210 647.840 ;
      LAYER met3 ;
        RECT 2900.365 1026.610 2900.695 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2900.365 1026.310 2924.800 1026.610 ;
        RECT 2900.365 1026.295 2900.695 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2186.905 647.850 2187.235 647.865 ;
        RECT 2169.670 647.550 2187.235 647.850 ;
        RECT 2169.670 646.880 2169.970 647.550 ;
        RECT 2186.905 647.535 2187.235 647.550 ;
        RECT 2166.000 646.280 2170.000 646.880 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2184.150 662.220 2184.470 662.280 ;
        RECT 2900.830 662.220 2901.150 662.280 ;
        RECT 2184.150 662.080 2901.150 662.220 ;
        RECT 2184.150 662.020 2184.470 662.080 ;
        RECT 2900.830 662.020 2901.150 662.080 ;
      LAYER via ;
        RECT 2184.180 662.020 2184.440 662.280 ;
        RECT 2900.860 662.020 2901.120 662.280 ;
      LAYER met2 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
        RECT 2900.920 662.310 2901.060 1260.875 ;
        RECT 2184.180 661.990 2184.440 662.310 ;
        RECT 2900.860 661.990 2901.120 662.310 ;
        RECT 2184.240 660.125 2184.380 661.990 ;
        RECT 2184.170 659.755 2184.450 660.125 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
        RECT 2184.170 659.800 2184.450 660.080 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2184.145 660.090 2184.475 660.105 ;
        RECT 2169.670 659.790 2184.475 660.090 ;
        RECT 2169.670 657.760 2169.970 659.790 ;
        RECT 2184.145 659.775 2184.475 659.790 ;
        RECT 2166.000 657.160 2170.000 657.760 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 669.360 2187.230 669.420 ;
        RECT 2904.050 669.360 2904.370 669.420 ;
        RECT 2186.910 669.220 2904.370 669.360 ;
        RECT 2186.910 669.160 2187.230 669.220 ;
        RECT 2904.050 669.160 2904.370 669.220 ;
      LAYER via ;
        RECT 2186.940 669.160 2187.200 669.420 ;
        RECT 2904.080 669.160 2904.340 669.420 ;
      LAYER met2 ;
        RECT 2904.070 1495.475 2904.350 1495.845 ;
        RECT 2904.140 669.450 2904.280 1495.475 ;
        RECT 2186.940 669.130 2187.200 669.450 ;
        RECT 2904.080 669.130 2904.340 669.450 ;
        RECT 2187.000 668.285 2187.140 669.130 ;
        RECT 2186.930 667.915 2187.210 668.285 ;
      LAYER via2 ;
        RECT 2904.070 1495.520 2904.350 1495.800 ;
        RECT 2186.930 667.960 2187.210 668.240 ;
      LAYER met3 ;
        RECT 2904.045 1495.810 2904.375 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2904.045 1495.510 2924.800 1495.810 ;
        RECT 2904.045 1495.495 2904.375 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2186.905 668.250 2187.235 668.265 ;
        RECT 2169.670 667.960 2187.235 668.250 ;
        RECT 2166.000 667.950 2187.235 667.960 ;
        RECT 2166.000 667.360 2170.000 667.950 ;
        RECT 2186.905 667.935 2187.235 667.950 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2524.090 1725.400 2524.410 1725.460 ;
        RECT 2899.910 1725.400 2900.230 1725.460 ;
        RECT 2524.090 1725.260 2900.230 1725.400 ;
        RECT 2524.090 1725.200 2524.410 1725.260 ;
        RECT 2899.910 1725.200 2900.230 1725.260 ;
        RECT 2521.790 1593.820 2522.110 1593.880 ;
        RECT 2522.250 1593.820 2522.570 1593.880 ;
        RECT 2521.790 1593.680 2522.570 1593.820 ;
        RECT 2521.790 1593.620 2522.110 1593.680 ;
        RECT 2522.250 1593.620 2522.570 1593.680 ;
        RECT 2521.790 1546.220 2522.110 1546.280 ;
        RECT 2522.250 1546.220 2522.570 1546.280 ;
        RECT 2521.790 1546.080 2522.570 1546.220 ;
        RECT 2521.790 1546.020 2522.110 1546.080 ;
        RECT 2522.250 1546.020 2522.570 1546.080 ;
        RECT 2520.870 1545.540 2521.190 1545.600 ;
        RECT 2521.790 1545.540 2522.110 1545.600 ;
        RECT 2520.870 1545.400 2522.110 1545.540 ;
        RECT 2520.870 1545.340 2521.190 1545.400 ;
        RECT 2521.790 1545.340 2522.110 1545.400 ;
        RECT 2520.870 1497.600 2521.190 1497.660 ;
        RECT 2522.250 1497.600 2522.570 1497.660 ;
        RECT 2520.870 1497.460 2522.570 1497.600 ;
        RECT 2520.870 1497.400 2521.190 1497.460 ;
        RECT 2522.250 1497.400 2522.570 1497.460 ;
        RECT 2522.250 1490.460 2522.570 1490.520 ;
        RECT 2523.630 1490.460 2523.950 1490.520 ;
        RECT 2522.250 1490.320 2523.950 1490.460 ;
        RECT 2522.250 1490.260 2522.570 1490.320 ;
        RECT 2523.630 1490.260 2523.950 1490.320 ;
        RECT 2522.710 1442.180 2523.030 1442.240 ;
        RECT 2523.630 1442.180 2523.950 1442.240 ;
        RECT 2522.710 1442.040 2523.950 1442.180 ;
        RECT 2522.710 1441.980 2523.030 1442.040 ;
        RECT 2523.630 1441.980 2523.950 1442.040 ;
        RECT 2522.250 1393.560 2522.570 1393.620 ;
        RECT 2522.710 1393.560 2523.030 1393.620 ;
        RECT 2522.250 1393.420 2523.030 1393.560 ;
        RECT 2522.250 1393.360 2522.570 1393.420 ;
        RECT 2522.710 1393.360 2523.030 1393.420 ;
        RECT 2521.330 1304.140 2521.650 1304.200 ;
        RECT 2522.710 1304.140 2523.030 1304.200 ;
        RECT 2521.330 1304.000 2523.030 1304.140 ;
        RECT 2521.330 1303.940 2521.650 1304.000 ;
        RECT 2522.710 1303.940 2523.030 1304.000 ;
        RECT 2521.330 1269.120 2521.650 1269.180 ;
        RECT 2522.710 1269.120 2523.030 1269.180 ;
        RECT 2521.330 1268.980 2523.030 1269.120 ;
        RECT 2521.330 1268.920 2521.650 1268.980 ;
        RECT 2522.710 1268.920 2523.030 1268.980 ;
        RECT 2520.410 1255.860 2520.730 1255.920 ;
        RECT 2521.330 1255.860 2521.650 1255.920 ;
        RECT 2520.410 1255.720 2521.650 1255.860 ;
        RECT 2520.410 1255.660 2520.730 1255.720 ;
        RECT 2521.330 1255.660 2521.650 1255.720 ;
        RECT 2520.410 1207.580 2520.730 1207.640 ;
        RECT 2522.250 1207.580 2522.570 1207.640 ;
        RECT 2520.410 1207.440 2522.570 1207.580 ;
        RECT 2520.410 1207.380 2520.730 1207.440 ;
        RECT 2522.250 1207.380 2522.570 1207.440 ;
        RECT 2522.250 1173.580 2522.570 1173.640 ;
        RECT 2521.880 1173.440 2522.570 1173.580 ;
        RECT 2521.880 1172.960 2522.020 1173.440 ;
        RECT 2522.250 1173.380 2522.570 1173.440 ;
        RECT 2521.790 1172.700 2522.110 1172.960 ;
        RECT 2520.870 1158.960 2521.190 1159.020 ;
        RECT 2521.790 1158.960 2522.110 1159.020 ;
        RECT 2520.870 1158.820 2522.110 1158.960 ;
        RECT 2520.870 1158.760 2521.190 1158.820 ;
        RECT 2521.790 1158.760 2522.110 1158.820 ;
        RECT 2520.870 1111.020 2521.190 1111.080 ;
        RECT 2522.250 1111.020 2522.570 1111.080 ;
        RECT 2520.870 1110.880 2522.570 1111.020 ;
        RECT 2520.870 1110.820 2521.190 1110.880 ;
        RECT 2522.250 1110.820 2522.570 1110.880 ;
        RECT 2522.250 1077.020 2522.570 1077.080 ;
        RECT 2521.420 1076.880 2522.570 1077.020 ;
        RECT 2521.420 1076.400 2521.560 1076.880 ;
        RECT 2522.250 1076.820 2522.570 1076.880 ;
        RECT 2521.330 1076.140 2521.650 1076.400 ;
        RECT 2520.870 1028.400 2521.190 1028.460 ;
        RECT 2520.870 1028.260 2521.560 1028.400 ;
        RECT 2520.870 1028.200 2521.190 1028.260 ;
        RECT 2521.420 1028.120 2521.560 1028.260 ;
        RECT 2521.330 1027.860 2521.650 1028.120 ;
        RECT 2520.870 1014.460 2521.190 1014.520 ;
        RECT 2521.330 1014.460 2521.650 1014.520 ;
        RECT 2520.870 1014.320 2521.650 1014.460 ;
        RECT 2520.870 1014.260 2521.190 1014.320 ;
        RECT 2521.330 1014.260 2521.650 1014.320 ;
        RECT 2520.870 1006.300 2521.190 1006.360 ;
        RECT 2522.250 1006.300 2522.570 1006.360 ;
        RECT 2520.870 1006.160 2522.570 1006.300 ;
        RECT 2520.870 1006.100 2521.190 1006.160 ;
        RECT 2522.250 1006.100 2522.570 1006.160 ;
        RECT 2522.250 869.620 2522.570 869.680 ;
        RECT 2523.170 869.620 2523.490 869.680 ;
        RECT 2522.250 869.480 2523.490 869.620 ;
        RECT 2522.250 869.420 2522.570 869.480 ;
        RECT 2523.170 869.420 2523.490 869.480 ;
        RECT 2520.870 821.000 2521.190 821.060 ;
        RECT 2521.790 821.000 2522.110 821.060 ;
        RECT 2520.870 820.860 2522.110 821.000 ;
        RECT 2520.870 820.800 2521.190 820.860 ;
        RECT 2521.790 820.800 2522.110 820.860 ;
        RECT 2185.070 682.960 2185.390 683.020 ;
        RECT 2522.250 682.960 2522.570 683.020 ;
        RECT 2185.070 682.820 2522.570 682.960 ;
        RECT 2185.070 682.760 2185.390 682.820 ;
        RECT 2522.250 682.760 2522.570 682.820 ;
      LAYER via ;
        RECT 2524.120 1725.200 2524.380 1725.460 ;
        RECT 2899.940 1725.200 2900.200 1725.460 ;
        RECT 2521.820 1593.620 2522.080 1593.880 ;
        RECT 2522.280 1593.620 2522.540 1593.880 ;
        RECT 2521.820 1546.020 2522.080 1546.280 ;
        RECT 2522.280 1546.020 2522.540 1546.280 ;
        RECT 2520.900 1545.340 2521.160 1545.600 ;
        RECT 2521.820 1545.340 2522.080 1545.600 ;
        RECT 2520.900 1497.400 2521.160 1497.660 ;
        RECT 2522.280 1497.400 2522.540 1497.660 ;
        RECT 2522.280 1490.260 2522.540 1490.520 ;
        RECT 2523.660 1490.260 2523.920 1490.520 ;
        RECT 2522.740 1441.980 2523.000 1442.240 ;
        RECT 2523.660 1441.980 2523.920 1442.240 ;
        RECT 2522.280 1393.360 2522.540 1393.620 ;
        RECT 2522.740 1393.360 2523.000 1393.620 ;
        RECT 2521.360 1303.940 2521.620 1304.200 ;
        RECT 2522.740 1303.940 2523.000 1304.200 ;
        RECT 2521.360 1268.920 2521.620 1269.180 ;
        RECT 2522.740 1268.920 2523.000 1269.180 ;
        RECT 2520.440 1255.660 2520.700 1255.920 ;
        RECT 2521.360 1255.660 2521.620 1255.920 ;
        RECT 2520.440 1207.380 2520.700 1207.640 ;
        RECT 2522.280 1207.380 2522.540 1207.640 ;
        RECT 2522.280 1173.380 2522.540 1173.640 ;
        RECT 2521.820 1172.700 2522.080 1172.960 ;
        RECT 2520.900 1158.760 2521.160 1159.020 ;
        RECT 2521.820 1158.760 2522.080 1159.020 ;
        RECT 2520.900 1110.820 2521.160 1111.080 ;
        RECT 2522.280 1110.820 2522.540 1111.080 ;
        RECT 2522.280 1076.820 2522.540 1077.080 ;
        RECT 2521.360 1076.140 2521.620 1076.400 ;
        RECT 2520.900 1028.200 2521.160 1028.460 ;
        RECT 2521.360 1027.860 2521.620 1028.120 ;
        RECT 2520.900 1014.260 2521.160 1014.520 ;
        RECT 2521.360 1014.260 2521.620 1014.520 ;
        RECT 2520.900 1006.100 2521.160 1006.360 ;
        RECT 2522.280 1006.100 2522.540 1006.360 ;
        RECT 2522.280 869.420 2522.540 869.680 ;
        RECT 2523.200 869.420 2523.460 869.680 ;
        RECT 2520.900 820.800 2521.160 821.060 ;
        RECT 2521.820 820.800 2522.080 821.060 ;
        RECT 2185.100 682.760 2185.360 683.020 ;
        RECT 2522.280 682.760 2522.540 683.020 ;
      LAYER met2 ;
        RECT 2899.930 1730.075 2900.210 1730.445 ;
        RECT 2900.000 1725.490 2900.140 1730.075 ;
        RECT 2524.120 1725.170 2524.380 1725.490 ;
        RECT 2899.940 1725.170 2900.200 1725.490 ;
        RECT 2524.180 1663.010 2524.320 1725.170 ;
        RECT 2522.340 1662.870 2524.320 1663.010 ;
        RECT 2522.340 1656.210 2522.480 1662.870 ;
        RECT 2521.880 1656.070 2522.480 1656.210 ;
        RECT 2521.880 1593.910 2522.020 1656.070 ;
        RECT 2521.820 1593.590 2522.080 1593.910 ;
        RECT 2522.280 1593.590 2522.540 1593.910 ;
        RECT 2522.340 1546.310 2522.480 1593.590 ;
        RECT 2521.820 1545.990 2522.080 1546.310 ;
        RECT 2522.280 1545.990 2522.540 1546.310 ;
        RECT 2521.880 1545.630 2522.020 1545.990 ;
        RECT 2520.900 1545.310 2521.160 1545.630 ;
        RECT 2521.820 1545.310 2522.080 1545.630 ;
        RECT 2520.960 1497.690 2521.100 1545.310 ;
        RECT 2520.900 1497.370 2521.160 1497.690 ;
        RECT 2522.280 1497.370 2522.540 1497.690 ;
        RECT 2522.340 1490.550 2522.480 1497.370 ;
        RECT 2522.280 1490.230 2522.540 1490.550 ;
        RECT 2523.660 1490.230 2523.920 1490.550 ;
        RECT 2523.720 1442.270 2523.860 1490.230 ;
        RECT 2522.740 1441.950 2523.000 1442.270 ;
        RECT 2523.660 1441.950 2523.920 1442.270 ;
        RECT 2522.800 1401.210 2522.940 1441.950 ;
        RECT 2522.340 1401.070 2522.940 1401.210 ;
        RECT 2522.340 1393.650 2522.480 1401.070 ;
        RECT 2522.280 1393.330 2522.540 1393.650 ;
        RECT 2522.740 1393.330 2523.000 1393.650 ;
        RECT 2522.800 1304.765 2522.940 1393.330 ;
        RECT 2521.350 1304.395 2521.630 1304.765 ;
        RECT 2522.730 1304.395 2523.010 1304.765 ;
        RECT 2521.420 1304.230 2521.560 1304.395 ;
        RECT 2521.360 1303.910 2521.620 1304.230 ;
        RECT 2522.740 1303.910 2523.000 1304.230 ;
        RECT 2522.800 1269.210 2522.940 1303.910 ;
        RECT 2521.360 1268.890 2521.620 1269.210 ;
        RECT 2522.740 1268.890 2523.000 1269.210 ;
        RECT 2521.420 1255.950 2521.560 1268.890 ;
        RECT 2520.440 1255.630 2520.700 1255.950 ;
        RECT 2521.360 1255.630 2521.620 1255.950 ;
        RECT 2520.500 1207.670 2520.640 1255.630 ;
        RECT 2520.440 1207.350 2520.700 1207.670 ;
        RECT 2522.280 1207.350 2522.540 1207.670 ;
        RECT 2522.340 1173.670 2522.480 1207.350 ;
        RECT 2522.280 1173.350 2522.540 1173.670 ;
        RECT 2521.820 1172.670 2522.080 1172.990 ;
        RECT 2521.880 1159.050 2522.020 1172.670 ;
        RECT 2520.900 1158.730 2521.160 1159.050 ;
        RECT 2521.820 1158.730 2522.080 1159.050 ;
        RECT 2520.960 1111.110 2521.100 1158.730 ;
        RECT 2520.900 1110.790 2521.160 1111.110 ;
        RECT 2522.280 1110.790 2522.540 1111.110 ;
        RECT 2522.340 1077.110 2522.480 1110.790 ;
        RECT 2522.280 1076.790 2522.540 1077.110 ;
        RECT 2521.360 1076.110 2521.620 1076.430 ;
        RECT 2521.420 1062.570 2521.560 1076.110 ;
        RECT 2520.960 1062.430 2521.560 1062.570 ;
        RECT 2520.960 1028.490 2521.100 1062.430 ;
        RECT 2520.900 1028.170 2521.160 1028.490 ;
        RECT 2521.360 1027.830 2521.620 1028.150 ;
        RECT 2521.420 1014.550 2521.560 1027.830 ;
        RECT 2520.900 1014.230 2521.160 1014.550 ;
        RECT 2521.360 1014.230 2521.620 1014.550 ;
        RECT 2520.960 1006.390 2521.100 1014.230 ;
        RECT 2520.900 1006.070 2521.160 1006.390 ;
        RECT 2522.280 1006.070 2522.540 1006.390 ;
        RECT 2522.340 931.330 2522.480 1006.070 ;
        RECT 2521.880 931.190 2522.480 931.330 ;
        RECT 2521.880 917.845 2522.020 931.190 ;
        RECT 2521.810 917.475 2522.090 917.845 ;
        RECT 2523.190 917.475 2523.470 917.845 ;
        RECT 2523.260 869.710 2523.400 917.475 ;
        RECT 2522.280 869.390 2522.540 869.710 ;
        RECT 2523.200 869.390 2523.460 869.710 ;
        RECT 2522.340 834.770 2522.480 869.390 ;
        RECT 2521.880 834.630 2522.480 834.770 ;
        RECT 2521.880 821.090 2522.020 834.630 ;
        RECT 2520.900 820.770 2521.160 821.090 ;
        RECT 2521.820 820.770 2522.080 821.090 ;
        RECT 2520.960 773.005 2521.100 820.770 ;
        RECT 2520.890 772.635 2521.170 773.005 ;
        RECT 2522.270 772.635 2522.550 773.005 ;
        RECT 2522.340 683.050 2522.480 772.635 ;
        RECT 2185.100 682.730 2185.360 683.050 ;
        RECT 2522.280 682.730 2522.540 683.050 ;
        RECT 2185.160 680.525 2185.300 682.730 ;
        RECT 2185.090 680.155 2185.370 680.525 ;
      LAYER via2 ;
        RECT 2899.930 1730.120 2900.210 1730.400 ;
        RECT 2521.350 1304.440 2521.630 1304.720 ;
        RECT 2522.730 1304.440 2523.010 1304.720 ;
        RECT 2521.810 917.520 2522.090 917.800 ;
        RECT 2523.190 917.520 2523.470 917.800 ;
        RECT 2520.890 772.680 2521.170 772.960 ;
        RECT 2522.270 772.680 2522.550 772.960 ;
        RECT 2185.090 680.200 2185.370 680.480 ;
      LAYER met3 ;
        RECT 2899.905 1730.410 2900.235 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2899.905 1730.110 2924.800 1730.410 ;
        RECT 2899.905 1730.095 2900.235 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2521.325 1304.730 2521.655 1304.745 ;
        RECT 2522.705 1304.730 2523.035 1304.745 ;
        RECT 2521.325 1304.430 2523.035 1304.730 ;
        RECT 2521.325 1304.415 2521.655 1304.430 ;
        RECT 2522.705 1304.415 2523.035 1304.430 ;
        RECT 2521.785 917.810 2522.115 917.825 ;
        RECT 2523.165 917.810 2523.495 917.825 ;
        RECT 2521.785 917.510 2523.495 917.810 ;
        RECT 2521.785 917.495 2522.115 917.510 ;
        RECT 2523.165 917.495 2523.495 917.510 ;
        RECT 2520.865 772.970 2521.195 772.985 ;
        RECT 2522.245 772.970 2522.575 772.985 ;
        RECT 2520.865 772.670 2522.575 772.970 ;
        RECT 2520.865 772.655 2521.195 772.670 ;
        RECT 2522.245 772.655 2522.575 772.670 ;
        RECT 2185.065 680.490 2185.395 680.505 ;
        RECT 2169.670 680.190 2185.395 680.490 ;
        RECT 2169.670 678.840 2169.970 680.190 ;
        RECT 2185.065 680.175 2185.395 680.190 ;
        RECT 2166.000 678.240 2170.000 678.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 689.760 2187.230 689.820 ;
        RECT 2902.670 689.760 2902.990 689.820 ;
        RECT 2186.910 689.620 2902.990 689.760 ;
        RECT 2186.910 689.560 2187.230 689.620 ;
        RECT 2902.670 689.560 2902.990 689.620 ;
      LAYER via ;
        RECT 2186.940 689.560 2187.200 689.820 ;
        RECT 2902.700 689.560 2902.960 689.820 ;
      LAYER met2 ;
        RECT 2902.690 1964.675 2902.970 1965.045 ;
        RECT 2902.760 689.850 2902.900 1964.675 ;
        RECT 2186.940 689.530 2187.200 689.850 ;
        RECT 2902.700 689.530 2902.960 689.850 ;
        RECT 2187.000 689.365 2187.140 689.530 ;
        RECT 2186.930 688.995 2187.210 689.365 ;
      LAYER via2 ;
        RECT 2902.690 1964.720 2902.970 1965.000 ;
        RECT 2186.930 689.040 2187.210 689.320 ;
      LAYER met3 ;
        RECT 2902.665 1965.010 2902.995 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2902.665 1964.710 2924.800 1965.010 ;
        RECT 2902.665 1964.695 2902.995 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2186.905 689.330 2187.235 689.345 ;
        RECT 2169.670 689.040 2187.235 689.330 ;
        RECT 2166.000 689.030 2187.235 689.040 ;
        RECT 2166.000 688.440 2170.000 689.030 ;
        RECT 2186.905 689.015 2187.235 689.030 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2186.910 703.700 2187.230 703.760 ;
        RECT 2902.210 703.700 2902.530 703.760 ;
        RECT 2186.910 703.560 2902.530 703.700 ;
        RECT 2186.910 703.500 2187.230 703.560 ;
        RECT 2902.210 703.500 2902.530 703.560 ;
      LAYER via ;
        RECT 2186.940 703.500 2187.200 703.760 ;
        RECT 2902.240 703.500 2902.500 703.760 ;
      LAYER met2 ;
        RECT 2902.230 2199.275 2902.510 2199.645 ;
        RECT 2902.300 703.790 2902.440 2199.275 ;
        RECT 2186.940 703.470 2187.200 703.790 ;
        RECT 2902.240 703.470 2902.500 703.790 ;
        RECT 2187.000 701.605 2187.140 703.470 ;
        RECT 2186.930 701.235 2187.210 701.605 ;
      LAYER via2 ;
        RECT 2902.230 2199.320 2902.510 2199.600 ;
        RECT 2186.930 701.280 2187.210 701.560 ;
      LAYER met3 ;
        RECT 2902.205 2199.610 2902.535 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2902.205 2199.310 2924.800 2199.610 ;
        RECT 2902.205 2199.295 2902.535 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2186.905 701.570 2187.235 701.585 ;
        RECT 2169.670 701.270 2187.235 701.570 ;
        RECT 2169.670 699.920 2169.970 701.270 ;
        RECT 2186.905 701.255 2187.235 701.270 ;
        RECT 2166.000 699.320 2170.000 699.920 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 917.860 207.160 919.380 207.300 ;
        RECT 660.170 206.960 660.490 207.020 ;
        RECT 917.860 206.960 918.000 207.160 ;
        RECT 660.170 206.820 918.000 206.960 ;
        RECT 919.240 206.960 919.380 207.160 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 919.240 206.820 2901.150 206.960 ;
        RECT 660.170 206.760 660.490 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 660.200 206.760 660.460 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 660.190 801.875 660.470 802.245 ;
        RECT 660.260 207.050 660.400 801.875 ;
        RECT 660.200 206.730 660.460 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 660.190 801.920 660.470 802.200 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 660.165 802.210 660.495 802.225 ;
        RECT 670.000 802.210 674.000 802.600 ;
        RECT 660.165 802.000 674.000 802.210 ;
        RECT 660.165 801.910 670.220 802.000 ;
        RECT 660.165 801.895 660.495 801.910 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 653.730 2501.280 654.050 2501.340 ;
        RECT 2902.670 2501.280 2902.990 2501.340 ;
        RECT 653.730 2501.140 2902.990 2501.280 ;
        RECT 653.730 2501.080 654.050 2501.140 ;
        RECT 2902.670 2501.080 2902.990 2501.140 ;
      LAYER via ;
        RECT 653.760 2501.080 654.020 2501.340 ;
        RECT 2902.700 2501.080 2902.960 2501.340 ;
      LAYER met2 ;
        RECT 2902.690 2551.515 2902.970 2551.885 ;
        RECT 2902.760 2501.370 2902.900 2551.515 ;
        RECT 653.760 2501.050 654.020 2501.370 ;
        RECT 2902.700 2501.050 2902.960 2501.370 ;
        RECT 653.820 854.605 653.960 2501.050 ;
        RECT 653.750 854.235 654.030 854.605 ;
      LAYER via2 ;
        RECT 2902.690 2551.560 2902.970 2551.840 ;
        RECT 653.750 854.280 654.030 854.560 ;
      LAYER met3 ;
        RECT 2902.665 2551.850 2902.995 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2902.665 2551.550 2924.800 2551.850 ;
        RECT 2902.665 2551.535 2902.995 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 653.725 854.570 654.055 854.585 ;
        RECT 670.000 854.570 674.000 854.960 ;
        RECT 653.725 854.360 674.000 854.570 ;
        RECT 653.725 854.270 670.220 854.360 ;
        RECT 653.725 854.255 654.055 854.270 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 653.270 2501.620 653.590 2501.680 ;
        RECT 2902.210 2501.620 2902.530 2501.680 ;
        RECT 653.270 2501.480 2902.530 2501.620 ;
        RECT 653.270 2501.420 653.590 2501.480 ;
        RECT 2902.210 2501.420 2902.530 2501.480 ;
      LAYER via ;
        RECT 653.300 2501.420 653.560 2501.680 ;
        RECT 2902.240 2501.420 2902.500 2501.680 ;
      LAYER met2 ;
        RECT 2902.230 2786.115 2902.510 2786.485 ;
        RECT 2902.300 2501.710 2902.440 2786.115 ;
        RECT 653.300 2501.390 653.560 2501.710 ;
        RECT 2902.240 2501.390 2902.500 2501.710 ;
        RECT 653.360 860.045 653.500 2501.390 ;
        RECT 653.290 859.675 653.570 860.045 ;
      LAYER via2 ;
        RECT 2902.230 2786.160 2902.510 2786.440 ;
        RECT 653.290 859.720 653.570 860.000 ;
      LAYER met3 ;
        RECT 2902.205 2786.450 2902.535 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2902.205 2786.150 2924.800 2786.450 ;
        RECT 2902.205 2786.135 2902.535 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 653.265 860.010 653.595 860.025 ;
        RECT 670.000 860.010 674.000 860.400 ;
        RECT 653.265 859.800 674.000 860.010 ;
        RECT 653.265 859.710 670.220 859.800 ;
        RECT 653.265 859.695 653.595 859.710 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 654.650 3015.700 654.970 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 654.650 3015.560 2901.150 3015.700 ;
        RECT 654.650 3015.500 654.970 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 654.680 3015.500 654.940 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 654.680 3015.470 654.940 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 654.740 864.805 654.880 3015.470 ;
        RECT 654.670 864.435 654.950 864.805 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 654.670 864.480 654.950 864.760 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 654.645 864.770 654.975 864.785 ;
        RECT 670.000 864.770 674.000 865.160 ;
        RECT 654.645 864.560 674.000 864.770 ;
        RECT 654.645 864.470 670.220 864.560 ;
        RECT 654.645 864.455 654.975 864.470 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 647.750 3250.300 648.070 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 647.750 3250.160 2901.150 3250.300 ;
        RECT 647.750 3250.100 648.070 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 647.750 875.740 648.070 875.800 ;
        RECT 660.170 875.740 660.490 875.800 ;
        RECT 647.750 875.600 660.490 875.740 ;
        RECT 647.750 875.540 648.070 875.600 ;
        RECT 660.170 875.540 660.490 875.600 ;
      LAYER via ;
        RECT 647.780 3250.100 648.040 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 647.780 875.540 648.040 875.800 ;
        RECT 660.200 875.540 660.460 875.800 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 647.780 3250.070 648.040 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 647.840 875.830 647.980 3250.070 ;
        RECT 647.780 875.510 648.040 875.830 ;
        RECT 660.200 875.510 660.460 875.830 ;
        RECT 660.260 870.245 660.400 875.510 ;
        RECT 660.190 869.875 660.470 870.245 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 660.190 869.920 660.470 870.200 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 660.165 870.210 660.495 870.225 ;
        RECT 670.000 870.210 674.000 870.600 ;
        RECT 660.165 870.000 674.000 870.210 ;
        RECT 660.165 869.910 670.220 870.000 ;
        RECT 660.165 869.895 660.495 869.910 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 648.210 3484.900 648.530 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 648.210 3484.760 2901.150 3484.900 ;
        RECT 648.210 3484.700 648.530 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 648.210 876.080 648.530 876.140 ;
        RECT 656.030 876.080 656.350 876.140 ;
        RECT 648.210 875.940 656.350 876.080 ;
        RECT 648.210 875.880 648.530 875.940 ;
        RECT 656.030 875.880 656.350 875.940 ;
      LAYER via ;
        RECT 648.240 3484.700 648.500 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 648.240 875.880 648.500 876.140 ;
        RECT 656.060 875.880 656.320 876.140 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 648.240 3484.670 648.500 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 648.300 876.170 648.440 3484.670 ;
        RECT 648.240 875.850 648.500 876.170 ;
        RECT 656.060 875.850 656.320 876.170 ;
        RECT 656.120 875.685 656.260 875.850 ;
        RECT 656.050 875.315 656.330 875.685 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 656.050 875.360 656.330 875.640 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 656.025 875.650 656.355 875.665 ;
        RECT 670.000 875.650 674.000 876.040 ;
        RECT 656.025 875.440 674.000 875.650 ;
        RECT 656.025 875.350 670.220 875.440 ;
        RECT 656.025 875.335 656.355 875.350 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.930 3501.900 663.250 3501.960 ;
        RECT 2635.870 3501.900 2636.190 3501.960 ;
        RECT 662.930 3501.760 2636.190 3501.900 ;
        RECT 662.930 3501.700 663.250 3501.760 ;
        RECT 2635.870 3501.700 2636.190 3501.760 ;
        RECT 662.930 906.340 663.250 906.400 ;
        RECT 666.150 906.340 666.470 906.400 ;
        RECT 662.930 906.200 666.470 906.340 ;
        RECT 662.930 906.140 663.250 906.200 ;
        RECT 666.150 906.140 666.470 906.200 ;
      LAYER via ;
        RECT 662.960 3501.700 663.220 3501.960 ;
        RECT 2635.900 3501.700 2636.160 3501.960 ;
        RECT 662.960 906.140 663.220 906.400 ;
        RECT 666.180 906.140 666.440 906.400 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.990 2636.100 3517.600 ;
        RECT 662.960 3501.670 663.220 3501.990 ;
        RECT 2635.900 3501.670 2636.160 3501.990 ;
        RECT 663.020 906.430 663.160 3501.670 ;
        RECT 662.960 906.110 663.220 906.430 ;
        RECT 666.180 906.110 666.440 906.430 ;
        RECT 666.240 881.125 666.380 906.110 ;
        RECT 666.170 880.755 666.450 881.125 ;
      LAYER via2 ;
        RECT 666.170 880.800 666.450 881.080 ;
      LAYER met3 ;
        RECT 666.145 881.090 666.475 881.105 ;
        RECT 670.000 881.090 674.000 881.480 ;
        RECT 666.145 880.880 674.000 881.090 ;
        RECT 666.145 880.790 670.220 880.880 ;
        RECT 666.145 880.775 666.475 880.790 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.070 3502.920 667.390 3502.980 ;
        RECT 2311.570 3502.920 2311.890 3502.980 ;
        RECT 667.070 3502.780 2311.890 3502.920 ;
        RECT 667.070 3502.720 667.390 3502.780 ;
        RECT 2311.570 3502.720 2311.890 3502.780 ;
      LAYER via ;
        RECT 667.100 3502.720 667.360 3502.980 ;
        RECT 2311.600 3502.720 2311.860 3502.980 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3503.010 2311.800 3517.600 ;
        RECT 667.100 3502.690 667.360 3503.010 ;
        RECT 2311.600 3502.690 2311.860 3503.010 ;
        RECT 667.160 885.885 667.300 3502.690 ;
        RECT 667.090 885.515 667.370 885.885 ;
      LAYER via2 ;
        RECT 667.090 885.560 667.370 885.840 ;
      LAYER met3 ;
        RECT 667.065 885.850 667.395 885.865 ;
        RECT 670.000 885.850 674.000 886.240 ;
        RECT 667.065 885.640 674.000 885.850 ;
        RECT 667.065 885.550 670.220 885.640 ;
        RECT 667.065 885.535 667.395 885.550 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 666.150 3504.280 666.470 3504.340 ;
        RECT 1987.270 3504.280 1987.590 3504.340 ;
        RECT 666.150 3504.140 1987.590 3504.280 ;
        RECT 666.150 3504.080 666.470 3504.140 ;
        RECT 1987.270 3504.080 1987.590 3504.140 ;
      LAYER via ;
        RECT 666.180 3504.080 666.440 3504.340 ;
        RECT 1987.300 3504.080 1987.560 3504.340 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3504.370 1987.500 3517.600 ;
        RECT 666.180 3504.050 666.440 3504.370 ;
        RECT 1987.300 3504.050 1987.560 3504.370 ;
        RECT 666.240 927.365 666.380 3504.050 ;
        RECT 666.170 926.995 666.450 927.365 ;
        RECT 664.330 911.355 664.610 911.725 ;
        RECT 664.400 891.325 664.540 911.355 ;
        RECT 664.330 890.955 664.610 891.325 ;
      LAYER via2 ;
        RECT 666.170 927.040 666.450 927.320 ;
        RECT 664.330 911.400 664.610 911.680 ;
        RECT 664.330 891.000 664.610 891.280 ;
      LAYER met3 ;
        RECT 664.510 927.330 664.890 927.340 ;
        RECT 666.145 927.330 666.475 927.345 ;
        RECT 664.510 927.030 666.475 927.330 ;
        RECT 664.510 927.020 664.890 927.030 ;
        RECT 666.145 927.015 666.475 927.030 ;
        RECT 664.305 911.700 664.635 911.705 ;
        RECT 664.305 911.690 664.890 911.700 ;
        RECT 664.305 911.390 665.090 911.690 ;
        RECT 664.305 911.380 664.890 911.390 ;
        RECT 664.305 911.375 664.635 911.380 ;
        RECT 664.305 891.290 664.635 891.305 ;
        RECT 670.000 891.290 674.000 891.680 ;
        RECT 664.305 891.080 674.000 891.290 ;
        RECT 664.305 890.990 670.220 891.080 ;
        RECT 664.305 890.975 664.635 890.990 ;
      LAYER via3 ;
        RECT 664.540 927.020 664.860 927.340 ;
        RECT 664.540 911.380 664.860 911.700 ;
      LAYER met4 ;
        RECT 664.535 927.015 664.865 927.345 ;
        RECT 664.550 911.705 664.850 927.015 ;
        RECT 664.535 911.375 664.865 911.705 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 666.610 3501.220 666.930 3501.280 ;
        RECT 1662.510 3501.220 1662.830 3501.280 ;
        RECT 666.610 3501.080 1662.830 3501.220 ;
        RECT 666.610 3501.020 666.930 3501.080 ;
        RECT 1662.510 3501.020 1662.830 3501.080 ;
      LAYER via ;
        RECT 666.640 3501.020 666.900 3501.280 ;
        RECT 1662.540 3501.020 1662.800 3501.280 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3501.310 1662.740 3517.600 ;
        RECT 666.640 3500.990 666.900 3501.310 ;
        RECT 1662.540 3500.990 1662.800 3501.310 ;
        RECT 666.700 896.765 666.840 3500.990 ;
        RECT 666.630 896.395 666.910 896.765 ;
      LAYER via2 ;
        RECT 666.630 896.440 666.910 896.720 ;
      LAYER met3 ;
        RECT 666.605 896.730 666.935 896.745 ;
        RECT 670.000 896.730 674.000 897.120 ;
        RECT 666.605 896.520 674.000 896.730 ;
        RECT 666.605 896.430 670.220 896.520 ;
        RECT 666.605 896.415 666.935 896.430 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 660.170 3500.540 660.490 3500.600 ;
        RECT 1338.210 3500.540 1338.530 3500.600 ;
        RECT 660.170 3500.400 1338.530 3500.540 ;
        RECT 660.170 3500.340 660.490 3500.400 ;
        RECT 1338.210 3500.340 1338.530 3500.400 ;
      LAYER via ;
        RECT 660.200 3500.340 660.460 3500.600 ;
        RECT 1338.240 3500.340 1338.500 3500.600 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3500.630 1338.440 3517.600 ;
        RECT 660.200 3500.310 660.460 3500.630 ;
        RECT 1338.240 3500.310 1338.500 3500.630 ;
        RECT 660.260 902.205 660.400 3500.310 ;
        RECT 660.190 901.835 660.470 902.205 ;
      LAYER via2 ;
        RECT 660.190 901.880 660.470 902.160 ;
      LAYER met3 ;
        RECT 660.165 902.170 660.495 902.185 ;
        RECT 670.000 902.170 674.000 902.560 ;
        RECT 660.165 901.960 674.000 902.170 ;
        RECT 660.165 901.870 670.220 901.960 ;
        RECT 660.165 901.855 660.495 901.870 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.530 441.560 667.850 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 667.530 441.420 2901.150 441.560 ;
        RECT 667.530 441.360 667.850 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 667.560 441.360 667.820 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 667.550 806.635 667.830 807.005 ;
        RECT 667.620 441.650 667.760 806.635 ;
        RECT 667.560 441.330 667.820 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 667.550 806.680 667.830 806.960 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 667.525 806.970 667.855 806.985 ;
        RECT 670.000 806.970 674.000 807.360 ;
        RECT 667.525 806.760 674.000 806.970 ;
        RECT 667.525 806.670 670.220 806.760 ;
        RECT 667.525 806.655 667.855 806.670 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 665.690 3500.200 666.010 3500.260 ;
        RECT 1013.910 3500.200 1014.230 3500.260 ;
        RECT 665.690 3500.060 1014.230 3500.200 ;
        RECT 665.690 3500.000 666.010 3500.060 ;
        RECT 1013.910 3500.000 1014.230 3500.060 ;
      LAYER via ;
        RECT 665.720 3500.000 665.980 3500.260 ;
        RECT 1013.940 3500.000 1014.200 3500.260 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3500.290 1014.140 3517.600 ;
        RECT 665.720 3499.970 665.980 3500.290 ;
        RECT 1013.940 3499.970 1014.200 3500.290 ;
        RECT 665.780 926.570 665.920 3499.970 ;
        RECT 665.780 926.430 666.380 926.570 ;
        RECT 666.240 906.965 666.380 926.430 ;
        RECT 666.170 906.595 666.450 906.965 ;
      LAYER via2 ;
        RECT 666.170 906.640 666.450 906.920 ;
      LAYER met3 ;
        RECT 666.145 906.930 666.475 906.945 ;
        RECT 670.000 906.930 674.000 907.320 ;
        RECT 666.145 906.720 674.000 906.930 ;
        RECT 666.145 906.630 670.220 906.720 ;
        RECT 666.145 906.615 666.475 906.630 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 665.230 3498.500 665.550 3498.560 ;
        RECT 689.150 3498.500 689.470 3498.560 ;
        RECT 665.230 3498.360 689.470 3498.500 ;
        RECT 665.230 3498.300 665.550 3498.360 ;
        RECT 689.150 3498.300 689.470 3498.360 ;
        RECT 664.310 925.040 664.630 925.100 ;
        RECT 665.230 925.040 665.550 925.100 ;
        RECT 664.310 924.900 665.550 925.040 ;
        RECT 664.310 924.840 664.630 924.900 ;
        RECT 665.230 924.840 665.550 924.900 ;
      LAYER via ;
        RECT 665.260 3498.300 665.520 3498.560 ;
        RECT 689.180 3498.300 689.440 3498.560 ;
        RECT 664.340 924.840 664.600 925.100 ;
        RECT 665.260 924.840 665.520 925.100 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3498.590 689.380 3517.600 ;
        RECT 665.260 3498.270 665.520 3498.590 ;
        RECT 689.180 3498.270 689.440 3498.590 ;
        RECT 665.320 925.130 665.460 3498.270 ;
        RECT 664.340 924.810 664.600 925.130 ;
        RECT 665.260 924.810 665.520 925.130 ;
        RECT 664.400 912.405 664.540 924.810 ;
        RECT 664.330 912.035 664.610 912.405 ;
      LAYER via2 ;
        RECT 664.330 912.080 664.610 912.360 ;
      LAYER met3 ;
        RECT 664.305 912.370 664.635 912.385 ;
        RECT 670.000 912.370 674.000 912.760 ;
        RECT 664.305 912.160 674.000 912.370 ;
        RECT 664.305 912.070 670.220 912.160 ;
        RECT 664.305 912.055 664.635 912.070 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 362.090 3498.500 362.410 3498.560 ;
        RECT 364.850 3498.500 365.170 3498.560 ;
        RECT 362.090 3498.360 365.170 3498.500 ;
        RECT 362.090 3498.300 362.410 3498.360 ;
        RECT 364.850 3498.300 365.170 3498.360 ;
        RECT 362.090 917.560 362.410 917.620 ;
        RECT 656.030 917.560 656.350 917.620 ;
        RECT 362.090 917.420 656.350 917.560 ;
        RECT 362.090 917.360 362.410 917.420 ;
        RECT 656.030 917.360 656.350 917.420 ;
      LAYER via ;
        RECT 362.120 3498.300 362.380 3498.560 ;
        RECT 364.880 3498.300 365.140 3498.560 ;
        RECT 362.120 917.360 362.380 917.620 ;
        RECT 656.060 917.360 656.320 917.620 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3498.590 365.080 3517.600 ;
        RECT 362.120 3498.270 362.380 3498.590 ;
        RECT 364.880 3498.270 365.140 3498.590 ;
        RECT 362.180 917.650 362.320 3498.270 ;
        RECT 362.120 917.330 362.380 917.650 ;
        RECT 656.050 917.475 656.330 917.845 ;
        RECT 656.060 917.330 656.320 917.475 ;
      LAYER via2 ;
        RECT 656.050 917.520 656.330 917.800 ;
      LAYER met3 ;
        RECT 656.025 917.810 656.355 917.825 ;
        RECT 670.000 917.810 674.000 918.200 ;
        RECT 656.025 917.600 674.000 917.810 ;
        RECT 656.025 917.510 670.220 917.600 ;
        RECT 656.025 917.495 656.355 917.510 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 39.630 3477.420 39.950 3477.480 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 39.630 3477.280 41.330 3477.420 ;
        RECT 39.630 3477.220 39.950 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 39.630 3429.480 39.950 3429.540 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 39.630 3429.340 40.870 3429.480 ;
        RECT 39.630 3429.280 39.950 3429.340 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3270.700 40.410 3270.760 ;
        RECT 41.010 3270.700 41.330 3270.760 ;
        RECT 40.090 3270.560 41.330 3270.700 ;
        RECT 40.090 3270.500 40.410 3270.560 ;
        RECT 41.010 3270.500 41.330 3270.560 ;
        RECT 40.090 3174.140 40.410 3174.200 ;
        RECT 41.010 3174.140 41.330 3174.200 ;
        RECT 40.090 3174.000 41.330 3174.140 ;
        RECT 40.090 3173.940 40.410 3174.000 ;
        RECT 41.010 3173.940 41.330 3174.000 ;
        RECT 40.090 3077.580 40.410 3077.640 ;
        RECT 41.010 3077.580 41.330 3077.640 ;
        RECT 40.090 3077.440 41.330 3077.580 ;
        RECT 40.090 3077.380 40.410 3077.440 ;
        RECT 41.010 3077.380 41.330 3077.440 ;
        RECT 40.090 2981.020 40.410 2981.080 ;
        RECT 41.010 2981.020 41.330 2981.080 ;
        RECT 40.090 2980.880 41.330 2981.020 ;
        RECT 40.090 2980.820 40.410 2980.880 ;
        RECT 41.010 2980.820 41.330 2980.880 ;
        RECT 38.250 2898.060 38.570 2898.120 ;
        RECT 39.630 2898.060 39.950 2898.120 ;
        RECT 38.250 2897.920 39.950 2898.060 ;
        RECT 38.250 2897.860 38.570 2897.920 ;
        RECT 39.630 2897.860 39.950 2897.920 ;
        RECT 38.250 2849.780 38.570 2849.840 ;
        RECT 39.170 2849.780 39.490 2849.840 ;
        RECT 38.250 2849.640 39.490 2849.780 ;
        RECT 38.250 2849.580 38.570 2849.640 ;
        RECT 39.170 2849.580 39.490 2849.640 ;
        RECT 39.170 2815.240 39.490 2815.500 ;
        RECT 39.260 2814.760 39.400 2815.240 ;
        RECT 39.630 2814.760 39.950 2814.820 ;
        RECT 39.260 2814.620 39.950 2814.760 ;
        RECT 39.630 2814.560 39.950 2814.620 ;
        RECT 40.090 2752.880 40.410 2752.940 ;
        RECT 40.550 2752.880 40.870 2752.940 ;
        RECT 40.090 2752.740 40.870 2752.880 ;
        RECT 40.090 2752.680 40.410 2752.740 ;
        RECT 40.550 2752.680 40.870 2752.740 ;
        RECT 40.550 2704.940 40.870 2705.000 ;
        RECT 41.010 2704.940 41.330 2705.000 ;
        RECT 40.550 2704.800 41.330 2704.940 ;
        RECT 40.550 2704.740 40.870 2704.800 ;
        RECT 41.010 2704.740 41.330 2704.800 ;
        RECT 41.010 2608.380 41.330 2608.440 ;
        RECT 41.930 2608.380 42.250 2608.440 ;
        RECT 41.010 2608.240 42.250 2608.380 ;
        RECT 41.010 2608.180 41.330 2608.240 ;
        RECT 41.930 2608.180 42.250 2608.240 ;
        RECT 41.010 2511.820 41.330 2511.880 ;
        RECT 41.930 2511.820 42.250 2511.880 ;
        RECT 41.010 2511.680 42.250 2511.820 ;
        RECT 41.010 2511.620 41.330 2511.680 ;
        RECT 41.930 2511.620 42.250 2511.680 ;
        RECT 40.550 2429.000 40.870 2429.260 ;
        RECT 40.640 2428.860 40.780 2429.000 ;
        RECT 41.010 2428.860 41.330 2428.920 ;
        RECT 40.640 2428.720 41.330 2428.860 ;
        RECT 41.010 2428.660 41.330 2428.720 ;
        RECT 39.630 2414.920 39.950 2414.980 ;
        RECT 41.010 2414.920 41.330 2414.980 ;
        RECT 39.630 2414.780 41.330 2414.920 ;
        RECT 39.630 2414.720 39.950 2414.780 ;
        RECT 41.010 2414.720 41.330 2414.780 ;
        RECT 40.550 2332.100 40.870 2332.360 ;
        RECT 40.640 2331.960 40.780 2332.100 ;
        RECT 41.010 2331.960 41.330 2332.020 ;
        RECT 40.640 2331.820 41.330 2331.960 ;
        RECT 41.010 2331.760 41.330 2331.820 ;
        RECT 39.170 2270.080 39.490 2270.140 ;
        RECT 40.090 2270.080 40.410 2270.140 ;
        RECT 39.170 2269.940 40.410 2270.080 ;
        RECT 39.170 2269.880 39.490 2269.940 ;
        RECT 40.090 2269.880 40.410 2269.940 ;
        RECT 39.170 2222.140 39.490 2222.200 ;
        RECT 39.630 2222.140 39.950 2222.200 ;
        RECT 39.170 2222.000 39.950 2222.140 ;
        RECT 39.170 2221.940 39.490 2222.000 ;
        RECT 39.630 2221.940 39.950 2222.000 ;
        RECT 40.550 2138.980 40.870 2139.240 ;
        RECT 40.640 2138.840 40.780 2138.980 ;
        RECT 41.010 2138.840 41.330 2138.900 ;
        RECT 40.640 2138.700 41.330 2138.840 ;
        RECT 41.010 2138.640 41.330 2138.700 ;
        RECT 39.630 2125.240 39.950 2125.300 ;
        RECT 41.010 2125.240 41.330 2125.300 ;
        RECT 39.630 2125.100 41.330 2125.240 ;
        RECT 39.630 2125.040 39.950 2125.100 ;
        RECT 41.010 2125.040 41.330 2125.100 ;
        RECT 39.630 2077.300 39.950 2077.360 ;
        RECT 40.550 2077.300 40.870 2077.360 ;
        RECT 39.630 2077.160 40.870 2077.300 ;
        RECT 39.630 2077.100 39.950 2077.160 ;
        RECT 40.550 2077.100 40.870 2077.160 ;
        RECT 40.550 2042.420 40.870 2042.680 ;
        RECT 40.640 2041.940 40.780 2042.420 ;
        RECT 41.010 2041.940 41.330 2042.000 ;
        RECT 40.640 2041.800 41.330 2041.940 ;
        RECT 41.010 2041.740 41.330 2041.800 ;
        RECT 41.010 2004.540 41.330 2004.600 ;
        RECT 41.930 2004.540 42.250 2004.600 ;
        RECT 41.010 2004.400 42.250 2004.540 ;
        RECT 41.010 2004.340 41.330 2004.400 ;
        RECT 41.930 2004.340 42.250 2004.400 ;
        RECT 40.090 1980.400 40.410 1980.460 ;
        RECT 41.930 1980.400 42.250 1980.460 ;
        RECT 40.090 1980.260 42.250 1980.400 ;
        RECT 40.090 1980.200 40.410 1980.260 ;
        RECT 41.930 1980.200 42.250 1980.260 ;
        RECT 40.090 1973.600 40.410 1973.660 ;
        RECT 40.550 1973.600 40.870 1973.660 ;
        RECT 40.090 1973.460 40.870 1973.600 ;
        RECT 40.090 1973.400 40.410 1973.460 ;
        RECT 40.550 1973.400 40.870 1973.460 ;
        RECT 40.550 1945.860 40.870 1946.120 ;
        RECT 40.640 1945.380 40.780 1945.860 ;
        RECT 41.010 1945.380 41.330 1945.440 ;
        RECT 40.640 1945.240 41.330 1945.380 ;
        RECT 41.010 1945.180 41.330 1945.240 ;
        RECT 41.010 1897.780 41.330 1897.840 ;
        RECT 40.180 1897.640 41.330 1897.780 ;
        RECT 40.180 1897.500 40.320 1897.640 ;
        RECT 41.010 1897.580 41.330 1897.640 ;
        RECT 40.090 1897.240 40.410 1897.500 ;
        RECT 39.170 1876.700 39.490 1876.760 ;
        RECT 40.090 1876.700 40.410 1876.760 ;
        RECT 39.170 1876.560 40.410 1876.700 ;
        RECT 39.170 1876.500 39.490 1876.560 ;
        RECT 40.090 1876.500 40.410 1876.560 ;
        RECT 39.170 1828.760 39.490 1828.820 ;
        RECT 40.550 1828.760 40.870 1828.820 ;
        RECT 39.170 1828.620 40.870 1828.760 ;
        RECT 39.170 1828.560 39.490 1828.620 ;
        RECT 40.550 1828.560 40.870 1828.620 ;
        RECT 40.550 1801.020 40.870 1801.280 ;
        RECT 40.640 1800.880 40.780 1801.020 ;
        RECT 41.010 1800.880 41.330 1800.940 ;
        RECT 40.640 1800.740 41.330 1800.880 ;
        RECT 41.010 1800.680 41.330 1800.740 ;
        RECT 41.010 1773.340 41.330 1773.400 ;
        RECT 41.930 1773.340 42.250 1773.400 ;
        RECT 41.010 1773.200 42.250 1773.340 ;
        RECT 41.010 1773.140 41.330 1773.200 ;
        RECT 41.930 1773.140 42.250 1773.200 ;
        RECT 41.010 1725.400 41.330 1725.460 ;
        RECT 41.930 1725.400 42.250 1725.460 ;
        RECT 41.010 1725.260 42.250 1725.400 ;
        RECT 41.010 1725.200 41.330 1725.260 ;
        RECT 41.930 1725.200 42.250 1725.260 ;
        RECT 40.090 1628.500 40.410 1628.560 ;
        RECT 41.010 1628.500 41.330 1628.560 ;
        RECT 40.090 1628.360 41.330 1628.500 ;
        RECT 40.090 1628.300 40.410 1628.360 ;
        RECT 41.010 1628.300 41.330 1628.360 ;
        RECT 40.090 1531.940 40.410 1532.000 ;
        RECT 41.010 1531.940 41.330 1532.000 ;
        RECT 40.090 1531.800 41.330 1531.940 ;
        RECT 40.090 1531.740 40.410 1531.800 ;
        RECT 41.010 1531.740 41.330 1531.800 ;
        RECT 40.090 1435.380 40.410 1435.440 ;
        RECT 41.010 1435.380 41.330 1435.440 ;
        RECT 40.090 1435.240 41.330 1435.380 ;
        RECT 40.090 1435.180 40.410 1435.240 ;
        RECT 41.010 1435.180 41.330 1435.240 ;
        RECT 40.090 1338.820 40.410 1338.880 ;
        RECT 41.010 1338.820 41.330 1338.880 ;
        RECT 40.090 1338.680 41.330 1338.820 ;
        RECT 40.090 1338.620 40.410 1338.680 ;
        RECT 41.010 1338.620 41.330 1338.680 ;
        RECT 38.710 1255.860 39.030 1255.920 ;
        RECT 39.630 1255.860 39.950 1255.920 ;
        RECT 38.710 1255.720 39.950 1255.860 ;
        RECT 38.710 1255.660 39.030 1255.720 ;
        RECT 39.630 1255.660 39.950 1255.720 ;
        RECT 38.710 1207.580 39.030 1207.640 ;
        RECT 40.090 1207.580 40.410 1207.640 ;
        RECT 38.710 1207.440 40.410 1207.580 ;
        RECT 38.710 1207.380 39.030 1207.440 ;
        RECT 40.090 1207.380 40.410 1207.440 ;
        RECT 40.090 1173.580 40.410 1173.640 ;
        RECT 39.720 1173.440 40.410 1173.580 ;
        RECT 39.720 1172.960 39.860 1173.440 ;
        RECT 40.090 1173.380 40.410 1173.440 ;
        RECT 39.630 1172.700 39.950 1172.960 ;
        RECT 38.710 1158.960 39.030 1159.020 ;
        RECT 39.630 1158.960 39.950 1159.020 ;
        RECT 38.710 1158.820 39.950 1158.960 ;
        RECT 38.710 1158.760 39.030 1158.820 ;
        RECT 39.630 1158.760 39.950 1158.820 ;
        RECT 38.710 1111.020 39.030 1111.080 ;
        RECT 40.090 1111.020 40.410 1111.080 ;
        RECT 38.710 1110.880 40.410 1111.020 ;
        RECT 38.710 1110.820 39.030 1110.880 ;
        RECT 40.090 1110.820 40.410 1110.880 ;
        RECT 40.090 1077.020 40.410 1077.080 ;
        RECT 39.720 1076.880 40.410 1077.020 ;
        RECT 39.720 1076.400 39.860 1076.880 ;
        RECT 40.090 1076.820 40.410 1076.880 ;
        RECT 39.630 1076.140 39.950 1076.400 ;
        RECT 40.090 1028.060 40.410 1028.120 ;
        RECT 40.090 1027.920 40.780 1028.060 ;
        RECT 40.090 1027.860 40.410 1027.920 ;
        RECT 40.640 1027.780 40.780 1027.920 ;
        RECT 40.550 1027.520 40.870 1027.780 ;
        RECT 40.090 1007.320 40.410 1007.380 ;
        RECT 40.550 1007.320 40.870 1007.380 ;
        RECT 40.090 1007.180 40.870 1007.320 ;
        RECT 40.090 1007.120 40.410 1007.180 ;
        RECT 40.550 1007.120 40.870 1007.180 ;
        RECT 41.470 924.360 41.790 924.420 ;
        RECT 656.030 924.360 656.350 924.420 ;
        RECT 41.470 924.220 656.350 924.360 ;
        RECT 41.470 924.160 41.790 924.220 ;
        RECT 656.030 924.160 656.350 924.220 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 39.660 3477.220 39.920 3477.480 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 39.660 3429.280 39.920 3429.540 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3270.500 40.380 3270.760 ;
        RECT 41.040 3270.500 41.300 3270.760 ;
        RECT 40.120 3173.940 40.380 3174.200 ;
        RECT 41.040 3173.940 41.300 3174.200 ;
        RECT 40.120 3077.380 40.380 3077.640 ;
        RECT 41.040 3077.380 41.300 3077.640 ;
        RECT 40.120 2980.820 40.380 2981.080 ;
        RECT 41.040 2980.820 41.300 2981.080 ;
        RECT 38.280 2897.860 38.540 2898.120 ;
        RECT 39.660 2897.860 39.920 2898.120 ;
        RECT 38.280 2849.580 38.540 2849.840 ;
        RECT 39.200 2849.580 39.460 2849.840 ;
        RECT 39.200 2815.240 39.460 2815.500 ;
        RECT 39.660 2814.560 39.920 2814.820 ;
        RECT 40.120 2752.680 40.380 2752.940 ;
        RECT 40.580 2752.680 40.840 2752.940 ;
        RECT 40.580 2704.740 40.840 2705.000 ;
        RECT 41.040 2704.740 41.300 2705.000 ;
        RECT 41.040 2608.180 41.300 2608.440 ;
        RECT 41.960 2608.180 42.220 2608.440 ;
        RECT 41.040 2511.620 41.300 2511.880 ;
        RECT 41.960 2511.620 42.220 2511.880 ;
        RECT 40.580 2429.000 40.840 2429.260 ;
        RECT 41.040 2428.660 41.300 2428.920 ;
        RECT 39.660 2414.720 39.920 2414.980 ;
        RECT 41.040 2414.720 41.300 2414.980 ;
        RECT 40.580 2332.100 40.840 2332.360 ;
        RECT 41.040 2331.760 41.300 2332.020 ;
        RECT 39.200 2269.880 39.460 2270.140 ;
        RECT 40.120 2269.880 40.380 2270.140 ;
        RECT 39.200 2221.940 39.460 2222.200 ;
        RECT 39.660 2221.940 39.920 2222.200 ;
        RECT 40.580 2138.980 40.840 2139.240 ;
        RECT 41.040 2138.640 41.300 2138.900 ;
        RECT 39.660 2125.040 39.920 2125.300 ;
        RECT 41.040 2125.040 41.300 2125.300 ;
        RECT 39.660 2077.100 39.920 2077.360 ;
        RECT 40.580 2077.100 40.840 2077.360 ;
        RECT 40.580 2042.420 40.840 2042.680 ;
        RECT 41.040 2041.740 41.300 2042.000 ;
        RECT 41.040 2004.340 41.300 2004.600 ;
        RECT 41.960 2004.340 42.220 2004.600 ;
        RECT 40.120 1980.200 40.380 1980.460 ;
        RECT 41.960 1980.200 42.220 1980.460 ;
        RECT 40.120 1973.400 40.380 1973.660 ;
        RECT 40.580 1973.400 40.840 1973.660 ;
        RECT 40.580 1945.860 40.840 1946.120 ;
        RECT 41.040 1945.180 41.300 1945.440 ;
        RECT 41.040 1897.580 41.300 1897.840 ;
        RECT 40.120 1897.240 40.380 1897.500 ;
        RECT 39.200 1876.500 39.460 1876.760 ;
        RECT 40.120 1876.500 40.380 1876.760 ;
        RECT 39.200 1828.560 39.460 1828.820 ;
        RECT 40.580 1828.560 40.840 1828.820 ;
        RECT 40.580 1801.020 40.840 1801.280 ;
        RECT 41.040 1800.680 41.300 1800.940 ;
        RECT 41.040 1773.140 41.300 1773.400 ;
        RECT 41.960 1773.140 42.220 1773.400 ;
        RECT 41.040 1725.200 41.300 1725.460 ;
        RECT 41.960 1725.200 42.220 1725.460 ;
        RECT 40.120 1628.300 40.380 1628.560 ;
        RECT 41.040 1628.300 41.300 1628.560 ;
        RECT 40.120 1531.740 40.380 1532.000 ;
        RECT 41.040 1531.740 41.300 1532.000 ;
        RECT 40.120 1435.180 40.380 1435.440 ;
        RECT 41.040 1435.180 41.300 1435.440 ;
        RECT 40.120 1338.620 40.380 1338.880 ;
        RECT 41.040 1338.620 41.300 1338.880 ;
        RECT 38.740 1255.660 39.000 1255.920 ;
        RECT 39.660 1255.660 39.920 1255.920 ;
        RECT 38.740 1207.380 39.000 1207.640 ;
        RECT 40.120 1207.380 40.380 1207.640 ;
        RECT 40.120 1173.380 40.380 1173.640 ;
        RECT 39.660 1172.700 39.920 1172.960 ;
        RECT 38.740 1158.760 39.000 1159.020 ;
        RECT 39.660 1158.760 39.920 1159.020 ;
        RECT 38.740 1110.820 39.000 1111.080 ;
        RECT 40.120 1110.820 40.380 1111.080 ;
        RECT 40.120 1076.820 40.380 1077.080 ;
        RECT 39.660 1076.140 39.920 1076.400 ;
        RECT 40.120 1027.860 40.380 1028.120 ;
        RECT 40.580 1027.520 40.840 1027.780 ;
        RECT 40.120 1007.120 40.380 1007.380 ;
        RECT 40.580 1007.120 40.840 1007.380 ;
        RECT 41.500 924.160 41.760 924.420 ;
        RECT 656.060 924.160 656.320 924.420 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 39.660 3477.190 39.920 3477.510 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 39.720 3429.570 39.860 3477.190 ;
        RECT 39.660 3429.250 39.920 3429.570 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3270.790 40.320 3318.670 ;
        RECT 40.120 3270.470 40.380 3270.790 ;
        RECT 41.040 3270.470 41.300 3270.790 ;
        RECT 41.100 3222.250 41.240 3270.470 ;
        RECT 40.180 3222.110 41.240 3222.250 ;
        RECT 40.180 3174.230 40.320 3222.110 ;
        RECT 40.120 3173.910 40.380 3174.230 ;
        RECT 41.040 3173.910 41.300 3174.230 ;
        RECT 41.100 3125.690 41.240 3173.910 ;
        RECT 40.180 3125.550 41.240 3125.690 ;
        RECT 40.180 3077.670 40.320 3125.550 ;
        RECT 40.120 3077.350 40.380 3077.670 ;
        RECT 41.040 3077.350 41.300 3077.670 ;
        RECT 41.100 3029.130 41.240 3077.350 ;
        RECT 40.180 3028.990 41.240 3029.130 ;
        RECT 40.180 2981.110 40.320 3028.990 ;
        RECT 40.120 2980.790 40.380 2981.110 ;
        RECT 41.040 2980.850 41.300 2981.110 ;
        RECT 40.640 2980.790 41.300 2980.850 ;
        RECT 40.640 2980.710 41.240 2980.790 ;
        RECT 40.640 2959.770 40.780 2980.710 ;
        RECT 40.180 2959.630 40.780 2959.770 ;
        RECT 40.180 2912.170 40.320 2959.630 ;
        RECT 39.720 2912.030 40.320 2912.170 ;
        RECT 39.720 2898.150 39.860 2912.030 ;
        RECT 38.280 2897.830 38.540 2898.150 ;
        RECT 39.660 2897.830 39.920 2898.150 ;
        RECT 38.340 2849.870 38.480 2897.830 ;
        RECT 38.280 2849.550 38.540 2849.870 ;
        RECT 39.200 2849.550 39.460 2849.870 ;
        RECT 39.260 2815.530 39.400 2849.550 ;
        RECT 39.200 2815.210 39.460 2815.530 ;
        RECT 39.660 2814.530 39.920 2814.850 ;
        RECT 39.720 2766.650 39.860 2814.530 ;
        RECT 39.720 2766.510 40.320 2766.650 ;
        RECT 40.180 2752.970 40.320 2766.510 ;
        RECT 40.120 2752.650 40.380 2752.970 ;
        RECT 40.580 2752.650 40.840 2752.970 ;
        RECT 40.640 2705.030 40.780 2752.650 ;
        RECT 40.580 2704.710 40.840 2705.030 ;
        RECT 41.040 2704.710 41.300 2705.030 ;
        RECT 41.100 2670.090 41.240 2704.710 ;
        RECT 40.640 2669.950 41.240 2670.090 ;
        RECT 40.640 2656.605 40.780 2669.950 ;
        RECT 40.570 2656.235 40.850 2656.605 ;
        RECT 41.950 2656.235 42.230 2656.605 ;
        RECT 42.020 2608.470 42.160 2656.235 ;
        RECT 41.040 2608.150 41.300 2608.470 ;
        RECT 41.960 2608.150 42.220 2608.470 ;
        RECT 41.100 2573.530 41.240 2608.150 ;
        RECT 40.640 2573.390 41.240 2573.530 ;
        RECT 40.640 2560.045 40.780 2573.390 ;
        RECT 40.570 2559.675 40.850 2560.045 ;
        RECT 41.950 2559.675 42.230 2560.045 ;
        RECT 42.020 2511.910 42.160 2559.675 ;
        RECT 41.040 2511.590 41.300 2511.910 ;
        RECT 41.960 2511.590 42.220 2511.910 ;
        RECT 41.100 2476.970 41.240 2511.590 ;
        RECT 40.640 2476.830 41.240 2476.970 ;
        RECT 40.640 2429.290 40.780 2476.830 ;
        RECT 40.580 2428.970 40.840 2429.290 ;
        RECT 41.040 2428.630 41.300 2428.950 ;
        RECT 41.100 2415.010 41.240 2428.630 ;
        RECT 39.660 2414.690 39.920 2415.010 ;
        RECT 41.040 2414.690 41.300 2415.010 ;
        RECT 39.720 2366.925 39.860 2414.690 ;
        RECT 39.650 2366.555 39.930 2366.925 ;
        RECT 40.570 2366.555 40.850 2366.925 ;
        RECT 40.640 2332.390 40.780 2366.555 ;
        RECT 40.580 2332.070 40.840 2332.390 ;
        RECT 41.040 2331.730 41.300 2332.050 ;
        RECT 41.100 2283.850 41.240 2331.730 ;
        RECT 40.180 2283.710 41.240 2283.850 ;
        RECT 40.180 2270.170 40.320 2283.710 ;
        RECT 39.200 2269.850 39.460 2270.170 ;
        RECT 40.120 2269.850 40.380 2270.170 ;
        RECT 39.260 2222.230 39.400 2269.850 ;
        RECT 39.200 2221.910 39.460 2222.230 ;
        RECT 39.660 2221.910 39.920 2222.230 ;
        RECT 39.720 2187.290 39.860 2221.910 ;
        RECT 39.720 2187.150 40.780 2187.290 ;
        RECT 40.640 2139.270 40.780 2187.150 ;
        RECT 40.580 2138.950 40.840 2139.270 ;
        RECT 41.040 2138.610 41.300 2138.930 ;
        RECT 41.100 2125.330 41.240 2138.610 ;
        RECT 39.660 2125.010 39.920 2125.330 ;
        RECT 41.040 2125.010 41.300 2125.330 ;
        RECT 39.720 2077.390 39.860 2125.010 ;
        RECT 39.660 2077.070 39.920 2077.390 ;
        RECT 40.580 2077.070 40.840 2077.390 ;
        RECT 40.640 2042.710 40.780 2077.070 ;
        RECT 40.580 2042.390 40.840 2042.710 ;
        RECT 41.040 2041.710 41.300 2042.030 ;
        RECT 41.100 2004.630 41.240 2041.710 ;
        RECT 41.040 2004.310 41.300 2004.630 ;
        RECT 41.960 2004.310 42.220 2004.630 ;
        RECT 42.020 1980.490 42.160 2004.310 ;
        RECT 40.120 1980.170 40.380 1980.490 ;
        RECT 41.960 1980.170 42.220 1980.490 ;
        RECT 40.180 1973.690 40.320 1980.170 ;
        RECT 40.120 1973.370 40.380 1973.690 ;
        RECT 40.580 1973.370 40.840 1973.690 ;
        RECT 40.640 1946.150 40.780 1973.370 ;
        RECT 40.580 1945.830 40.840 1946.150 ;
        RECT 41.040 1945.150 41.300 1945.470 ;
        RECT 41.100 1897.870 41.240 1945.150 ;
        RECT 41.040 1897.550 41.300 1897.870 ;
        RECT 40.120 1897.210 40.380 1897.530 ;
        RECT 40.180 1876.790 40.320 1897.210 ;
        RECT 39.200 1876.470 39.460 1876.790 ;
        RECT 40.120 1876.470 40.380 1876.790 ;
        RECT 39.260 1828.850 39.400 1876.470 ;
        RECT 39.200 1828.530 39.460 1828.850 ;
        RECT 40.580 1828.530 40.840 1828.850 ;
        RECT 40.640 1801.310 40.780 1828.530 ;
        RECT 40.580 1800.990 40.840 1801.310 ;
        RECT 41.040 1800.650 41.300 1800.970 ;
        RECT 41.100 1773.430 41.240 1800.650 ;
        RECT 41.040 1773.110 41.300 1773.430 ;
        RECT 41.960 1773.110 42.220 1773.430 ;
        RECT 42.020 1725.490 42.160 1773.110 ;
        RECT 41.040 1725.170 41.300 1725.490 ;
        RECT 41.960 1725.170 42.220 1725.490 ;
        RECT 41.100 1676.610 41.240 1725.170 ;
        RECT 40.180 1676.470 41.240 1676.610 ;
        RECT 40.180 1628.590 40.320 1676.470 ;
        RECT 40.120 1628.270 40.380 1628.590 ;
        RECT 41.040 1628.270 41.300 1628.590 ;
        RECT 41.100 1580.050 41.240 1628.270 ;
        RECT 40.180 1579.910 41.240 1580.050 ;
        RECT 40.180 1532.030 40.320 1579.910 ;
        RECT 40.120 1531.710 40.380 1532.030 ;
        RECT 41.040 1531.710 41.300 1532.030 ;
        RECT 41.100 1483.490 41.240 1531.710 ;
        RECT 40.180 1483.350 41.240 1483.490 ;
        RECT 40.180 1435.470 40.320 1483.350 ;
        RECT 40.120 1435.150 40.380 1435.470 ;
        RECT 41.040 1435.150 41.300 1435.470 ;
        RECT 41.100 1386.930 41.240 1435.150 ;
        RECT 40.180 1386.790 41.240 1386.930 ;
        RECT 40.180 1338.910 40.320 1386.790 ;
        RECT 40.120 1338.590 40.380 1338.910 ;
        RECT 41.040 1338.650 41.300 1338.910 ;
        RECT 40.640 1338.590 41.300 1338.650 ;
        RECT 40.640 1338.510 41.240 1338.590 ;
        RECT 40.640 1317.570 40.780 1338.510 ;
        RECT 40.180 1317.430 40.780 1317.570 ;
        RECT 40.180 1269.970 40.320 1317.430 ;
        RECT 39.720 1269.830 40.320 1269.970 ;
        RECT 39.720 1255.950 39.860 1269.830 ;
        RECT 38.740 1255.630 39.000 1255.950 ;
        RECT 39.660 1255.630 39.920 1255.950 ;
        RECT 38.800 1207.670 38.940 1255.630 ;
        RECT 38.740 1207.350 39.000 1207.670 ;
        RECT 40.120 1207.350 40.380 1207.670 ;
        RECT 40.180 1173.670 40.320 1207.350 ;
        RECT 40.120 1173.350 40.380 1173.670 ;
        RECT 39.660 1172.670 39.920 1172.990 ;
        RECT 39.720 1159.050 39.860 1172.670 ;
        RECT 38.740 1158.730 39.000 1159.050 ;
        RECT 39.660 1158.730 39.920 1159.050 ;
        RECT 38.800 1111.110 38.940 1158.730 ;
        RECT 38.740 1110.790 39.000 1111.110 ;
        RECT 40.120 1110.790 40.380 1111.110 ;
        RECT 40.180 1077.110 40.320 1110.790 ;
        RECT 40.120 1076.790 40.380 1077.110 ;
        RECT 39.660 1076.110 39.920 1076.430 ;
        RECT 39.720 1062.570 39.860 1076.110 ;
        RECT 39.720 1062.430 40.320 1062.570 ;
        RECT 40.180 1028.150 40.320 1062.430 ;
        RECT 40.120 1027.830 40.380 1028.150 ;
        RECT 40.580 1027.490 40.840 1027.810 ;
        RECT 40.640 1007.410 40.780 1027.490 ;
        RECT 40.120 1007.090 40.380 1007.410 ;
        RECT 40.580 1007.090 40.840 1007.410 ;
        RECT 40.180 966.125 40.320 1007.090 ;
        RECT 40.110 965.755 40.390 966.125 ;
        RECT 41.490 965.755 41.770 966.125 ;
        RECT 41.560 924.450 41.700 965.755 ;
        RECT 41.500 924.130 41.760 924.450 ;
        RECT 656.060 924.130 656.320 924.450 ;
        RECT 656.120 922.605 656.260 924.130 ;
        RECT 656.050 922.235 656.330 922.605 ;
      LAYER via2 ;
        RECT 40.570 2656.280 40.850 2656.560 ;
        RECT 41.950 2656.280 42.230 2656.560 ;
        RECT 40.570 2559.720 40.850 2560.000 ;
        RECT 41.950 2559.720 42.230 2560.000 ;
        RECT 39.650 2366.600 39.930 2366.880 ;
        RECT 40.570 2366.600 40.850 2366.880 ;
        RECT 40.110 965.800 40.390 966.080 ;
        RECT 41.490 965.800 41.770 966.080 ;
        RECT 656.050 922.280 656.330 922.560 ;
      LAYER met3 ;
        RECT 40.545 2656.570 40.875 2656.585 ;
        RECT 41.925 2656.570 42.255 2656.585 ;
        RECT 40.545 2656.270 42.255 2656.570 ;
        RECT 40.545 2656.255 40.875 2656.270 ;
        RECT 41.925 2656.255 42.255 2656.270 ;
        RECT 40.545 2560.010 40.875 2560.025 ;
        RECT 41.925 2560.010 42.255 2560.025 ;
        RECT 40.545 2559.710 42.255 2560.010 ;
        RECT 40.545 2559.695 40.875 2559.710 ;
        RECT 41.925 2559.695 42.255 2559.710 ;
        RECT 39.625 2366.890 39.955 2366.905 ;
        RECT 40.545 2366.890 40.875 2366.905 ;
        RECT 39.625 2366.590 40.875 2366.890 ;
        RECT 39.625 2366.575 39.955 2366.590 ;
        RECT 40.545 2366.575 40.875 2366.590 ;
        RECT 40.085 966.090 40.415 966.105 ;
        RECT 41.465 966.090 41.795 966.105 ;
        RECT 40.085 965.790 41.795 966.090 ;
        RECT 40.085 965.775 40.415 965.790 ;
        RECT 41.465 965.775 41.795 965.790 ;
        RECT 656.025 922.570 656.355 922.585 ;
        RECT 670.000 922.570 674.000 922.960 ;
        RECT 656.025 922.360 674.000 922.570 ;
        RECT 656.025 922.270 670.220 922.360 ;
        RECT 656.025 922.255 656.355 922.270 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 931.500 17.870 931.560 ;
        RECT 656.030 931.500 656.350 931.560 ;
        RECT 17.550 931.360 656.350 931.500 ;
        RECT 17.550 931.300 17.870 931.360 ;
        RECT 656.030 931.300 656.350 931.360 ;
      LAYER via ;
        RECT 17.580 931.300 17.840 931.560 ;
        RECT 656.060 931.300 656.320 931.560 ;
      LAYER met2 ;
        RECT 17.570 3267.555 17.850 3267.925 ;
        RECT 17.640 931.590 17.780 3267.555 ;
        RECT 17.580 931.270 17.840 931.590 ;
        RECT 656.060 931.270 656.320 931.590 ;
        RECT 656.120 928.045 656.260 931.270 ;
        RECT 656.050 927.675 656.330 928.045 ;
      LAYER via2 ;
        RECT 17.570 3267.600 17.850 3267.880 ;
        RECT 656.050 927.720 656.330 928.000 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 17.545 3267.890 17.875 3267.905 ;
        RECT -4.800 3267.590 17.875 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 17.545 3267.575 17.875 3267.590 ;
        RECT 656.025 928.010 656.355 928.025 ;
        RECT 670.000 928.010 674.000 928.400 ;
        RECT 656.025 927.800 674.000 928.010 ;
        RECT 656.025 927.710 670.220 927.800 ;
        RECT 656.025 927.695 656.355 927.710 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 938.300 18.790 938.360 ;
        RECT 656.030 938.300 656.350 938.360 ;
        RECT 18.470 938.160 656.350 938.300 ;
        RECT 18.470 938.100 18.790 938.160 ;
        RECT 656.030 938.100 656.350 938.160 ;
      LAYER via ;
        RECT 18.500 938.100 18.760 938.360 ;
        RECT 656.060 938.100 656.320 938.360 ;
      LAYER met2 ;
        RECT 18.490 2979.915 18.770 2980.285 ;
        RECT 18.560 938.390 18.700 2979.915 ;
        RECT 18.500 938.070 18.760 938.390 ;
        RECT 656.060 938.070 656.320 938.390 ;
        RECT 656.120 933.485 656.260 938.070 ;
        RECT 656.050 933.115 656.330 933.485 ;
      LAYER via2 ;
        RECT 18.490 2979.960 18.770 2980.240 ;
        RECT 656.050 933.160 656.330 933.440 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 18.465 2980.250 18.795 2980.265 ;
        RECT -4.800 2979.950 18.795 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 18.465 2979.935 18.795 2979.950 ;
        RECT 656.025 933.450 656.355 933.465 ;
        RECT 670.000 933.450 674.000 933.840 ;
        RECT 656.025 933.240 674.000 933.450 ;
        RECT 656.025 933.150 670.220 933.240 ;
        RECT 656.025 933.135 656.355 933.150 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 2692.360 20.170 2692.420 ;
        RECT 23.990 2692.360 24.310 2692.420 ;
        RECT 19.850 2692.220 24.310 2692.360 ;
        RECT 19.850 2692.160 20.170 2692.220 ;
        RECT 23.990 2692.160 24.310 2692.220 ;
        RECT 23.990 944.420 24.310 944.480 ;
        RECT 23.990 944.280 48.140 944.420 ;
        RECT 23.990 944.220 24.310 944.280 ;
        RECT 48.000 944.080 48.140 944.280 ;
        RECT 48.370 944.220 48.690 944.480 ;
        RECT 96.210 944.420 96.530 944.480 ;
        RECT 110.470 944.420 110.790 944.480 ;
        RECT 96.210 944.280 110.790 944.420 ;
        RECT 96.210 944.220 96.530 944.280 ;
        RECT 110.470 944.220 110.790 944.280 ;
        RECT 110.930 944.420 111.250 944.480 ;
        RECT 110.930 944.280 144.740 944.420 ;
        RECT 110.930 944.220 111.250 944.280 ;
        RECT 48.460 944.080 48.600 944.220 ;
        RECT 48.000 943.940 48.600 944.080 ;
        RECT 144.600 944.080 144.740 944.280 ;
        RECT 338.170 944.080 338.490 944.140 ;
        RECT 434.770 944.080 435.090 944.140 ;
        RECT 579.670 944.080 579.990 944.140 ;
        RECT 144.600 943.940 158.540 944.080 ;
        RECT 158.400 943.400 158.540 943.940 ;
        RECT 304.220 943.940 338.490 944.080 ;
        RECT 207.530 943.740 207.850 943.800 ;
        RECT 303.670 943.740 303.990 943.800 ;
        RECT 304.220 943.740 304.360 943.940 ;
        RECT 338.170 943.880 338.490 943.940 ;
        RECT 406.340 943.940 435.090 944.080 ;
        RECT 207.530 943.600 241.800 943.740 ;
        RECT 207.530 943.540 207.850 943.600 ;
        RECT 241.660 943.460 241.800 943.600 ;
        RECT 303.670 943.600 304.360 943.740 ;
        RECT 386.010 943.740 386.330 943.800 ;
        RECT 399.810 943.740 400.130 943.800 ;
        RECT 386.010 943.600 400.130 943.740 ;
        RECT 303.670 943.540 303.990 943.600 ;
        RECT 386.010 943.540 386.330 943.600 ;
        RECT 399.810 943.540 400.130 943.600 ;
        RECT 400.270 943.740 400.590 943.800 ;
        RECT 406.340 943.740 406.480 943.940 ;
        RECT 434.770 943.880 435.090 943.940 ;
        RECT 544.800 943.940 579.990 944.080 ;
        RECT 544.800 943.740 544.940 943.940 ;
        RECT 579.670 943.880 579.990 943.940 ;
        RECT 400.270 943.600 406.480 943.740 ;
        RECT 531.000 943.600 544.940 943.740 ;
        RECT 400.270 943.540 400.590 943.600 ;
        RECT 206.610 943.400 206.930 943.460 ;
        RECT 158.400 943.260 206.930 943.400 ;
        RECT 206.610 943.200 206.930 943.260 ;
        RECT 241.570 943.200 241.890 943.460 ;
        RECT 289.410 943.400 289.730 943.460 ;
        RECT 303.210 943.400 303.530 943.460 ;
        RECT 289.410 943.260 303.530 943.400 ;
        RECT 289.410 943.200 289.730 943.260 ;
        RECT 303.210 943.200 303.530 943.260 ;
        RECT 482.610 943.400 482.930 943.460 ;
        RECT 496.870 943.400 497.190 943.460 ;
        RECT 482.610 943.260 497.190 943.400 ;
        RECT 482.610 943.200 482.930 943.260 ;
        RECT 496.870 943.200 497.190 943.260 ;
        RECT 497.330 943.400 497.650 943.460 ;
        RECT 531.000 943.400 531.140 943.600 ;
        RECT 627.510 943.540 627.830 943.800 ;
        RECT 497.330 943.260 531.140 943.400 ;
        RECT 627.600 943.400 627.740 943.540 ;
        RECT 627.600 943.260 656.260 943.400 ;
        RECT 497.330 943.200 497.650 943.260 ;
        RECT 656.120 943.120 656.260 943.260 ;
        RECT 656.030 942.860 656.350 943.120 ;
        RECT 241.570 942.720 241.890 942.780 ;
        RECT 289.410 942.720 289.730 942.780 ;
        RECT 241.570 942.580 289.730 942.720 ;
        RECT 241.570 942.520 241.890 942.580 ;
        RECT 289.410 942.520 289.730 942.580 ;
      LAYER via ;
        RECT 19.880 2692.160 20.140 2692.420 ;
        RECT 24.020 2692.160 24.280 2692.420 ;
        RECT 24.020 944.220 24.280 944.480 ;
        RECT 48.400 944.220 48.660 944.480 ;
        RECT 96.240 944.220 96.500 944.480 ;
        RECT 110.500 944.220 110.760 944.480 ;
        RECT 110.960 944.220 111.220 944.480 ;
        RECT 207.560 943.540 207.820 943.800 ;
        RECT 303.700 943.540 303.960 943.800 ;
        RECT 338.200 943.880 338.460 944.140 ;
        RECT 386.040 943.540 386.300 943.800 ;
        RECT 399.840 943.540 400.100 943.800 ;
        RECT 400.300 943.540 400.560 943.800 ;
        RECT 434.800 943.880 435.060 944.140 ;
        RECT 579.700 943.880 579.960 944.140 ;
        RECT 206.640 943.200 206.900 943.460 ;
        RECT 241.600 943.200 241.860 943.460 ;
        RECT 289.440 943.200 289.700 943.460 ;
        RECT 303.240 943.200 303.500 943.460 ;
        RECT 482.640 943.200 482.900 943.460 ;
        RECT 496.900 943.200 497.160 943.460 ;
        RECT 497.360 943.200 497.620 943.460 ;
        RECT 627.540 943.540 627.800 943.800 ;
        RECT 656.060 942.860 656.320 943.120 ;
        RECT 241.600 942.520 241.860 942.780 ;
        RECT 289.440 942.520 289.700 942.780 ;
      LAYER met2 ;
        RECT 19.870 2692.955 20.150 2693.325 ;
        RECT 19.940 2692.450 20.080 2692.955 ;
        RECT 19.880 2692.130 20.140 2692.450 ;
        RECT 24.020 2692.130 24.280 2692.450 ;
        RECT 24.080 944.510 24.220 2692.130 ;
        RECT 48.390 944.675 48.670 945.045 ;
        RECT 96.230 944.675 96.510 945.045 ;
        RECT 48.460 944.510 48.600 944.675 ;
        RECT 96.300 944.510 96.440 944.675 ;
        RECT 24.020 944.190 24.280 944.510 ;
        RECT 48.400 944.190 48.660 944.510 ;
        RECT 96.240 944.190 96.500 944.510 ;
        RECT 110.500 944.250 110.760 944.510 ;
        RECT 110.960 944.250 111.220 944.510 ;
        RECT 110.500 944.190 111.220 944.250 ;
        RECT 110.560 944.110 111.160 944.190 ;
        RECT 338.190 943.995 338.470 944.365 ;
        RECT 386.030 943.995 386.310 944.365 ;
        RECT 434.790 943.995 435.070 944.365 ;
        RECT 481.710 943.995 481.990 944.365 ;
        RECT 579.690 943.995 579.970 944.365 ;
        RECT 627.530 943.995 627.810 944.365 ;
        RECT 338.200 943.850 338.460 943.995 ;
        RECT 386.100 943.830 386.240 943.995 ;
        RECT 434.800 943.850 435.060 943.995 ;
        RECT 207.560 943.570 207.820 943.830 ;
        RECT 303.700 943.570 303.960 943.830 ;
        RECT 206.700 943.510 207.820 943.570 ;
        RECT 303.300 943.510 303.960 943.570 ;
        RECT 386.040 943.510 386.300 943.830 ;
        RECT 399.840 943.570 400.100 943.830 ;
        RECT 400.300 943.570 400.560 943.830 ;
        RECT 399.840 943.510 400.560 943.570 ;
        RECT 206.700 943.490 207.760 943.510 ;
        RECT 303.300 943.490 303.900 943.510 ;
        RECT 206.640 943.430 207.760 943.490 ;
        RECT 206.640 943.170 206.900 943.430 ;
        RECT 241.600 943.170 241.860 943.490 ;
        RECT 289.440 943.170 289.700 943.490 ;
        RECT 303.240 943.430 303.900 943.490 ;
        RECT 399.900 943.430 400.500 943.510 ;
        RECT 303.240 943.170 303.500 943.430 ;
        RECT 241.660 942.810 241.800 943.170 ;
        RECT 289.500 942.810 289.640 943.170 ;
        RECT 481.780 942.890 481.920 943.995 ;
        RECT 579.700 943.850 579.960 943.995 ;
        RECT 627.600 943.830 627.740 943.995 ;
        RECT 496.960 943.490 497.560 943.570 ;
        RECT 627.540 943.510 627.800 943.830 ;
        RECT 482.640 943.170 482.900 943.490 ;
        RECT 496.900 943.430 497.620 943.490 ;
        RECT 496.900 943.170 497.160 943.430 ;
        RECT 497.360 943.170 497.620 943.430 ;
        RECT 482.700 942.890 482.840 943.170 ;
        RECT 241.600 942.490 241.860 942.810 ;
        RECT 289.440 942.490 289.700 942.810 ;
        RECT 481.780 942.750 482.840 942.890 ;
        RECT 656.060 942.830 656.320 943.150 ;
        RECT 656.120 938.925 656.260 942.830 ;
        RECT 656.050 938.555 656.330 938.925 ;
      LAYER via2 ;
        RECT 19.870 2693.000 20.150 2693.280 ;
        RECT 48.390 944.720 48.670 945.000 ;
        RECT 96.230 944.720 96.510 945.000 ;
        RECT 338.190 944.040 338.470 944.320 ;
        RECT 386.030 944.040 386.310 944.320 ;
        RECT 434.790 944.040 435.070 944.320 ;
        RECT 481.710 944.040 481.990 944.320 ;
        RECT 579.690 944.040 579.970 944.320 ;
        RECT 627.530 944.040 627.810 944.320 ;
        RECT 656.050 938.600 656.330 938.880 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 19.845 2693.290 20.175 2693.305 ;
        RECT -4.800 2692.990 20.175 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 19.845 2692.975 20.175 2692.990 ;
        RECT 48.365 945.010 48.695 945.025 ;
        RECT 96.205 945.010 96.535 945.025 ;
        RECT 48.365 944.710 96.535 945.010 ;
        RECT 48.365 944.695 48.695 944.710 ;
        RECT 96.205 944.695 96.535 944.710 ;
        RECT 338.165 944.330 338.495 944.345 ;
        RECT 386.005 944.330 386.335 944.345 ;
        RECT 338.165 944.030 386.335 944.330 ;
        RECT 338.165 944.015 338.495 944.030 ;
        RECT 386.005 944.015 386.335 944.030 ;
        RECT 434.765 944.330 435.095 944.345 ;
        RECT 481.685 944.330 482.015 944.345 ;
        RECT 434.765 944.030 482.015 944.330 ;
        RECT 434.765 944.015 435.095 944.030 ;
        RECT 481.685 944.015 482.015 944.030 ;
        RECT 579.665 944.330 579.995 944.345 ;
        RECT 627.505 944.330 627.835 944.345 ;
        RECT 579.665 944.030 627.835 944.330 ;
        RECT 579.665 944.015 579.995 944.030 ;
        RECT 627.505 944.015 627.835 944.030 ;
        RECT 656.025 938.890 656.355 938.905 ;
        RECT 670.000 938.890 674.000 939.280 ;
        RECT 656.025 938.680 674.000 938.890 ;
        RECT 656.025 938.590 670.220 938.680 ;
        RECT 656.025 938.575 656.355 938.590 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2405.400 16.030 2405.460 ;
        RECT 24.450 2405.400 24.770 2405.460 ;
        RECT 15.710 2405.260 24.770 2405.400 ;
        RECT 15.710 2405.200 16.030 2405.260 ;
        RECT 24.450 2405.200 24.770 2405.260 ;
        RECT 24.450 945.100 24.770 945.160 ;
        RECT 656.030 945.100 656.350 945.160 ;
        RECT 24.450 944.960 656.350 945.100 ;
        RECT 24.450 944.900 24.770 944.960 ;
        RECT 656.030 944.900 656.350 944.960 ;
      LAYER via ;
        RECT 15.740 2405.200 16.000 2405.460 ;
        RECT 24.480 2405.200 24.740 2405.460 ;
        RECT 24.480 944.900 24.740 945.160 ;
        RECT 656.060 944.900 656.320 945.160 ;
      LAYER met2 ;
        RECT 15.730 2405.315 16.010 2405.685 ;
        RECT 15.740 2405.170 16.000 2405.315 ;
        RECT 24.480 2405.170 24.740 2405.490 ;
        RECT 24.540 945.190 24.680 2405.170 ;
        RECT 24.480 944.870 24.740 945.190 ;
        RECT 656.060 944.870 656.320 945.190 ;
        RECT 656.120 943.685 656.260 944.870 ;
        RECT 656.050 943.315 656.330 943.685 ;
      LAYER via2 ;
        RECT 15.730 2405.360 16.010 2405.640 ;
        RECT 656.050 943.360 656.330 943.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 15.705 2405.650 16.035 2405.665 ;
        RECT -4.800 2405.350 16.035 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 15.705 2405.335 16.035 2405.350 ;
        RECT 656.025 943.650 656.355 943.665 ;
        RECT 670.000 943.650 674.000 944.040 ;
        RECT 656.025 943.440 674.000 943.650 ;
        RECT 656.025 943.350 670.220 943.440 ;
        RECT 656.025 943.335 656.355 943.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 952.240 16.490 952.300 ;
        RECT 656.030 952.240 656.350 952.300 ;
        RECT 16.170 952.100 656.350 952.240 ;
        RECT 16.170 952.040 16.490 952.100 ;
        RECT 656.030 952.040 656.350 952.100 ;
      LAYER via ;
        RECT 16.200 952.040 16.460 952.300 ;
        RECT 656.060 952.040 656.320 952.300 ;
      LAYER met2 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
        RECT 16.260 952.330 16.400 2118.355 ;
        RECT 16.200 952.010 16.460 952.330 ;
        RECT 656.060 952.010 656.320 952.330 ;
        RECT 656.120 949.125 656.260 952.010 ;
        RECT 656.050 948.755 656.330 949.125 ;
      LAYER via2 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
        RECT 656.050 948.800 656.330 949.080 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
        RECT 656.025 949.090 656.355 949.105 ;
        RECT 670.000 949.090 674.000 949.480 ;
        RECT 656.025 948.880 674.000 949.090 ;
        RECT 656.025 948.790 670.220 948.880 ;
        RECT 656.025 948.775 656.355 948.790 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 1830.800 15.110 1830.860 ;
        RECT 24.910 1830.800 25.230 1830.860 ;
        RECT 14.790 1830.660 25.230 1830.800 ;
        RECT 14.790 1830.600 15.110 1830.660 ;
        RECT 24.910 1830.600 25.230 1830.660 ;
        RECT 24.910 959.040 25.230 959.100 ;
        RECT 656.030 959.040 656.350 959.100 ;
        RECT 24.910 958.900 656.350 959.040 ;
        RECT 24.910 958.840 25.230 958.900 ;
        RECT 656.030 958.840 656.350 958.900 ;
      LAYER via ;
        RECT 14.820 1830.600 15.080 1830.860 ;
        RECT 24.940 1830.600 25.200 1830.860 ;
        RECT 24.940 958.840 25.200 959.100 ;
        RECT 656.060 958.840 656.320 959.100 ;
      LAYER met2 ;
        RECT 14.810 1830.715 15.090 1831.085 ;
        RECT 14.820 1830.570 15.080 1830.715 ;
        RECT 24.940 1830.570 25.200 1830.890 ;
        RECT 25.000 959.130 25.140 1830.570 ;
        RECT 24.940 958.810 25.200 959.130 ;
        RECT 656.060 958.810 656.320 959.130 ;
        RECT 656.120 954.565 656.260 958.810 ;
        RECT 656.050 954.195 656.330 954.565 ;
      LAYER via2 ;
        RECT 14.810 1830.760 15.090 1831.040 ;
        RECT 656.050 954.240 656.330 954.520 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 14.785 1831.050 15.115 1831.065 ;
        RECT -4.800 1830.750 15.115 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 14.785 1830.735 15.115 1830.750 ;
        RECT 656.025 954.530 656.355 954.545 ;
        RECT 670.000 954.530 674.000 954.920 ;
        RECT 656.025 954.320 674.000 954.530 ;
        RECT 656.025 954.230 670.220 954.320 ;
        RECT 656.025 954.215 656.355 954.230 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 603.400 662.330 603.460 ;
        RECT 2901.290 603.400 2901.610 603.460 ;
        RECT 662.010 603.260 2901.610 603.400 ;
        RECT 662.010 603.200 662.330 603.260 ;
        RECT 2901.290 603.200 2901.610 603.260 ;
      LAYER via ;
        RECT 662.040 603.200 662.300 603.460 ;
        RECT 2901.320 603.200 2901.580 603.460 ;
      LAYER met2 ;
        RECT 662.030 812.075 662.310 812.445 ;
        RECT 662.100 603.490 662.240 812.075 ;
        RECT 2901.310 674.035 2901.590 674.405 ;
        RECT 2901.380 603.490 2901.520 674.035 ;
        RECT 662.040 603.170 662.300 603.490 ;
        RECT 2901.320 603.170 2901.580 603.490 ;
      LAYER via2 ;
        RECT 662.030 812.120 662.310 812.400 ;
        RECT 2901.310 674.080 2901.590 674.360 ;
      LAYER met3 ;
        RECT 662.005 812.410 662.335 812.425 ;
        RECT 670.000 812.410 674.000 812.800 ;
        RECT 662.005 812.200 674.000 812.410 ;
        RECT 662.005 812.110 670.220 812.200 ;
        RECT 662.005 812.095 662.335 812.110 ;
        RECT 2901.285 674.370 2901.615 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2901.285 674.070 2924.800 674.370 ;
        RECT 2901.285 674.055 2901.615 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 1539.080 15.110 1539.140 ;
        RECT 25.830 1539.080 26.150 1539.140 ;
        RECT 14.790 1538.940 26.150 1539.080 ;
        RECT 14.790 1538.880 15.110 1538.940 ;
        RECT 25.830 1538.880 26.150 1538.940 ;
        RECT 25.830 965.840 26.150 965.900 ;
        RECT 25.830 965.700 656.720 965.840 ;
        RECT 25.830 965.640 26.150 965.700 ;
        RECT 656.030 964.140 656.350 964.200 ;
        RECT 656.580 964.140 656.720 965.700 ;
        RECT 656.030 964.000 656.720 964.140 ;
        RECT 656.030 963.940 656.350 964.000 ;
      LAYER via ;
        RECT 14.820 1538.880 15.080 1539.140 ;
        RECT 25.860 1538.880 26.120 1539.140 ;
        RECT 25.860 965.640 26.120 965.900 ;
        RECT 656.060 963.940 656.320 964.200 ;
      LAYER met2 ;
        RECT 14.810 1543.755 15.090 1544.125 ;
        RECT 14.880 1539.170 15.020 1543.755 ;
        RECT 14.820 1538.850 15.080 1539.170 ;
        RECT 25.860 1538.850 26.120 1539.170 ;
        RECT 25.920 965.930 26.060 1538.850 ;
        RECT 25.860 965.610 26.120 965.930 ;
        RECT 656.060 963.910 656.320 964.230 ;
        RECT 656.120 960.005 656.260 963.910 ;
        RECT 656.050 959.635 656.330 960.005 ;
      LAYER via2 ;
        RECT 14.810 1543.800 15.090 1544.080 ;
        RECT 656.050 959.680 656.330 959.960 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 14.785 1544.090 15.115 1544.105 ;
        RECT -4.800 1543.790 15.115 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 14.785 1543.775 15.115 1543.790 ;
        RECT 656.025 959.970 656.355 959.985 ;
        RECT 670.000 959.970 674.000 960.360 ;
        RECT 656.025 959.760 674.000 959.970 ;
        RECT 656.025 959.670 670.220 959.760 ;
        RECT 656.025 959.655 656.355 959.670 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 1324.880 14.650 1324.940 ;
        RECT 26.290 1324.880 26.610 1324.940 ;
        RECT 14.330 1324.740 26.610 1324.880 ;
        RECT 14.330 1324.680 14.650 1324.740 ;
        RECT 26.290 1324.680 26.610 1324.740 ;
        RECT 26.290 965.500 26.610 965.560 ;
        RECT 656.030 965.500 656.350 965.560 ;
        RECT 26.290 965.360 656.350 965.500 ;
        RECT 26.290 965.300 26.610 965.360 ;
        RECT 656.030 965.300 656.350 965.360 ;
      LAYER via ;
        RECT 14.360 1324.680 14.620 1324.940 ;
        RECT 26.320 1324.680 26.580 1324.940 ;
        RECT 26.320 965.300 26.580 965.560 ;
        RECT 656.060 965.300 656.320 965.560 ;
      LAYER met2 ;
        RECT 14.350 1328.195 14.630 1328.565 ;
        RECT 14.420 1324.970 14.560 1328.195 ;
        RECT 14.360 1324.650 14.620 1324.970 ;
        RECT 26.320 1324.650 26.580 1324.970 ;
        RECT 26.380 965.590 26.520 1324.650 ;
        RECT 26.320 965.270 26.580 965.590 ;
        RECT 656.060 965.270 656.320 965.590 ;
        RECT 656.120 964.765 656.260 965.270 ;
        RECT 656.050 964.395 656.330 964.765 ;
      LAYER via2 ;
        RECT 14.350 1328.240 14.630 1328.520 ;
        RECT 656.050 964.440 656.330 964.720 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 14.325 1328.530 14.655 1328.545 ;
        RECT -4.800 1328.230 14.655 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 14.325 1328.215 14.655 1328.230 ;
        RECT 656.025 964.730 656.355 964.745 ;
        RECT 670.000 964.730 674.000 965.120 ;
        RECT 656.025 964.520 674.000 964.730 ;
        RECT 656.025 964.430 670.220 964.520 ;
        RECT 656.025 964.415 656.355 964.430 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 1112.720 14.190 1112.780 ;
        RECT 30.890 1112.720 31.210 1112.780 ;
        RECT 13.870 1112.580 31.210 1112.720 ;
        RECT 13.870 1112.520 14.190 1112.580 ;
        RECT 30.890 1112.520 31.210 1112.580 ;
        RECT 30.890 972.300 31.210 972.360 ;
        RECT 656.030 972.300 656.350 972.360 ;
        RECT 30.890 972.160 656.350 972.300 ;
        RECT 30.890 972.100 31.210 972.160 ;
        RECT 656.030 972.100 656.350 972.160 ;
      LAYER via ;
        RECT 13.900 1112.520 14.160 1112.780 ;
        RECT 30.920 1112.520 31.180 1112.780 ;
        RECT 30.920 972.100 31.180 972.360 ;
        RECT 656.060 972.100 656.320 972.360 ;
      LAYER met2 ;
        RECT 13.890 1112.635 14.170 1113.005 ;
        RECT 13.900 1112.490 14.160 1112.635 ;
        RECT 30.920 1112.490 31.180 1112.810 ;
        RECT 30.980 972.390 31.120 1112.490 ;
        RECT 30.920 972.070 31.180 972.390 ;
        RECT 656.060 972.070 656.320 972.390 ;
        RECT 656.120 970.205 656.260 972.070 ;
        RECT 656.050 969.835 656.330 970.205 ;
      LAYER via2 ;
        RECT 13.890 1112.680 14.170 1112.960 ;
        RECT 656.050 969.880 656.330 970.160 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 13.865 1112.970 14.195 1112.985 ;
        RECT -4.800 1112.670 14.195 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 13.865 1112.655 14.195 1112.670 ;
        RECT 656.025 970.170 656.355 970.185 ;
        RECT 670.000 970.170 674.000 970.560 ;
        RECT 656.025 969.960 674.000 970.170 ;
        RECT 656.025 969.870 670.220 969.960 ;
        RECT 656.025 969.855 656.355 969.870 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 44.690 972.980 45.010 973.040 ;
        RECT 656.030 972.980 656.350 973.040 ;
        RECT 44.690 972.840 656.350 972.980 ;
        RECT 44.690 972.780 45.010 972.840 ;
        RECT 656.030 972.780 656.350 972.840 ;
        RECT 18.470 897.500 18.790 897.560 ;
        RECT 44.690 897.500 45.010 897.560 ;
        RECT 18.470 897.360 45.010 897.500 ;
        RECT 18.470 897.300 18.790 897.360 ;
        RECT 44.690 897.300 45.010 897.360 ;
      LAYER via ;
        RECT 44.720 972.780 44.980 973.040 ;
        RECT 656.060 972.780 656.320 973.040 ;
        RECT 18.500 897.300 18.760 897.560 ;
        RECT 44.720 897.300 44.980 897.560 ;
      LAYER met2 ;
        RECT 656.050 975.275 656.330 975.645 ;
        RECT 656.120 973.070 656.260 975.275 ;
        RECT 44.720 972.750 44.980 973.070 ;
        RECT 656.060 972.750 656.320 973.070 ;
        RECT 44.780 897.590 44.920 972.750 ;
        RECT 18.500 897.445 18.760 897.590 ;
        RECT 18.490 897.075 18.770 897.445 ;
        RECT 44.720 897.270 44.980 897.590 ;
      LAYER via2 ;
        RECT 656.050 975.320 656.330 975.600 ;
        RECT 18.490 897.120 18.770 897.400 ;
      LAYER met3 ;
        RECT 656.025 975.610 656.355 975.625 ;
        RECT 670.000 975.610 674.000 976.000 ;
        RECT 656.025 975.400 674.000 975.610 ;
        RECT 656.025 975.310 670.220 975.400 ;
        RECT 656.025 975.295 656.355 975.310 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 18.465 897.410 18.795 897.425 ;
        RECT -4.800 897.110 18.795 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 18.465 897.095 18.795 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.750 980.120 27.070 980.180 ;
        RECT 656.030 980.120 656.350 980.180 ;
        RECT 26.750 979.980 656.350 980.120 ;
        RECT 26.750 979.920 27.070 979.980 ;
        RECT 656.030 979.920 656.350 979.980 ;
        RECT 13.870 681.940 14.190 682.000 ;
        RECT 26.750 681.940 27.070 682.000 ;
        RECT 13.870 681.800 27.070 681.940 ;
        RECT 13.870 681.740 14.190 681.800 ;
        RECT 26.750 681.740 27.070 681.800 ;
      LAYER via ;
        RECT 26.780 979.920 27.040 980.180 ;
        RECT 656.060 979.920 656.320 980.180 ;
        RECT 13.900 681.740 14.160 682.000 ;
        RECT 26.780 681.740 27.040 682.000 ;
      LAYER met2 ;
        RECT 26.780 979.890 27.040 980.210 ;
        RECT 656.050 980.035 656.330 980.405 ;
        RECT 656.060 979.890 656.320 980.035 ;
        RECT 26.840 682.030 26.980 979.890 ;
        RECT 13.900 681.885 14.160 682.030 ;
        RECT 13.890 681.515 14.170 681.885 ;
        RECT 26.780 681.710 27.040 682.030 ;
      LAYER via2 ;
        RECT 656.050 980.080 656.330 980.360 ;
        RECT 13.890 681.560 14.170 681.840 ;
      LAYER met3 ;
        RECT 670.000 981.050 674.000 981.440 ;
        RECT 656.270 980.840 674.000 981.050 ;
        RECT 656.270 980.750 670.220 980.840 ;
        RECT 656.270 980.385 656.570 980.750 ;
        RECT 656.025 980.070 656.570 980.385 ;
        RECT 656.025 980.055 656.355 980.070 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 13.865 681.850 14.195 681.865 ;
        RECT -4.800 681.550 14.195 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 13.865 681.535 14.195 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.490 981.820 656.810 981.880 ;
        RECT 656.490 981.680 657.180 981.820 ;
        RECT 656.490 981.620 656.810 981.680 ;
        RECT 72.290 980.460 72.610 980.520 ;
        RECT 657.040 980.460 657.180 981.680 ;
        RECT 72.290 980.320 657.180 980.460 ;
        RECT 72.290 980.260 72.610 980.320 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 72.290 469.100 72.610 469.160 ;
        RECT 17.090 468.960 72.610 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 72.290 468.900 72.610 468.960 ;
      LAYER via ;
        RECT 656.520 981.620 656.780 981.880 ;
        RECT 72.320 980.260 72.580 980.520 ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 72.320 468.900 72.580 469.160 ;
      LAYER met2 ;
        RECT 656.510 985.475 656.790 985.845 ;
        RECT 656.580 981.910 656.720 985.475 ;
        RECT 656.520 981.590 656.780 981.910 ;
        RECT 72.320 980.230 72.580 980.550 ;
        RECT 72.380 469.190 72.520 980.230 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 72.320 468.870 72.580 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 656.510 985.520 656.790 985.800 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 656.485 985.810 656.815 985.825 ;
        RECT 670.000 985.810 674.000 986.200 ;
        RECT 656.485 985.600 674.000 985.810 ;
        RECT 656.485 985.510 670.220 985.600 ;
        RECT 656.485 985.495 656.815 985.510 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 986.920 20.630 986.980 ;
        RECT 656.030 986.920 656.350 986.980 ;
        RECT 20.310 986.780 656.350 986.920 ;
        RECT 20.310 986.720 20.630 986.780 ;
        RECT 656.030 986.720 656.350 986.780 ;
      LAYER via ;
        RECT 20.340 986.720 20.600 986.980 ;
        RECT 656.060 986.720 656.320 986.980 ;
      LAYER met2 ;
        RECT 656.050 990.915 656.330 991.285 ;
        RECT 656.120 987.010 656.260 990.915 ;
        RECT 20.340 986.690 20.600 987.010 ;
        RECT 656.060 986.690 656.320 987.010 ;
        RECT 20.400 250.765 20.540 986.690 ;
        RECT 20.330 250.395 20.610 250.765 ;
      LAYER via2 ;
        RECT 656.050 990.960 656.330 991.240 ;
        RECT 20.330 250.440 20.610 250.720 ;
      LAYER met3 ;
        RECT 656.025 991.250 656.355 991.265 ;
        RECT 670.000 991.250 674.000 991.640 ;
        RECT 656.025 991.040 674.000 991.250 ;
        RECT 656.025 990.950 670.220 991.040 ;
        RECT 656.025 990.935 656.355 990.950 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 20.305 250.730 20.635 250.745 ;
        RECT -4.800 250.430 20.635 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 20.305 250.415 20.635 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.390 993.720 19.710 993.780 ;
        RECT 656.030 993.720 656.350 993.780 ;
        RECT 19.390 993.580 656.350 993.720 ;
        RECT 19.390 993.520 19.710 993.580 ;
        RECT 656.030 993.520 656.350 993.580 ;
      LAYER via ;
        RECT 19.420 993.520 19.680 993.780 ;
        RECT 656.060 993.520 656.320 993.780 ;
      LAYER met2 ;
        RECT 656.050 996.355 656.330 996.725 ;
        RECT 656.120 993.810 656.260 996.355 ;
        RECT 19.420 993.490 19.680 993.810 ;
        RECT 656.060 993.490 656.320 993.810 ;
        RECT 19.480 35.885 19.620 993.490 ;
        RECT 19.410 35.515 19.690 35.885 ;
      LAYER via2 ;
        RECT 656.050 996.400 656.330 996.680 ;
        RECT 19.410 35.560 19.690 35.840 ;
      LAYER met3 ;
        RECT 656.025 996.690 656.355 996.705 ;
        RECT 670.000 996.690 674.000 997.080 ;
        RECT 656.025 996.480 674.000 996.690 ;
        RECT 656.025 996.390 670.220 996.480 ;
        RECT 656.025 996.375 656.355 996.390 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 19.385 35.850 19.715 35.865 ;
        RECT -4.800 35.550 19.715 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 19.385 35.535 19.715 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 668.910 1000.860 669.230 1000.920 ;
        RECT 2899.910 1000.860 2900.230 1000.920 ;
        RECT 668.910 1000.720 2900.230 1000.860 ;
        RECT 668.910 1000.660 669.230 1000.720 ;
        RECT 2899.910 1000.660 2900.230 1000.720 ;
        RECT 667.530 948.840 667.850 948.900 ;
        RECT 668.910 948.840 669.230 948.900 ;
        RECT 667.530 948.700 669.230 948.840 ;
        RECT 667.530 948.640 667.850 948.700 ;
        RECT 668.910 948.640 669.230 948.700 ;
      LAYER via ;
        RECT 668.940 1000.660 669.200 1000.920 ;
        RECT 2899.940 1000.660 2900.200 1000.920 ;
        RECT 667.560 948.640 667.820 948.900 ;
        RECT 668.940 948.640 669.200 948.900 ;
      LAYER met2 ;
        RECT 668.940 1000.630 669.200 1000.950 ;
        RECT 2899.940 1000.630 2900.200 1000.950 ;
        RECT 669.000 948.930 669.140 1000.630 ;
        RECT 667.560 948.610 667.820 948.930 ;
        RECT 668.940 948.610 669.200 948.930 ;
        RECT 667.620 817.885 667.760 948.610 ;
        RECT 2900.000 909.685 2900.140 1000.630 ;
        RECT 2899.930 909.315 2900.210 909.685 ;
        RECT 667.550 817.515 667.830 817.885 ;
      LAYER via2 ;
        RECT 2899.930 909.360 2900.210 909.640 ;
        RECT 667.550 817.560 667.830 817.840 ;
      LAYER met3 ;
        RECT 2899.905 909.650 2900.235 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2899.905 909.350 2924.800 909.650 ;
        RECT 2899.905 909.335 2900.235 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT 667.525 817.850 667.855 817.865 ;
        RECT 670.000 817.850 674.000 818.240 ;
        RECT 667.525 817.640 674.000 817.850 ;
        RECT 667.525 817.550 670.220 817.640 ;
        RECT 667.525 817.535 667.855 817.550 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 663.390 1138.900 663.710 1138.960 ;
        RECT 2900.370 1138.900 2900.690 1138.960 ;
        RECT 663.390 1138.760 2900.690 1138.900 ;
        RECT 663.390 1138.700 663.710 1138.760 ;
        RECT 2900.370 1138.700 2900.690 1138.760 ;
      LAYER via ;
        RECT 663.420 1138.700 663.680 1138.960 ;
        RECT 2900.400 1138.700 2900.660 1138.960 ;
      LAYER met2 ;
        RECT 2900.390 1143.915 2900.670 1144.285 ;
        RECT 2900.460 1138.990 2900.600 1143.915 ;
        RECT 663.420 1138.670 663.680 1138.990 ;
        RECT 2900.400 1138.670 2900.660 1138.990 ;
        RECT 663.480 822.645 663.620 1138.670 ;
        RECT 663.410 822.275 663.690 822.645 ;
      LAYER via2 ;
        RECT 2900.390 1143.960 2900.670 1144.240 ;
        RECT 663.410 822.320 663.690 822.600 ;
      LAYER met3 ;
        RECT 2900.365 1144.250 2900.695 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.365 1143.950 2924.800 1144.250 ;
        RECT 2900.365 1143.935 2900.695 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 663.385 822.610 663.715 822.625 ;
        RECT 670.000 822.610 674.000 823.000 ;
        RECT 663.385 822.400 674.000 822.610 ;
        RECT 663.385 822.310 670.220 822.400 ;
        RECT 663.385 822.295 663.715 822.310 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 657.870 1373.500 658.190 1373.560 ;
        RECT 2899.910 1373.500 2900.230 1373.560 ;
        RECT 657.870 1373.360 2900.230 1373.500 ;
        RECT 657.870 1373.300 658.190 1373.360 ;
        RECT 2899.910 1373.300 2900.230 1373.360 ;
      LAYER via ;
        RECT 657.900 1373.300 658.160 1373.560 ;
        RECT 2899.940 1373.300 2900.200 1373.560 ;
      LAYER met2 ;
        RECT 2899.930 1378.515 2900.210 1378.885 ;
        RECT 2900.000 1373.590 2900.140 1378.515 ;
        RECT 657.900 1373.270 658.160 1373.590 ;
        RECT 2899.940 1373.270 2900.200 1373.590 ;
        RECT 657.960 828.085 658.100 1373.270 ;
        RECT 657.890 827.715 658.170 828.085 ;
      LAYER via2 ;
        RECT 2899.930 1378.560 2900.210 1378.840 ;
        RECT 657.890 827.760 658.170 828.040 ;
      LAYER met3 ;
        RECT 2899.905 1378.850 2900.235 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2899.905 1378.550 2924.800 1378.850 ;
        RECT 2899.905 1378.535 2900.235 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 657.865 828.050 658.195 828.065 ;
        RECT 670.000 828.050 674.000 828.440 ;
        RECT 657.865 827.840 674.000 828.050 ;
        RECT 657.865 827.750 670.220 827.840 ;
        RECT 657.865 827.735 658.195 827.750 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 650.050 1608.100 650.370 1608.160 ;
        RECT 2900.830 1608.100 2901.150 1608.160 ;
        RECT 650.050 1607.960 2901.150 1608.100 ;
        RECT 650.050 1607.900 650.370 1607.960 ;
        RECT 2900.830 1607.900 2901.150 1607.960 ;
        RECT 650.050 834.260 650.370 834.320 ;
        RECT 660.170 834.260 660.490 834.320 ;
        RECT 650.050 834.120 660.490 834.260 ;
        RECT 650.050 834.060 650.370 834.120 ;
        RECT 660.170 834.060 660.490 834.120 ;
      LAYER via ;
        RECT 650.080 1607.900 650.340 1608.160 ;
        RECT 2900.860 1607.900 2901.120 1608.160 ;
        RECT 650.080 834.060 650.340 834.320 ;
        RECT 660.200 834.060 660.460 834.320 ;
      LAYER met2 ;
        RECT 2900.850 1613.115 2901.130 1613.485 ;
        RECT 2900.920 1608.190 2901.060 1613.115 ;
        RECT 650.080 1607.870 650.340 1608.190 ;
        RECT 2900.860 1607.870 2901.120 1608.190 ;
        RECT 650.140 834.350 650.280 1607.870 ;
        RECT 650.080 834.030 650.340 834.350 ;
        RECT 660.200 834.030 660.460 834.350 ;
        RECT 660.260 833.525 660.400 834.030 ;
        RECT 660.190 833.155 660.470 833.525 ;
      LAYER via2 ;
        RECT 2900.850 1613.160 2901.130 1613.440 ;
        RECT 660.190 833.200 660.470 833.480 ;
      LAYER met3 ;
        RECT 2900.825 1613.450 2901.155 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.825 1613.150 2924.800 1613.450 ;
        RECT 2900.825 1613.135 2901.155 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 660.165 833.490 660.495 833.505 ;
        RECT 670.000 833.490 674.000 833.880 ;
        RECT 660.165 833.280 674.000 833.490 ;
        RECT 660.165 833.190 670.220 833.280 ;
        RECT 660.165 833.175 660.495 833.190 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 1004.940 662.330 1005.000 ;
        RECT 2903.590 1004.940 2903.910 1005.000 ;
        RECT 662.010 1004.800 2903.910 1004.940 ;
        RECT 662.010 1004.740 662.330 1004.800 ;
        RECT 2903.590 1004.740 2903.910 1004.800 ;
      LAYER via ;
        RECT 662.040 1004.740 662.300 1005.000 ;
        RECT 2903.620 1004.740 2903.880 1005.000 ;
      LAYER met2 ;
        RECT 2903.610 1847.715 2903.890 1848.085 ;
        RECT 2903.680 1005.030 2903.820 1847.715 ;
        RECT 662.040 1004.710 662.300 1005.030 ;
        RECT 2903.620 1004.710 2903.880 1005.030 ;
        RECT 662.100 838.965 662.240 1004.710 ;
        RECT 662.030 838.595 662.310 838.965 ;
      LAYER via2 ;
        RECT 2903.610 1847.760 2903.890 1848.040 ;
        RECT 662.030 838.640 662.310 838.920 ;
      LAYER met3 ;
        RECT 2903.585 1848.050 2903.915 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2903.585 1847.750 2924.800 1848.050 ;
        RECT 2903.585 1847.735 2903.915 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 662.005 838.930 662.335 838.945 ;
        RECT 670.000 838.930 674.000 839.320 ;
        RECT 662.005 838.720 674.000 838.930 ;
        RECT 662.005 838.630 670.220 838.720 ;
        RECT 662.005 838.615 662.335 838.630 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 664.770 2077.300 665.090 2077.360 ;
        RECT 2898.990 2077.300 2899.310 2077.360 ;
        RECT 664.770 2077.160 2899.310 2077.300 ;
        RECT 664.770 2077.100 665.090 2077.160 ;
        RECT 2898.990 2077.100 2899.310 2077.160 ;
      LAYER via ;
        RECT 664.800 2077.100 665.060 2077.360 ;
        RECT 2899.020 2077.100 2899.280 2077.360 ;
      LAYER met2 ;
        RECT 2899.010 2082.315 2899.290 2082.685 ;
        RECT 2899.080 2077.390 2899.220 2082.315 ;
        RECT 664.800 2077.070 665.060 2077.390 ;
        RECT 2899.020 2077.070 2899.280 2077.390 ;
        RECT 664.860 843.725 665.000 2077.070 ;
        RECT 664.790 843.355 665.070 843.725 ;
      LAYER via2 ;
        RECT 2899.010 2082.360 2899.290 2082.640 ;
        RECT 664.790 843.400 665.070 843.680 ;
      LAYER met3 ;
        RECT 2898.985 2082.650 2899.315 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2898.985 2082.350 2924.800 2082.650 ;
        RECT 2898.985 2082.335 2899.315 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 664.765 843.690 665.095 843.705 ;
        RECT 670.000 843.690 674.000 844.080 ;
        RECT 664.765 843.480 674.000 843.690 ;
        RECT 664.765 843.390 670.220 843.480 ;
        RECT 664.765 843.375 665.095 843.390 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 652.810 2311.900 653.130 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 652.810 2311.760 2901.150 2311.900 ;
        RECT 652.810 2311.700 653.130 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
      LAYER via ;
        RECT 652.840 2311.700 653.100 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 652.840 2311.670 653.100 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 652.900 849.165 653.040 2311.670 ;
        RECT 652.830 848.795 653.110 849.165 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 652.830 848.840 653.110 849.120 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 652.805 849.130 653.135 849.145 ;
        RECT 670.000 849.130 674.000 849.520 ;
        RECT 652.805 848.920 674.000 849.130 ;
        RECT 652.805 848.830 670.220 848.920 ;
        RECT 652.805 848.815 653.135 848.830 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 660.630 151.540 660.950 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 660.630 151.400 2901.150 151.540 ;
        RECT 660.630 151.340 660.950 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 660.660 151.340 660.920 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 660.650 601.955 660.930 602.325 ;
        RECT 660.720 151.630 660.860 601.955 ;
        RECT 660.660 151.310 660.920 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 660.650 602.000 660.930 602.280 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 660.625 602.290 660.955 602.305 ;
        RECT 670.000 602.290 674.000 602.680 ;
        RECT 660.625 602.080 674.000 602.290 ;
        RECT 660.625 601.990 670.220 602.080 ;
        RECT 660.625 601.975 660.955 601.990 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 659.250 2491.080 659.570 2491.140 ;
        RECT 2899.450 2491.080 2899.770 2491.140 ;
        RECT 659.250 2490.940 2899.770 2491.080 ;
        RECT 659.250 2490.880 659.570 2490.940 ;
        RECT 2899.450 2490.880 2899.770 2490.940 ;
      LAYER via ;
        RECT 659.280 2490.880 659.540 2491.140 ;
        RECT 2899.480 2490.880 2899.740 2491.140 ;
      LAYER met2 ;
        RECT 2899.470 2493.035 2899.750 2493.405 ;
        RECT 2899.540 2491.170 2899.680 2493.035 ;
        RECT 659.280 2490.850 659.540 2491.170 ;
        RECT 2899.480 2490.850 2899.740 2491.170 ;
        RECT 659.340 654.685 659.480 2490.850 ;
        RECT 659.270 654.315 659.550 654.685 ;
      LAYER via2 ;
        RECT 2899.470 2493.080 2899.750 2493.360 ;
        RECT 659.270 654.360 659.550 654.640 ;
      LAYER met3 ;
        RECT 2899.445 2493.370 2899.775 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2899.445 2493.070 2924.800 2493.370 ;
        RECT 2899.445 2493.055 2899.775 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 659.245 654.650 659.575 654.665 ;
        RECT 670.000 654.650 674.000 655.040 ;
        RECT 659.245 654.440 674.000 654.650 ;
        RECT 659.245 654.350 670.220 654.440 ;
        RECT 659.245 654.335 659.575 654.350 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.490 1004.600 656.810 1004.660 ;
        RECT 2901.750 1004.600 2902.070 1004.660 ;
        RECT 656.490 1004.460 2902.070 1004.600 ;
        RECT 656.490 1004.400 656.810 1004.460 ;
        RECT 2901.750 1004.400 2902.070 1004.460 ;
      LAYER via ;
        RECT 656.520 1004.400 656.780 1004.660 ;
        RECT 2901.780 1004.400 2902.040 1004.660 ;
      LAYER met2 ;
        RECT 2901.770 2727.635 2902.050 2728.005 ;
        RECT 2901.840 1004.690 2901.980 2727.635 ;
        RECT 656.520 1004.370 656.780 1004.690 ;
        RECT 2901.780 1004.370 2902.040 1004.690 ;
        RECT 656.580 986.410 656.720 1004.370 ;
        RECT 656.120 986.270 656.720 986.410 ;
        RECT 656.120 980.970 656.260 986.270 ;
        RECT 656.120 980.830 656.720 980.970 ;
        RECT 656.580 660.125 656.720 980.830 ;
        RECT 656.510 659.755 656.790 660.125 ;
      LAYER via2 ;
        RECT 2901.770 2727.680 2902.050 2727.960 ;
        RECT 656.510 659.800 656.790 660.080 ;
      LAYER met3 ;
        RECT 2901.745 2727.970 2902.075 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2901.745 2727.670 2924.800 2727.970 ;
        RECT 2901.745 2727.655 2902.075 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 656.485 660.090 656.815 660.105 ;
        RECT 670.000 660.090 674.000 660.480 ;
        RECT 656.485 659.880 674.000 660.090 ;
        RECT 656.485 659.790 670.220 659.880 ;
        RECT 656.485 659.775 656.815 659.790 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 669.830 2960.280 670.150 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 669.830 2960.140 2901.150 2960.280 ;
        RECT 669.830 2960.080 670.150 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 669.860 2960.080 670.120 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 669.860 2960.050 670.120 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 669.920 667.605 670.060 2960.050 ;
        RECT 669.850 667.235 670.130 667.605 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
        RECT 669.850 667.280 670.130 667.560 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 669.825 667.570 670.155 667.585 ;
        RECT 669.825 667.255 670.370 667.570 ;
        RECT 670.070 665.240 670.370 667.255 ;
        RECT 670.000 664.640 674.000 665.240 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 659.710 3194.880 660.030 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 659.710 3194.740 2901.150 3194.880 ;
        RECT 659.710 3194.680 660.030 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 659.740 3194.680 660.000 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 659.740 3194.650 660.000 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 659.800 670.325 659.940 3194.650 ;
        RECT 659.730 669.955 660.010 670.325 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 659.730 670.000 660.010 670.280 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 659.705 670.290 660.035 670.305 ;
        RECT 670.000 670.290 674.000 670.680 ;
        RECT 659.705 670.080 674.000 670.290 ;
        RECT 659.705 669.990 670.220 670.080 ;
        RECT 659.705 669.975 660.035 669.990 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 660.630 3429.480 660.950 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 660.630 3429.340 2901.150 3429.480 ;
        RECT 660.630 3429.280 660.950 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 660.660 3429.280 660.920 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 660.660 3429.250 660.920 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 660.720 675.765 660.860 3429.250 ;
        RECT 660.650 675.395 660.930 675.765 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 660.650 675.440 660.930 675.720 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 660.625 675.730 660.955 675.745 ;
        RECT 670.000 675.730 674.000 676.120 ;
        RECT 660.625 675.520 674.000 675.730 ;
        RECT 660.625 675.430 670.220 675.520 ;
        RECT 660.625 675.415 660.955 675.430 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.470 3501.560 662.790 3501.620 ;
        RECT 2717.290 3501.560 2717.610 3501.620 ;
        RECT 662.470 3501.420 2717.610 3501.560 ;
        RECT 662.470 3501.360 662.790 3501.420 ;
        RECT 2717.290 3501.360 2717.610 3501.420 ;
      LAYER via ;
        RECT 662.500 3501.360 662.760 3501.620 ;
        RECT 2717.320 3501.360 2717.580 3501.620 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.650 2717.520 3517.600 ;
        RECT 662.500 3501.330 662.760 3501.650 ;
        RECT 2717.320 3501.330 2717.580 3501.650 ;
        RECT 662.560 681.205 662.700 3501.330 ;
        RECT 662.490 680.835 662.770 681.205 ;
      LAYER via2 ;
        RECT 662.490 680.880 662.770 681.160 ;
      LAYER met3 ;
        RECT 662.465 681.170 662.795 681.185 ;
        RECT 670.000 681.170 674.000 681.560 ;
        RECT 662.465 680.960 674.000 681.170 ;
        RECT 662.465 680.870 670.220 680.960 ;
        RECT 662.465 680.855 662.795 680.870 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 668.450 3502.580 668.770 3502.640 ;
        RECT 2392.530 3502.580 2392.850 3502.640 ;
        RECT 668.450 3502.440 2392.850 3502.580 ;
        RECT 668.450 3502.380 668.770 3502.440 ;
        RECT 2392.530 3502.380 2392.850 3502.440 ;
      LAYER via ;
        RECT 668.480 3502.380 668.740 3502.640 ;
        RECT 2392.560 3502.380 2392.820 3502.640 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3502.670 2392.760 3517.600 ;
        RECT 668.480 3502.350 668.740 3502.670 ;
        RECT 2392.560 3502.350 2392.820 3502.670 ;
        RECT 668.540 685.965 668.680 3502.350 ;
        RECT 668.470 685.595 668.750 685.965 ;
      LAYER via2 ;
        RECT 668.470 685.640 668.750 685.920 ;
      LAYER met3 ;
        RECT 668.445 685.930 668.775 685.945 ;
        RECT 670.000 685.930 674.000 686.320 ;
        RECT 668.445 685.720 674.000 685.930 ;
        RECT 668.445 685.630 670.220 685.720 ;
        RECT 668.445 685.615 668.775 685.630 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 655.570 3503.600 655.890 3503.660 ;
        RECT 2068.230 3503.600 2068.550 3503.660 ;
        RECT 655.570 3503.460 2068.550 3503.600 ;
        RECT 655.570 3503.400 655.890 3503.460 ;
        RECT 2068.230 3503.400 2068.550 3503.460 ;
        RECT 654.650 731.920 654.970 731.980 ;
        RECT 655.570 731.920 655.890 731.980 ;
        RECT 654.650 731.780 655.890 731.920 ;
        RECT 654.650 731.720 654.970 731.780 ;
        RECT 655.570 731.720 655.890 731.780 ;
      LAYER via ;
        RECT 655.600 3503.400 655.860 3503.660 ;
        RECT 2068.260 3503.400 2068.520 3503.660 ;
        RECT 654.680 731.720 654.940 731.980 ;
        RECT 655.600 731.720 655.860 731.980 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3503.690 2068.460 3517.600 ;
        RECT 655.600 3503.370 655.860 3503.690 ;
        RECT 2068.260 3503.370 2068.520 3503.690 ;
        RECT 655.660 732.010 655.800 3503.370 ;
        RECT 654.680 731.690 654.940 732.010 ;
        RECT 655.600 731.690 655.860 732.010 ;
        RECT 654.740 721.890 654.880 731.690 ;
        RECT 654.740 721.750 655.800 721.890 ;
        RECT 655.660 691.405 655.800 721.750 ;
        RECT 655.590 691.035 655.870 691.405 ;
      LAYER via2 ;
        RECT 655.590 691.080 655.870 691.360 ;
      LAYER met3 ;
        RECT 655.565 691.370 655.895 691.385 ;
        RECT 670.000 691.370 674.000 691.760 ;
        RECT 655.565 691.160 674.000 691.370 ;
        RECT 655.565 691.070 670.220 691.160 ;
        RECT 655.565 691.055 655.895 691.070 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 667.990 3504.620 668.310 3504.680 ;
        RECT 1743.930 3504.620 1744.250 3504.680 ;
        RECT 667.990 3504.480 1744.250 3504.620 ;
        RECT 667.990 3504.420 668.310 3504.480 ;
        RECT 1743.930 3504.420 1744.250 3504.480 ;
      LAYER via ;
        RECT 668.020 3504.420 668.280 3504.680 ;
        RECT 1743.960 3504.420 1744.220 3504.680 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3504.710 1744.160 3517.600 ;
        RECT 668.020 3504.390 668.280 3504.710 ;
        RECT 1743.960 3504.390 1744.220 3504.710 ;
        RECT 668.080 696.845 668.220 3504.390 ;
        RECT 668.010 696.475 668.290 696.845 ;
      LAYER via2 ;
        RECT 668.010 696.520 668.290 696.800 ;
      LAYER met3 ;
        RECT 667.985 696.810 668.315 696.825 ;
        RECT 670.000 696.810 674.000 697.200 ;
        RECT 667.985 696.600 674.000 696.810 ;
        RECT 667.985 696.510 670.220 696.600 ;
        RECT 667.985 696.495 668.315 696.510 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 661.550 3500.880 661.870 3500.940 ;
        RECT 1419.170 3500.880 1419.490 3500.940 ;
        RECT 661.550 3500.740 1419.490 3500.880 ;
        RECT 661.550 3500.680 661.870 3500.740 ;
        RECT 1419.170 3500.680 1419.490 3500.740 ;
        RECT 661.550 737.840 661.870 738.100 ;
        RECT 661.640 737.700 661.780 737.840 ;
        RECT 661.180 737.560 661.780 737.700 ;
        RECT 661.180 733.000 661.320 737.560 ;
        RECT 661.090 732.740 661.410 733.000 ;
      LAYER via ;
        RECT 661.580 3500.680 661.840 3500.940 ;
        RECT 1419.200 3500.680 1419.460 3500.940 ;
        RECT 661.580 737.840 661.840 738.100 ;
        RECT 661.120 732.740 661.380 733.000 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3500.970 1419.400 3517.600 ;
        RECT 661.580 3500.650 661.840 3500.970 ;
        RECT 1419.200 3500.650 1419.460 3500.970 ;
        RECT 661.640 738.130 661.780 3500.650 ;
        RECT 661.580 737.810 661.840 738.130 ;
        RECT 661.120 732.710 661.380 733.030 ;
        RECT 661.180 702.285 661.320 732.710 ;
        RECT 661.110 701.915 661.390 702.285 ;
      LAYER via2 ;
        RECT 661.110 701.960 661.390 702.240 ;
      LAYER met3 ;
        RECT 661.085 702.250 661.415 702.265 ;
        RECT 670.000 702.250 674.000 702.640 ;
        RECT 661.085 702.040 674.000 702.250 ;
        RECT 661.085 701.950 670.220 702.040 ;
        RECT 661.085 701.935 661.415 701.950 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 661.550 386.140 661.870 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 661.550 386.000 2901.150 386.140 ;
        RECT 661.550 385.940 661.870 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 661.580 385.940 661.840 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 661.570 606.715 661.850 607.085 ;
        RECT 661.640 386.230 661.780 606.715 ;
        RECT 661.580 385.910 661.840 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 661.570 606.760 661.850 607.040 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 661.545 607.050 661.875 607.065 ;
        RECT 670.000 607.050 674.000 607.440 ;
        RECT 661.545 606.840 674.000 607.050 ;
        RECT 661.545 606.750 670.220 606.840 ;
        RECT 661.545 606.735 661.875 606.750 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 669.370 3504.960 669.690 3505.020 ;
        RECT 1094.870 3504.960 1095.190 3505.020 ;
        RECT 669.370 3504.820 1095.190 3504.960 ;
        RECT 669.370 3504.760 669.690 3504.820 ;
        RECT 1094.870 3504.760 1095.190 3504.820 ;
      LAYER via ;
        RECT 669.400 3504.760 669.660 3505.020 ;
        RECT 1094.900 3504.760 1095.160 3505.020 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3505.050 1095.100 3517.600 ;
        RECT 669.400 3504.730 669.660 3505.050 ;
        RECT 1094.900 3504.730 1095.160 3505.050 ;
        RECT 669.460 707.045 669.600 3504.730 ;
        RECT 669.390 706.675 669.670 707.045 ;
      LAYER via2 ;
        RECT 669.390 706.720 669.670 707.000 ;
      LAYER met3 ;
        RECT 669.365 707.010 669.695 707.025 ;
        RECT 670.000 707.010 674.000 707.400 ;
        RECT 669.365 706.800 674.000 707.010 ;
        RECT 669.365 706.710 670.220 706.800 ;
        RECT 669.365 706.695 669.695 706.710 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 661.090 3503.940 661.410 3504.000 ;
        RECT 770.570 3503.940 770.890 3504.000 ;
        RECT 661.090 3503.800 770.890 3503.940 ;
        RECT 661.090 3503.740 661.410 3503.800 ;
        RECT 770.570 3503.740 770.890 3503.800 ;
      LAYER via ;
        RECT 661.120 3503.740 661.380 3504.000 ;
        RECT 770.600 3503.740 770.860 3504.000 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3504.030 770.800 3517.600 ;
        RECT 661.120 3503.710 661.380 3504.030 ;
        RECT 770.600 3503.710 770.860 3504.030 ;
        RECT 661.180 739.005 661.320 3503.710 ;
        RECT 661.110 738.635 661.390 739.005 ;
        RECT 661.570 737.275 661.850 737.645 ;
        RECT 661.640 712.485 661.780 737.275 ;
        RECT 661.570 712.115 661.850 712.485 ;
      LAYER via2 ;
        RECT 661.110 738.680 661.390 738.960 ;
        RECT 661.570 737.320 661.850 737.600 ;
        RECT 661.570 712.160 661.850 712.440 ;
      LAYER met3 ;
        RECT 661.085 738.980 661.415 738.985 ;
        RECT 660.830 738.970 661.415 738.980 ;
        RECT 660.630 738.670 661.415 738.970 ;
        RECT 660.830 738.660 661.415 738.670 ;
        RECT 661.085 738.655 661.415 738.660 ;
        RECT 660.830 737.610 661.210 737.620 ;
        RECT 661.545 737.610 661.875 737.625 ;
        RECT 660.830 737.310 661.875 737.610 ;
        RECT 660.830 737.300 661.210 737.310 ;
        RECT 661.545 737.295 661.875 737.310 ;
        RECT 661.545 712.450 661.875 712.465 ;
        RECT 670.000 712.450 674.000 712.840 ;
        RECT 661.545 712.240 674.000 712.450 ;
        RECT 661.545 712.150 670.220 712.240 ;
        RECT 661.545 712.135 661.875 712.150 ;
      LAYER via3 ;
        RECT 660.860 738.660 661.180 738.980 ;
        RECT 660.860 737.300 661.180 737.620 ;
      LAYER met4 ;
        RECT 660.855 738.655 661.185 738.985 ;
        RECT 660.870 737.625 661.170 738.655 ;
        RECT 660.855 737.295 661.185 737.625 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 2763.420 448.430 2763.480 ;
        RECT 644.990 2763.420 645.310 2763.480 ;
        RECT 448.110 2763.280 645.310 2763.420 ;
        RECT 448.110 2763.220 448.430 2763.280 ;
        RECT 644.990 2763.220 645.310 2763.280 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 2763.220 448.400 2763.480 ;
        RECT 645.020 2763.220 645.280 2763.480 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 2763.510 448.340 3498.270 ;
        RECT 448.140 2763.190 448.400 2763.510 ;
        RECT 645.020 2763.190 645.280 2763.510 ;
        RECT 645.080 717.925 645.220 2763.190 ;
        RECT 645.010 717.555 645.290 717.925 ;
      LAYER via2 ;
        RECT 645.010 717.600 645.290 717.880 ;
      LAYER met3 ;
        RECT 644.985 717.890 645.315 717.905 ;
        RECT 670.000 717.890 674.000 718.280 ;
        RECT 644.985 717.680 674.000 717.890 ;
        RECT 644.985 717.590 670.220 717.680 ;
        RECT 644.985 717.575 645.315 717.590 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 724.440 124.130 724.500 ;
        RECT 655.570 724.440 655.890 724.500 ;
        RECT 123.810 724.300 579.900 724.440 ;
        RECT 123.810 724.240 124.130 724.300 ;
        RECT 579.760 724.100 579.900 724.300 ;
        RECT 613.340 724.300 655.890 724.440 ;
        RECT 613.340 724.100 613.480 724.300 ;
        RECT 655.570 724.240 655.890 724.300 ;
        RECT 579.760 723.960 613.480 724.100 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 724.240 124.100 724.500 ;
        RECT 655.600 724.240 655.860 724.500 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 724.530 124.040 3498.270 ;
        RECT 123.840 724.210 124.100 724.530 ;
        RECT 655.600 724.210 655.860 724.530 ;
        RECT 655.660 722.685 655.800 724.210 ;
        RECT 655.590 722.315 655.870 722.685 ;
      LAYER via2 ;
        RECT 655.590 722.360 655.870 722.640 ;
      LAYER met3 ;
        RECT 655.565 722.650 655.895 722.665 ;
        RECT 670.000 722.650 674.000 723.040 ;
        RECT 655.565 722.440 674.000 722.650 ;
        RECT 655.565 722.350 670.220 722.440 ;
        RECT 655.565 722.335 655.895 722.350 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 731.240 17.410 731.300 ;
        RECT 655.570 731.240 655.890 731.300 ;
        RECT 17.090 731.100 655.890 731.240 ;
        RECT 17.090 731.040 17.410 731.100 ;
        RECT 655.570 731.040 655.890 731.100 ;
      LAYER via ;
        RECT 17.120 731.040 17.380 731.300 ;
        RECT 655.600 731.040 655.860 731.300 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.180 731.330 17.320 3339.635 ;
        RECT 17.120 731.010 17.380 731.330 ;
        RECT 655.600 731.010 655.860 731.330 ;
        RECT 655.660 728.125 655.800 731.010 ;
        RECT 655.590 727.755 655.870 728.125 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 655.590 727.800 655.870 728.080 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 655.565 728.090 655.895 728.105 ;
        RECT 670.000 728.090 674.000 728.480 ;
        RECT 655.565 727.880 674.000 728.090 ;
        RECT 655.565 727.790 670.220 727.880 ;
        RECT 655.565 727.775 655.895 727.790 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 738.040 18.330 738.100 ;
        RECT 661.090 738.040 661.410 738.100 ;
        RECT 18.010 737.900 661.410 738.040 ;
        RECT 18.010 737.840 18.330 737.900 ;
        RECT 661.090 737.840 661.410 737.900 ;
      LAYER via ;
        RECT 18.040 737.840 18.300 738.100 ;
        RECT 661.120 737.840 661.380 738.100 ;
      LAYER met2 ;
        RECT 18.030 3051.995 18.310 3052.365 ;
        RECT 18.100 738.130 18.240 3051.995 ;
        RECT 18.040 737.810 18.300 738.130 ;
        RECT 661.120 737.810 661.380 738.130 ;
        RECT 661.180 733.565 661.320 737.810 ;
        RECT 661.110 733.195 661.390 733.565 ;
      LAYER via2 ;
        RECT 18.030 3052.040 18.310 3052.320 ;
        RECT 661.110 733.240 661.390 733.520 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 18.005 3052.330 18.335 3052.345 ;
        RECT -4.800 3052.030 18.335 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 18.005 3052.015 18.335 3052.030 ;
        RECT 661.085 733.530 661.415 733.545 ;
        RECT 670.000 733.530 674.000 733.920 ;
        RECT 661.085 733.320 674.000 733.530 ;
        RECT 661.085 733.230 670.220 733.320 ;
        RECT 661.085 733.215 661.415 733.230 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 579.670 744.300 579.990 744.560 ;
        RECT 351.970 744.160 352.290 744.220 ;
        RECT 420.970 744.160 421.290 744.220 ;
        RECT 579.760 744.160 579.900 744.300 ;
        RECT 351.970 744.020 372.440 744.160 ;
        RECT 351.970 743.960 352.290 744.020 ;
        RECT 110.930 743.820 111.250 743.880 ;
        RECT 207.530 743.820 207.850 743.880 ;
        RECT 254.910 743.820 255.230 743.880 ;
        RECT 110.930 743.680 131.400 743.820 ;
        RECT 110.930 743.620 111.250 743.680 ;
        RECT 131.260 743.540 131.400 743.680 ;
        RECT 207.530 743.680 255.230 743.820 ;
        RECT 207.530 743.620 207.850 743.680 ;
        RECT 254.910 743.620 255.230 743.680 ;
        RECT 282.970 743.820 283.290 743.880 ;
        RECT 324.370 743.820 324.690 743.880 ;
        RECT 282.970 743.680 324.690 743.820 ;
        RECT 372.300 743.820 372.440 744.020 ;
        RECT 400.820 744.020 421.290 744.160 ;
        RECT 399.810 743.820 400.130 743.880 ;
        RECT 372.300 743.680 400.130 743.820 ;
        RECT 282.970 743.620 283.290 743.680 ;
        RECT 324.370 743.620 324.690 743.680 ;
        RECT 399.810 743.620 400.130 743.680 ;
        RECT 400.270 743.820 400.590 743.880 ;
        RECT 400.820 743.820 400.960 744.020 ;
        RECT 420.970 743.960 421.290 744.020 ;
        RECT 544.800 744.020 579.900 744.160 ;
        RECT 544.800 743.820 544.940 744.020 ;
        RECT 400.270 743.680 400.960 743.820 ;
        RECT 517.200 743.680 544.940 743.820 ;
        RECT 400.270 743.620 400.590 743.680 ;
        RECT 18.930 743.480 19.250 743.540 ;
        RECT 110.010 743.480 110.330 743.540 ;
        RECT 18.930 743.340 110.330 743.480 ;
        RECT 18.930 743.280 19.250 743.340 ;
        RECT 110.010 743.280 110.330 743.340 ;
        RECT 131.170 743.280 131.490 743.540 ;
        RECT 179.010 743.480 179.330 743.540 ;
        RECT 206.610 743.480 206.930 743.540 ;
        RECT 179.010 743.340 206.930 743.480 ;
        RECT 179.010 743.280 179.330 743.340 ;
        RECT 206.610 743.280 206.930 743.340 ;
        RECT 255.370 743.480 255.690 743.540 ;
        RECT 282.510 743.480 282.830 743.540 ;
        RECT 255.370 743.340 282.830 743.480 ;
        RECT 255.370 743.280 255.690 743.340 ;
        RECT 282.510 743.280 282.830 743.340 ;
        RECT 468.810 743.480 469.130 743.540 ;
        RECT 496.870 743.480 497.190 743.540 ;
        RECT 468.810 743.340 497.190 743.480 ;
        RECT 468.810 743.280 469.130 743.340 ;
        RECT 496.870 743.280 497.190 743.340 ;
        RECT 497.330 743.480 497.650 743.540 ;
        RECT 517.200 743.480 517.340 743.680 ;
        RECT 497.330 743.340 517.340 743.480 ;
        RECT 497.330 743.280 497.650 743.340 ;
        RECT 580.130 743.140 580.450 743.200 ;
        RECT 656.030 743.140 656.350 743.200 ;
        RECT 580.130 743.000 656.350 743.140 ;
        RECT 580.130 742.940 580.450 743.000 ;
        RECT 656.030 742.940 656.350 743.000 ;
        RECT 131.170 742.800 131.490 742.860 ;
        RECT 179.010 742.800 179.330 742.860 ;
        RECT 131.170 742.660 179.330 742.800 ;
        RECT 131.170 742.600 131.490 742.660 ;
        RECT 179.010 742.600 179.330 742.660 ;
      LAYER via ;
        RECT 579.700 744.300 579.960 744.560 ;
        RECT 352.000 743.960 352.260 744.220 ;
        RECT 110.960 743.620 111.220 743.880 ;
        RECT 207.560 743.620 207.820 743.880 ;
        RECT 254.940 743.620 255.200 743.880 ;
        RECT 283.000 743.620 283.260 743.880 ;
        RECT 324.400 743.620 324.660 743.880 ;
        RECT 399.840 743.620 400.100 743.880 ;
        RECT 400.300 743.620 400.560 743.880 ;
        RECT 421.000 743.960 421.260 744.220 ;
        RECT 18.960 743.280 19.220 743.540 ;
        RECT 110.040 743.280 110.300 743.540 ;
        RECT 131.200 743.280 131.460 743.540 ;
        RECT 179.040 743.280 179.300 743.540 ;
        RECT 206.640 743.280 206.900 743.540 ;
        RECT 255.400 743.280 255.660 743.540 ;
        RECT 282.540 743.280 282.800 743.540 ;
        RECT 468.840 743.280 469.100 743.540 ;
        RECT 496.900 743.280 497.160 743.540 ;
        RECT 497.360 743.280 497.620 743.540 ;
        RECT 580.160 742.940 580.420 743.200 ;
        RECT 656.060 742.940 656.320 743.200 ;
        RECT 131.200 742.600 131.460 742.860 ;
        RECT 179.040 742.600 179.300 742.860 ;
      LAYER met2 ;
        RECT 18.950 2765.035 19.230 2765.405 ;
        RECT 19.020 743.570 19.160 2765.035 ;
        RECT 579.760 744.870 580.360 745.010 ;
        RECT 579.760 744.590 579.900 744.870 ;
        RECT 352.000 743.930 352.260 744.250 ;
        RECT 420.990 744.075 421.270 744.445 ;
        RECT 467.910 744.075 468.190 744.445 ;
        RECT 579.700 744.270 579.960 744.590 ;
        RECT 421.000 743.930 421.260 744.075 ;
        RECT 110.960 743.650 111.220 743.910 ;
        RECT 207.560 743.650 207.820 743.910 ;
        RECT 110.100 743.590 111.220 743.650 ;
        RECT 206.700 743.590 207.820 743.650 ;
        RECT 254.940 743.650 255.200 743.910 ;
        RECT 283.000 743.650 283.260 743.910 ;
        RECT 324.400 743.765 324.660 743.910 ;
        RECT 352.060 743.765 352.200 743.930 ;
        RECT 254.940 743.590 255.600 743.650 ;
        RECT 110.100 743.570 111.160 743.590 ;
        RECT 206.700 743.570 207.760 743.590 ;
        RECT 18.960 743.250 19.220 743.570 ;
        RECT 110.040 743.510 111.160 743.570 ;
        RECT 110.040 743.250 110.300 743.510 ;
        RECT 131.200 743.250 131.460 743.570 ;
        RECT 179.040 743.250 179.300 743.570 ;
        RECT 206.640 743.510 207.760 743.570 ;
        RECT 255.000 743.570 255.600 743.590 ;
        RECT 282.600 743.590 283.260 743.650 ;
        RECT 282.600 743.570 283.200 743.590 ;
        RECT 255.000 743.510 255.660 743.570 ;
        RECT 206.640 743.250 206.900 743.510 ;
        RECT 255.400 743.250 255.660 743.510 ;
        RECT 282.540 743.510 283.200 743.570 ;
        RECT 282.540 743.250 282.800 743.510 ;
        RECT 324.390 743.395 324.670 743.765 ;
        RECT 351.990 743.395 352.270 743.765 ;
        RECT 399.840 743.650 400.100 743.910 ;
        RECT 400.300 743.650 400.560 743.910 ;
        RECT 399.840 743.590 400.560 743.650 ;
        RECT 399.900 743.510 400.500 743.590 ;
        RECT 131.260 742.890 131.400 743.250 ;
        RECT 179.100 742.890 179.240 743.250 ;
        RECT 467.980 742.970 468.120 744.075 ;
        RECT 496.960 743.570 497.560 743.650 ;
        RECT 468.840 743.250 469.100 743.570 ;
        RECT 496.900 743.510 497.620 743.570 ;
        RECT 496.900 743.250 497.160 743.510 ;
        RECT 497.360 743.250 497.620 743.510 ;
        RECT 468.900 742.970 469.040 743.250 ;
        RECT 580.220 743.230 580.360 744.870 ;
        RECT 131.200 742.570 131.460 742.890 ;
        RECT 179.040 742.570 179.300 742.890 ;
        RECT 467.980 742.830 469.040 742.970 ;
        RECT 580.160 742.910 580.420 743.230 ;
        RECT 656.060 742.910 656.320 743.230 ;
        RECT 656.120 741.725 656.260 742.910 ;
        RECT 656.050 741.355 656.330 741.725 ;
      LAYER via2 ;
        RECT 18.950 2765.080 19.230 2765.360 ;
        RECT 420.990 744.120 421.270 744.400 ;
        RECT 467.910 744.120 468.190 744.400 ;
        RECT 324.390 743.440 324.670 743.720 ;
        RECT 351.990 743.440 352.270 743.720 ;
        RECT 656.050 741.400 656.330 741.680 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 18.925 2765.370 19.255 2765.385 ;
        RECT -4.800 2765.070 19.255 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 18.925 2765.055 19.255 2765.070 ;
        RECT 420.965 744.410 421.295 744.425 ;
        RECT 467.885 744.410 468.215 744.425 ;
        RECT 420.965 744.110 468.215 744.410 ;
        RECT 420.965 744.095 421.295 744.110 ;
        RECT 467.885 744.095 468.215 744.110 ;
        RECT 324.365 743.730 324.695 743.745 ;
        RECT 351.965 743.730 352.295 743.745 ;
        RECT 324.365 743.430 352.295 743.730 ;
        RECT 324.365 743.415 324.695 743.430 ;
        RECT 351.965 743.415 352.295 743.430 ;
        RECT 656.025 741.690 656.355 741.705 ;
        RECT 656.025 741.390 670.370 741.690 ;
        RECT 656.025 741.375 656.355 741.390 ;
        RECT 670.070 739.360 670.370 741.390 ;
        RECT 670.000 738.760 674.000 739.360 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 745.180 20.170 745.240 ;
        RECT 656.030 745.180 656.350 745.240 ;
        RECT 19.850 745.040 656.350 745.180 ;
        RECT 19.850 744.980 20.170 745.040 ;
        RECT 656.030 744.980 656.350 745.040 ;
      LAYER via ;
        RECT 19.880 744.980 20.140 745.240 ;
        RECT 656.060 744.980 656.320 745.240 ;
      LAYER met2 ;
        RECT 19.870 2477.395 20.150 2477.765 ;
        RECT 19.940 745.270 20.080 2477.395 ;
        RECT 19.880 744.950 20.140 745.270 ;
        RECT 656.060 744.950 656.320 745.270 ;
        RECT 656.120 743.765 656.260 744.950 ;
        RECT 656.050 743.395 656.330 743.765 ;
      LAYER via2 ;
        RECT 19.870 2477.440 20.150 2477.720 ;
        RECT 656.050 743.440 656.330 743.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 19.845 2477.730 20.175 2477.745 ;
        RECT -4.800 2477.430 20.175 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 19.845 2477.415 20.175 2477.430 ;
        RECT 656.025 743.730 656.355 743.745 ;
        RECT 670.000 743.730 674.000 744.120 ;
        RECT 656.025 743.520 674.000 743.730 ;
        RECT 656.025 743.430 670.220 743.520 ;
        RECT 656.025 743.415 656.355 743.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 751.980 16.950 752.040 ;
        RECT 656.030 751.980 656.350 752.040 ;
        RECT 16.630 751.840 656.350 751.980 ;
        RECT 16.630 751.780 16.950 751.840 ;
        RECT 656.030 751.780 656.350 751.840 ;
      LAYER via ;
        RECT 16.660 751.780 16.920 752.040 ;
        RECT 656.060 751.780 656.320 752.040 ;
      LAYER met2 ;
        RECT 16.650 2189.755 16.930 2190.125 ;
        RECT 16.720 752.070 16.860 2189.755 ;
        RECT 16.660 751.750 16.920 752.070 ;
        RECT 656.060 751.750 656.320 752.070 ;
        RECT 656.120 749.205 656.260 751.750 ;
        RECT 656.050 748.835 656.330 749.205 ;
      LAYER via2 ;
        RECT 16.650 2189.800 16.930 2190.080 ;
        RECT 656.050 748.880 656.330 749.160 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 16.625 2190.090 16.955 2190.105 ;
        RECT -4.800 2189.790 16.955 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 16.625 2189.775 16.955 2189.790 ;
        RECT 656.025 749.170 656.355 749.185 ;
        RECT 670.000 749.170 674.000 749.560 ;
        RECT 656.025 748.960 674.000 749.170 ;
        RECT 656.025 748.870 670.220 748.960 ;
        RECT 656.025 748.855 656.355 748.870 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 656.030 758.780 656.350 758.840 ;
        RECT 15.710 758.640 656.350 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 656.030 758.580 656.350 758.640 ;
      LAYER via ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 656.060 758.580 656.320 758.840 ;
      LAYER met2 ;
        RECT 15.730 1902.795 16.010 1903.165 ;
        RECT 15.800 758.870 15.940 1902.795 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 656.060 758.550 656.320 758.870 ;
        RECT 656.120 754.645 656.260 758.550 ;
        RECT 656.050 754.275 656.330 754.645 ;
      LAYER via2 ;
        RECT 15.730 1902.840 16.010 1903.120 ;
        RECT 656.050 754.320 656.330 754.600 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 15.705 1903.130 16.035 1903.145 ;
        RECT -4.800 1902.830 16.035 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 15.705 1902.815 16.035 1902.830 ;
        RECT 656.025 754.610 656.355 754.625 ;
        RECT 670.000 754.610 674.000 755.000 ;
        RECT 656.025 754.400 674.000 754.610 ;
        RECT 656.025 754.310 670.220 754.400 ;
        RECT 656.025 754.295 656.355 754.310 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 670.290 604.080 670.610 604.140 ;
        RECT 2904.510 604.080 2904.830 604.140 ;
        RECT 670.290 603.940 2904.830 604.080 ;
        RECT 670.290 603.880 670.610 603.940 ;
        RECT 2904.510 603.880 2904.830 603.940 ;
      LAYER via ;
        RECT 670.320 603.880 670.580 604.140 ;
        RECT 2904.540 603.880 2904.800 604.140 ;
      LAYER met2 ;
        RECT 2904.530 615.555 2904.810 615.925 ;
        RECT 670.310 609.435 670.590 609.805 ;
        RECT 670.380 604.170 670.520 609.435 ;
        RECT 2904.600 604.170 2904.740 615.555 ;
        RECT 670.320 603.850 670.580 604.170 ;
        RECT 2904.540 603.850 2904.800 604.170 ;
      LAYER via2 ;
        RECT 2904.530 615.600 2904.810 615.880 ;
        RECT 670.310 609.480 670.590 609.760 ;
      LAYER met3 ;
        RECT 2904.505 615.890 2904.835 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2904.505 615.590 2924.800 615.890 ;
        RECT 2904.505 615.575 2904.835 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
        RECT 670.000 612.280 674.000 612.880 ;
        RECT 670.070 609.785 670.370 612.280 ;
        RECT 670.070 609.470 670.615 609.785 ;
        RECT 670.285 609.455 670.615 609.470 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 1614.900 15.110 1614.960 ;
        RECT 25.370 1614.900 25.690 1614.960 ;
        RECT 14.790 1614.760 25.690 1614.900 ;
        RECT 14.790 1614.700 15.110 1614.760 ;
        RECT 25.370 1614.700 25.690 1614.760 ;
        RECT 25.370 765.580 25.690 765.640 ;
        RECT 25.370 765.440 34.340 765.580 ;
        RECT 25.370 765.380 25.690 765.440 ;
        RECT 34.200 765.240 34.340 765.440 ;
        RECT 34.570 765.380 34.890 765.640 ;
        RECT 158.400 765.440 351.740 765.580 ;
        RECT 34.660 765.240 34.800 765.380 ;
        RECT 158.400 765.240 158.540 765.440 ;
        RECT 34.200 765.100 34.800 765.240 ;
        RECT 111.020 765.100 158.540 765.240 ;
        RECT 351.600 765.240 351.740 765.440 ;
        RECT 414.070 765.380 414.390 765.640 ;
        RECT 414.530 765.580 414.850 765.640 ;
        RECT 414.530 765.440 469.500 765.580 ;
        RECT 414.530 765.380 414.850 765.440 ;
        RECT 414.160 765.240 414.300 765.380 ;
        RECT 351.600 765.100 359.560 765.240 ;
        RECT 82.410 764.900 82.730 764.960 ;
        RECT 82.410 764.760 105.180 764.900 ;
        RECT 82.410 764.700 82.730 764.760 ;
        RECT 105.040 764.560 105.180 764.760 ;
        RECT 111.020 764.560 111.160 765.100 ;
        RECT 359.420 764.900 359.560 765.100 ;
        RECT 400.820 765.100 414.300 765.240 ;
        RECT 469.360 765.240 469.500 765.440 ;
        RECT 469.360 765.100 544.940 765.240 ;
        RECT 400.820 764.900 400.960 765.100 ;
        RECT 359.420 764.760 400.960 764.900 ;
        RECT 544.800 764.900 544.940 765.100 ;
        RECT 581.510 764.900 581.830 764.960 ;
        RECT 544.800 764.760 581.830 764.900 ;
        RECT 581.510 764.700 581.830 764.760 ;
        RECT 105.040 764.420 111.160 764.560 ;
        RECT 581.510 764.220 581.830 764.280 ;
        RECT 656.030 764.220 656.350 764.280 ;
        RECT 581.510 764.080 656.350 764.220 ;
        RECT 581.510 764.020 581.830 764.080 ;
        RECT 656.030 764.020 656.350 764.080 ;
      LAYER via ;
        RECT 14.820 1614.700 15.080 1614.960 ;
        RECT 25.400 1614.700 25.660 1614.960 ;
        RECT 25.400 765.380 25.660 765.640 ;
        RECT 34.600 765.380 34.860 765.640 ;
        RECT 414.100 765.380 414.360 765.640 ;
        RECT 414.560 765.380 414.820 765.640 ;
        RECT 82.440 764.700 82.700 764.960 ;
        RECT 581.540 764.700 581.800 764.960 ;
        RECT 581.540 764.020 581.800 764.280 ;
        RECT 656.060 764.020 656.320 764.280 ;
      LAYER met2 ;
        RECT 14.810 1615.155 15.090 1615.525 ;
        RECT 14.880 1614.990 15.020 1615.155 ;
        RECT 14.820 1614.670 15.080 1614.990 ;
        RECT 25.400 1614.670 25.660 1614.990 ;
        RECT 25.460 765.670 25.600 1614.670 ;
        RECT 25.400 765.350 25.660 765.670 ;
        RECT 34.600 765.525 34.860 765.670 ;
        RECT 34.590 765.155 34.870 765.525 ;
        RECT 82.430 765.155 82.710 765.525 ;
        RECT 414.100 765.410 414.360 765.670 ;
        RECT 414.560 765.410 414.820 765.670 ;
        RECT 414.100 765.350 414.820 765.410 ;
        RECT 414.160 765.270 414.760 765.350 ;
        RECT 82.500 764.990 82.640 765.155 ;
        RECT 82.440 764.670 82.700 764.990 ;
        RECT 581.540 764.670 581.800 764.990 ;
        RECT 581.600 764.310 581.740 764.670 ;
        RECT 581.540 763.990 581.800 764.310 ;
        RECT 656.060 763.990 656.320 764.310 ;
        RECT 656.120 760.085 656.260 763.990 ;
        RECT 656.050 759.715 656.330 760.085 ;
      LAYER via2 ;
        RECT 14.810 1615.200 15.090 1615.480 ;
        RECT 34.590 765.200 34.870 765.480 ;
        RECT 82.430 765.200 82.710 765.480 ;
        RECT 656.050 759.760 656.330 760.040 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 14.785 1615.490 15.115 1615.505 ;
        RECT -4.800 1615.190 15.115 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 14.785 1615.175 15.115 1615.190 ;
        RECT 34.565 765.490 34.895 765.505 ;
        RECT 82.405 765.490 82.735 765.505 ;
        RECT 34.565 765.190 82.735 765.490 ;
        RECT 34.565 765.175 34.895 765.190 ;
        RECT 82.405 765.175 82.735 765.190 ;
        RECT 656.025 760.050 656.355 760.065 ;
        RECT 670.000 760.050 674.000 760.440 ;
        RECT 656.025 759.840 674.000 760.050 ;
        RECT 656.025 759.750 670.220 759.840 ;
        RECT 656.025 759.735 656.355 759.750 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 765.920 15.110 765.980 ;
        RECT 656.030 765.920 656.350 765.980 ;
        RECT 14.790 765.780 656.350 765.920 ;
        RECT 14.790 765.720 15.110 765.780 ;
        RECT 656.030 765.720 656.350 765.780 ;
      LAYER via ;
        RECT 14.820 765.720 15.080 765.980 ;
        RECT 656.060 765.720 656.320 765.980 ;
      LAYER met2 ;
        RECT 14.810 1400.275 15.090 1400.645 ;
        RECT 14.880 766.010 15.020 1400.275 ;
        RECT 14.820 765.690 15.080 766.010 ;
        RECT 656.060 765.690 656.320 766.010 ;
        RECT 656.120 764.845 656.260 765.690 ;
        RECT 656.050 764.475 656.330 764.845 ;
      LAYER via2 ;
        RECT 14.810 1400.320 15.090 1400.600 ;
        RECT 656.050 764.520 656.330 764.800 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 14.785 1400.610 15.115 1400.625 ;
        RECT -4.800 1400.310 15.115 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 14.785 1400.295 15.115 1400.310 ;
        RECT 656.025 764.810 656.355 764.825 ;
        RECT 670.000 764.810 674.000 765.200 ;
        RECT 656.025 764.600 674.000 764.810 ;
        RECT 656.025 764.510 670.220 764.600 ;
        RECT 656.025 764.495 656.355 764.510 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 772.720 14.650 772.780 ;
        RECT 656.030 772.720 656.350 772.780 ;
        RECT 14.330 772.580 656.350 772.720 ;
        RECT 14.330 772.520 14.650 772.580 ;
        RECT 656.030 772.520 656.350 772.580 ;
      LAYER via ;
        RECT 14.360 772.520 14.620 772.780 ;
        RECT 656.060 772.520 656.320 772.780 ;
      LAYER met2 ;
        RECT 14.350 1184.715 14.630 1185.085 ;
        RECT 14.420 772.810 14.560 1184.715 ;
        RECT 14.360 772.490 14.620 772.810 ;
        RECT 656.060 772.490 656.320 772.810 ;
        RECT 656.120 770.285 656.260 772.490 ;
        RECT 656.050 769.915 656.330 770.285 ;
      LAYER via2 ;
        RECT 14.350 1184.760 14.630 1185.040 ;
        RECT 656.050 769.960 656.330 770.240 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 14.325 1185.050 14.655 1185.065 ;
        RECT -4.800 1184.750 14.655 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 14.325 1184.735 14.655 1184.750 ;
        RECT 656.025 770.250 656.355 770.265 ;
        RECT 670.000 770.250 674.000 770.640 ;
        RECT 656.025 770.040 674.000 770.250 ;
        RECT 656.025 769.950 670.220 770.040 ;
        RECT 656.025 769.935 656.355 769.950 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 779.520 15.570 779.580 ;
        RECT 15.250 779.380 656.260 779.520 ;
        RECT 15.250 779.320 15.570 779.380 ;
        RECT 656.120 779.240 656.260 779.380 ;
        RECT 656.030 778.980 656.350 779.240 ;
      LAYER via ;
        RECT 15.280 779.320 15.540 779.580 ;
        RECT 656.060 778.980 656.320 779.240 ;
      LAYER met2 ;
        RECT 15.270 969.155 15.550 969.525 ;
        RECT 15.340 779.610 15.480 969.155 ;
        RECT 15.280 779.290 15.540 779.610 ;
        RECT 656.060 778.950 656.320 779.270 ;
        RECT 656.120 775.725 656.260 778.950 ;
        RECT 656.050 775.355 656.330 775.725 ;
      LAYER via2 ;
        RECT 15.270 969.200 15.550 969.480 ;
        RECT 656.050 775.400 656.330 775.680 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.245 969.490 15.575 969.505 ;
        RECT -4.800 969.190 15.575 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.245 969.175 15.575 969.190 ;
        RECT 656.025 775.690 656.355 775.705 ;
        RECT 670.000 775.690 674.000 776.080 ;
        RECT 656.025 775.480 674.000 775.690 ;
        RECT 656.025 775.390 670.220 775.480 ;
        RECT 656.025 775.375 656.355 775.390 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.770 779.860 21.090 779.920 ;
        RECT 656.030 779.860 656.350 779.920 ;
        RECT 20.770 779.720 656.350 779.860 ;
        RECT 20.770 779.660 21.090 779.720 ;
        RECT 656.030 779.660 656.350 779.720 ;
      LAYER via ;
        RECT 20.800 779.660 21.060 779.920 ;
        RECT 656.060 779.660 656.320 779.920 ;
      LAYER met2 ;
        RECT 656.050 780.795 656.330 781.165 ;
        RECT 656.120 779.950 656.260 780.795 ;
        RECT 20.800 779.630 21.060 779.950 ;
        RECT 656.060 779.630 656.320 779.950 ;
        RECT 20.860 753.965 21.000 779.630 ;
        RECT 20.790 753.595 21.070 753.965 ;
      LAYER via2 ;
        RECT 656.050 780.840 656.330 781.120 ;
        RECT 20.790 753.640 21.070 753.920 ;
      LAYER met3 ;
        RECT 656.025 781.130 656.355 781.145 ;
        RECT 670.000 781.130 674.000 781.520 ;
        RECT 656.025 780.920 674.000 781.130 ;
        RECT 656.025 780.830 670.220 780.920 ;
        RECT 656.025 780.815 656.355 780.830 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 20.765 753.930 21.095 753.945 ;
        RECT -4.800 753.630 21.095 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 20.765 753.615 21.095 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 654.650 741.100 654.970 741.160 ;
        RECT 656.030 741.100 656.350 741.160 ;
        RECT 654.650 740.960 656.350 741.100 ;
        RECT 654.650 740.900 654.970 740.960 ;
        RECT 656.030 740.900 656.350 740.960 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 656.030 544.920 656.350 544.980 ;
        RECT 16.170 544.780 656.350 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 656.030 544.720 656.350 544.780 ;
      LAYER via ;
        RECT 654.680 740.900 654.940 741.160 ;
        RECT 656.060 740.900 656.320 741.160 ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 656.060 544.720 656.320 544.980 ;
      LAYER met2 ;
        RECT 654.670 782.835 654.950 783.205 ;
        RECT 654.740 741.190 654.880 782.835 ;
        RECT 654.680 740.870 654.940 741.190 ;
        RECT 656.060 740.870 656.320 741.190 ;
        RECT 656.120 545.010 656.260 740.870 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 656.060 544.690 656.320 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 654.670 782.880 654.950 783.160 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 670.000 785.680 674.000 786.280 ;
        RECT 654.645 783.170 654.975 783.185 ;
        RECT 670.070 783.170 670.370 785.680 ;
        RECT 654.645 782.870 670.370 783.170 ;
        RECT 654.645 782.855 654.975 782.870 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 657.870 324.260 658.190 324.320 ;
        RECT 16.630 324.120 658.190 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 657.870 324.060 658.190 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 657.900 324.060 658.160 324.320 ;
      LAYER met2 ;
        RECT 657.890 790.995 658.170 791.365 ;
        RECT 657.960 324.350 658.100 790.995 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 657.900 324.030 658.160 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 657.890 791.040 658.170 791.320 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 657.865 791.330 658.195 791.345 ;
        RECT 670.000 791.330 674.000 791.720 ;
        RECT 657.865 791.120 674.000 791.330 ;
        RECT 657.865 791.030 670.220 791.120 ;
        RECT 657.865 791.015 658.195 791.030 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 23.990 793.800 24.310 793.860 ;
        RECT 656.030 793.800 656.350 793.860 ;
        RECT 23.990 793.660 656.350 793.800 ;
        RECT 23.990 793.600 24.310 793.660 ;
        RECT 656.030 793.600 656.350 793.660 ;
        RECT 13.870 107.340 14.190 107.400 ;
        RECT 23.990 107.340 24.310 107.400 ;
        RECT 13.870 107.200 24.310 107.340 ;
        RECT 13.870 107.140 14.190 107.200 ;
        RECT 23.990 107.140 24.310 107.200 ;
      LAYER via ;
        RECT 24.020 793.600 24.280 793.860 ;
        RECT 656.060 793.600 656.320 793.860 ;
        RECT 13.900 107.140 14.160 107.400 ;
        RECT 24.020 107.140 24.280 107.400 ;
      LAYER met2 ;
        RECT 656.050 796.435 656.330 796.805 ;
        RECT 656.120 793.890 656.260 796.435 ;
        RECT 24.020 793.570 24.280 793.890 ;
        RECT 656.060 793.570 656.320 793.890 ;
        RECT 24.080 107.430 24.220 793.570 ;
        RECT 13.900 107.285 14.160 107.430 ;
        RECT 13.890 106.915 14.170 107.285 ;
        RECT 24.020 107.110 24.280 107.430 ;
      LAYER via2 ;
        RECT 656.050 796.480 656.330 796.760 ;
        RECT 13.890 106.960 14.170 107.240 ;
      LAYER met3 ;
        RECT 656.025 796.770 656.355 796.785 ;
        RECT 670.000 796.770 674.000 797.160 ;
        RECT 656.025 796.560 674.000 796.770 ;
        RECT 656.025 796.470 670.220 796.560 ;
        RECT 656.025 796.455 656.355 796.470 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 13.865 107.250 14.195 107.265 ;
        RECT -4.800 106.950 14.195 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 13.865 106.935 14.195 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 669.830 603.740 670.150 603.800 ;
        RECT 2901.750 603.740 2902.070 603.800 ;
        RECT 669.830 603.600 2902.070 603.740 ;
        RECT 669.830 603.540 670.150 603.600 ;
        RECT 2901.750 603.540 2902.070 603.600 ;
      LAYER via ;
        RECT 669.860 603.540 670.120 603.800 ;
        RECT 2901.780 603.540 2902.040 603.800 ;
      LAYER met2 ;
        RECT 2901.770 850.155 2902.050 850.525 ;
        RECT 669.850 614.875 670.130 615.245 ;
        RECT 669.920 603.830 670.060 614.875 ;
        RECT 2901.840 603.830 2901.980 850.155 ;
        RECT 669.860 603.510 670.120 603.830 ;
        RECT 2901.780 603.510 2902.040 603.830 ;
      LAYER via2 ;
        RECT 2901.770 850.200 2902.050 850.480 ;
        RECT 669.850 614.920 670.130 615.200 ;
      LAYER met3 ;
        RECT 2901.745 850.490 2902.075 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2901.745 850.190 2924.800 850.490 ;
        RECT 2901.745 850.175 2902.075 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT 670.000 617.720 674.000 618.320 ;
        RECT 670.070 615.225 670.370 617.720 ;
        RECT 669.825 614.910 670.370 615.225 ;
        RECT 669.825 614.895 670.155 614.910 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 663.850 1083.480 664.170 1083.540 ;
        RECT 2898.990 1083.480 2899.310 1083.540 ;
        RECT 663.850 1083.340 2899.310 1083.480 ;
        RECT 663.850 1083.280 664.170 1083.340 ;
        RECT 2898.990 1083.280 2899.310 1083.340 ;
      LAYER via ;
        RECT 663.880 1083.280 664.140 1083.540 ;
        RECT 2899.020 1083.280 2899.280 1083.540 ;
      LAYER met2 ;
        RECT 2899.010 1084.755 2899.290 1085.125 ;
        RECT 2899.080 1083.570 2899.220 1084.755 ;
        RECT 663.880 1083.250 664.140 1083.570 ;
        RECT 2899.020 1083.250 2899.280 1083.570 ;
        RECT 663.940 622.725 664.080 1083.250 ;
        RECT 663.870 622.355 664.150 622.725 ;
      LAYER via2 ;
        RECT 2899.010 1084.800 2899.290 1085.080 ;
        RECT 663.870 622.400 664.150 622.680 ;
      LAYER met3 ;
        RECT 2898.985 1085.090 2899.315 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2898.985 1084.790 2924.800 1085.090 ;
        RECT 2898.985 1084.775 2899.315 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
        RECT 663.845 622.690 664.175 622.705 ;
        RECT 670.000 622.690 674.000 623.080 ;
        RECT 663.845 622.480 674.000 622.690 ;
        RECT 663.845 622.390 670.220 622.480 ;
        RECT 663.845 622.375 664.175 622.390 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 658.330 1318.080 658.650 1318.140 ;
        RECT 2900.830 1318.080 2901.150 1318.140 ;
        RECT 658.330 1317.940 2901.150 1318.080 ;
        RECT 658.330 1317.880 658.650 1317.940 ;
        RECT 2900.830 1317.880 2901.150 1317.940 ;
      LAYER via ;
        RECT 658.360 1317.880 658.620 1318.140 ;
        RECT 2900.860 1317.880 2901.120 1318.140 ;
      LAYER met2 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
        RECT 2900.920 1318.170 2901.060 1319.355 ;
        RECT 658.360 1317.850 658.620 1318.170 ;
        RECT 2900.860 1317.850 2901.120 1318.170 ;
        RECT 658.420 628.165 658.560 1317.850 ;
        RECT 658.350 627.795 658.630 628.165 ;
      LAYER via2 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
        RECT 658.350 627.840 658.630 628.120 ;
      LAYER met3 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 658.325 628.130 658.655 628.145 ;
        RECT 670.000 628.130 674.000 628.520 ;
        RECT 658.325 627.920 674.000 628.130 ;
        RECT 658.325 627.830 670.220 627.920 ;
        RECT 658.325 627.815 658.655 627.830 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 658.790 1552.680 659.110 1552.740 ;
        RECT 2900.830 1552.680 2901.150 1552.740 ;
        RECT 658.790 1552.540 2901.150 1552.680 ;
        RECT 658.790 1552.480 659.110 1552.540 ;
        RECT 2900.830 1552.480 2901.150 1552.540 ;
      LAYER via ;
        RECT 658.820 1552.480 659.080 1552.740 ;
        RECT 2900.860 1552.480 2901.120 1552.740 ;
      LAYER met2 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
        RECT 2900.920 1552.770 2901.060 1553.955 ;
        RECT 658.820 1552.450 659.080 1552.770 ;
        RECT 2900.860 1552.450 2901.120 1552.770 ;
        RECT 658.880 633.605 659.020 1552.450 ;
        RECT 658.810 633.235 659.090 633.605 ;
      LAYER via2 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
        RECT 658.810 633.280 659.090 633.560 ;
      LAYER met3 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 658.785 633.570 659.115 633.585 ;
        RECT 670.000 633.570 674.000 633.960 ;
        RECT 658.785 633.360 674.000 633.570 ;
        RECT 658.785 633.270 670.220 633.360 ;
        RECT 658.785 633.255 659.115 633.270 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 657.410 1003.920 657.730 1003.980 ;
        RECT 2904.510 1003.920 2904.830 1003.980 ;
        RECT 657.410 1003.780 2904.830 1003.920 ;
        RECT 657.410 1003.720 657.730 1003.780 ;
        RECT 2904.510 1003.720 2904.830 1003.780 ;
      LAYER via ;
        RECT 657.440 1003.720 657.700 1003.980 ;
        RECT 2904.540 1003.720 2904.800 1003.980 ;
      LAYER met2 ;
        RECT 2904.530 1789.235 2904.810 1789.605 ;
        RECT 2904.600 1004.010 2904.740 1789.235 ;
        RECT 657.440 1003.690 657.700 1004.010 ;
        RECT 2904.540 1003.690 2904.800 1004.010 ;
        RECT 657.500 639.045 657.640 1003.690 ;
        RECT 657.430 638.675 657.710 639.045 ;
      LAYER via2 ;
        RECT 2904.530 1789.280 2904.810 1789.560 ;
        RECT 657.430 638.720 657.710 639.000 ;
      LAYER met3 ;
        RECT 2904.505 1789.570 2904.835 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2904.505 1789.270 2924.800 1789.570 ;
        RECT 2904.505 1789.255 2904.835 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 657.405 639.010 657.735 639.025 ;
        RECT 670.000 639.010 674.000 639.400 ;
        RECT 657.405 638.800 674.000 639.010 ;
        RECT 657.405 638.710 670.220 638.800 ;
        RECT 657.405 638.695 657.735 638.710 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 1004.260 657.270 1004.320 ;
        RECT 2903.130 1004.260 2903.450 1004.320 ;
        RECT 656.950 1004.120 2903.450 1004.260 ;
        RECT 656.950 1004.060 657.270 1004.120 ;
        RECT 2903.130 1004.060 2903.450 1004.120 ;
      LAYER via ;
        RECT 656.980 1004.060 657.240 1004.320 ;
        RECT 2903.160 1004.060 2903.420 1004.320 ;
      LAYER met2 ;
        RECT 2903.150 2023.835 2903.430 2024.205 ;
        RECT 2903.220 1004.350 2903.360 2023.835 ;
        RECT 656.980 1004.030 657.240 1004.350 ;
        RECT 2903.160 1004.030 2903.420 1004.350 ;
        RECT 657.040 643.805 657.180 1004.030 ;
        RECT 656.970 643.435 657.250 643.805 ;
      LAYER via2 ;
        RECT 2903.150 2023.880 2903.430 2024.160 ;
        RECT 656.970 643.480 657.250 643.760 ;
      LAYER met3 ;
        RECT 2903.125 2024.170 2903.455 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2903.125 2023.870 2924.800 2024.170 ;
        RECT 2903.125 2023.855 2903.455 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 656.945 643.770 657.275 643.785 ;
        RECT 670.000 643.770 674.000 644.160 ;
        RECT 656.945 643.560 674.000 643.770 ;
        RECT 656.945 643.470 670.220 643.560 ;
        RECT 656.945 643.455 657.275 643.470 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 670.290 2256.480 670.610 2256.540 ;
        RECT 2899.450 2256.480 2899.770 2256.540 ;
        RECT 670.290 2256.340 2899.770 2256.480 ;
        RECT 670.290 2256.280 670.610 2256.340 ;
        RECT 2899.450 2256.280 2899.770 2256.340 ;
      LAYER via ;
        RECT 670.320 2256.280 670.580 2256.540 ;
        RECT 2899.480 2256.280 2899.740 2256.540 ;
      LAYER met2 ;
        RECT 2899.470 2258.435 2899.750 2258.805 ;
        RECT 2899.540 2256.570 2899.680 2258.435 ;
        RECT 670.320 2256.250 670.580 2256.570 ;
        RECT 2899.480 2256.250 2899.740 2256.570 ;
        RECT 670.380 651.965 670.520 2256.250 ;
        RECT 670.310 651.595 670.590 651.965 ;
      LAYER via2 ;
        RECT 2899.470 2258.480 2899.750 2258.760 ;
        RECT 670.310 651.640 670.590 651.920 ;
      LAYER met3 ;
        RECT 2899.445 2258.770 2899.775 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2899.445 2258.470 2924.800 2258.770 ;
        RECT 2899.445 2258.455 2899.775 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 670.285 651.930 670.615 651.945 ;
        RECT 670.070 651.615 670.615 651.930 ;
        RECT 670.070 649.600 670.370 651.615 ;
        RECT 670.000 649.000 674.000 649.600 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 36.960 633.350 37.020 ;
        RECT 994.130 36.960 994.450 37.020 ;
        RECT 633.030 36.820 994.450 36.960 ;
        RECT 633.030 36.760 633.350 36.820 ;
        RECT 994.130 36.760 994.450 36.820 ;
      LAYER via ;
        RECT 633.060 36.760 633.320 37.020 ;
        RECT 994.160 36.760 994.420 37.020 ;
      LAYER met2 ;
        RECT 995.770 600.170 996.050 604.000 ;
        RECT 994.220 600.030 996.050 600.170 ;
        RECT 994.220 37.050 994.360 600.030 ;
        RECT 995.770 600.000 996.050 600.030 ;
        RECT 633.060 36.730 633.320 37.050 ;
        RECT 994.160 36.730 994.420 37.050 ;
        RECT 633.120 2.400 633.260 36.730 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1914.590 572.800 1914.910 572.860 ;
        RECT 1915.510 572.800 1915.830 572.860 ;
        RECT 1914.590 572.660 1915.830 572.800 ;
        RECT 1914.590 572.600 1914.910 572.660 ;
        RECT 1915.510 572.600 1915.830 572.660 ;
        RECT 1915.510 545.400 1915.830 545.660 ;
        RECT 1915.600 544.980 1915.740 545.400 ;
        RECT 1915.510 544.720 1915.830 544.980 ;
        RECT 1916.430 497.320 1916.750 497.380 ;
        RECT 1916.060 497.180 1916.750 497.320 ;
        RECT 1916.060 496.700 1916.200 497.180 ;
        RECT 1916.430 497.120 1916.750 497.180 ;
        RECT 1915.970 496.440 1916.290 496.700 ;
        RECT 1914.590 483.040 1914.910 483.100 ;
        RECT 1915.970 483.040 1916.290 483.100 ;
        RECT 1914.590 482.900 1916.290 483.040 ;
        RECT 1914.590 482.840 1914.910 482.900 ;
        RECT 1915.970 482.840 1916.290 482.900 ;
        RECT 1914.590 435.100 1914.910 435.160 ;
        RECT 1915.510 435.100 1915.830 435.160 ;
        RECT 1914.590 434.960 1915.830 435.100 ;
        RECT 1914.590 434.900 1914.910 434.960 ;
        RECT 1915.510 434.900 1915.830 434.960 ;
        RECT 1916.430 338.200 1916.750 338.260 ;
        RECT 1918.270 338.200 1918.590 338.260 ;
        RECT 1916.430 338.060 1918.590 338.200 ;
        RECT 1916.430 338.000 1916.750 338.060 ;
        RECT 1918.270 338.000 1918.590 338.060 ;
        RECT 1916.430 304.200 1916.750 304.260 ;
        RECT 1916.060 304.060 1916.750 304.200 ;
        RECT 1916.060 303.580 1916.200 304.060 ;
        RECT 1916.430 304.000 1916.750 304.060 ;
        RECT 1915.970 303.320 1916.290 303.580 ;
        RECT 1915.050 289.580 1915.370 289.640 ;
        RECT 1915.970 289.580 1916.290 289.640 ;
        RECT 1915.050 289.440 1916.290 289.580 ;
        RECT 1915.050 289.380 1915.370 289.440 ;
        RECT 1915.970 289.380 1916.290 289.440 ;
        RECT 1915.050 241.640 1915.370 241.700 ;
        RECT 1916.430 241.640 1916.750 241.700 ;
        RECT 1915.050 241.500 1916.750 241.640 ;
        RECT 1915.050 241.440 1915.370 241.500 ;
        RECT 1916.430 241.440 1916.750 241.500 ;
        RECT 1915.050 193.020 1915.370 193.080 ;
        RECT 1915.970 193.020 1916.290 193.080 ;
        RECT 1915.050 192.880 1916.290 193.020 ;
        RECT 1915.050 192.820 1915.370 192.880 ;
        RECT 1915.970 192.820 1916.290 192.880 ;
        RECT 1915.050 145.080 1915.370 145.140 ;
        RECT 1916.430 145.080 1916.750 145.140 ;
        RECT 1915.050 144.940 1916.750 145.080 ;
        RECT 1915.050 144.880 1915.370 144.940 ;
        RECT 1916.430 144.880 1916.750 144.940 ;
        RECT 1916.890 36.960 1917.210 37.020 ;
        RECT 2417.370 36.960 2417.690 37.020 ;
        RECT 1916.890 36.820 2417.690 36.960 ;
        RECT 1916.890 36.760 1917.210 36.820 ;
        RECT 2417.370 36.760 2417.690 36.820 ;
      LAYER via ;
        RECT 1914.620 572.600 1914.880 572.860 ;
        RECT 1915.540 572.600 1915.800 572.860 ;
        RECT 1915.540 545.400 1915.800 545.660 ;
        RECT 1915.540 544.720 1915.800 544.980 ;
        RECT 1916.460 497.120 1916.720 497.380 ;
        RECT 1916.000 496.440 1916.260 496.700 ;
        RECT 1914.620 482.840 1914.880 483.100 ;
        RECT 1916.000 482.840 1916.260 483.100 ;
        RECT 1914.620 434.900 1914.880 435.160 ;
        RECT 1915.540 434.900 1915.800 435.160 ;
        RECT 1916.460 338.000 1916.720 338.260 ;
        RECT 1918.300 338.000 1918.560 338.260 ;
        RECT 1916.460 304.000 1916.720 304.260 ;
        RECT 1916.000 303.320 1916.260 303.580 ;
        RECT 1915.080 289.380 1915.340 289.640 ;
        RECT 1916.000 289.380 1916.260 289.640 ;
        RECT 1915.080 241.440 1915.340 241.700 ;
        RECT 1916.460 241.440 1916.720 241.700 ;
        RECT 1915.080 192.820 1915.340 193.080 ;
        RECT 1916.000 192.820 1916.260 193.080 ;
        RECT 1915.080 144.880 1915.340 145.140 ;
        RECT 1916.460 144.880 1916.720 145.140 ;
        RECT 1916.920 36.760 1917.180 37.020 ;
        RECT 2417.400 36.760 2417.660 37.020 ;
      LAYER met2 ;
        RECT 1913.930 600.170 1914.210 604.000 ;
        RECT 1913.930 600.030 1914.820 600.170 ;
        RECT 1913.930 600.000 1914.210 600.030 ;
        RECT 1914.680 572.890 1914.820 600.030 ;
        RECT 1914.620 572.570 1914.880 572.890 ;
        RECT 1915.540 572.570 1915.800 572.890 ;
        RECT 1915.600 545.690 1915.740 572.570 ;
        RECT 1915.540 545.370 1915.800 545.690 ;
        RECT 1915.540 544.690 1915.800 545.010 ;
        RECT 1915.600 531.605 1915.740 544.690 ;
        RECT 1915.530 531.235 1915.810 531.605 ;
        RECT 1916.450 531.235 1916.730 531.605 ;
        RECT 1916.520 497.410 1916.660 531.235 ;
        RECT 1916.460 497.090 1916.720 497.410 ;
        RECT 1916.000 496.410 1916.260 496.730 ;
        RECT 1916.060 483.130 1916.200 496.410 ;
        RECT 1914.620 482.810 1914.880 483.130 ;
        RECT 1916.000 482.810 1916.260 483.130 ;
        RECT 1914.680 435.190 1914.820 482.810 ;
        RECT 1914.620 434.870 1914.880 435.190 ;
        RECT 1915.540 434.870 1915.800 435.190 ;
        RECT 1915.600 399.570 1915.740 434.870 ;
        RECT 1915.600 399.430 1916.200 399.570 ;
        RECT 1916.060 386.085 1916.200 399.430 ;
        RECT 1915.990 385.715 1916.270 386.085 ;
        RECT 1918.290 385.715 1918.570 386.085 ;
        RECT 1918.360 338.290 1918.500 385.715 ;
        RECT 1916.460 337.970 1916.720 338.290 ;
        RECT 1918.300 337.970 1918.560 338.290 ;
        RECT 1916.520 304.290 1916.660 337.970 ;
        RECT 1916.460 303.970 1916.720 304.290 ;
        RECT 1916.000 303.290 1916.260 303.610 ;
        RECT 1916.060 289.670 1916.200 303.290 ;
        RECT 1915.080 289.350 1915.340 289.670 ;
        RECT 1916.000 289.350 1916.260 289.670 ;
        RECT 1915.140 241.730 1915.280 289.350 ;
        RECT 1915.080 241.410 1915.340 241.730 ;
        RECT 1916.460 241.410 1916.720 241.730 ;
        RECT 1916.520 217.330 1916.660 241.410 ;
        RECT 1916.060 217.190 1916.660 217.330 ;
        RECT 1916.060 193.110 1916.200 217.190 ;
        RECT 1915.080 192.790 1915.340 193.110 ;
        RECT 1916.000 192.790 1916.260 193.110 ;
        RECT 1915.140 145.170 1915.280 192.790 ;
        RECT 1915.080 144.850 1915.340 145.170 ;
        RECT 1916.460 144.850 1916.720 145.170 ;
        RECT 1916.520 144.685 1916.660 144.850 ;
        RECT 1916.450 144.315 1916.730 144.685 ;
        RECT 1916.910 109.635 1917.190 110.005 ;
        RECT 1916.980 37.050 1917.120 109.635 ;
        RECT 1916.920 36.730 1917.180 37.050 ;
        RECT 2417.400 36.730 2417.660 37.050 ;
        RECT 2417.460 2.400 2417.600 36.730 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
      LAYER via2 ;
        RECT 1915.530 531.280 1915.810 531.560 ;
        RECT 1916.450 531.280 1916.730 531.560 ;
        RECT 1915.990 385.760 1916.270 386.040 ;
        RECT 1918.290 385.760 1918.570 386.040 ;
        RECT 1916.450 144.360 1916.730 144.640 ;
        RECT 1916.910 109.680 1917.190 109.960 ;
      LAYER met3 ;
        RECT 1915.505 531.570 1915.835 531.585 ;
        RECT 1916.425 531.570 1916.755 531.585 ;
        RECT 1915.505 531.270 1916.755 531.570 ;
        RECT 1915.505 531.255 1915.835 531.270 ;
        RECT 1916.425 531.255 1916.755 531.270 ;
        RECT 1915.965 386.050 1916.295 386.065 ;
        RECT 1918.265 386.050 1918.595 386.065 ;
        RECT 1915.965 385.750 1918.595 386.050 ;
        RECT 1915.965 385.735 1916.295 385.750 ;
        RECT 1918.265 385.735 1918.595 385.750 ;
        RECT 1916.425 144.660 1916.755 144.665 ;
        RECT 1916.425 144.650 1917.010 144.660 ;
        RECT 1916.425 144.350 1917.210 144.650 ;
        RECT 1916.425 144.340 1917.010 144.350 ;
        RECT 1916.425 144.335 1916.755 144.340 ;
        RECT 1916.885 109.980 1917.215 109.985 ;
        RECT 1916.630 109.970 1917.215 109.980 ;
        RECT 1916.430 109.670 1917.215 109.970 ;
        RECT 1916.630 109.660 1917.215 109.670 ;
        RECT 1916.885 109.655 1917.215 109.660 ;
      LAYER via3 ;
        RECT 1916.660 144.340 1916.980 144.660 ;
        RECT 1916.660 109.660 1916.980 109.980 ;
      LAYER met4 ;
        RECT 1916.655 144.335 1916.985 144.665 ;
        RECT 1916.670 109.985 1916.970 144.335 ;
        RECT 1916.655 109.655 1916.985 109.985 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1924.710 37.300 1925.030 37.360 ;
        RECT 2434.850 37.300 2435.170 37.360 ;
        RECT 1924.710 37.160 2435.170 37.300 ;
        RECT 1924.710 37.100 1925.030 37.160 ;
        RECT 2434.850 37.100 2435.170 37.160 ;
      LAYER via ;
        RECT 1924.740 37.100 1925.000 37.360 ;
        RECT 2434.880 37.100 2435.140 37.360 ;
      LAYER met2 ;
        RECT 1923.130 600.170 1923.410 604.000 ;
        RECT 1923.130 600.030 1924.020 600.170 ;
        RECT 1923.130 600.000 1923.410 600.030 ;
        RECT 1923.880 587.250 1924.020 600.030 ;
        RECT 1923.880 587.110 1924.940 587.250 ;
        RECT 1924.800 37.390 1924.940 587.110 ;
        RECT 1924.740 37.070 1925.000 37.390 ;
        RECT 2434.880 37.070 2435.140 37.390 ;
        RECT 2434.940 2.400 2435.080 37.070 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1933.910 586.740 1934.230 586.800 ;
        RECT 1938.050 586.740 1938.370 586.800 ;
        RECT 1933.910 586.600 1938.370 586.740 ;
        RECT 1933.910 586.540 1934.230 586.600 ;
        RECT 1938.050 586.540 1938.370 586.600 ;
        RECT 1938.050 37.640 1938.370 37.700 ;
        RECT 2452.790 37.640 2453.110 37.700 ;
        RECT 1938.050 37.500 2453.110 37.640 ;
        RECT 1938.050 37.440 1938.370 37.500 ;
        RECT 2452.790 37.440 2453.110 37.500 ;
      LAYER via ;
        RECT 1933.940 586.540 1934.200 586.800 ;
        RECT 1938.080 586.540 1938.340 586.800 ;
        RECT 1938.080 37.440 1938.340 37.700 ;
        RECT 2452.820 37.440 2453.080 37.700 ;
      LAYER met2 ;
        RECT 1932.330 600.170 1932.610 604.000 ;
        RECT 1932.330 600.030 1934.140 600.170 ;
        RECT 1932.330 600.000 1932.610 600.030 ;
        RECT 1934.000 586.830 1934.140 600.030 ;
        RECT 1933.940 586.510 1934.200 586.830 ;
        RECT 1938.080 586.510 1938.340 586.830 ;
        RECT 1938.140 37.730 1938.280 586.510 ;
        RECT 1938.080 37.410 1938.340 37.730 ;
        RECT 2452.820 37.410 2453.080 37.730 ;
        RECT 2452.880 2.400 2453.020 37.410 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1944.030 545.260 1944.350 545.320 ;
        RECT 1944.950 545.260 1945.270 545.320 ;
        RECT 1944.030 545.120 1945.270 545.260 ;
        RECT 1944.030 545.060 1944.350 545.120 ;
        RECT 1944.950 545.060 1945.270 545.120 ;
        RECT 1944.950 41.380 1945.270 41.440 ;
        RECT 2470.730 41.380 2471.050 41.440 ;
        RECT 1944.950 41.240 2471.050 41.380 ;
        RECT 1944.950 41.180 1945.270 41.240 ;
        RECT 2470.730 41.180 2471.050 41.240 ;
      LAYER via ;
        RECT 1944.060 545.060 1944.320 545.320 ;
        RECT 1944.980 545.060 1945.240 545.320 ;
        RECT 1944.980 41.180 1945.240 41.440 ;
        RECT 2470.760 41.180 2471.020 41.440 ;
      LAYER met2 ;
        RECT 1941.530 600.170 1941.810 604.000 ;
        RECT 1941.530 600.030 1944.260 600.170 ;
        RECT 1941.530 600.000 1941.810 600.030 ;
        RECT 1944.120 545.350 1944.260 600.030 ;
        RECT 1944.060 545.030 1944.320 545.350 ;
        RECT 1944.980 545.030 1945.240 545.350 ;
        RECT 1945.040 41.470 1945.180 545.030 ;
        RECT 1944.980 41.150 1945.240 41.470 ;
        RECT 2470.760 41.150 2471.020 41.470 ;
        RECT 2470.820 2.400 2470.960 41.150 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1952.310 41.040 1952.630 41.100 ;
        RECT 2488.670 41.040 2488.990 41.100 ;
        RECT 1952.310 40.900 2488.990 41.040 ;
        RECT 1952.310 40.840 1952.630 40.900 ;
        RECT 2488.670 40.840 2488.990 40.900 ;
      LAYER via ;
        RECT 1952.340 40.840 1952.600 41.100 ;
        RECT 2488.700 40.840 2488.960 41.100 ;
      LAYER met2 ;
        RECT 1950.730 600.170 1951.010 604.000 ;
        RECT 1950.730 600.030 1952.540 600.170 ;
        RECT 1950.730 600.000 1951.010 600.030 ;
        RECT 1952.400 41.130 1952.540 600.030 ;
        RECT 1952.340 40.810 1952.600 41.130 ;
        RECT 2488.700 40.810 2488.960 41.130 ;
        RECT 2488.760 2.400 2488.900 40.810 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1961.510 586.740 1961.830 586.800 ;
        RECT 1965.650 586.740 1965.970 586.800 ;
        RECT 1961.510 586.600 1965.970 586.740 ;
        RECT 1961.510 586.540 1961.830 586.600 ;
        RECT 1965.650 586.540 1965.970 586.600 ;
        RECT 1965.650 47.160 1965.970 47.220 ;
        RECT 2506.150 47.160 2506.470 47.220 ;
        RECT 1965.650 47.020 2506.470 47.160 ;
        RECT 1965.650 46.960 1965.970 47.020 ;
        RECT 2506.150 46.960 2506.470 47.020 ;
      LAYER via ;
        RECT 1961.540 586.540 1961.800 586.800 ;
        RECT 1965.680 586.540 1965.940 586.800 ;
        RECT 1965.680 46.960 1965.940 47.220 ;
        RECT 2506.180 46.960 2506.440 47.220 ;
      LAYER met2 ;
        RECT 1959.930 600.170 1960.210 604.000 ;
        RECT 1959.930 600.030 1961.740 600.170 ;
        RECT 1959.930 600.000 1960.210 600.030 ;
        RECT 1961.600 586.830 1961.740 600.030 ;
        RECT 1961.540 586.510 1961.800 586.830 ;
        RECT 1965.680 586.510 1965.940 586.830 ;
        RECT 1965.740 47.250 1965.880 586.510 ;
        RECT 1965.680 46.930 1965.940 47.250 ;
        RECT 2506.180 46.930 2506.440 47.250 ;
        RECT 2506.240 2.400 2506.380 46.930 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1971.630 545.260 1971.950 545.320 ;
        RECT 1972.550 545.260 1972.870 545.320 ;
        RECT 1971.630 545.120 1972.870 545.260 ;
        RECT 1971.630 545.060 1971.950 545.120 ;
        RECT 1972.550 545.060 1972.870 545.120 ;
        RECT 1972.550 46.820 1972.870 46.880 ;
        RECT 2524.090 46.820 2524.410 46.880 ;
        RECT 1972.550 46.680 2524.410 46.820 ;
        RECT 1972.550 46.620 1972.870 46.680 ;
        RECT 2524.090 46.620 2524.410 46.680 ;
      LAYER via ;
        RECT 1971.660 545.060 1971.920 545.320 ;
        RECT 1972.580 545.060 1972.840 545.320 ;
        RECT 1972.580 46.620 1972.840 46.880 ;
        RECT 2524.120 46.620 2524.380 46.880 ;
      LAYER met2 ;
        RECT 1969.130 600.170 1969.410 604.000 ;
        RECT 1969.130 600.030 1971.860 600.170 ;
        RECT 1969.130 600.000 1969.410 600.030 ;
        RECT 1971.720 545.350 1971.860 600.030 ;
        RECT 1971.660 545.030 1971.920 545.350 ;
        RECT 1972.580 545.030 1972.840 545.350 ;
        RECT 1972.640 46.910 1972.780 545.030 ;
        RECT 1972.580 46.590 1972.840 46.910 ;
        RECT 2524.120 46.590 2524.380 46.910 ;
        RECT 2524.180 2.400 2524.320 46.590 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1979.910 46.480 1980.230 46.540 ;
        RECT 2542.030 46.480 2542.350 46.540 ;
        RECT 1979.910 46.340 2542.350 46.480 ;
        RECT 1979.910 46.280 1980.230 46.340 ;
        RECT 2542.030 46.280 2542.350 46.340 ;
      LAYER via ;
        RECT 1979.940 46.280 1980.200 46.540 ;
        RECT 2542.060 46.280 2542.320 46.540 ;
      LAYER met2 ;
        RECT 1978.330 600.170 1978.610 604.000 ;
        RECT 1978.330 600.030 1980.140 600.170 ;
        RECT 1978.330 600.000 1978.610 600.030 ;
        RECT 1980.000 46.570 1980.140 600.030 ;
        RECT 1979.940 46.250 1980.200 46.570 ;
        RECT 2542.060 46.250 2542.320 46.570 ;
        RECT 2542.120 2.400 2542.260 46.250 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1989.110 586.740 1989.430 586.800 ;
        RECT 1993.250 586.740 1993.570 586.800 ;
        RECT 1989.110 586.600 1993.570 586.740 ;
        RECT 1989.110 586.540 1989.430 586.600 ;
        RECT 1993.250 586.540 1993.570 586.600 ;
        RECT 1993.250 46.140 1993.570 46.200 ;
        RECT 2559.970 46.140 2560.290 46.200 ;
        RECT 1993.250 46.000 2560.290 46.140 ;
        RECT 1993.250 45.940 1993.570 46.000 ;
        RECT 2559.970 45.940 2560.290 46.000 ;
      LAYER via ;
        RECT 1989.140 586.540 1989.400 586.800 ;
        RECT 1993.280 586.540 1993.540 586.800 ;
        RECT 1993.280 45.940 1993.540 46.200 ;
        RECT 2560.000 45.940 2560.260 46.200 ;
      LAYER met2 ;
        RECT 1987.530 600.170 1987.810 604.000 ;
        RECT 1987.530 600.030 1989.340 600.170 ;
        RECT 1987.530 600.000 1987.810 600.030 ;
        RECT 1989.200 586.830 1989.340 600.030 ;
        RECT 1989.140 586.510 1989.400 586.830 ;
        RECT 1993.280 586.510 1993.540 586.830 ;
        RECT 1993.340 46.230 1993.480 586.510 ;
        RECT 1993.280 45.910 1993.540 46.230 ;
        RECT 2560.000 45.910 2560.260 46.230 ;
        RECT 2560.060 2.400 2560.200 45.910 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1998.310 587.080 1998.630 587.140 ;
        RECT 2000.610 587.080 2000.930 587.140 ;
        RECT 1998.310 586.940 2000.930 587.080 ;
        RECT 1998.310 586.880 1998.630 586.940 ;
        RECT 2000.610 586.880 2000.930 586.940 ;
        RECT 2000.610 21.320 2000.930 21.380 ;
        RECT 2577.910 21.320 2578.230 21.380 ;
        RECT 2000.610 21.180 2578.230 21.320 ;
        RECT 2000.610 21.120 2000.930 21.180 ;
        RECT 2577.910 21.120 2578.230 21.180 ;
      LAYER via ;
        RECT 1998.340 586.880 1998.600 587.140 ;
        RECT 2000.640 586.880 2000.900 587.140 ;
        RECT 2000.640 21.120 2000.900 21.380 ;
        RECT 2577.940 21.120 2578.200 21.380 ;
      LAYER met2 ;
        RECT 1996.730 600.170 1997.010 604.000 ;
        RECT 1996.730 600.030 1998.540 600.170 ;
        RECT 1996.730 600.000 1997.010 600.030 ;
        RECT 1998.400 587.170 1998.540 600.030 ;
        RECT 1998.340 586.850 1998.600 587.170 ;
        RECT 2000.640 586.850 2000.900 587.170 ;
        RECT 2000.700 21.410 2000.840 586.850 ;
        RECT 2000.640 21.090 2000.900 21.410 ;
        RECT 2577.940 21.090 2578.200 21.410 ;
        RECT 2578.000 2.400 2578.140 21.090 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1085.210 532.340 1085.530 532.400 ;
        RECT 1084.840 532.200 1085.530 532.340 ;
        RECT 1084.840 531.720 1084.980 532.200 ;
        RECT 1085.210 532.140 1085.530 532.200 ;
        RECT 1084.750 531.460 1085.070 531.720 ;
        RECT 1084.750 497.120 1085.070 497.380 ;
        RECT 1084.840 496.700 1084.980 497.120 ;
        RECT 1084.750 496.440 1085.070 496.700 ;
        RECT 1084.750 476.240 1085.070 476.300 ;
        RECT 1085.210 476.240 1085.530 476.300 ;
        RECT 1084.750 476.100 1085.530 476.240 ;
        RECT 1084.750 476.040 1085.070 476.100 ;
        RECT 1085.210 476.040 1085.530 476.100 ;
        RECT 1084.750 434.760 1085.070 434.820 ;
        RECT 1085.210 434.760 1085.530 434.820 ;
        RECT 1084.750 434.620 1085.530 434.760 ;
        RECT 1084.750 434.560 1085.070 434.620 ;
        RECT 1085.210 434.560 1085.530 434.620 ;
        RECT 811.510 17.240 811.830 17.300 ;
        RECT 1084.750 17.240 1085.070 17.300 ;
        RECT 811.510 17.100 1085.070 17.240 ;
        RECT 811.510 17.040 811.830 17.100 ;
        RECT 1084.750 17.040 1085.070 17.100 ;
      LAYER via ;
        RECT 1085.240 532.140 1085.500 532.400 ;
        RECT 1084.780 531.460 1085.040 531.720 ;
        RECT 1084.780 497.120 1085.040 497.380 ;
        RECT 1084.780 496.440 1085.040 496.700 ;
        RECT 1084.780 476.040 1085.040 476.300 ;
        RECT 1085.240 476.040 1085.500 476.300 ;
        RECT 1084.780 434.560 1085.040 434.820 ;
        RECT 1085.240 434.560 1085.500 434.820 ;
        RECT 811.540 17.040 811.800 17.300 ;
        RECT 1084.780 17.040 1085.040 17.300 ;
      LAYER met2 ;
        RECT 1087.770 600.170 1088.050 604.000 ;
        RECT 1087.140 600.030 1088.050 600.170 ;
        RECT 1087.140 579.885 1087.280 600.030 ;
        RECT 1087.770 600.000 1088.050 600.030 ;
        RECT 1085.230 579.515 1085.510 579.885 ;
        RECT 1087.070 579.515 1087.350 579.885 ;
        RECT 1085.300 532.430 1085.440 579.515 ;
        RECT 1085.240 532.110 1085.500 532.430 ;
        RECT 1084.780 531.430 1085.040 531.750 ;
        RECT 1084.840 497.410 1084.980 531.430 ;
        RECT 1084.780 497.090 1085.040 497.410 ;
        RECT 1084.780 496.410 1085.040 496.730 ;
        RECT 1084.840 476.330 1084.980 496.410 ;
        RECT 1084.780 476.010 1085.040 476.330 ;
        RECT 1085.240 476.010 1085.500 476.330 ;
        RECT 1085.300 434.850 1085.440 476.010 ;
        RECT 1084.780 434.530 1085.040 434.850 ;
        RECT 1085.240 434.530 1085.500 434.850 ;
        RECT 1084.840 17.330 1084.980 434.530 ;
        RECT 811.540 17.010 811.800 17.330 ;
        RECT 1084.780 17.010 1085.040 17.330 ;
        RECT 811.600 2.400 811.740 17.010 ;
        RECT 811.390 -4.800 811.950 2.400 ;
      LAYER via2 ;
        RECT 1085.230 579.560 1085.510 579.840 ;
        RECT 1087.070 579.560 1087.350 579.840 ;
      LAYER met3 ;
        RECT 1085.205 579.850 1085.535 579.865 ;
        RECT 1087.045 579.850 1087.375 579.865 ;
        RECT 1085.205 579.550 1087.375 579.850 ;
        RECT 1085.205 579.535 1085.535 579.550 ;
        RECT 1087.045 579.535 1087.375 579.550 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.510 21.660 2007.830 21.720 ;
        RECT 2595.390 21.660 2595.710 21.720 ;
        RECT 2007.510 21.520 2595.710 21.660 ;
        RECT 2007.510 21.460 2007.830 21.520 ;
        RECT 2595.390 21.460 2595.710 21.520 ;
      LAYER via ;
        RECT 2007.540 21.460 2007.800 21.720 ;
        RECT 2595.420 21.460 2595.680 21.720 ;
      LAYER met2 ;
        RECT 2005.930 600.170 2006.210 604.000 ;
        RECT 2005.930 600.030 2007.740 600.170 ;
        RECT 2005.930 600.000 2006.210 600.030 ;
        RECT 2007.600 21.750 2007.740 600.030 ;
        RECT 2007.540 21.430 2007.800 21.750 ;
        RECT 2595.420 21.430 2595.680 21.750 ;
        RECT 2595.480 2.400 2595.620 21.430 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2016.710 586.740 2017.030 586.800 ;
        RECT 2021.310 586.740 2021.630 586.800 ;
        RECT 2016.710 586.600 2021.630 586.740 ;
        RECT 2016.710 586.540 2017.030 586.600 ;
        RECT 2021.310 586.540 2021.630 586.600 ;
        RECT 2021.310 22.000 2021.630 22.060 ;
        RECT 2613.330 22.000 2613.650 22.060 ;
        RECT 2021.310 21.860 2613.650 22.000 ;
        RECT 2021.310 21.800 2021.630 21.860 ;
        RECT 2613.330 21.800 2613.650 21.860 ;
      LAYER via ;
        RECT 2016.740 586.540 2017.000 586.800 ;
        RECT 2021.340 586.540 2021.600 586.800 ;
        RECT 2021.340 21.800 2021.600 22.060 ;
        RECT 2613.360 21.800 2613.620 22.060 ;
      LAYER met2 ;
        RECT 2015.130 600.170 2015.410 604.000 ;
        RECT 2015.130 600.030 2016.940 600.170 ;
        RECT 2015.130 600.000 2015.410 600.030 ;
        RECT 2016.800 586.830 2016.940 600.030 ;
        RECT 2016.740 586.510 2017.000 586.830 ;
        RECT 2021.340 586.510 2021.600 586.830 ;
        RECT 2021.400 22.090 2021.540 586.510 ;
        RECT 2021.340 21.770 2021.600 22.090 ;
        RECT 2613.360 21.770 2613.620 22.090 ;
        RECT 2613.420 2.400 2613.560 21.770 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2025.910 586.740 2026.230 586.800 ;
        RECT 2028.210 586.740 2028.530 586.800 ;
        RECT 2025.910 586.600 2028.530 586.740 ;
        RECT 2025.910 586.540 2026.230 586.600 ;
        RECT 2028.210 586.540 2028.530 586.600 ;
        RECT 2028.210 22.340 2028.530 22.400 ;
        RECT 2631.270 22.340 2631.590 22.400 ;
        RECT 2028.210 22.200 2631.590 22.340 ;
        RECT 2028.210 22.140 2028.530 22.200 ;
        RECT 2631.270 22.140 2631.590 22.200 ;
      LAYER via ;
        RECT 2025.940 586.540 2026.200 586.800 ;
        RECT 2028.240 586.540 2028.500 586.800 ;
        RECT 2028.240 22.140 2028.500 22.400 ;
        RECT 2631.300 22.140 2631.560 22.400 ;
      LAYER met2 ;
        RECT 2024.330 600.170 2024.610 604.000 ;
        RECT 2024.330 600.030 2026.140 600.170 ;
        RECT 2024.330 600.000 2024.610 600.030 ;
        RECT 2026.000 586.830 2026.140 600.030 ;
        RECT 2025.940 586.510 2026.200 586.830 ;
        RECT 2028.240 586.510 2028.500 586.830 ;
        RECT 2028.300 22.430 2028.440 586.510 ;
        RECT 2028.240 22.110 2028.500 22.430 ;
        RECT 2631.300 22.110 2631.560 22.430 ;
        RECT 2631.360 2.400 2631.500 22.110 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2034.650 22.680 2034.970 22.740 ;
        RECT 2649.210 22.680 2649.530 22.740 ;
        RECT 2034.650 22.540 2649.530 22.680 ;
        RECT 2034.650 22.480 2034.970 22.540 ;
        RECT 2649.210 22.480 2649.530 22.540 ;
      LAYER via ;
        RECT 2034.680 22.480 2034.940 22.740 ;
        RECT 2649.240 22.480 2649.500 22.740 ;
      LAYER met2 ;
        RECT 2033.530 600.170 2033.810 604.000 ;
        RECT 2033.530 600.030 2034.880 600.170 ;
        RECT 2033.530 600.000 2033.810 600.030 ;
        RECT 2034.740 22.770 2034.880 600.030 ;
        RECT 2034.680 22.450 2034.940 22.770 ;
        RECT 2649.240 22.450 2649.500 22.770 ;
        RECT 2649.300 2.400 2649.440 22.450 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2044.310 586.740 2044.630 586.800 ;
        RECT 2048.450 586.740 2048.770 586.800 ;
        RECT 2044.310 586.600 2048.770 586.740 ;
        RECT 2044.310 586.540 2044.630 586.600 ;
        RECT 2048.450 586.540 2048.770 586.600 ;
        RECT 2048.910 23.020 2049.230 23.080 ;
        RECT 2667.150 23.020 2667.470 23.080 ;
        RECT 2048.910 22.880 2667.470 23.020 ;
        RECT 2048.910 22.820 2049.230 22.880 ;
        RECT 2667.150 22.820 2667.470 22.880 ;
      LAYER via ;
        RECT 2044.340 586.540 2044.600 586.800 ;
        RECT 2048.480 586.540 2048.740 586.800 ;
        RECT 2048.940 22.820 2049.200 23.080 ;
        RECT 2667.180 22.820 2667.440 23.080 ;
      LAYER met2 ;
        RECT 2042.730 600.170 2043.010 604.000 ;
        RECT 2042.730 600.030 2044.540 600.170 ;
        RECT 2042.730 600.000 2043.010 600.030 ;
        RECT 2044.400 586.830 2044.540 600.030 ;
        RECT 2044.340 586.510 2044.600 586.830 ;
        RECT 2048.480 586.510 2048.740 586.830 ;
        RECT 2048.540 42.570 2048.680 586.510 ;
        RECT 2048.540 42.430 2049.140 42.570 ;
        RECT 2049.000 23.110 2049.140 42.430 ;
        RECT 2048.940 22.790 2049.200 23.110 ;
        RECT 2667.180 22.790 2667.440 23.110 ;
        RECT 2667.240 2.400 2667.380 22.790 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2053.510 586.740 2053.830 586.800 ;
        RECT 2055.810 586.740 2056.130 586.800 ;
        RECT 2053.510 586.600 2056.130 586.740 ;
        RECT 2053.510 586.540 2053.830 586.600 ;
        RECT 2055.810 586.540 2056.130 586.600 ;
        RECT 2055.810 23.360 2056.130 23.420 ;
        RECT 2684.630 23.360 2684.950 23.420 ;
        RECT 2055.810 23.220 2684.950 23.360 ;
        RECT 2055.810 23.160 2056.130 23.220 ;
        RECT 2684.630 23.160 2684.950 23.220 ;
      LAYER via ;
        RECT 2053.540 586.540 2053.800 586.800 ;
        RECT 2055.840 586.540 2056.100 586.800 ;
        RECT 2055.840 23.160 2056.100 23.420 ;
        RECT 2684.660 23.160 2684.920 23.420 ;
      LAYER met2 ;
        RECT 2051.930 600.170 2052.210 604.000 ;
        RECT 2051.930 600.030 2053.740 600.170 ;
        RECT 2051.930 600.000 2052.210 600.030 ;
        RECT 2053.600 586.830 2053.740 600.030 ;
        RECT 2053.540 586.510 2053.800 586.830 ;
        RECT 2055.840 586.510 2056.100 586.830 ;
        RECT 2055.900 23.450 2056.040 586.510 ;
        RECT 2055.840 23.130 2056.100 23.450 ;
        RECT 2684.660 23.130 2684.920 23.450 ;
        RECT 2684.720 2.400 2684.860 23.130 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2062.710 23.700 2063.030 23.760 ;
        RECT 2702.570 23.700 2702.890 23.760 ;
        RECT 2062.710 23.560 2702.890 23.700 ;
        RECT 2062.710 23.500 2063.030 23.560 ;
        RECT 2702.570 23.500 2702.890 23.560 ;
      LAYER via ;
        RECT 2062.740 23.500 2063.000 23.760 ;
        RECT 2702.600 23.500 2702.860 23.760 ;
      LAYER met2 ;
        RECT 2061.130 600.170 2061.410 604.000 ;
        RECT 2061.130 600.030 2062.940 600.170 ;
        RECT 2061.130 600.000 2061.410 600.030 ;
        RECT 2062.800 23.790 2062.940 600.030 ;
        RECT 2062.740 23.470 2063.000 23.790 ;
        RECT 2702.600 23.470 2702.860 23.790 ;
        RECT 2702.660 2.400 2702.800 23.470 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2071.910 586.740 2072.230 586.800 ;
        RECT 2076.510 586.740 2076.830 586.800 ;
        RECT 2071.910 586.600 2076.830 586.740 ;
        RECT 2071.910 586.540 2072.230 586.600 ;
        RECT 2076.510 586.540 2076.830 586.600 ;
        RECT 2076.510 27.440 2076.830 27.500 ;
        RECT 2720.510 27.440 2720.830 27.500 ;
        RECT 2076.510 27.300 2720.830 27.440 ;
        RECT 2076.510 27.240 2076.830 27.300 ;
        RECT 2720.510 27.240 2720.830 27.300 ;
      LAYER via ;
        RECT 2071.940 586.540 2072.200 586.800 ;
        RECT 2076.540 586.540 2076.800 586.800 ;
        RECT 2076.540 27.240 2076.800 27.500 ;
        RECT 2720.540 27.240 2720.800 27.500 ;
      LAYER met2 ;
        RECT 2070.330 600.170 2070.610 604.000 ;
        RECT 2070.330 600.030 2072.140 600.170 ;
        RECT 2070.330 600.000 2070.610 600.030 ;
        RECT 2072.000 586.830 2072.140 600.030 ;
        RECT 2071.940 586.510 2072.200 586.830 ;
        RECT 2076.540 586.510 2076.800 586.830 ;
        RECT 2076.600 27.530 2076.740 586.510 ;
        RECT 2076.540 27.210 2076.800 27.530 ;
        RECT 2720.540 27.210 2720.800 27.530 ;
        RECT 2720.600 2.400 2720.740 27.210 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2081.110 586.740 2081.430 586.800 ;
        RECT 2083.410 586.740 2083.730 586.800 ;
        RECT 2081.110 586.600 2083.730 586.740 ;
        RECT 2081.110 586.540 2081.430 586.600 ;
        RECT 2083.410 586.540 2083.730 586.600 ;
        RECT 2083.410 27.100 2083.730 27.160 ;
        RECT 2738.450 27.100 2738.770 27.160 ;
        RECT 2083.410 26.960 2738.770 27.100 ;
        RECT 2083.410 26.900 2083.730 26.960 ;
        RECT 2738.450 26.900 2738.770 26.960 ;
      LAYER via ;
        RECT 2081.140 586.540 2081.400 586.800 ;
        RECT 2083.440 586.540 2083.700 586.800 ;
        RECT 2083.440 26.900 2083.700 27.160 ;
        RECT 2738.480 26.900 2738.740 27.160 ;
      LAYER met2 ;
        RECT 2079.530 600.170 2079.810 604.000 ;
        RECT 2079.530 600.030 2081.340 600.170 ;
        RECT 2079.530 600.000 2079.810 600.030 ;
        RECT 2081.200 586.830 2081.340 600.030 ;
        RECT 2081.140 586.510 2081.400 586.830 ;
        RECT 2083.440 586.510 2083.700 586.830 ;
        RECT 2083.500 27.190 2083.640 586.510 ;
        RECT 2083.440 26.870 2083.700 27.190 ;
        RECT 2738.480 26.870 2738.740 27.190 ;
        RECT 2738.540 2.400 2738.680 26.870 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 26.760 2090.630 26.820 ;
        RECT 2755.930 26.760 2756.250 26.820 ;
        RECT 2090.310 26.620 2756.250 26.760 ;
        RECT 2090.310 26.560 2090.630 26.620 ;
        RECT 2755.930 26.560 2756.250 26.620 ;
      LAYER via ;
        RECT 2090.340 26.560 2090.600 26.820 ;
        RECT 2755.960 26.560 2756.220 26.820 ;
      LAYER met2 ;
        RECT 2088.730 600.170 2089.010 604.000 ;
        RECT 2088.730 600.030 2090.540 600.170 ;
        RECT 2088.730 600.000 2089.010 600.030 ;
        RECT 2090.400 26.850 2090.540 600.030 ;
        RECT 2090.340 26.530 2090.600 26.850 ;
        RECT 2755.960 26.530 2756.220 26.850 ;
        RECT 2756.020 2.400 2756.160 26.530 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 829.450 17.580 829.770 17.640 ;
        RECT 1097.170 17.580 1097.490 17.640 ;
        RECT 829.450 17.440 1097.490 17.580 ;
        RECT 829.450 17.380 829.770 17.440 ;
        RECT 1097.170 17.380 1097.490 17.440 ;
      LAYER via ;
        RECT 829.480 17.380 829.740 17.640 ;
        RECT 1097.200 17.380 1097.460 17.640 ;
      LAYER met2 ;
        RECT 1096.970 600.000 1097.250 604.000 ;
        RECT 1097.030 598.810 1097.170 600.000 ;
        RECT 1097.030 598.670 1097.400 598.810 ;
        RECT 1097.260 17.670 1097.400 598.670 ;
        RECT 829.480 17.350 829.740 17.670 ;
        RECT 1097.200 17.350 1097.460 17.670 ;
        RECT 829.540 2.400 829.680 17.350 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2099.510 586.740 2099.830 586.800 ;
        RECT 2104.110 586.740 2104.430 586.800 ;
        RECT 2099.510 586.600 2104.430 586.740 ;
        RECT 2099.510 586.540 2099.830 586.600 ;
        RECT 2104.110 586.540 2104.430 586.600 ;
        RECT 2104.110 26.420 2104.430 26.480 ;
        RECT 2773.870 26.420 2774.190 26.480 ;
        RECT 2104.110 26.280 2774.190 26.420 ;
        RECT 2104.110 26.220 2104.430 26.280 ;
        RECT 2773.870 26.220 2774.190 26.280 ;
      LAYER via ;
        RECT 2099.540 586.540 2099.800 586.800 ;
        RECT 2104.140 586.540 2104.400 586.800 ;
        RECT 2104.140 26.220 2104.400 26.480 ;
        RECT 2773.900 26.220 2774.160 26.480 ;
      LAYER met2 ;
        RECT 2097.930 600.170 2098.210 604.000 ;
        RECT 2097.930 600.030 2099.740 600.170 ;
        RECT 2097.930 600.000 2098.210 600.030 ;
        RECT 2099.600 586.830 2099.740 600.030 ;
        RECT 2099.540 586.510 2099.800 586.830 ;
        RECT 2104.140 586.510 2104.400 586.830 ;
        RECT 2104.200 26.510 2104.340 586.510 ;
        RECT 2104.140 26.190 2104.400 26.510 ;
        RECT 2773.900 26.190 2774.160 26.510 ;
        RECT 2773.960 2.400 2774.100 26.190 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2108.710 587.080 2109.030 587.140 ;
        RECT 2111.010 587.080 2111.330 587.140 ;
        RECT 2108.710 586.940 2111.330 587.080 ;
        RECT 2108.710 586.880 2109.030 586.940 ;
        RECT 2111.010 586.880 2111.330 586.940 ;
        RECT 2111.010 26.080 2111.330 26.140 ;
        RECT 2791.810 26.080 2792.130 26.140 ;
        RECT 2111.010 25.940 2792.130 26.080 ;
        RECT 2111.010 25.880 2111.330 25.940 ;
        RECT 2791.810 25.880 2792.130 25.940 ;
      LAYER via ;
        RECT 2108.740 586.880 2109.000 587.140 ;
        RECT 2111.040 586.880 2111.300 587.140 ;
        RECT 2111.040 25.880 2111.300 26.140 ;
        RECT 2791.840 25.880 2792.100 26.140 ;
      LAYER met2 ;
        RECT 2107.130 600.170 2107.410 604.000 ;
        RECT 2107.130 600.030 2108.940 600.170 ;
        RECT 2107.130 600.000 2107.410 600.030 ;
        RECT 2108.800 587.170 2108.940 600.030 ;
        RECT 2108.740 586.850 2109.000 587.170 ;
        RECT 2111.040 586.850 2111.300 587.170 ;
        RECT 2111.100 26.170 2111.240 586.850 ;
        RECT 2111.040 25.850 2111.300 26.170 ;
        RECT 2791.840 25.850 2792.100 26.170 ;
        RECT 2791.900 2.400 2792.040 25.850 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2117.450 25.400 2117.770 25.460 ;
        RECT 2809.750 25.400 2810.070 25.460 ;
        RECT 2117.450 25.260 2810.070 25.400 ;
        RECT 2117.450 25.200 2117.770 25.260 ;
        RECT 2809.750 25.200 2810.070 25.260 ;
      LAYER via ;
        RECT 2117.480 25.200 2117.740 25.460 ;
        RECT 2809.780 25.200 2810.040 25.460 ;
      LAYER met2 ;
        RECT 2116.330 600.170 2116.610 604.000 ;
        RECT 2116.330 600.030 2117.680 600.170 ;
        RECT 2116.330 600.000 2116.610 600.030 ;
        RECT 2117.540 25.490 2117.680 600.030 ;
        RECT 2117.480 25.170 2117.740 25.490 ;
        RECT 2809.780 25.170 2810.040 25.490 ;
        RECT 2809.840 2.400 2809.980 25.170 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2127.110 586.740 2127.430 586.800 ;
        RECT 2131.710 586.740 2132.030 586.800 ;
        RECT 2127.110 586.600 2132.030 586.740 ;
        RECT 2127.110 586.540 2127.430 586.600 ;
        RECT 2131.710 586.540 2132.030 586.600 ;
        RECT 2131.710 25.740 2132.030 25.800 ;
        RECT 2827.690 25.740 2828.010 25.800 ;
        RECT 2131.710 25.600 2828.010 25.740 ;
        RECT 2131.710 25.540 2132.030 25.600 ;
        RECT 2827.690 25.540 2828.010 25.600 ;
      LAYER via ;
        RECT 2127.140 586.540 2127.400 586.800 ;
        RECT 2131.740 586.540 2132.000 586.800 ;
        RECT 2131.740 25.540 2132.000 25.800 ;
        RECT 2827.720 25.540 2827.980 25.800 ;
      LAYER met2 ;
        RECT 2125.530 600.170 2125.810 604.000 ;
        RECT 2125.530 600.030 2127.340 600.170 ;
        RECT 2125.530 600.000 2125.810 600.030 ;
        RECT 2127.200 586.830 2127.340 600.030 ;
        RECT 2127.140 586.510 2127.400 586.830 ;
        RECT 2131.740 586.510 2132.000 586.830 ;
        RECT 2131.800 25.830 2131.940 586.510 ;
        RECT 2131.740 25.510 2132.000 25.830 ;
        RECT 2827.720 25.510 2827.980 25.830 ;
        RECT 2827.780 2.400 2827.920 25.510 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2136.310 586.740 2136.630 586.800 ;
        RECT 2138.610 586.740 2138.930 586.800 ;
        RECT 2136.310 586.600 2138.930 586.740 ;
        RECT 2136.310 586.540 2136.630 586.600 ;
        RECT 2138.610 586.540 2138.930 586.600 ;
        RECT 2138.610 25.060 2138.930 25.120 ;
        RECT 2845.170 25.060 2845.490 25.120 ;
        RECT 2138.610 24.920 2845.490 25.060 ;
        RECT 2138.610 24.860 2138.930 24.920 ;
        RECT 2845.170 24.860 2845.490 24.920 ;
      LAYER via ;
        RECT 2136.340 586.540 2136.600 586.800 ;
        RECT 2138.640 586.540 2138.900 586.800 ;
        RECT 2138.640 24.860 2138.900 25.120 ;
        RECT 2845.200 24.860 2845.460 25.120 ;
      LAYER met2 ;
        RECT 2134.730 600.170 2135.010 604.000 ;
        RECT 2134.730 600.030 2136.540 600.170 ;
        RECT 2134.730 600.000 2135.010 600.030 ;
        RECT 2136.400 586.830 2136.540 600.030 ;
        RECT 2136.340 586.510 2136.600 586.830 ;
        RECT 2138.640 586.510 2138.900 586.830 ;
        RECT 2138.700 25.150 2138.840 586.510 ;
        RECT 2138.640 24.830 2138.900 25.150 ;
        RECT 2845.200 24.830 2845.460 25.150 ;
        RECT 2845.260 2.400 2845.400 24.830 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.510 24.720 2145.830 24.780 ;
        RECT 2863.110 24.720 2863.430 24.780 ;
        RECT 2145.510 24.580 2863.430 24.720 ;
        RECT 2145.510 24.520 2145.830 24.580 ;
        RECT 2863.110 24.520 2863.430 24.580 ;
      LAYER via ;
        RECT 2145.540 24.520 2145.800 24.780 ;
        RECT 2863.140 24.520 2863.400 24.780 ;
      LAYER met2 ;
        RECT 2143.930 600.170 2144.210 604.000 ;
        RECT 2143.930 600.030 2145.740 600.170 ;
        RECT 2143.930 600.000 2144.210 600.030 ;
        RECT 2145.600 24.810 2145.740 600.030 ;
        RECT 2145.540 24.490 2145.800 24.810 ;
        RECT 2863.140 24.490 2863.400 24.810 ;
        RECT 2863.200 2.400 2863.340 24.490 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2154.710 586.740 2155.030 586.800 ;
        RECT 2159.310 586.740 2159.630 586.800 ;
        RECT 2154.710 586.600 2159.630 586.740 ;
        RECT 2154.710 586.540 2155.030 586.600 ;
        RECT 2159.310 586.540 2159.630 586.600 ;
        RECT 2159.310 24.380 2159.630 24.440 ;
        RECT 2881.050 24.380 2881.370 24.440 ;
        RECT 2159.310 24.240 2881.370 24.380 ;
        RECT 2159.310 24.180 2159.630 24.240 ;
        RECT 2881.050 24.180 2881.370 24.240 ;
      LAYER via ;
        RECT 2154.740 586.540 2155.000 586.800 ;
        RECT 2159.340 586.540 2159.600 586.800 ;
        RECT 2159.340 24.180 2159.600 24.440 ;
        RECT 2881.080 24.180 2881.340 24.440 ;
      LAYER met2 ;
        RECT 2153.130 600.170 2153.410 604.000 ;
        RECT 2153.130 600.030 2154.940 600.170 ;
        RECT 2153.130 600.000 2153.410 600.030 ;
        RECT 2154.800 586.830 2154.940 600.030 ;
        RECT 2154.740 586.510 2155.000 586.830 ;
        RECT 2159.340 586.510 2159.600 586.830 ;
        RECT 2159.400 24.470 2159.540 586.510 ;
        RECT 2159.340 24.150 2159.600 24.470 ;
        RECT 2881.080 24.150 2881.340 24.470 ;
        RECT 2881.140 2.400 2881.280 24.150 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2163.910 586.740 2164.230 586.800 ;
        RECT 2166.210 586.740 2166.530 586.800 ;
        RECT 2163.910 586.600 2166.530 586.740 ;
        RECT 2163.910 586.540 2164.230 586.600 ;
        RECT 2166.210 586.540 2166.530 586.600 ;
        RECT 2166.210 24.040 2166.530 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 2166.210 23.900 2899.310 24.040 ;
        RECT 2166.210 23.840 2166.530 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 2163.940 586.540 2164.200 586.800 ;
        RECT 2166.240 586.540 2166.500 586.800 ;
        RECT 2166.240 23.840 2166.500 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 2162.330 600.170 2162.610 604.000 ;
        RECT 2162.330 600.030 2164.140 600.170 ;
        RECT 2162.330 600.000 2162.610 600.030 ;
        RECT 2164.000 586.830 2164.140 600.030 ;
        RECT 2163.940 586.510 2164.200 586.830 ;
        RECT 2166.240 586.510 2166.500 586.830 ;
        RECT 2166.300 24.130 2166.440 586.510 ;
        RECT 2166.240 23.810 2166.500 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.400 2899.220 23.810 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 846.930 17.920 847.250 17.980 ;
        RECT 1104.070 17.920 1104.390 17.980 ;
        RECT 846.930 17.780 1104.390 17.920 ;
        RECT 846.930 17.720 847.250 17.780 ;
        RECT 1104.070 17.720 1104.390 17.780 ;
      LAYER via ;
        RECT 846.960 17.720 847.220 17.980 ;
        RECT 1104.100 17.720 1104.360 17.980 ;
      LAYER met2 ;
        RECT 1106.170 600.170 1106.450 604.000 ;
        RECT 1104.160 600.030 1106.450 600.170 ;
        RECT 1104.160 18.010 1104.300 600.030 ;
        RECT 1106.170 600.000 1106.450 600.030 ;
        RECT 846.960 17.690 847.220 18.010 ;
        RECT 1104.100 17.690 1104.360 18.010 ;
        RECT 847.020 2.400 847.160 17.690 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.970 568.720 1111.290 568.780 ;
        RECT 1113.270 568.720 1113.590 568.780 ;
        RECT 1110.970 568.580 1113.590 568.720 ;
        RECT 1110.970 568.520 1111.290 568.580 ;
        RECT 1113.270 568.520 1113.590 568.580 ;
        RECT 864.870 18.940 865.190 19.000 ;
        RECT 900.290 18.940 900.610 19.000 ;
        RECT 864.870 18.800 900.610 18.940 ;
        RECT 864.870 18.740 865.190 18.800 ;
        RECT 900.290 18.740 900.610 18.800 ;
        RECT 931.110 18.260 931.430 18.320 ;
        RECT 1110.970 18.260 1111.290 18.320 ;
        RECT 931.110 18.120 1111.290 18.260 ;
        RECT 931.110 18.060 931.430 18.120 ;
        RECT 1110.970 18.060 1111.290 18.120 ;
        RECT 900.290 15.880 900.610 15.940 ;
        RECT 930.650 15.880 930.970 15.940 ;
        RECT 900.290 15.740 930.970 15.880 ;
        RECT 900.290 15.680 900.610 15.740 ;
        RECT 930.650 15.680 930.970 15.740 ;
      LAYER via ;
        RECT 1111.000 568.520 1111.260 568.780 ;
        RECT 1113.300 568.520 1113.560 568.780 ;
        RECT 864.900 18.740 865.160 19.000 ;
        RECT 900.320 18.740 900.580 19.000 ;
        RECT 931.140 18.060 931.400 18.320 ;
        RECT 1111.000 18.060 1111.260 18.320 ;
        RECT 900.320 15.680 900.580 15.940 ;
        RECT 930.680 15.680 930.940 15.940 ;
      LAYER met2 ;
        RECT 1114.910 600.170 1115.190 604.000 ;
        RECT 1113.360 600.030 1115.190 600.170 ;
        RECT 1113.360 568.810 1113.500 600.030 ;
        RECT 1114.910 600.000 1115.190 600.030 ;
        RECT 1111.000 568.490 1111.260 568.810 ;
        RECT 1113.300 568.490 1113.560 568.810 ;
        RECT 864.900 18.710 865.160 19.030 ;
        RECT 900.320 18.710 900.580 19.030 ;
        RECT 864.960 2.400 865.100 18.710 ;
        RECT 900.380 15.970 900.520 18.710 ;
        RECT 1111.060 18.350 1111.200 568.490 ;
        RECT 931.140 18.090 931.400 18.350 ;
        RECT 930.740 18.030 931.400 18.090 ;
        RECT 1111.000 18.030 1111.260 18.350 ;
        RECT 930.740 17.950 931.340 18.030 ;
        RECT 930.740 15.970 930.880 17.950 ;
        RECT 900.320 15.650 900.580 15.970 ;
        RECT 930.680 15.650 930.940 15.970 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 883.730 18.600 884.050 18.660 ;
        RECT 1118.790 18.600 1119.110 18.660 ;
        RECT 883.730 18.460 1119.110 18.600 ;
        RECT 883.730 18.400 884.050 18.460 ;
        RECT 1118.790 18.400 1119.110 18.460 ;
      LAYER via ;
        RECT 883.760 18.400 884.020 18.660 ;
        RECT 1118.820 18.400 1119.080 18.660 ;
      LAYER met2 ;
        RECT 1124.110 600.170 1124.390 604.000 ;
        RECT 1122.100 600.030 1124.390 600.170 ;
        RECT 1122.100 588.610 1122.240 600.030 ;
        RECT 1124.110 600.000 1124.390 600.030 ;
        RECT 1118.880 588.470 1122.240 588.610 ;
        RECT 1118.880 18.690 1119.020 588.470 ;
        RECT 883.760 18.370 884.020 18.690 ;
        RECT 1118.820 18.370 1119.080 18.690 ;
        RECT 883.820 17.410 883.960 18.370 ;
        RECT 882.900 17.270 883.960 17.410 ;
        RECT 882.900 2.400 883.040 17.270 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 900.750 18.940 901.070 19.000 ;
        RECT 1110.510 18.940 1110.830 19.000 ;
        RECT 900.750 18.800 1110.830 18.940 ;
        RECT 900.750 18.740 901.070 18.800 ;
        RECT 1110.510 18.740 1110.830 18.800 ;
        RECT 1114.190 18.940 1114.510 19.000 ;
        RECT 1132.130 18.940 1132.450 19.000 ;
        RECT 1114.190 18.800 1132.450 18.940 ;
        RECT 1114.190 18.740 1114.510 18.800 ;
        RECT 1132.130 18.740 1132.450 18.800 ;
        RECT 1110.510 17.580 1110.830 17.640 ;
        RECT 1114.190 17.580 1114.510 17.640 ;
        RECT 1110.510 17.440 1114.510 17.580 ;
        RECT 1110.510 17.380 1110.830 17.440 ;
        RECT 1114.190 17.380 1114.510 17.440 ;
      LAYER via ;
        RECT 900.780 18.740 901.040 19.000 ;
        RECT 1110.540 18.740 1110.800 19.000 ;
        RECT 1114.220 18.740 1114.480 19.000 ;
        RECT 1132.160 18.740 1132.420 19.000 ;
        RECT 1110.540 17.380 1110.800 17.640 ;
        RECT 1114.220 17.380 1114.480 17.640 ;
      LAYER met2 ;
        RECT 1133.310 600.170 1133.590 604.000 ;
        RECT 1132.220 600.030 1133.590 600.170 ;
        RECT 1132.220 19.030 1132.360 600.030 ;
        RECT 1133.310 600.000 1133.590 600.030 ;
        RECT 900.780 18.710 901.040 19.030 ;
        RECT 1110.540 18.710 1110.800 19.030 ;
        RECT 1114.220 18.710 1114.480 19.030 ;
        RECT 1132.160 18.710 1132.420 19.030 ;
        RECT 900.840 2.400 900.980 18.710 ;
        RECT 1110.600 17.670 1110.740 18.710 ;
        RECT 1114.280 17.670 1114.420 18.710 ;
        RECT 1110.540 17.350 1110.800 17.670 ;
        RECT 1114.220 17.350 1114.480 17.670 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1139.490 497.320 1139.810 497.380 ;
        RECT 1139.120 497.180 1139.810 497.320 ;
        RECT 1139.120 496.700 1139.260 497.180 ;
        RECT 1139.490 497.120 1139.810 497.180 ;
        RECT 1139.030 496.440 1139.350 496.700 ;
        RECT 1139.030 448.500 1139.350 448.760 ;
        RECT 1139.120 448.020 1139.260 448.500 ;
        RECT 1139.490 448.020 1139.810 448.080 ;
        RECT 1139.120 447.880 1139.810 448.020 ;
        RECT 1139.490 447.820 1139.810 447.880 ;
        RECT 1137.650 427.620 1137.970 427.680 ;
        RECT 1139.490 427.620 1139.810 427.680 ;
        RECT 1137.650 427.480 1139.810 427.620 ;
        RECT 1137.650 427.420 1137.970 427.480 ;
        RECT 1139.490 427.420 1139.810 427.480 ;
        RECT 1137.650 379.680 1137.970 379.740 ;
        RECT 1138.570 379.680 1138.890 379.740 ;
        RECT 1137.650 379.540 1138.890 379.680 ;
        RECT 1137.650 379.480 1137.970 379.540 ;
        RECT 1138.570 379.480 1138.890 379.540 ;
        RECT 1139.030 303.520 1139.350 303.580 ;
        RECT 1139.950 303.520 1140.270 303.580 ;
        RECT 1139.030 303.380 1140.270 303.520 ;
        RECT 1139.030 303.320 1139.350 303.380 ;
        RECT 1139.950 303.320 1140.270 303.380 ;
        RECT 1138.570 289.580 1138.890 289.640 ;
        RECT 1139.950 289.580 1140.270 289.640 ;
        RECT 1138.570 289.440 1140.270 289.580 ;
        RECT 1138.570 289.380 1138.890 289.440 ;
        RECT 1139.950 289.380 1140.270 289.440 ;
        RECT 1138.570 241.640 1138.890 241.700 ;
        RECT 1139.490 241.640 1139.810 241.700 ;
        RECT 1138.570 241.500 1139.810 241.640 ;
        RECT 1138.570 241.440 1138.890 241.500 ;
        RECT 1139.490 241.440 1139.810 241.500 ;
        RECT 1139.490 207.780 1139.810 208.040 ;
        RECT 1139.580 207.360 1139.720 207.780 ;
        RECT 1139.490 207.100 1139.810 207.360 ;
        RECT 1139.490 158.820 1139.810 159.080 ;
        RECT 1139.580 158.400 1139.720 158.820 ;
        RECT 1139.490 158.140 1139.810 158.400 ;
        RECT 1139.030 145.080 1139.350 145.140 ;
        RECT 1139.490 145.080 1139.810 145.140 ;
        RECT 1139.030 144.940 1139.810 145.080 ;
        RECT 1139.030 144.880 1139.350 144.940 ;
        RECT 1139.490 144.880 1139.810 144.940 ;
        RECT 1014.370 22.000 1014.690 22.060 ;
        RECT 1139.950 22.000 1140.270 22.060 ;
        RECT 1014.370 21.860 1140.270 22.000 ;
        RECT 1014.370 21.800 1014.690 21.860 ;
        RECT 1139.950 21.800 1140.270 21.860 ;
        RECT 918.690 16.900 919.010 16.960 ;
        RECT 1014.370 16.900 1014.690 16.960 ;
        RECT 918.690 16.760 1014.690 16.900 ;
        RECT 918.690 16.700 919.010 16.760 ;
        RECT 1014.370 16.700 1014.690 16.760 ;
      LAYER via ;
        RECT 1139.520 497.120 1139.780 497.380 ;
        RECT 1139.060 496.440 1139.320 496.700 ;
        RECT 1139.060 448.500 1139.320 448.760 ;
        RECT 1139.520 447.820 1139.780 448.080 ;
        RECT 1137.680 427.420 1137.940 427.680 ;
        RECT 1139.520 427.420 1139.780 427.680 ;
        RECT 1137.680 379.480 1137.940 379.740 ;
        RECT 1138.600 379.480 1138.860 379.740 ;
        RECT 1139.060 303.320 1139.320 303.580 ;
        RECT 1139.980 303.320 1140.240 303.580 ;
        RECT 1138.600 289.380 1138.860 289.640 ;
        RECT 1139.980 289.380 1140.240 289.640 ;
        RECT 1138.600 241.440 1138.860 241.700 ;
        RECT 1139.520 241.440 1139.780 241.700 ;
        RECT 1139.520 207.780 1139.780 208.040 ;
        RECT 1139.520 207.100 1139.780 207.360 ;
        RECT 1139.520 158.820 1139.780 159.080 ;
        RECT 1139.520 158.140 1139.780 158.400 ;
        RECT 1139.060 144.880 1139.320 145.140 ;
        RECT 1139.520 144.880 1139.780 145.140 ;
        RECT 1014.400 21.800 1014.660 22.060 ;
        RECT 1139.980 21.800 1140.240 22.060 ;
        RECT 918.720 16.700 918.980 16.960 ;
        RECT 1014.400 16.700 1014.660 16.960 ;
      LAYER met2 ;
        RECT 1142.510 600.170 1142.790 604.000 ;
        RECT 1141.420 600.030 1142.790 600.170 ;
        RECT 1141.420 579.885 1141.560 600.030 ;
        RECT 1142.510 600.000 1142.790 600.030 ;
        RECT 1139.970 579.515 1140.250 579.885 ;
        RECT 1141.350 579.515 1141.630 579.885 ;
        RECT 1140.040 545.090 1140.180 579.515 ;
        RECT 1139.580 544.950 1140.180 545.090 ;
        RECT 1139.580 497.410 1139.720 544.950 ;
        RECT 1139.520 497.090 1139.780 497.410 ;
        RECT 1139.060 496.410 1139.320 496.730 ;
        RECT 1139.120 448.790 1139.260 496.410 ;
        RECT 1139.060 448.470 1139.320 448.790 ;
        RECT 1139.520 447.790 1139.780 448.110 ;
        RECT 1139.580 427.710 1139.720 447.790 ;
        RECT 1137.680 427.390 1137.940 427.710 ;
        RECT 1139.520 427.390 1139.780 427.710 ;
        RECT 1137.740 379.770 1137.880 427.390 ;
        RECT 1137.680 379.450 1137.940 379.770 ;
        RECT 1138.600 379.450 1138.860 379.770 ;
        RECT 1138.660 351.290 1138.800 379.450 ;
        RECT 1138.660 351.150 1139.260 351.290 ;
        RECT 1139.120 303.610 1139.260 351.150 ;
        RECT 1139.060 303.290 1139.320 303.610 ;
        RECT 1139.980 303.290 1140.240 303.610 ;
        RECT 1140.040 289.670 1140.180 303.290 ;
        RECT 1138.600 289.350 1138.860 289.670 ;
        RECT 1139.980 289.350 1140.240 289.670 ;
        RECT 1138.660 241.730 1138.800 289.350 ;
        RECT 1138.600 241.410 1138.860 241.730 ;
        RECT 1139.520 241.410 1139.780 241.730 ;
        RECT 1139.580 208.070 1139.720 241.410 ;
        RECT 1139.520 207.750 1139.780 208.070 ;
        RECT 1139.520 207.070 1139.780 207.390 ;
        RECT 1139.580 159.110 1139.720 207.070 ;
        RECT 1139.520 158.790 1139.780 159.110 ;
        RECT 1139.520 158.110 1139.780 158.430 ;
        RECT 1139.580 145.170 1139.720 158.110 ;
        RECT 1139.060 144.850 1139.320 145.170 ;
        RECT 1139.520 144.850 1139.780 145.170 ;
        RECT 1139.120 144.685 1139.260 144.850 ;
        RECT 1139.050 144.315 1139.330 144.685 ;
        RECT 1139.970 144.315 1140.250 144.685 ;
        RECT 1140.040 22.090 1140.180 144.315 ;
        RECT 1014.400 21.770 1014.660 22.090 ;
        RECT 1139.980 21.770 1140.240 22.090 ;
        RECT 1014.460 16.990 1014.600 21.770 ;
        RECT 918.720 16.670 918.980 16.990 ;
        RECT 1014.400 16.670 1014.660 16.990 ;
        RECT 918.780 2.400 918.920 16.670 ;
        RECT 918.570 -4.800 919.130 2.400 ;
      LAYER via2 ;
        RECT 1139.970 579.560 1140.250 579.840 ;
        RECT 1141.350 579.560 1141.630 579.840 ;
        RECT 1139.050 144.360 1139.330 144.640 ;
        RECT 1139.970 144.360 1140.250 144.640 ;
      LAYER met3 ;
        RECT 1139.945 579.850 1140.275 579.865 ;
        RECT 1141.325 579.850 1141.655 579.865 ;
        RECT 1139.945 579.550 1141.655 579.850 ;
        RECT 1139.945 579.535 1140.275 579.550 ;
        RECT 1141.325 579.535 1141.655 579.550 ;
        RECT 1139.025 144.650 1139.355 144.665 ;
        RECT 1139.945 144.650 1140.275 144.665 ;
        RECT 1139.025 144.350 1140.275 144.650 ;
        RECT 1139.025 144.335 1139.355 144.350 ;
        RECT 1139.945 144.335 1140.275 144.350 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1014.830 22.340 1015.150 22.400 ;
        RECT 1145.930 22.340 1146.250 22.400 ;
        RECT 1014.830 22.200 1146.250 22.340 ;
        RECT 1014.830 22.140 1015.150 22.200 ;
        RECT 1145.930 22.140 1146.250 22.200 ;
        RECT 972.970 16.560 973.290 16.620 ;
        RECT 1014.830 16.560 1015.150 16.620 ;
        RECT 972.970 16.420 1015.150 16.560 ;
        RECT 972.970 16.360 973.290 16.420 ;
        RECT 1014.830 16.360 1015.150 16.420 ;
        RECT 936.170 14.180 936.490 14.240 ;
        RECT 972.970 14.180 973.290 14.240 ;
        RECT 936.170 14.040 973.290 14.180 ;
        RECT 936.170 13.980 936.490 14.040 ;
        RECT 972.970 13.980 973.290 14.040 ;
      LAYER via ;
        RECT 1014.860 22.140 1015.120 22.400 ;
        RECT 1145.960 22.140 1146.220 22.400 ;
        RECT 973.000 16.360 973.260 16.620 ;
        RECT 1014.860 16.360 1015.120 16.620 ;
        RECT 936.200 13.980 936.460 14.240 ;
        RECT 973.000 13.980 973.260 14.240 ;
      LAYER met2 ;
        RECT 1151.710 600.170 1151.990 604.000 ;
        RECT 1149.700 600.030 1151.990 600.170 ;
        RECT 1149.700 587.930 1149.840 600.030 ;
        RECT 1151.710 600.000 1151.990 600.030 ;
        RECT 1146.020 587.790 1149.840 587.930 ;
        RECT 1146.020 22.430 1146.160 587.790 ;
        RECT 1014.860 22.110 1015.120 22.430 ;
        RECT 1145.960 22.110 1146.220 22.430 ;
        RECT 1014.920 16.650 1015.060 22.110 ;
        RECT 973.000 16.330 973.260 16.650 ;
        RECT 1014.860 16.330 1015.120 16.650 ;
        RECT 973.060 14.270 973.200 16.330 ;
        RECT 936.200 13.950 936.460 14.270 ;
        RECT 973.000 13.950 973.260 14.270 ;
        RECT 936.260 2.400 936.400 13.950 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1021.270 23.020 1021.590 23.080 ;
        RECT 1159.730 23.020 1160.050 23.080 ;
        RECT 1021.270 22.880 1160.050 23.020 ;
        RECT 1021.270 22.820 1021.590 22.880 ;
        RECT 1159.730 22.820 1160.050 22.880 ;
        RECT 954.110 15.540 954.430 15.600 ;
        RECT 1021.270 15.540 1021.590 15.600 ;
        RECT 954.110 15.400 1021.590 15.540 ;
        RECT 954.110 15.340 954.430 15.400 ;
        RECT 1021.270 15.340 1021.590 15.400 ;
      LAYER via ;
        RECT 1021.300 22.820 1021.560 23.080 ;
        RECT 1159.760 22.820 1160.020 23.080 ;
        RECT 954.140 15.340 954.400 15.600 ;
        RECT 1021.300 15.340 1021.560 15.600 ;
      LAYER met2 ;
        RECT 1160.910 600.170 1161.190 604.000 ;
        RECT 1159.820 600.030 1161.190 600.170 ;
        RECT 1159.820 23.110 1159.960 600.030 ;
        RECT 1160.910 600.000 1161.190 600.030 ;
        RECT 1021.300 22.790 1021.560 23.110 ;
        RECT 1159.760 22.790 1160.020 23.110 ;
        RECT 1021.360 15.630 1021.500 22.790 ;
        RECT 954.140 15.310 954.400 15.630 ;
        RECT 1021.300 15.310 1021.560 15.630 ;
        RECT 954.200 2.400 954.340 15.310 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1167.090 566.000 1167.410 566.060 ;
        RECT 1168.470 566.000 1168.790 566.060 ;
        RECT 1167.090 565.860 1168.790 566.000 ;
        RECT 1167.090 565.800 1167.410 565.860 ;
        RECT 1168.470 565.800 1168.790 565.860 ;
        RECT 1166.630 524.520 1166.950 524.580 ;
        RECT 1167.550 524.520 1167.870 524.580 ;
        RECT 1166.630 524.380 1167.870 524.520 ;
        RECT 1166.630 524.320 1166.950 524.380 ;
        RECT 1167.550 524.320 1167.870 524.380 ;
        RECT 1166.630 517.380 1166.950 517.440 ;
        RECT 1167.550 517.380 1167.870 517.440 ;
        RECT 1166.630 517.240 1167.870 517.380 ;
        RECT 1166.630 517.180 1166.950 517.240 ;
        RECT 1167.550 517.180 1167.870 517.240 ;
        RECT 1167.550 476.040 1167.870 476.300 ;
        RECT 1167.640 475.620 1167.780 476.040 ;
        RECT 1167.550 475.360 1167.870 475.620 ;
        RECT 1166.170 373.220 1166.490 373.280 ;
        RECT 1168.470 373.220 1168.790 373.280 ;
        RECT 1166.170 373.080 1168.790 373.220 ;
        RECT 1166.170 373.020 1166.490 373.080 ;
        RECT 1168.470 373.020 1168.790 373.080 ;
        RECT 1166.630 289.580 1166.950 289.640 ;
        RECT 1167.550 289.580 1167.870 289.640 ;
        RECT 1166.630 289.440 1167.870 289.580 ;
        RECT 1166.630 289.380 1166.950 289.440 ;
        RECT 1167.550 289.380 1167.870 289.440 ;
        RECT 1166.630 241.640 1166.950 241.700 ;
        RECT 1168.010 241.640 1168.330 241.700 ;
        RECT 1166.630 241.500 1168.330 241.640 ;
        RECT 1166.630 241.440 1166.950 241.500 ;
        RECT 1168.010 241.440 1168.330 241.500 ;
        RECT 1166.170 193.360 1166.490 193.420 ;
        RECT 1168.010 193.360 1168.330 193.420 ;
        RECT 1166.170 193.220 1168.330 193.360 ;
        RECT 1166.170 193.160 1166.490 193.220 ;
        RECT 1168.010 193.160 1168.330 193.220 ;
        RECT 1166.630 144.400 1166.950 144.460 ;
        RECT 1167.550 144.400 1167.870 144.460 ;
        RECT 1166.630 144.260 1167.870 144.400 ;
        RECT 1166.630 144.200 1166.950 144.260 ;
        RECT 1167.550 144.200 1167.870 144.260 ;
        RECT 1021.730 23.360 1022.050 23.420 ;
        RECT 1167.550 23.360 1167.870 23.420 ;
        RECT 1021.730 23.220 1167.870 23.360 ;
        RECT 1021.730 23.160 1022.050 23.220 ;
        RECT 1167.550 23.160 1167.870 23.220 ;
        RECT 972.050 15.200 972.370 15.260 ;
        RECT 1021.730 15.200 1022.050 15.260 ;
        RECT 972.050 15.060 1022.050 15.200 ;
        RECT 972.050 15.000 972.370 15.060 ;
        RECT 1021.730 15.000 1022.050 15.060 ;
      LAYER via ;
        RECT 1167.120 565.800 1167.380 566.060 ;
        RECT 1168.500 565.800 1168.760 566.060 ;
        RECT 1166.660 524.320 1166.920 524.580 ;
        RECT 1167.580 524.320 1167.840 524.580 ;
        RECT 1166.660 517.180 1166.920 517.440 ;
        RECT 1167.580 517.180 1167.840 517.440 ;
        RECT 1167.580 476.040 1167.840 476.300 ;
        RECT 1167.580 475.360 1167.840 475.620 ;
        RECT 1166.200 373.020 1166.460 373.280 ;
        RECT 1168.500 373.020 1168.760 373.280 ;
        RECT 1166.660 289.380 1166.920 289.640 ;
        RECT 1167.580 289.380 1167.840 289.640 ;
        RECT 1166.660 241.440 1166.920 241.700 ;
        RECT 1168.040 241.440 1168.300 241.700 ;
        RECT 1166.200 193.160 1166.460 193.420 ;
        RECT 1168.040 193.160 1168.300 193.420 ;
        RECT 1166.660 144.200 1166.920 144.460 ;
        RECT 1167.580 144.200 1167.840 144.460 ;
        RECT 1021.760 23.160 1022.020 23.420 ;
        RECT 1167.580 23.160 1167.840 23.420 ;
        RECT 972.080 15.000 972.340 15.260 ;
        RECT 1021.760 15.000 1022.020 15.260 ;
      LAYER met2 ;
        RECT 1170.110 600.170 1170.390 604.000 ;
        RECT 1168.560 600.030 1170.390 600.170 ;
        RECT 1168.560 566.090 1168.700 600.030 ;
        RECT 1170.110 600.000 1170.390 600.030 ;
        RECT 1167.120 565.770 1167.380 566.090 ;
        RECT 1168.500 565.770 1168.760 566.090 ;
        RECT 1167.180 532.170 1167.320 565.770 ;
        RECT 1167.180 532.030 1167.780 532.170 ;
        RECT 1167.640 524.610 1167.780 532.030 ;
        RECT 1166.660 524.290 1166.920 524.610 ;
        RECT 1167.580 524.290 1167.840 524.610 ;
        RECT 1166.720 517.470 1166.860 524.290 ;
        RECT 1166.660 517.150 1166.920 517.470 ;
        RECT 1167.580 517.150 1167.840 517.470 ;
        RECT 1167.640 476.330 1167.780 517.150 ;
        RECT 1167.580 476.010 1167.840 476.330 ;
        RECT 1167.580 475.330 1167.840 475.650 ;
        RECT 1167.640 447.850 1167.780 475.330 ;
        RECT 1167.180 447.710 1167.780 447.850 ;
        RECT 1167.180 401.045 1167.320 447.710 ;
        RECT 1167.110 400.675 1167.390 401.045 ;
        RECT 1166.190 399.315 1166.470 399.685 ;
        RECT 1166.260 373.310 1166.400 399.315 ;
        RECT 1166.200 372.990 1166.460 373.310 ;
        RECT 1168.500 372.990 1168.760 373.310 ;
        RECT 1168.560 290.090 1168.700 372.990 ;
        RECT 1167.640 289.950 1168.700 290.090 ;
        RECT 1167.640 289.670 1167.780 289.950 ;
        RECT 1166.660 289.350 1166.920 289.670 ;
        RECT 1167.580 289.350 1167.840 289.670 ;
        RECT 1166.720 241.730 1166.860 289.350 ;
        RECT 1166.660 241.410 1166.920 241.730 ;
        RECT 1168.040 241.410 1168.300 241.730 ;
        RECT 1168.100 193.450 1168.240 241.410 ;
        RECT 1166.200 193.130 1166.460 193.450 ;
        RECT 1168.040 193.130 1168.300 193.450 ;
        RECT 1166.260 158.170 1166.400 193.130 ;
        RECT 1166.260 158.030 1166.860 158.170 ;
        RECT 1166.720 144.490 1166.860 158.030 ;
        RECT 1166.660 144.170 1166.920 144.490 ;
        RECT 1167.580 144.170 1167.840 144.490 ;
        RECT 1167.640 23.450 1167.780 144.170 ;
        RECT 1021.760 23.130 1022.020 23.450 ;
        RECT 1167.580 23.130 1167.840 23.450 ;
        RECT 1021.820 15.290 1021.960 23.130 ;
        RECT 972.080 14.970 972.340 15.290 ;
        RECT 1021.760 14.970 1022.020 15.290 ;
        RECT 972.140 2.400 972.280 14.970 ;
        RECT 971.930 -4.800 972.490 2.400 ;
      LAYER via2 ;
        RECT 1167.110 400.720 1167.390 401.000 ;
        RECT 1166.190 399.360 1166.470 399.640 ;
      LAYER met3 ;
        RECT 1167.085 401.010 1167.415 401.025 ;
        RECT 1166.870 400.695 1167.415 401.010 ;
        RECT 1166.165 399.650 1166.495 399.665 ;
        RECT 1166.870 399.650 1167.170 400.695 ;
        RECT 1166.165 399.350 1167.170 399.650 ;
        RECT 1166.165 399.335 1166.495 399.350 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1000.570 557.500 1000.890 557.560 ;
        RECT 1003.330 557.500 1003.650 557.560 ;
        RECT 1000.570 557.360 1003.650 557.500 ;
        RECT 1000.570 557.300 1000.890 557.360 ;
        RECT 1003.330 557.300 1003.650 557.360 ;
        RECT 650.970 35.940 651.290 36.000 ;
        RECT 1000.570 35.940 1000.890 36.000 ;
        RECT 650.970 35.800 1000.890 35.940 ;
        RECT 650.970 35.740 651.290 35.800 ;
        RECT 1000.570 35.740 1000.890 35.800 ;
      LAYER via ;
        RECT 1000.600 557.300 1000.860 557.560 ;
        RECT 1003.360 557.300 1003.620 557.560 ;
        RECT 651.000 35.740 651.260 36.000 ;
        RECT 1000.600 35.740 1000.860 36.000 ;
      LAYER met2 ;
        RECT 1004.970 600.170 1005.250 604.000 ;
        RECT 1003.420 600.030 1005.250 600.170 ;
        RECT 1003.420 557.590 1003.560 600.030 ;
        RECT 1004.970 600.000 1005.250 600.030 ;
        RECT 1000.600 557.270 1000.860 557.590 ;
        RECT 1003.360 557.270 1003.620 557.590 ;
        RECT 1000.660 36.030 1000.800 557.270 ;
        RECT 651.000 35.710 651.260 36.030 ;
        RECT 1000.600 35.710 1000.860 36.030 ;
        RECT 651.060 2.400 651.200 35.710 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1034.610 23.700 1034.930 23.760 ;
        RECT 1173.530 23.700 1173.850 23.760 ;
        RECT 1034.610 23.560 1173.850 23.700 ;
        RECT 1034.610 23.500 1034.930 23.560 ;
        RECT 1173.530 23.500 1173.850 23.560 ;
        RECT 989.990 19.280 990.310 19.340 ;
        RECT 1034.610 19.280 1034.930 19.340 ;
        RECT 989.990 19.140 1034.930 19.280 ;
        RECT 989.990 19.080 990.310 19.140 ;
        RECT 1034.610 19.080 1034.930 19.140 ;
      LAYER via ;
        RECT 1034.640 23.500 1034.900 23.760 ;
        RECT 1173.560 23.500 1173.820 23.760 ;
        RECT 990.020 19.080 990.280 19.340 ;
        RECT 1034.640 19.080 1034.900 19.340 ;
      LAYER met2 ;
        RECT 1179.310 600.170 1179.590 604.000 ;
        RECT 1177.300 600.030 1179.590 600.170 ;
        RECT 1177.300 588.440 1177.440 600.030 ;
        RECT 1179.310 600.000 1179.590 600.030 ;
        RECT 1173.620 588.300 1177.440 588.440 ;
        RECT 1173.620 23.790 1173.760 588.300 ;
        RECT 1034.640 23.470 1034.900 23.790 ;
        RECT 1173.560 23.470 1173.820 23.790 ;
        RECT 1034.700 19.370 1034.840 23.470 ;
        RECT 990.020 19.050 990.280 19.370 ;
        RECT 1034.640 19.050 1034.900 19.370 ;
        RECT 990.080 2.400 990.220 19.050 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.510 27.100 1041.830 27.160 ;
        RECT 1187.330 27.100 1187.650 27.160 ;
        RECT 1041.510 26.960 1187.650 27.100 ;
        RECT 1041.510 26.900 1041.830 26.960 ;
        RECT 1187.330 26.900 1187.650 26.960 ;
        RECT 1007.470 14.520 1007.790 14.580 ;
        RECT 1041.510 14.520 1041.830 14.580 ;
        RECT 1007.470 14.380 1041.830 14.520 ;
        RECT 1007.470 14.320 1007.790 14.380 ;
        RECT 1041.510 14.320 1041.830 14.380 ;
      LAYER via ;
        RECT 1041.540 26.900 1041.800 27.160 ;
        RECT 1187.360 26.900 1187.620 27.160 ;
        RECT 1007.500 14.320 1007.760 14.580 ;
        RECT 1041.540 14.320 1041.800 14.580 ;
      LAYER met2 ;
        RECT 1188.510 600.170 1188.790 604.000 ;
        RECT 1187.420 600.030 1188.790 600.170 ;
        RECT 1187.420 27.190 1187.560 600.030 ;
        RECT 1188.510 600.000 1188.790 600.030 ;
        RECT 1041.540 26.870 1041.800 27.190 ;
        RECT 1187.360 26.870 1187.620 27.190 ;
        RECT 1041.600 14.610 1041.740 26.870 ;
        RECT 1007.500 14.290 1007.760 14.610 ;
        RECT 1041.540 14.290 1041.800 14.610 ;
        RECT 1007.560 2.400 1007.700 14.290 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1194.690 579.600 1195.010 579.660 ;
        RECT 1195.610 579.600 1195.930 579.660 ;
        RECT 1194.690 579.460 1195.930 579.600 ;
        RECT 1194.690 579.400 1195.010 579.460 ;
        RECT 1195.610 579.400 1195.930 579.460 ;
        RECT 1194.690 337.860 1195.010 337.920 ;
        RECT 1195.610 337.860 1195.930 337.920 ;
        RECT 1194.690 337.720 1195.930 337.860 ;
        RECT 1194.690 337.660 1195.010 337.720 ;
        RECT 1195.610 337.660 1195.930 337.720 ;
        RECT 1194.690 289.920 1195.010 289.980 ;
        RECT 1195.610 289.920 1195.930 289.980 ;
        RECT 1194.690 289.780 1195.930 289.920 ;
        RECT 1194.690 289.720 1195.010 289.780 ;
        RECT 1195.610 289.720 1195.930 289.780 ;
        RECT 1193.770 241.300 1194.090 241.360 ;
        RECT 1194.690 241.300 1195.010 241.360 ;
        RECT 1193.770 241.160 1195.010 241.300 ;
        RECT 1193.770 241.100 1194.090 241.160 ;
        RECT 1194.690 241.100 1195.010 241.160 ;
        RECT 1194.690 120.940 1195.010 121.000 ;
        RECT 1195.610 120.940 1195.930 121.000 ;
        RECT 1194.690 120.800 1195.930 120.940 ;
        RECT 1194.690 120.740 1195.010 120.800 ;
        RECT 1195.610 120.740 1195.930 120.800 ;
        RECT 1194.690 96.800 1195.010 96.860 ;
        RECT 1195.610 96.800 1195.930 96.860 ;
        RECT 1194.690 96.660 1195.930 96.800 ;
        RECT 1194.690 96.600 1195.010 96.660 ;
        RECT 1195.610 96.600 1195.930 96.660 ;
        RECT 1164.330 48.180 1164.650 48.240 ;
        RECT 1194.690 48.180 1195.010 48.240 ;
        RECT 1164.330 48.040 1195.010 48.180 ;
        RECT 1164.330 47.980 1164.650 48.040 ;
        RECT 1194.690 47.980 1195.010 48.040 ;
        RECT 1046.110 27.440 1046.430 27.500 ;
        RECT 1164.330 27.440 1164.650 27.500 ;
        RECT 1046.110 27.300 1164.650 27.440 ;
        RECT 1046.110 27.240 1046.430 27.300 ;
        RECT 1164.330 27.240 1164.650 27.300 ;
        RECT 1025.410 14.180 1025.730 14.240 ;
        RECT 1046.110 14.180 1046.430 14.240 ;
        RECT 1025.410 14.040 1046.430 14.180 ;
        RECT 1025.410 13.980 1025.730 14.040 ;
        RECT 1046.110 13.980 1046.430 14.040 ;
      LAYER via ;
        RECT 1194.720 579.400 1194.980 579.660 ;
        RECT 1195.640 579.400 1195.900 579.660 ;
        RECT 1194.720 337.660 1194.980 337.920 ;
        RECT 1195.640 337.660 1195.900 337.920 ;
        RECT 1194.720 289.720 1194.980 289.980 ;
        RECT 1195.640 289.720 1195.900 289.980 ;
        RECT 1193.800 241.100 1194.060 241.360 ;
        RECT 1194.720 241.100 1194.980 241.360 ;
        RECT 1194.720 120.740 1194.980 121.000 ;
        RECT 1195.640 120.740 1195.900 121.000 ;
        RECT 1194.720 96.600 1194.980 96.860 ;
        RECT 1195.640 96.600 1195.900 96.860 ;
        RECT 1164.360 47.980 1164.620 48.240 ;
        RECT 1194.720 47.980 1194.980 48.240 ;
        RECT 1046.140 27.240 1046.400 27.500 ;
        RECT 1164.360 27.240 1164.620 27.500 ;
        RECT 1025.440 13.980 1025.700 14.240 ;
        RECT 1046.140 13.980 1046.400 14.240 ;
      LAYER met2 ;
        RECT 1197.710 600.170 1197.990 604.000 ;
        RECT 1196.620 600.030 1197.990 600.170 ;
        RECT 1196.620 596.770 1196.760 600.030 ;
        RECT 1197.710 600.000 1197.990 600.030 ;
        RECT 1194.780 596.630 1196.760 596.770 ;
        RECT 1194.780 579.690 1194.920 596.630 ;
        RECT 1194.720 579.370 1194.980 579.690 ;
        RECT 1195.640 579.370 1195.900 579.690 ;
        RECT 1195.700 531.605 1195.840 579.370 ;
        RECT 1194.710 531.235 1194.990 531.605 ;
        RECT 1195.630 531.235 1195.910 531.605 ;
        RECT 1194.780 400.930 1194.920 531.235 ;
        RECT 1194.320 400.790 1194.920 400.930 ;
        RECT 1194.320 400.250 1194.460 400.790 ;
        RECT 1194.320 400.110 1194.920 400.250 ;
        RECT 1194.780 337.950 1194.920 400.110 ;
        RECT 1194.720 337.630 1194.980 337.950 ;
        RECT 1195.640 337.630 1195.900 337.950 ;
        RECT 1195.700 290.010 1195.840 337.630 ;
        RECT 1194.720 289.690 1194.980 290.010 ;
        RECT 1195.640 289.690 1195.900 290.010 ;
        RECT 1194.780 241.390 1194.920 289.690 ;
        RECT 1193.800 241.070 1194.060 241.390 ;
        RECT 1194.720 241.070 1194.980 241.390 ;
        RECT 1193.860 216.650 1194.000 241.070 ;
        RECT 1193.860 216.510 1194.920 216.650 ;
        RECT 1194.780 121.030 1194.920 216.510 ;
        RECT 1194.720 120.710 1194.980 121.030 ;
        RECT 1195.640 120.710 1195.900 121.030 ;
        RECT 1195.700 96.890 1195.840 120.710 ;
        RECT 1194.720 96.570 1194.980 96.890 ;
        RECT 1195.640 96.570 1195.900 96.890 ;
        RECT 1194.780 48.270 1194.920 96.570 ;
        RECT 1164.360 47.950 1164.620 48.270 ;
        RECT 1194.720 47.950 1194.980 48.270 ;
        RECT 1164.420 27.530 1164.560 47.950 ;
        RECT 1046.140 27.210 1046.400 27.530 ;
        RECT 1164.360 27.210 1164.620 27.530 ;
        RECT 1046.200 14.270 1046.340 27.210 ;
        RECT 1025.440 13.950 1025.700 14.270 ;
        RECT 1046.140 13.950 1046.400 14.270 ;
        RECT 1025.500 2.400 1025.640 13.950 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
      LAYER via2 ;
        RECT 1194.710 531.280 1194.990 531.560 ;
        RECT 1195.630 531.280 1195.910 531.560 ;
      LAYER met3 ;
        RECT 1194.685 531.570 1195.015 531.585 ;
        RECT 1195.605 531.570 1195.935 531.585 ;
        RECT 1194.685 531.270 1195.935 531.570 ;
        RECT 1194.685 531.255 1195.015 531.270 ;
        RECT 1195.605 531.255 1195.935 531.270 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1201.590 400.760 1201.910 400.820 ;
        RECT 1201.220 400.620 1201.910 400.760 ;
        RECT 1201.220 400.480 1201.360 400.620 ;
        RECT 1201.590 400.560 1201.910 400.620 ;
        RECT 1201.130 400.220 1201.450 400.480 ;
        RECT 1043.350 24.380 1043.670 24.440 ;
        RECT 1200.670 24.380 1200.990 24.440 ;
        RECT 1043.350 24.240 1200.990 24.380 ;
        RECT 1043.350 24.180 1043.670 24.240 ;
        RECT 1200.670 24.180 1200.990 24.240 ;
      LAYER via ;
        RECT 1201.620 400.560 1201.880 400.820 ;
        RECT 1201.160 400.220 1201.420 400.480 ;
        RECT 1043.380 24.180 1043.640 24.440 ;
        RECT 1200.700 24.180 1200.960 24.440 ;
      LAYER met2 ;
        RECT 1206.910 600.170 1207.190 604.000 ;
        RECT 1204.440 600.030 1207.190 600.170 ;
        RECT 1204.440 596.770 1204.580 600.030 ;
        RECT 1206.910 600.000 1207.190 600.030 ;
        RECT 1202.600 596.630 1204.580 596.770 ;
        RECT 1202.600 569.570 1202.740 596.630 ;
        RECT 1201.220 569.430 1202.740 569.570 ;
        RECT 1201.220 507.010 1201.360 569.430 ;
        RECT 1201.220 506.870 1202.280 507.010 ;
        RECT 1202.140 496.130 1202.280 506.870 ;
        RECT 1201.680 495.990 1202.280 496.130 ;
        RECT 1201.680 400.850 1201.820 495.990 ;
        RECT 1201.620 400.530 1201.880 400.850 ;
        RECT 1201.160 400.190 1201.420 400.510 ;
        RECT 1201.220 351.970 1201.360 400.190 ;
        RECT 1200.760 351.830 1201.360 351.970 ;
        RECT 1200.760 351.290 1200.900 351.830 ;
        RECT 1200.760 351.150 1201.360 351.290 ;
        RECT 1201.220 255.410 1201.360 351.150 ;
        RECT 1200.760 255.270 1201.360 255.410 ;
        RECT 1200.760 254.730 1200.900 255.270 ;
        RECT 1200.760 254.590 1201.360 254.730 ;
        RECT 1201.220 158.850 1201.360 254.590 ;
        RECT 1200.760 158.710 1201.360 158.850 ;
        RECT 1200.760 158.170 1200.900 158.710 ;
        RECT 1200.760 158.030 1201.360 158.170 ;
        RECT 1201.220 62.290 1201.360 158.030 ;
        RECT 1200.760 62.150 1201.360 62.290 ;
        RECT 1200.760 24.470 1200.900 62.150 ;
        RECT 1043.380 24.150 1043.640 24.470 ;
        RECT 1200.700 24.150 1200.960 24.470 ;
        RECT 1043.440 2.400 1043.580 24.150 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1061.290 24.040 1061.610 24.100 ;
        RECT 1214.930 24.040 1215.250 24.100 ;
        RECT 1061.290 23.900 1215.250 24.040 ;
        RECT 1061.290 23.840 1061.610 23.900 ;
        RECT 1214.930 23.840 1215.250 23.900 ;
      LAYER via ;
        RECT 1061.320 23.840 1061.580 24.100 ;
        RECT 1214.960 23.840 1215.220 24.100 ;
      LAYER met2 ;
        RECT 1216.110 600.170 1216.390 604.000 ;
        RECT 1215.020 600.030 1216.390 600.170 ;
        RECT 1215.020 24.130 1215.160 600.030 ;
        RECT 1216.110 600.000 1216.390 600.030 ;
        RECT 1061.320 23.810 1061.580 24.130 ;
        RECT 1214.960 23.810 1215.220 24.130 ;
        RECT 1061.380 2.400 1061.520 23.810 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1221.370 379.680 1221.690 379.740 ;
        RECT 1222.290 379.680 1222.610 379.740 ;
        RECT 1221.370 379.540 1222.610 379.680 ;
        RECT 1221.370 379.480 1221.690 379.540 ;
        RECT 1222.290 379.480 1222.610 379.540 ;
        RECT 1221.830 331.400 1222.150 331.460 ;
        RECT 1223.210 331.400 1223.530 331.460 ;
        RECT 1221.830 331.260 1223.530 331.400 ;
        RECT 1221.830 331.200 1222.150 331.260 ;
        RECT 1223.210 331.200 1223.530 331.260 ;
        RECT 1221.370 283.120 1221.690 283.180 ;
        RECT 1222.750 283.120 1223.070 283.180 ;
        RECT 1221.370 282.980 1223.070 283.120 ;
        RECT 1221.370 282.920 1221.690 282.980 ;
        RECT 1222.750 282.920 1223.070 282.980 ;
        RECT 1221.370 193.360 1221.690 193.420 ;
        RECT 1222.750 193.360 1223.070 193.420 ;
        RECT 1221.370 193.220 1223.070 193.360 ;
        RECT 1221.370 193.160 1221.690 193.220 ;
        RECT 1222.750 193.160 1223.070 193.220 ;
        RECT 1220.450 186.220 1220.770 186.280 ;
        RECT 1221.370 186.220 1221.690 186.280 ;
        RECT 1220.450 186.080 1221.690 186.220 ;
        RECT 1220.450 186.020 1220.770 186.080 ;
        RECT 1221.370 186.020 1221.690 186.080 ;
        RECT 1220.450 138.280 1220.770 138.340 ;
        RECT 1221.830 138.280 1222.150 138.340 ;
        RECT 1220.450 138.140 1222.150 138.280 ;
        RECT 1220.450 138.080 1220.770 138.140 ;
        RECT 1221.830 138.080 1222.150 138.140 ;
        RECT 1221.830 110.400 1222.150 110.460 ;
        RECT 1222.750 110.400 1223.070 110.460 ;
        RECT 1221.830 110.260 1223.070 110.400 ;
        RECT 1221.830 110.200 1222.150 110.260 ;
        RECT 1222.750 110.200 1223.070 110.260 ;
        RECT 1079.230 24.720 1079.550 24.780 ;
        RECT 1222.750 24.720 1223.070 24.780 ;
        RECT 1079.230 24.580 1223.070 24.720 ;
        RECT 1079.230 24.520 1079.550 24.580 ;
        RECT 1222.750 24.520 1223.070 24.580 ;
      LAYER via ;
        RECT 1221.400 379.480 1221.660 379.740 ;
        RECT 1222.320 379.480 1222.580 379.740 ;
        RECT 1221.860 331.200 1222.120 331.460 ;
        RECT 1223.240 331.200 1223.500 331.460 ;
        RECT 1221.400 282.920 1221.660 283.180 ;
        RECT 1222.780 282.920 1223.040 283.180 ;
        RECT 1221.400 193.160 1221.660 193.420 ;
        RECT 1222.780 193.160 1223.040 193.420 ;
        RECT 1220.480 186.020 1220.740 186.280 ;
        RECT 1221.400 186.020 1221.660 186.280 ;
        RECT 1220.480 138.080 1220.740 138.340 ;
        RECT 1221.860 138.080 1222.120 138.340 ;
        RECT 1221.860 110.200 1222.120 110.460 ;
        RECT 1222.780 110.200 1223.040 110.460 ;
        RECT 1079.260 24.520 1079.520 24.780 ;
        RECT 1222.780 24.520 1223.040 24.780 ;
      LAYER met2 ;
        RECT 1225.310 600.170 1225.590 604.000 ;
        RECT 1222.840 600.030 1225.590 600.170 ;
        RECT 1222.840 596.770 1222.980 600.030 ;
        RECT 1225.310 600.000 1225.590 600.030 ;
        RECT 1222.380 596.630 1222.980 596.770 ;
        RECT 1222.380 555.290 1222.520 596.630 ;
        RECT 1221.460 555.150 1222.520 555.290 ;
        RECT 1221.460 496.810 1221.600 555.150 ;
        RECT 1221.460 496.670 1222.520 496.810 ;
        RECT 1222.380 379.770 1222.520 496.670 ;
        RECT 1221.400 379.450 1221.660 379.770 ;
        RECT 1222.320 379.450 1222.580 379.770 ;
        RECT 1221.460 379.285 1221.600 379.450 ;
        RECT 1221.390 378.915 1221.670 379.285 ;
        RECT 1223.230 378.915 1223.510 379.285 ;
        RECT 1223.300 331.490 1223.440 378.915 ;
        RECT 1221.860 331.170 1222.120 331.490 ;
        RECT 1223.240 331.170 1223.500 331.490 ;
        RECT 1221.920 330.890 1222.060 331.170 ;
        RECT 1221.460 330.750 1222.060 330.890 ;
        RECT 1221.460 283.210 1221.600 330.750 ;
        RECT 1221.400 282.890 1221.660 283.210 ;
        RECT 1222.780 282.890 1223.040 283.210 ;
        RECT 1222.840 193.450 1222.980 282.890 ;
        RECT 1221.400 193.130 1221.660 193.450 ;
        RECT 1222.780 193.130 1223.040 193.450 ;
        RECT 1221.460 186.310 1221.600 193.130 ;
        RECT 1220.480 185.990 1220.740 186.310 ;
        RECT 1221.400 185.990 1221.660 186.310 ;
        RECT 1220.540 138.370 1220.680 185.990 ;
        RECT 1220.480 138.050 1220.740 138.370 ;
        RECT 1221.860 138.050 1222.120 138.370 ;
        RECT 1221.920 110.490 1222.060 138.050 ;
        RECT 1221.860 110.170 1222.120 110.490 ;
        RECT 1222.780 110.170 1223.040 110.490 ;
        RECT 1222.840 60.250 1222.980 110.170 ;
        RECT 1222.840 60.110 1223.440 60.250 ;
        RECT 1223.300 58.890 1223.440 60.110 ;
        RECT 1222.840 58.750 1223.440 58.890 ;
        RECT 1222.840 24.810 1222.980 58.750 ;
        RECT 1079.260 24.490 1079.520 24.810 ;
        RECT 1222.780 24.490 1223.040 24.810 ;
        RECT 1079.320 2.400 1079.460 24.490 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
      LAYER via2 ;
        RECT 1221.390 378.960 1221.670 379.240 ;
        RECT 1223.230 378.960 1223.510 379.240 ;
      LAYER met3 ;
        RECT 1221.365 379.250 1221.695 379.265 ;
        RECT 1223.205 379.250 1223.535 379.265 ;
        RECT 1221.365 378.950 1223.535 379.250 ;
        RECT 1221.365 378.935 1221.695 378.950 ;
        RECT 1223.205 378.935 1223.535 378.950 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1228.730 550.020 1229.050 550.080 ;
        RECT 1232.870 550.020 1233.190 550.080 ;
        RECT 1228.730 549.880 1233.190 550.020 ;
        RECT 1228.730 549.820 1229.050 549.880 ;
        RECT 1232.870 549.820 1233.190 549.880 ;
        RECT 1096.710 25.060 1097.030 25.120 ;
        RECT 1228.730 25.060 1229.050 25.120 ;
        RECT 1096.710 24.920 1229.050 25.060 ;
        RECT 1096.710 24.860 1097.030 24.920 ;
        RECT 1228.730 24.860 1229.050 24.920 ;
      LAYER via ;
        RECT 1228.760 549.820 1229.020 550.080 ;
        RECT 1232.900 549.820 1233.160 550.080 ;
        RECT 1096.740 24.860 1097.000 25.120 ;
        RECT 1228.760 24.860 1229.020 25.120 ;
      LAYER met2 ;
        RECT 1234.510 600.170 1234.790 604.000 ;
        RECT 1232.960 600.030 1234.790 600.170 ;
        RECT 1232.960 550.110 1233.100 600.030 ;
        RECT 1234.510 600.000 1234.790 600.030 ;
        RECT 1228.760 549.790 1229.020 550.110 ;
        RECT 1232.900 549.790 1233.160 550.110 ;
        RECT 1228.820 25.150 1228.960 549.790 ;
        RECT 1096.740 24.830 1097.000 25.150 ;
        RECT 1228.760 24.830 1229.020 25.150 ;
        RECT 1096.800 2.400 1096.940 24.830 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1114.650 17.580 1114.970 17.640 ;
        RECT 1242.530 17.580 1242.850 17.640 ;
        RECT 1114.650 17.440 1242.850 17.580 ;
        RECT 1114.650 17.380 1114.970 17.440 ;
        RECT 1242.530 17.380 1242.850 17.440 ;
      LAYER via ;
        RECT 1114.680 17.380 1114.940 17.640 ;
        RECT 1242.560 17.380 1242.820 17.640 ;
      LAYER met2 ;
        RECT 1243.710 600.170 1243.990 604.000 ;
        RECT 1242.620 600.030 1243.990 600.170 ;
        RECT 1242.620 17.670 1242.760 600.030 ;
        RECT 1243.710 600.000 1243.990 600.030 ;
        RECT 1114.680 17.350 1114.940 17.670 ;
        RECT 1242.560 17.350 1242.820 17.670 ;
        RECT 1114.740 2.400 1114.880 17.350 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1250.350 572.800 1250.670 572.860 ;
        RECT 1251.730 572.800 1252.050 572.860 ;
        RECT 1250.350 572.660 1252.050 572.800 ;
        RECT 1250.350 572.600 1250.670 572.660 ;
        RECT 1251.730 572.600 1252.050 572.660 ;
        RECT 1249.430 496.780 1249.750 497.040 ;
        RECT 1249.520 496.640 1249.660 496.780 ;
        RECT 1249.890 496.640 1250.210 496.700 ;
        RECT 1249.520 496.500 1250.210 496.640 ;
        RECT 1249.890 496.440 1250.210 496.500 ;
        RECT 1249.430 400.760 1249.750 400.820 ;
        RECT 1249.060 400.620 1249.750 400.760 ;
        RECT 1249.060 400.480 1249.200 400.620 ;
        RECT 1249.430 400.560 1249.750 400.620 ;
        RECT 1248.970 400.220 1249.290 400.480 ;
        RECT 1248.970 379.340 1249.290 379.400 ;
        RECT 1249.430 379.340 1249.750 379.400 ;
        RECT 1248.970 379.200 1249.750 379.340 ;
        RECT 1248.970 379.140 1249.290 379.200 ;
        RECT 1249.430 379.140 1249.750 379.200 ;
        RECT 1249.430 351.940 1249.750 352.200 ;
        RECT 1249.520 351.800 1249.660 351.940 ;
        RECT 1249.890 351.800 1250.210 351.860 ;
        RECT 1249.520 351.660 1250.210 351.800 ;
        RECT 1249.890 351.600 1250.210 351.660 ;
        RECT 1249.430 330.860 1249.750 331.120 ;
        RECT 1249.520 330.720 1249.660 330.860 ;
        RECT 1250.810 330.720 1251.130 330.780 ;
        RECT 1249.520 330.580 1251.130 330.720 ;
        RECT 1250.810 330.520 1251.130 330.580 ;
        RECT 1250.350 283.120 1250.670 283.180 ;
        RECT 1250.810 283.120 1251.130 283.180 ;
        RECT 1250.350 282.980 1251.130 283.120 ;
        RECT 1250.350 282.920 1250.670 282.980 ;
        RECT 1250.810 282.920 1251.130 282.980 ;
        RECT 1248.970 193.360 1249.290 193.420 ;
        RECT 1250.350 193.360 1250.670 193.420 ;
        RECT 1248.970 193.220 1250.670 193.360 ;
        RECT 1248.970 193.160 1249.290 193.220 ;
        RECT 1250.350 193.160 1250.670 193.220 ;
        RECT 1248.970 186.220 1249.290 186.280 ;
        RECT 1250.810 186.220 1251.130 186.280 ;
        RECT 1248.970 186.080 1251.130 186.220 ;
        RECT 1248.970 186.020 1249.290 186.080 ;
        RECT 1250.810 186.020 1251.130 186.080 ;
        RECT 1249.430 138.280 1249.750 138.340 ;
        RECT 1250.810 138.280 1251.130 138.340 ;
        RECT 1249.430 138.140 1251.130 138.280 ;
        RECT 1249.430 138.080 1249.750 138.140 ;
        RECT 1250.810 138.080 1251.130 138.140 ;
        RECT 1249.430 110.400 1249.750 110.460 ;
        RECT 1250.350 110.400 1250.670 110.460 ;
        RECT 1249.430 110.260 1250.670 110.400 ;
        RECT 1249.430 110.200 1249.750 110.260 ;
        RECT 1250.350 110.200 1250.670 110.260 ;
        RECT 1132.590 18.600 1132.910 18.660 ;
        RECT 1132.590 18.460 1146.160 18.600 ;
        RECT 1132.590 18.400 1132.910 18.460 ;
        RECT 1146.020 17.920 1146.160 18.460 ;
        RECT 1250.350 17.920 1250.670 17.980 ;
        RECT 1146.020 17.780 1250.670 17.920 ;
        RECT 1250.350 17.720 1250.670 17.780 ;
      LAYER via ;
        RECT 1250.380 572.600 1250.640 572.860 ;
        RECT 1251.760 572.600 1252.020 572.860 ;
        RECT 1249.460 496.780 1249.720 497.040 ;
        RECT 1249.920 496.440 1250.180 496.700 ;
        RECT 1249.460 400.560 1249.720 400.820 ;
        RECT 1249.000 400.220 1249.260 400.480 ;
        RECT 1249.000 379.140 1249.260 379.400 ;
        RECT 1249.460 379.140 1249.720 379.400 ;
        RECT 1249.460 351.940 1249.720 352.200 ;
        RECT 1249.920 351.600 1250.180 351.860 ;
        RECT 1249.460 330.860 1249.720 331.120 ;
        RECT 1250.840 330.520 1251.100 330.780 ;
        RECT 1250.380 282.920 1250.640 283.180 ;
        RECT 1250.840 282.920 1251.100 283.180 ;
        RECT 1249.000 193.160 1249.260 193.420 ;
        RECT 1250.380 193.160 1250.640 193.420 ;
        RECT 1249.000 186.020 1249.260 186.280 ;
        RECT 1250.840 186.020 1251.100 186.280 ;
        RECT 1249.460 138.080 1249.720 138.340 ;
        RECT 1250.840 138.080 1251.100 138.340 ;
        RECT 1249.460 110.200 1249.720 110.460 ;
        RECT 1250.380 110.200 1250.640 110.460 ;
        RECT 1132.620 18.400 1132.880 18.660 ;
        RECT 1250.380 17.720 1250.640 17.980 ;
      LAYER met2 ;
        RECT 1252.910 600.170 1253.190 604.000 ;
        RECT 1251.820 600.030 1253.190 600.170 ;
        RECT 1251.820 572.890 1251.960 600.030 ;
        RECT 1252.910 600.000 1253.190 600.030 ;
        RECT 1250.380 572.570 1250.640 572.890 ;
        RECT 1251.760 572.570 1252.020 572.890 ;
        RECT 1250.440 545.090 1250.580 572.570 ;
        RECT 1249.980 544.950 1250.580 545.090 ;
        RECT 1249.980 531.320 1250.120 544.950 ;
        RECT 1249.520 531.180 1250.120 531.320 ;
        RECT 1249.520 497.070 1249.660 531.180 ;
        RECT 1249.460 496.750 1249.720 497.070 ;
        RECT 1249.920 496.410 1250.180 496.730 ;
        RECT 1249.980 483.210 1250.120 496.410 ;
        RECT 1249.520 483.070 1250.120 483.210 ;
        RECT 1249.520 400.850 1249.660 483.070 ;
        RECT 1249.460 400.530 1249.720 400.850 ;
        RECT 1249.000 400.190 1249.260 400.510 ;
        RECT 1249.060 379.430 1249.200 400.190 ;
        RECT 1249.000 379.110 1249.260 379.430 ;
        RECT 1249.460 379.110 1249.720 379.430 ;
        RECT 1249.520 352.230 1249.660 379.110 ;
        RECT 1249.460 351.910 1249.720 352.230 ;
        RECT 1249.920 351.570 1250.180 351.890 ;
        RECT 1249.980 331.570 1250.120 351.570 ;
        RECT 1249.520 331.430 1250.120 331.570 ;
        RECT 1249.520 331.150 1249.660 331.430 ;
        RECT 1249.460 330.830 1249.720 331.150 ;
        RECT 1250.840 330.490 1251.100 330.810 ;
        RECT 1250.900 283.210 1251.040 330.490 ;
        RECT 1250.380 282.890 1250.640 283.210 ;
        RECT 1250.840 282.890 1251.100 283.210 ;
        RECT 1250.440 193.450 1250.580 282.890 ;
        RECT 1249.000 193.130 1249.260 193.450 ;
        RECT 1250.380 193.130 1250.640 193.450 ;
        RECT 1249.060 186.310 1249.200 193.130 ;
        RECT 1249.000 185.990 1249.260 186.310 ;
        RECT 1250.840 185.990 1251.100 186.310 ;
        RECT 1250.900 138.370 1251.040 185.990 ;
        RECT 1249.460 138.050 1249.720 138.370 ;
        RECT 1250.840 138.050 1251.100 138.370 ;
        RECT 1249.520 110.490 1249.660 138.050 ;
        RECT 1249.460 110.170 1249.720 110.490 ;
        RECT 1250.380 110.170 1250.640 110.490 ;
        RECT 1132.620 18.370 1132.880 18.690 ;
        RECT 1132.680 2.400 1132.820 18.370 ;
        RECT 1250.440 18.010 1250.580 110.170 ;
        RECT 1250.380 17.690 1250.640 18.010 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1256.330 531.320 1256.650 531.380 ;
        RECT 1257.250 531.320 1257.570 531.380 ;
        RECT 1256.330 531.180 1257.570 531.320 ;
        RECT 1256.330 531.120 1256.650 531.180 ;
        RECT 1257.250 531.120 1257.570 531.180 ;
        RECT 1256.330 483.380 1256.650 483.440 ;
        RECT 1257.250 483.380 1257.570 483.440 ;
        RECT 1256.330 483.240 1257.570 483.380 ;
        RECT 1256.330 483.180 1256.650 483.240 ;
        RECT 1257.250 483.180 1257.570 483.240 ;
        RECT 1256.330 448.160 1256.650 448.420 ;
        RECT 1256.420 448.020 1256.560 448.160 ;
        RECT 1256.790 448.020 1257.110 448.080 ;
        RECT 1256.420 447.880 1257.110 448.020 ;
        RECT 1256.790 447.820 1257.110 447.880 ;
        RECT 1256.330 331.400 1256.650 331.460 ;
        RECT 1256.790 331.400 1257.110 331.460 ;
        RECT 1256.330 331.260 1257.110 331.400 ;
        RECT 1256.330 331.200 1256.650 331.260 ;
        RECT 1256.790 331.200 1257.110 331.260 ;
        RECT 1255.870 193.020 1256.190 193.080 ;
        RECT 1256.790 193.020 1257.110 193.080 ;
        RECT 1255.870 192.880 1257.110 193.020 ;
        RECT 1255.870 192.820 1256.190 192.880 ;
        RECT 1256.790 192.820 1257.110 192.880 ;
        RECT 1255.870 159.020 1256.190 159.080 ;
        RECT 1255.870 158.880 1256.560 159.020 ;
        RECT 1255.870 158.820 1256.190 158.880 ;
        RECT 1256.420 158.740 1256.560 158.880 ;
        RECT 1256.330 158.480 1256.650 158.740 ;
        RECT 1150.530 18.600 1150.850 18.660 ;
        RECT 1255.870 18.600 1256.190 18.660 ;
        RECT 1150.530 18.460 1256.190 18.600 ;
        RECT 1150.530 18.400 1150.850 18.460 ;
        RECT 1255.870 18.400 1256.190 18.460 ;
      LAYER via ;
        RECT 1256.360 531.120 1256.620 531.380 ;
        RECT 1257.280 531.120 1257.540 531.380 ;
        RECT 1256.360 483.180 1256.620 483.440 ;
        RECT 1257.280 483.180 1257.540 483.440 ;
        RECT 1256.360 448.160 1256.620 448.420 ;
        RECT 1256.820 447.820 1257.080 448.080 ;
        RECT 1256.360 331.200 1256.620 331.460 ;
        RECT 1256.820 331.200 1257.080 331.460 ;
        RECT 1255.900 192.820 1256.160 193.080 ;
        RECT 1256.820 192.820 1257.080 193.080 ;
        RECT 1255.900 158.820 1256.160 159.080 ;
        RECT 1256.360 158.480 1256.620 158.740 ;
        RECT 1150.560 18.400 1150.820 18.660 ;
        RECT 1255.900 18.400 1256.160 18.660 ;
      LAYER met2 ;
        RECT 1262.110 600.170 1262.390 604.000 ;
        RECT 1259.640 600.030 1262.390 600.170 ;
        RECT 1259.640 596.770 1259.780 600.030 ;
        RECT 1262.110 600.000 1262.390 600.030 ;
        RECT 1257.800 596.630 1259.780 596.770 ;
        RECT 1257.800 569.570 1257.940 596.630 ;
        RECT 1256.880 569.430 1257.940 569.570 ;
        RECT 1256.880 545.090 1257.020 569.430 ;
        RECT 1256.420 544.950 1257.020 545.090 ;
        RECT 1256.420 531.410 1256.560 544.950 ;
        RECT 1256.360 531.090 1256.620 531.410 ;
        RECT 1257.280 531.090 1257.540 531.410 ;
        RECT 1257.340 483.470 1257.480 531.090 ;
        RECT 1256.360 483.150 1256.620 483.470 ;
        RECT 1257.280 483.150 1257.540 483.470 ;
        RECT 1256.420 448.450 1256.560 483.150 ;
        RECT 1256.360 448.130 1256.620 448.450 ;
        RECT 1256.820 447.790 1257.080 448.110 ;
        RECT 1256.880 331.490 1257.020 447.790 ;
        RECT 1256.360 331.170 1256.620 331.490 ;
        RECT 1256.820 331.170 1257.080 331.490 ;
        RECT 1256.420 303.690 1256.560 331.170 ;
        RECT 1256.420 303.550 1257.020 303.690 ;
        RECT 1256.880 193.110 1257.020 303.550 ;
        RECT 1255.900 192.790 1256.160 193.110 ;
        RECT 1256.820 192.790 1257.080 193.110 ;
        RECT 1255.960 159.110 1256.100 192.790 ;
        RECT 1255.900 158.790 1256.160 159.110 ;
        RECT 1256.360 158.450 1256.620 158.770 ;
        RECT 1256.420 110.570 1256.560 158.450 ;
        RECT 1256.420 110.430 1257.020 110.570 ;
        RECT 1256.880 62.290 1257.020 110.430 ;
        RECT 1255.960 62.150 1257.020 62.290 ;
        RECT 1255.960 18.690 1256.100 62.150 ;
        RECT 1150.560 18.370 1150.820 18.690 ;
        RECT 1255.900 18.370 1256.160 18.690 ;
        RECT 1150.620 2.400 1150.760 18.370 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 36.280 669.230 36.340 ;
        RECT 1014.370 36.280 1014.690 36.340 ;
        RECT 668.910 36.140 1014.690 36.280 ;
        RECT 668.910 36.080 669.230 36.140 ;
        RECT 1014.370 36.080 1014.690 36.140 ;
      LAYER via ;
        RECT 668.940 36.080 669.200 36.340 ;
        RECT 1014.400 36.080 1014.660 36.340 ;
      LAYER met2 ;
        RECT 1014.170 600.000 1014.450 604.000 ;
        RECT 1014.230 598.810 1014.370 600.000 ;
        RECT 1014.230 598.670 1014.600 598.810 ;
        RECT 1014.460 36.370 1014.600 598.670 ;
        RECT 668.940 36.050 669.200 36.370 ;
        RECT 1014.400 36.050 1014.660 36.370 ;
        RECT 669.000 2.400 669.140 36.050 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1172.610 590.820 1172.930 590.880 ;
        RECT 1269.670 590.820 1269.990 590.880 ;
        RECT 1172.610 590.680 1269.990 590.820 ;
        RECT 1172.610 590.620 1172.930 590.680 ;
        RECT 1269.670 590.620 1269.990 590.680 ;
        RECT 1168.470 20.640 1168.790 20.700 ;
        RECT 1172.610 20.640 1172.930 20.700 ;
        RECT 1168.470 20.500 1172.930 20.640 ;
        RECT 1168.470 20.440 1168.790 20.500 ;
        RECT 1172.610 20.440 1172.930 20.500 ;
      LAYER via ;
        RECT 1172.640 590.620 1172.900 590.880 ;
        RECT 1269.700 590.620 1269.960 590.880 ;
        RECT 1168.500 20.440 1168.760 20.700 ;
        RECT 1172.640 20.440 1172.900 20.700 ;
      LAYER met2 ;
        RECT 1271.310 600.170 1271.590 604.000 ;
        RECT 1269.760 600.030 1271.590 600.170 ;
        RECT 1269.760 590.910 1269.900 600.030 ;
        RECT 1271.310 600.000 1271.590 600.030 ;
        RECT 1172.640 590.590 1172.900 590.910 ;
        RECT 1269.700 590.590 1269.960 590.910 ;
        RECT 1172.700 20.730 1172.840 590.590 ;
        RECT 1168.500 20.410 1168.760 20.730 ;
        RECT 1172.640 20.410 1172.900 20.730 ;
        RECT 1168.560 2.400 1168.700 20.410 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1185.950 591.500 1186.270 591.560 ;
        RECT 1278.870 591.500 1279.190 591.560 ;
        RECT 1185.950 591.360 1279.190 591.500 ;
        RECT 1185.950 591.300 1186.270 591.360 ;
        RECT 1278.870 591.300 1279.190 591.360 ;
      LAYER via ;
        RECT 1185.980 591.300 1186.240 591.560 ;
        RECT 1278.900 591.300 1279.160 591.560 ;
      LAYER met2 ;
        RECT 1280.510 600.170 1280.790 604.000 ;
        RECT 1278.960 600.030 1280.790 600.170 ;
        RECT 1278.960 591.590 1279.100 600.030 ;
        RECT 1280.510 600.000 1280.790 600.030 ;
        RECT 1185.980 591.270 1186.240 591.590 ;
        RECT 1278.900 591.270 1279.160 591.590 ;
        RECT 1186.040 2.400 1186.180 591.270 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.110 589.460 1207.430 589.520 ;
        RECT 1288.070 589.460 1288.390 589.520 ;
        RECT 1207.110 589.320 1288.390 589.460 ;
        RECT 1207.110 589.260 1207.430 589.320 ;
        RECT 1288.070 589.260 1288.390 589.320 ;
        RECT 1203.890 20.640 1204.210 20.700 ;
        RECT 1207.110 20.640 1207.430 20.700 ;
        RECT 1203.890 20.500 1207.430 20.640 ;
        RECT 1203.890 20.440 1204.210 20.500 ;
        RECT 1207.110 20.440 1207.430 20.500 ;
      LAYER via ;
        RECT 1207.140 589.260 1207.400 589.520 ;
        RECT 1288.100 589.260 1288.360 589.520 ;
        RECT 1203.920 20.440 1204.180 20.700 ;
        RECT 1207.140 20.440 1207.400 20.700 ;
      LAYER met2 ;
        RECT 1289.710 600.170 1289.990 604.000 ;
        RECT 1288.160 600.030 1289.990 600.170 ;
        RECT 1288.160 589.550 1288.300 600.030 ;
        RECT 1289.710 600.000 1289.990 600.030 ;
        RECT 1207.140 589.230 1207.400 589.550 ;
        RECT 1288.100 589.230 1288.360 589.550 ;
        RECT 1207.200 20.730 1207.340 589.230 ;
        RECT 1203.920 20.410 1204.180 20.730 ;
        RECT 1207.140 20.410 1207.400 20.730 ;
        RECT 1203.980 2.400 1204.120 20.410 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1227.810 588.440 1228.130 588.500 ;
        RECT 1297.270 588.440 1297.590 588.500 ;
        RECT 1227.810 588.300 1297.590 588.440 ;
        RECT 1227.810 588.240 1228.130 588.300 ;
        RECT 1297.270 588.240 1297.590 588.300 ;
        RECT 1221.830 20.640 1222.150 20.700 ;
        RECT 1227.810 20.640 1228.130 20.700 ;
        RECT 1221.830 20.500 1228.130 20.640 ;
        RECT 1221.830 20.440 1222.150 20.500 ;
        RECT 1227.810 20.440 1228.130 20.500 ;
      LAYER via ;
        RECT 1227.840 588.240 1228.100 588.500 ;
        RECT 1297.300 588.240 1297.560 588.500 ;
        RECT 1221.860 20.440 1222.120 20.700 ;
        RECT 1227.840 20.440 1228.100 20.700 ;
      LAYER met2 ;
        RECT 1298.910 600.170 1299.190 604.000 ;
        RECT 1297.360 600.030 1299.190 600.170 ;
        RECT 1297.360 588.530 1297.500 600.030 ;
        RECT 1298.910 600.000 1299.190 600.030 ;
        RECT 1227.840 588.210 1228.100 588.530 ;
        RECT 1297.300 588.210 1297.560 588.530 ;
        RECT 1227.900 20.730 1228.040 588.210 ;
        RECT 1221.860 20.410 1222.120 20.730 ;
        RECT 1227.840 20.410 1228.100 20.730 ;
        RECT 1221.920 2.400 1222.060 20.410 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.610 587.760 1241.930 587.820 ;
        RECT 1306.470 587.760 1306.790 587.820 ;
        RECT 1241.610 587.620 1306.790 587.760 ;
        RECT 1241.610 587.560 1241.930 587.620 ;
        RECT 1306.470 587.560 1306.790 587.620 ;
        RECT 1241.150 579.600 1241.470 579.660 ;
        RECT 1241.610 579.600 1241.930 579.660 ;
        RECT 1241.150 579.460 1241.930 579.600 ;
        RECT 1241.150 579.400 1241.470 579.460 ;
        RECT 1241.610 579.400 1241.930 579.460 ;
        RECT 1241.150 531.660 1241.470 531.720 ;
        RECT 1241.610 531.660 1241.930 531.720 ;
        RECT 1241.150 531.520 1241.930 531.660 ;
        RECT 1241.150 531.460 1241.470 531.520 ;
        RECT 1241.610 531.460 1241.930 531.520 ;
        RECT 1239.770 90.000 1240.090 90.060 ;
        RECT 1241.610 90.000 1241.930 90.060 ;
        RECT 1239.770 89.860 1241.930 90.000 ;
        RECT 1239.770 89.800 1240.090 89.860 ;
        RECT 1241.610 89.800 1241.930 89.860 ;
        RECT 1239.770 47.980 1240.090 48.240 ;
        RECT 1239.860 47.560 1240.000 47.980 ;
        RECT 1239.770 47.300 1240.090 47.560 ;
      LAYER via ;
        RECT 1241.640 587.560 1241.900 587.820 ;
        RECT 1306.500 587.560 1306.760 587.820 ;
        RECT 1241.180 579.400 1241.440 579.660 ;
        RECT 1241.640 579.400 1241.900 579.660 ;
        RECT 1241.180 531.460 1241.440 531.720 ;
        RECT 1241.640 531.460 1241.900 531.720 ;
        RECT 1239.800 89.800 1240.060 90.060 ;
        RECT 1241.640 89.800 1241.900 90.060 ;
        RECT 1239.800 47.980 1240.060 48.240 ;
        RECT 1239.800 47.300 1240.060 47.560 ;
      LAYER met2 ;
        RECT 1308.110 600.170 1308.390 604.000 ;
        RECT 1306.560 600.030 1308.390 600.170 ;
        RECT 1306.560 587.850 1306.700 600.030 ;
        RECT 1308.110 600.000 1308.390 600.030 ;
        RECT 1241.640 587.530 1241.900 587.850 ;
        RECT 1306.500 587.530 1306.760 587.850 ;
        RECT 1241.700 579.690 1241.840 587.530 ;
        RECT 1241.180 579.370 1241.440 579.690 ;
        RECT 1241.640 579.370 1241.900 579.690 ;
        RECT 1241.240 531.750 1241.380 579.370 ;
        RECT 1241.180 531.430 1241.440 531.750 ;
        RECT 1241.640 531.430 1241.900 531.750 ;
        RECT 1241.700 90.090 1241.840 531.430 ;
        RECT 1239.800 89.770 1240.060 90.090 ;
        RECT 1241.640 89.770 1241.900 90.090 ;
        RECT 1239.860 48.270 1240.000 89.770 ;
        RECT 1239.800 47.950 1240.060 48.270 ;
        RECT 1239.800 47.270 1240.060 47.590 ;
        RECT 1239.860 2.400 1240.000 47.270 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.350 588.100 1296.670 588.160 ;
        RECT 1315.670 588.100 1315.990 588.160 ;
        RECT 1296.350 587.960 1315.990 588.100 ;
        RECT 1296.350 587.900 1296.670 587.960 ;
        RECT 1315.670 587.900 1315.990 587.960 ;
        RECT 1262.310 586.740 1262.630 586.800 ;
        RECT 1296.350 586.740 1296.670 586.800 ;
        RECT 1262.310 586.600 1296.670 586.740 ;
        RECT 1262.310 586.540 1262.630 586.600 ;
        RECT 1296.350 586.540 1296.670 586.600 ;
        RECT 1257.250 20.640 1257.570 20.700 ;
        RECT 1262.310 20.640 1262.630 20.700 ;
        RECT 1257.250 20.500 1262.630 20.640 ;
        RECT 1257.250 20.440 1257.570 20.500 ;
        RECT 1262.310 20.440 1262.630 20.500 ;
      LAYER via ;
        RECT 1296.380 587.900 1296.640 588.160 ;
        RECT 1315.700 587.900 1315.960 588.160 ;
        RECT 1262.340 586.540 1262.600 586.800 ;
        RECT 1296.380 586.540 1296.640 586.800 ;
        RECT 1257.280 20.440 1257.540 20.700 ;
        RECT 1262.340 20.440 1262.600 20.700 ;
      LAYER met2 ;
        RECT 1317.310 600.170 1317.590 604.000 ;
        RECT 1315.760 600.030 1317.590 600.170 ;
        RECT 1315.760 588.190 1315.900 600.030 ;
        RECT 1317.310 600.000 1317.590 600.030 ;
        RECT 1296.380 587.870 1296.640 588.190 ;
        RECT 1315.700 587.870 1315.960 588.190 ;
        RECT 1296.440 586.830 1296.580 587.870 ;
        RECT 1262.340 586.510 1262.600 586.830 ;
        RECT 1296.380 586.510 1296.640 586.830 ;
        RECT 1262.400 20.730 1262.540 586.510 ;
        RECT 1257.280 20.410 1257.540 20.730 ;
        RECT 1262.340 20.410 1262.600 20.730 ;
        RECT 1257.340 2.400 1257.480 20.410 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.110 590.480 1276.430 590.540 ;
        RECT 1324.870 590.480 1325.190 590.540 ;
        RECT 1276.110 590.340 1325.190 590.480 ;
        RECT 1276.110 590.280 1276.430 590.340 ;
        RECT 1324.870 590.280 1325.190 590.340 ;
      LAYER via ;
        RECT 1276.140 590.280 1276.400 590.540 ;
        RECT 1324.900 590.280 1325.160 590.540 ;
      LAYER met2 ;
        RECT 1326.510 600.170 1326.790 604.000 ;
        RECT 1324.960 600.030 1326.790 600.170 ;
        RECT 1324.960 590.570 1325.100 600.030 ;
        RECT 1326.510 600.000 1326.790 600.030 ;
        RECT 1276.140 590.250 1276.400 590.570 ;
        RECT 1324.900 590.250 1325.160 590.570 ;
        RECT 1276.200 16.730 1276.340 590.250 ;
        RECT 1275.280 16.590 1276.340 16.730 ;
        RECT 1275.280 2.400 1275.420 16.590 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 586.740 1297.130 586.800 ;
        RECT 1334.070 586.740 1334.390 586.800 ;
        RECT 1296.810 586.600 1334.390 586.740 ;
        RECT 1296.810 586.540 1297.130 586.600 ;
        RECT 1334.070 586.540 1334.390 586.600 ;
        RECT 1293.130 15.540 1293.450 15.600 ;
        RECT 1296.810 15.540 1297.130 15.600 ;
        RECT 1293.130 15.400 1297.130 15.540 ;
        RECT 1293.130 15.340 1293.450 15.400 ;
        RECT 1296.810 15.340 1297.130 15.400 ;
      LAYER via ;
        RECT 1296.840 586.540 1297.100 586.800 ;
        RECT 1334.100 586.540 1334.360 586.800 ;
        RECT 1293.160 15.340 1293.420 15.600 ;
        RECT 1296.840 15.340 1297.100 15.600 ;
      LAYER met2 ;
        RECT 1335.710 600.170 1335.990 604.000 ;
        RECT 1334.160 600.030 1335.990 600.170 ;
        RECT 1334.160 586.830 1334.300 600.030 ;
        RECT 1335.710 600.000 1335.990 600.030 ;
        RECT 1296.840 586.510 1297.100 586.830 ;
        RECT 1334.100 586.510 1334.360 586.830 ;
        RECT 1296.900 15.630 1297.040 586.510 ;
        RECT 1293.160 15.310 1293.420 15.630 ;
        RECT 1296.840 15.310 1297.100 15.630 ;
        RECT 1293.220 2.400 1293.360 15.310 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1317.510 589.460 1317.830 589.520 ;
        RECT 1343.270 589.460 1343.590 589.520 ;
        RECT 1317.510 589.320 1343.590 589.460 ;
        RECT 1317.510 589.260 1317.830 589.320 ;
        RECT 1343.270 589.260 1343.590 589.320 ;
        RECT 1311.070 17.580 1311.390 17.640 ;
        RECT 1317.510 17.580 1317.830 17.640 ;
        RECT 1311.070 17.440 1317.830 17.580 ;
        RECT 1311.070 17.380 1311.390 17.440 ;
        RECT 1317.510 17.380 1317.830 17.440 ;
      LAYER via ;
        RECT 1317.540 589.260 1317.800 589.520 ;
        RECT 1343.300 589.260 1343.560 589.520 ;
        RECT 1311.100 17.380 1311.360 17.640 ;
        RECT 1317.540 17.380 1317.800 17.640 ;
      LAYER met2 ;
        RECT 1344.910 600.170 1345.190 604.000 ;
        RECT 1343.360 600.030 1345.190 600.170 ;
        RECT 1343.360 589.550 1343.500 600.030 ;
        RECT 1344.910 600.000 1345.190 600.030 ;
        RECT 1317.540 589.230 1317.800 589.550 ;
        RECT 1343.300 589.230 1343.560 589.550 ;
        RECT 1317.600 17.670 1317.740 589.230 ;
        RECT 1311.100 17.350 1311.360 17.670 ;
        RECT 1317.540 17.350 1317.800 17.670 ;
        RECT 1311.160 2.400 1311.300 17.350 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.310 590.140 1331.630 590.200 ;
        RECT 1352.470 590.140 1352.790 590.200 ;
        RECT 1331.310 590.000 1352.790 590.140 ;
        RECT 1331.310 589.940 1331.630 590.000 ;
        RECT 1352.470 589.940 1352.790 590.000 ;
        RECT 1329.010 17.580 1329.330 17.640 ;
        RECT 1331.310 17.580 1331.630 17.640 ;
        RECT 1329.010 17.440 1331.630 17.580 ;
        RECT 1329.010 17.380 1329.330 17.440 ;
        RECT 1331.310 17.380 1331.630 17.440 ;
      LAYER via ;
        RECT 1331.340 589.940 1331.600 590.200 ;
        RECT 1352.500 589.940 1352.760 590.200 ;
        RECT 1329.040 17.380 1329.300 17.640 ;
        RECT 1331.340 17.380 1331.600 17.640 ;
      LAYER met2 ;
        RECT 1354.110 600.170 1354.390 604.000 ;
        RECT 1352.560 600.030 1354.390 600.170 ;
        RECT 1352.560 590.230 1352.700 600.030 ;
        RECT 1354.110 600.000 1354.390 600.030 ;
        RECT 1331.340 589.910 1331.600 590.230 ;
        RECT 1352.500 589.910 1352.760 590.230 ;
        RECT 1331.400 17.670 1331.540 589.910 ;
        RECT 1329.040 17.350 1329.300 17.670 ;
        RECT 1331.340 17.350 1331.600 17.670 ;
        RECT 1329.100 2.400 1329.240 17.350 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 37.980 686.710 38.040 ;
        RECT 1021.270 37.980 1021.590 38.040 ;
        RECT 686.390 37.840 1021.590 37.980 ;
        RECT 686.390 37.780 686.710 37.840 ;
        RECT 1021.270 37.780 1021.590 37.840 ;
      LAYER via ;
        RECT 686.420 37.780 686.680 38.040 ;
        RECT 1021.300 37.780 1021.560 38.040 ;
      LAYER met2 ;
        RECT 1023.370 600.170 1023.650 604.000 ;
        RECT 1021.360 600.030 1023.650 600.170 ;
        RECT 1021.360 38.070 1021.500 600.030 ;
        RECT 1023.370 600.000 1023.650 600.030 ;
        RECT 686.420 37.750 686.680 38.070 ;
        RECT 1021.300 37.750 1021.560 38.070 ;
        RECT 686.480 2.400 686.620 37.750 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1355.690 586.740 1356.010 586.800 ;
        RECT 1361.670 586.740 1361.990 586.800 ;
        RECT 1355.690 586.600 1361.990 586.740 ;
        RECT 1355.690 586.540 1356.010 586.600 ;
        RECT 1361.670 586.540 1361.990 586.600 ;
        RECT 1346.490 15.200 1346.810 15.260 ;
        RECT 1355.690 15.200 1356.010 15.260 ;
        RECT 1346.490 15.060 1356.010 15.200 ;
        RECT 1346.490 15.000 1346.810 15.060 ;
        RECT 1355.690 15.000 1356.010 15.060 ;
      LAYER via ;
        RECT 1355.720 586.540 1355.980 586.800 ;
        RECT 1361.700 586.540 1361.960 586.800 ;
        RECT 1346.520 15.000 1346.780 15.260 ;
        RECT 1355.720 15.000 1355.980 15.260 ;
      LAYER met2 ;
        RECT 1363.310 600.170 1363.590 604.000 ;
        RECT 1361.760 600.030 1363.590 600.170 ;
        RECT 1361.760 586.830 1361.900 600.030 ;
        RECT 1363.310 600.000 1363.590 600.030 ;
        RECT 1355.720 586.510 1355.980 586.830 ;
        RECT 1361.700 586.510 1361.960 586.830 ;
        RECT 1355.780 15.290 1355.920 586.510 ;
        RECT 1346.520 14.970 1346.780 15.290 ;
        RECT 1355.720 14.970 1355.980 15.290 ;
        RECT 1346.580 2.400 1346.720 14.970 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 586.740 1366.130 586.800 ;
        RECT 1370.870 586.740 1371.190 586.800 ;
        RECT 1365.810 586.600 1371.190 586.740 ;
        RECT 1365.810 586.540 1366.130 586.600 ;
        RECT 1370.870 586.540 1371.190 586.600 ;
      LAYER via ;
        RECT 1365.840 586.540 1366.100 586.800 ;
        RECT 1370.900 586.540 1371.160 586.800 ;
      LAYER met2 ;
        RECT 1372.510 600.170 1372.790 604.000 ;
        RECT 1370.960 600.030 1372.790 600.170 ;
        RECT 1370.960 586.830 1371.100 600.030 ;
        RECT 1372.510 600.000 1372.790 600.030 ;
        RECT 1365.840 586.510 1366.100 586.830 ;
        RECT 1370.900 586.510 1371.160 586.830 ;
        RECT 1365.900 17.410 1366.040 586.510 ;
        RECT 1364.520 17.270 1366.040 17.410 ;
        RECT 1364.520 2.400 1364.660 17.270 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.530 572.800 1380.850 572.860 ;
        RECT 1380.990 572.800 1381.310 572.860 ;
        RECT 1380.530 572.660 1381.310 572.800 ;
        RECT 1380.530 572.600 1380.850 572.660 ;
        RECT 1380.990 572.600 1381.310 572.660 ;
        RECT 1379.610 524.180 1379.930 524.240 ;
        RECT 1380.530 524.180 1380.850 524.240 ;
        RECT 1379.610 524.040 1380.850 524.180 ;
        RECT 1379.610 523.980 1379.930 524.040 ;
        RECT 1380.530 523.980 1380.850 524.040 ;
        RECT 1379.610 476.240 1379.930 476.300 ;
        RECT 1380.070 476.240 1380.390 476.300 ;
        RECT 1379.610 476.100 1380.390 476.240 ;
        RECT 1379.610 476.040 1379.930 476.100 ;
        RECT 1380.070 476.040 1380.390 476.100 ;
        RECT 1380.070 475.560 1380.390 475.620 ;
        RECT 1381.450 475.560 1381.770 475.620 ;
        RECT 1380.070 475.420 1381.770 475.560 ;
        RECT 1380.070 475.360 1380.390 475.420 ;
        RECT 1381.450 475.360 1381.770 475.420 ;
        RECT 1380.530 427.620 1380.850 427.680 ;
        RECT 1380.990 427.620 1381.310 427.680 ;
        RECT 1380.530 427.480 1381.310 427.620 ;
        RECT 1380.530 427.420 1380.850 427.480 ;
        RECT 1380.990 427.420 1381.310 427.480 ;
        RECT 1380.070 420.820 1380.390 420.880 ;
        RECT 1380.990 420.820 1381.310 420.880 ;
        RECT 1380.070 420.680 1381.310 420.820 ;
        RECT 1380.070 420.620 1380.390 420.680 ;
        RECT 1380.990 420.620 1381.310 420.680 ;
        RECT 1379.610 372.880 1379.930 372.940 ;
        RECT 1380.070 372.880 1380.390 372.940 ;
        RECT 1379.610 372.740 1380.390 372.880 ;
        RECT 1379.610 372.680 1379.930 372.740 ;
        RECT 1380.070 372.680 1380.390 372.740 ;
        RECT 1380.530 289.580 1380.850 289.640 ;
        RECT 1380.990 289.580 1381.310 289.640 ;
        RECT 1380.530 289.440 1381.310 289.580 ;
        RECT 1380.530 289.380 1380.850 289.440 ;
        RECT 1380.990 289.380 1381.310 289.440 ;
        RECT 1380.530 241.980 1380.850 242.040 ;
        RECT 1380.990 241.980 1381.310 242.040 ;
        RECT 1380.530 241.840 1381.310 241.980 ;
        RECT 1380.530 241.780 1380.850 241.840 ;
        RECT 1380.990 241.780 1381.310 241.840 ;
        RECT 1380.530 234.500 1380.850 234.560 ;
        RECT 1380.990 234.500 1381.310 234.560 ;
        RECT 1380.530 234.360 1381.310 234.500 ;
        RECT 1380.530 234.300 1380.850 234.360 ;
        RECT 1380.990 234.300 1381.310 234.360 ;
        RECT 1380.530 145.420 1380.850 145.480 ;
        RECT 1380.990 145.420 1381.310 145.480 ;
        RECT 1380.530 145.280 1381.310 145.420 ;
        RECT 1380.530 145.220 1380.850 145.280 ;
        RECT 1380.990 145.220 1381.310 145.280 ;
        RECT 1379.610 137.940 1379.930 138.000 ;
        RECT 1380.530 137.940 1380.850 138.000 ;
        RECT 1379.610 137.800 1380.850 137.940 ;
        RECT 1379.610 137.740 1379.930 137.800 ;
        RECT 1380.530 137.740 1380.850 137.800 ;
        RECT 1379.610 90.000 1379.930 90.060 ;
        RECT 1380.530 90.000 1380.850 90.060 ;
        RECT 1379.610 89.860 1380.850 90.000 ;
        RECT 1379.610 89.800 1379.930 89.860 ;
        RECT 1380.530 89.800 1380.850 89.860 ;
        RECT 1380.530 62.260 1380.850 62.520 ;
        RECT 1380.620 61.780 1380.760 62.260 ;
        RECT 1382.370 61.780 1382.690 61.840 ;
        RECT 1380.620 61.640 1382.690 61.780 ;
        RECT 1382.370 61.580 1382.690 61.640 ;
      LAYER via ;
        RECT 1380.560 572.600 1380.820 572.860 ;
        RECT 1381.020 572.600 1381.280 572.860 ;
        RECT 1379.640 523.980 1379.900 524.240 ;
        RECT 1380.560 523.980 1380.820 524.240 ;
        RECT 1379.640 476.040 1379.900 476.300 ;
        RECT 1380.100 476.040 1380.360 476.300 ;
        RECT 1380.100 475.360 1380.360 475.620 ;
        RECT 1381.480 475.360 1381.740 475.620 ;
        RECT 1380.560 427.420 1380.820 427.680 ;
        RECT 1381.020 427.420 1381.280 427.680 ;
        RECT 1380.100 420.620 1380.360 420.880 ;
        RECT 1381.020 420.620 1381.280 420.880 ;
        RECT 1379.640 372.680 1379.900 372.940 ;
        RECT 1380.100 372.680 1380.360 372.940 ;
        RECT 1380.560 289.380 1380.820 289.640 ;
        RECT 1381.020 289.380 1381.280 289.640 ;
        RECT 1380.560 241.780 1380.820 242.040 ;
        RECT 1381.020 241.780 1381.280 242.040 ;
        RECT 1380.560 234.300 1380.820 234.560 ;
        RECT 1381.020 234.300 1381.280 234.560 ;
        RECT 1380.560 145.220 1380.820 145.480 ;
        RECT 1381.020 145.220 1381.280 145.480 ;
        RECT 1379.640 137.740 1379.900 138.000 ;
        RECT 1380.560 137.740 1380.820 138.000 ;
        RECT 1379.640 89.800 1379.900 90.060 ;
        RECT 1380.560 89.800 1380.820 90.060 ;
        RECT 1380.560 62.260 1380.820 62.520 ;
        RECT 1382.400 61.580 1382.660 61.840 ;
      LAYER met2 ;
        RECT 1381.250 600.000 1381.530 604.000 ;
        RECT 1381.310 598.810 1381.450 600.000 ;
        RECT 1381.080 598.670 1381.450 598.810 ;
        RECT 1381.080 572.890 1381.220 598.670 ;
        RECT 1380.560 572.570 1380.820 572.890 ;
        RECT 1381.020 572.570 1381.280 572.890 ;
        RECT 1380.620 524.270 1380.760 572.570 ;
        RECT 1379.640 523.950 1379.900 524.270 ;
        RECT 1380.560 523.950 1380.820 524.270 ;
        RECT 1379.700 476.330 1379.840 523.950 ;
        RECT 1379.640 476.010 1379.900 476.330 ;
        RECT 1380.100 476.010 1380.360 476.330 ;
        RECT 1380.160 475.650 1380.300 476.010 ;
        RECT 1380.100 475.330 1380.360 475.650 ;
        RECT 1381.480 475.330 1381.740 475.650 ;
        RECT 1381.540 428.245 1381.680 475.330 ;
        RECT 1380.550 427.875 1380.830 428.245 ;
        RECT 1381.470 427.875 1381.750 428.245 ;
        RECT 1380.620 427.710 1380.760 427.875 ;
        RECT 1380.560 427.390 1380.820 427.710 ;
        RECT 1381.020 427.390 1381.280 427.710 ;
        RECT 1381.080 420.910 1381.220 427.390 ;
        RECT 1380.100 420.590 1380.360 420.910 ;
        RECT 1381.020 420.590 1381.280 420.910 ;
        RECT 1380.160 372.970 1380.300 420.590 ;
        RECT 1379.640 372.650 1379.900 372.970 ;
        RECT 1380.100 372.650 1380.360 372.970 ;
        RECT 1379.700 337.010 1379.840 372.650 ;
        RECT 1379.700 336.870 1380.760 337.010 ;
        RECT 1380.620 289.670 1380.760 336.870 ;
        RECT 1380.560 289.350 1380.820 289.670 ;
        RECT 1381.020 289.350 1381.280 289.670 ;
        RECT 1381.080 242.070 1381.220 289.350 ;
        RECT 1380.560 241.750 1380.820 242.070 ;
        RECT 1381.020 241.750 1381.280 242.070 ;
        RECT 1380.620 234.590 1380.760 241.750 ;
        RECT 1380.560 234.270 1380.820 234.590 ;
        RECT 1381.020 234.270 1381.280 234.590 ;
        RECT 1381.080 145.510 1381.220 234.270 ;
        RECT 1380.560 145.190 1380.820 145.510 ;
        RECT 1381.020 145.190 1381.280 145.510 ;
        RECT 1380.620 138.030 1380.760 145.190 ;
        RECT 1379.640 137.710 1379.900 138.030 ;
        RECT 1380.560 137.710 1380.820 138.030 ;
        RECT 1379.700 90.090 1379.840 137.710 ;
        RECT 1379.640 89.770 1379.900 90.090 ;
        RECT 1380.560 89.770 1380.820 90.090 ;
        RECT 1380.620 62.550 1380.760 89.770 ;
        RECT 1380.560 62.230 1380.820 62.550 ;
        RECT 1382.400 61.550 1382.660 61.870 ;
        RECT 1382.460 2.400 1382.600 61.550 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
      LAYER via2 ;
        RECT 1380.550 427.920 1380.830 428.200 ;
        RECT 1381.470 427.920 1381.750 428.200 ;
      LAYER met3 ;
        RECT 1380.525 428.210 1380.855 428.225 ;
        RECT 1381.445 428.210 1381.775 428.225 ;
        RECT 1380.525 427.910 1381.775 428.210 ;
        RECT 1380.525 427.895 1380.855 427.910 ;
        RECT 1381.445 427.895 1381.775 427.910 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1392.950 20.640 1393.270 20.700 ;
        RECT 1400.310 20.640 1400.630 20.700 ;
        RECT 1392.950 20.500 1400.630 20.640 ;
        RECT 1392.950 20.440 1393.270 20.500 ;
        RECT 1400.310 20.440 1400.630 20.500 ;
      LAYER via ;
        RECT 1392.980 20.440 1393.240 20.700 ;
        RECT 1400.340 20.440 1400.600 20.700 ;
      LAYER met2 ;
        RECT 1390.450 600.170 1390.730 604.000 ;
        RECT 1390.450 600.030 1393.180 600.170 ;
        RECT 1390.450 600.000 1390.730 600.030 ;
        RECT 1393.040 20.730 1393.180 600.030 ;
        RECT 1392.980 20.410 1393.240 20.730 ;
        RECT 1400.340 20.410 1400.600 20.730 ;
        RECT 1400.400 2.400 1400.540 20.410 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1398.930 17.920 1399.250 17.980 ;
        RECT 1418.250 17.920 1418.570 17.980 ;
        RECT 1398.930 17.780 1418.570 17.920 ;
        RECT 1398.930 17.720 1399.250 17.780 ;
        RECT 1418.250 17.720 1418.570 17.780 ;
      LAYER via ;
        RECT 1398.960 17.720 1399.220 17.980 ;
        RECT 1418.280 17.720 1418.540 17.980 ;
      LAYER met2 ;
        RECT 1399.650 600.000 1399.930 604.000 ;
        RECT 1399.710 598.810 1399.850 600.000 ;
        RECT 1399.710 598.670 1400.080 598.810 ;
        RECT 1399.940 56.850 1400.080 598.670 ;
        RECT 1399.020 56.710 1400.080 56.850 ;
        RECT 1399.020 18.010 1399.160 56.710 ;
        RECT 1398.960 17.690 1399.220 18.010 ;
        RECT 1418.280 17.690 1418.540 18.010 ;
        RECT 1418.340 2.400 1418.480 17.690 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1410.430 586.740 1410.750 586.800 ;
        RECT 1414.110 586.740 1414.430 586.800 ;
        RECT 1410.430 586.600 1414.430 586.740 ;
        RECT 1410.430 586.540 1410.750 586.600 ;
        RECT 1414.110 586.540 1414.430 586.600 ;
        RECT 1414.110 16.900 1414.430 16.960 ;
        RECT 1435.730 16.900 1436.050 16.960 ;
        RECT 1414.110 16.760 1436.050 16.900 ;
        RECT 1414.110 16.700 1414.430 16.760 ;
        RECT 1435.730 16.700 1436.050 16.760 ;
      LAYER via ;
        RECT 1410.460 586.540 1410.720 586.800 ;
        RECT 1414.140 586.540 1414.400 586.800 ;
        RECT 1414.140 16.700 1414.400 16.960 ;
        RECT 1435.760 16.700 1436.020 16.960 ;
      LAYER met2 ;
        RECT 1408.850 600.170 1409.130 604.000 ;
        RECT 1408.850 600.030 1410.660 600.170 ;
        RECT 1408.850 600.000 1409.130 600.030 ;
        RECT 1410.520 586.830 1410.660 600.030 ;
        RECT 1410.460 586.510 1410.720 586.830 ;
        RECT 1414.140 586.510 1414.400 586.830 ;
        RECT 1414.200 16.990 1414.340 586.510 ;
        RECT 1414.140 16.670 1414.400 16.990 ;
        RECT 1435.760 16.670 1436.020 16.990 ;
        RECT 1435.820 2.400 1435.960 16.670 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.010 18.260 1421.330 18.320 ;
        RECT 1453.670 18.260 1453.990 18.320 ;
        RECT 1421.010 18.120 1453.990 18.260 ;
        RECT 1421.010 18.060 1421.330 18.120 ;
        RECT 1453.670 18.060 1453.990 18.120 ;
      LAYER via ;
        RECT 1421.040 18.060 1421.300 18.320 ;
        RECT 1453.700 18.060 1453.960 18.320 ;
      LAYER met2 ;
        RECT 1418.050 600.170 1418.330 604.000 ;
        RECT 1418.050 600.030 1420.780 600.170 ;
        RECT 1418.050 600.000 1418.330 600.030 ;
        RECT 1420.640 583.170 1420.780 600.030 ;
        RECT 1420.640 583.030 1421.240 583.170 ;
        RECT 1421.100 18.350 1421.240 583.030 ;
        RECT 1421.040 18.030 1421.300 18.350 ;
        RECT 1453.700 18.030 1453.960 18.350 ;
        RECT 1453.760 2.400 1453.900 18.030 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1426.990 17.580 1427.310 17.640 ;
        RECT 1471.610 17.580 1471.930 17.640 ;
        RECT 1426.990 17.440 1471.930 17.580 ;
        RECT 1426.990 17.380 1427.310 17.440 ;
        RECT 1471.610 17.380 1471.930 17.440 ;
      LAYER via ;
        RECT 1427.020 17.380 1427.280 17.640 ;
        RECT 1471.640 17.380 1471.900 17.640 ;
      LAYER met2 ;
        RECT 1427.250 600.000 1427.530 604.000 ;
        RECT 1427.310 598.810 1427.450 600.000 ;
        RECT 1427.080 598.670 1427.450 598.810 ;
        RECT 1427.080 17.670 1427.220 598.670 ;
        RECT 1427.020 17.350 1427.280 17.670 ;
        RECT 1471.640 17.350 1471.900 17.670 ;
        RECT 1471.700 2.400 1471.840 17.350 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1438.030 586.740 1438.350 586.800 ;
        RECT 1441.710 586.740 1442.030 586.800 ;
        RECT 1438.030 586.600 1442.030 586.740 ;
        RECT 1438.030 586.540 1438.350 586.600 ;
        RECT 1441.710 586.540 1442.030 586.600 ;
        RECT 1441.710 16.560 1442.030 16.620 ;
        RECT 1489.550 16.560 1489.870 16.620 ;
        RECT 1441.710 16.420 1489.870 16.560 ;
        RECT 1441.710 16.360 1442.030 16.420 ;
        RECT 1489.550 16.360 1489.870 16.420 ;
      LAYER via ;
        RECT 1438.060 586.540 1438.320 586.800 ;
        RECT 1441.740 586.540 1442.000 586.800 ;
        RECT 1441.740 16.360 1442.000 16.620 ;
        RECT 1489.580 16.360 1489.840 16.620 ;
      LAYER met2 ;
        RECT 1436.450 600.170 1436.730 604.000 ;
        RECT 1436.450 600.030 1438.260 600.170 ;
        RECT 1436.450 600.000 1436.730 600.030 ;
        RECT 1438.120 586.830 1438.260 600.030 ;
        RECT 1438.060 586.510 1438.320 586.830 ;
        RECT 1441.740 586.510 1442.000 586.830 ;
        RECT 1441.800 16.650 1441.940 586.510 ;
        RECT 1441.740 16.330 1442.000 16.650 ;
        RECT 1489.580 16.330 1489.840 16.650 ;
        RECT 1489.640 2.400 1489.780 16.330 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1448.610 20.640 1448.930 20.700 ;
        RECT 1507.030 20.640 1507.350 20.700 ;
        RECT 1448.610 20.500 1507.350 20.640 ;
        RECT 1448.610 20.440 1448.930 20.500 ;
        RECT 1507.030 20.440 1507.350 20.500 ;
      LAYER via ;
        RECT 1448.640 20.440 1448.900 20.700 ;
        RECT 1507.060 20.440 1507.320 20.700 ;
      LAYER met2 ;
        RECT 1445.650 600.170 1445.930 604.000 ;
        RECT 1445.650 600.030 1448.380 600.170 ;
        RECT 1445.650 600.000 1445.930 600.030 ;
        RECT 1448.240 583.170 1448.380 600.030 ;
        RECT 1448.240 583.030 1448.840 583.170 ;
        RECT 1448.700 20.730 1448.840 583.030 ;
        RECT 1448.640 20.410 1448.900 20.730 ;
        RECT 1507.060 20.410 1507.320 20.730 ;
        RECT 1507.120 2.400 1507.260 20.410 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1028.170 583.000 1028.490 583.060 ;
        RECT 1030.930 583.000 1031.250 583.060 ;
        RECT 1028.170 582.860 1031.250 583.000 ;
        RECT 1028.170 582.800 1028.490 582.860 ;
        RECT 1030.930 582.800 1031.250 582.860 ;
        RECT 704.330 38.660 704.650 38.720 ;
        RECT 1028.170 38.660 1028.490 38.720 ;
        RECT 704.330 38.520 1028.490 38.660 ;
        RECT 704.330 38.460 704.650 38.520 ;
        RECT 1028.170 38.460 1028.490 38.520 ;
      LAYER via ;
        RECT 1028.200 582.800 1028.460 583.060 ;
        RECT 1030.960 582.800 1031.220 583.060 ;
        RECT 704.360 38.460 704.620 38.720 ;
        RECT 1028.200 38.460 1028.460 38.720 ;
      LAYER met2 ;
        RECT 1032.570 600.170 1032.850 604.000 ;
        RECT 1031.020 600.030 1032.850 600.170 ;
        RECT 1031.020 583.090 1031.160 600.030 ;
        RECT 1032.570 600.000 1032.850 600.030 ;
        RECT 1028.200 582.770 1028.460 583.090 ;
        RECT 1030.960 582.770 1031.220 583.090 ;
        RECT 1028.260 38.750 1028.400 582.770 ;
        RECT 704.360 38.430 704.620 38.750 ;
        RECT 1028.200 38.430 1028.460 38.750 ;
        RECT 704.420 2.400 704.560 38.430 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.510 590.820 1455.830 590.880 ;
        RECT 1525.890 590.820 1526.210 590.880 ;
        RECT 1455.510 590.680 1526.210 590.820 ;
        RECT 1455.510 590.620 1455.830 590.680 ;
        RECT 1525.890 590.620 1526.210 590.680 ;
        RECT 1524.970 2.960 1525.290 3.020 ;
        RECT 1525.890 2.960 1526.210 3.020 ;
        RECT 1524.970 2.820 1526.210 2.960 ;
        RECT 1524.970 2.760 1525.290 2.820 ;
        RECT 1525.890 2.760 1526.210 2.820 ;
      LAYER via ;
        RECT 1455.540 590.620 1455.800 590.880 ;
        RECT 1525.920 590.620 1526.180 590.880 ;
        RECT 1525.000 2.760 1525.260 3.020 ;
        RECT 1525.920 2.760 1526.180 3.020 ;
      LAYER met2 ;
        RECT 1454.850 600.170 1455.130 604.000 ;
        RECT 1454.850 600.030 1455.740 600.170 ;
        RECT 1454.850 600.000 1455.130 600.030 ;
        RECT 1455.600 590.910 1455.740 600.030 ;
        RECT 1455.540 590.590 1455.800 590.910 ;
        RECT 1525.920 590.590 1526.180 590.910 ;
        RECT 1525.980 3.050 1526.120 590.590 ;
        RECT 1525.000 2.730 1525.260 3.050 ;
        RECT 1525.920 2.730 1526.180 3.050 ;
        RECT 1525.060 2.400 1525.200 2.730 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1465.630 590.480 1465.950 590.540 ;
        RECT 1539.690 590.480 1540.010 590.540 ;
        RECT 1465.630 590.340 1540.010 590.480 ;
        RECT 1465.630 590.280 1465.950 590.340 ;
        RECT 1539.690 590.280 1540.010 590.340 ;
        RECT 1539.690 2.960 1540.010 3.020 ;
        RECT 1542.910 2.960 1543.230 3.020 ;
        RECT 1539.690 2.820 1543.230 2.960 ;
        RECT 1539.690 2.760 1540.010 2.820 ;
        RECT 1542.910 2.760 1543.230 2.820 ;
      LAYER via ;
        RECT 1465.660 590.280 1465.920 590.540 ;
        RECT 1539.720 590.280 1539.980 590.540 ;
        RECT 1539.720 2.760 1539.980 3.020 ;
        RECT 1542.940 2.760 1543.200 3.020 ;
      LAYER met2 ;
        RECT 1464.050 600.170 1464.330 604.000 ;
        RECT 1464.050 600.030 1465.860 600.170 ;
        RECT 1464.050 600.000 1464.330 600.030 ;
        RECT 1465.720 590.570 1465.860 600.030 ;
        RECT 1465.660 590.250 1465.920 590.570 ;
        RECT 1539.720 590.250 1539.980 590.570 ;
        RECT 1539.780 3.050 1539.920 590.250 ;
        RECT 1539.720 2.730 1539.980 3.050 ;
        RECT 1542.940 2.730 1543.200 3.050 ;
        RECT 1543.000 2.400 1543.140 2.730 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1474.830 590.140 1475.150 590.200 ;
        RECT 1474.830 590.000 1530.720 590.140 ;
        RECT 1474.830 589.940 1475.150 590.000 ;
        RECT 1530.580 589.460 1530.720 590.000 ;
        RECT 1559.470 589.460 1559.790 589.520 ;
        RECT 1530.580 589.320 1559.790 589.460 ;
        RECT 1559.470 589.260 1559.790 589.320 ;
      LAYER via ;
        RECT 1474.860 589.940 1475.120 590.200 ;
        RECT 1559.500 589.260 1559.760 589.520 ;
      LAYER met2 ;
        RECT 1473.250 600.170 1473.530 604.000 ;
        RECT 1473.250 600.030 1475.060 600.170 ;
        RECT 1473.250 600.000 1473.530 600.030 ;
        RECT 1474.920 590.230 1475.060 600.030 ;
        RECT 1474.860 589.910 1475.120 590.230 ;
        RECT 1559.500 589.230 1559.760 589.550 ;
        RECT 1559.560 3.130 1559.700 589.230 ;
        RECT 1559.560 2.990 1561.080 3.130 ;
        RECT 1560.940 2.400 1561.080 2.990 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1482.650 589.460 1482.970 589.520 ;
        RECT 1482.650 589.320 1511.860 589.460 ;
        RECT 1482.650 589.260 1482.970 589.320 ;
        RECT 1511.720 588.780 1511.860 589.320 ;
        RECT 1573.270 588.780 1573.590 588.840 ;
        RECT 1511.720 588.640 1573.590 588.780 ;
        RECT 1573.270 588.580 1573.590 588.640 ;
        RECT 1573.270 62.120 1573.590 62.180 ;
        RECT 1578.790 62.120 1579.110 62.180 ;
        RECT 1573.270 61.980 1579.110 62.120 ;
        RECT 1573.270 61.920 1573.590 61.980 ;
        RECT 1578.790 61.920 1579.110 61.980 ;
      LAYER via ;
        RECT 1482.680 589.260 1482.940 589.520 ;
        RECT 1573.300 588.580 1573.560 588.840 ;
        RECT 1573.300 61.920 1573.560 62.180 ;
        RECT 1578.820 61.920 1579.080 62.180 ;
      LAYER met2 ;
        RECT 1482.450 600.000 1482.730 604.000 ;
        RECT 1482.510 598.810 1482.650 600.000 ;
        RECT 1482.510 598.670 1482.880 598.810 ;
        RECT 1482.740 589.550 1482.880 598.670 ;
        RECT 1482.680 589.230 1482.940 589.550 ;
        RECT 1573.300 588.550 1573.560 588.870 ;
        RECT 1573.360 62.210 1573.500 588.550 ;
        RECT 1573.300 61.890 1573.560 62.210 ;
        RECT 1578.820 61.890 1579.080 62.210 ;
        RECT 1578.880 2.400 1579.020 61.890 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1493.230 593.200 1493.550 593.260 ;
        RECT 1594.890 593.200 1595.210 593.260 ;
        RECT 1493.230 593.060 1595.210 593.200 ;
        RECT 1493.230 593.000 1493.550 593.060 ;
        RECT 1594.890 593.000 1595.210 593.060 ;
      LAYER via ;
        RECT 1493.260 593.000 1493.520 593.260 ;
        RECT 1594.920 593.000 1595.180 593.260 ;
      LAYER met2 ;
        RECT 1491.650 600.170 1491.930 604.000 ;
        RECT 1491.650 600.030 1493.460 600.170 ;
        RECT 1491.650 600.000 1491.930 600.030 ;
        RECT 1493.320 593.290 1493.460 600.030 ;
        RECT 1493.260 592.970 1493.520 593.290 ;
        RECT 1594.920 592.970 1595.180 593.290 ;
        RECT 1594.980 2.960 1595.120 592.970 ;
        RECT 1594.980 2.820 1596.500 2.960 ;
        RECT 1596.360 2.400 1596.500 2.820 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1502.430 591.160 1502.750 591.220 ;
        RECT 1502.430 591.020 1535.320 591.160 ;
        RECT 1502.430 590.960 1502.750 591.020 ;
        RECT 1535.180 590.820 1535.320 591.020 ;
        RECT 1535.180 590.680 1540.840 590.820 ;
        RECT 1540.700 589.800 1540.840 590.680 ;
        RECT 1608.690 589.800 1609.010 589.860 ;
        RECT 1540.700 589.660 1609.010 589.800 ;
        RECT 1608.690 589.600 1609.010 589.660 ;
      LAYER via ;
        RECT 1502.460 590.960 1502.720 591.220 ;
        RECT 1608.720 589.600 1608.980 589.860 ;
      LAYER met2 ;
        RECT 1500.850 600.170 1501.130 604.000 ;
        RECT 1500.850 600.030 1502.660 600.170 ;
        RECT 1500.850 600.000 1501.130 600.030 ;
        RECT 1502.520 591.250 1502.660 600.030 ;
        RECT 1502.460 590.930 1502.720 591.250 ;
        RECT 1608.720 589.570 1608.980 589.890 ;
        RECT 1608.780 14.010 1608.920 589.570 ;
        RECT 1608.780 13.870 1614.440 14.010 ;
        RECT 1614.300 2.400 1614.440 13.870 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1510.710 592.180 1511.030 592.240 ;
        RECT 1629.390 592.180 1629.710 592.240 ;
        RECT 1510.710 592.040 1629.710 592.180 ;
        RECT 1510.710 591.980 1511.030 592.040 ;
        RECT 1629.390 591.980 1629.710 592.040 ;
        RECT 1629.390 2.960 1629.710 3.020 ;
        RECT 1632.150 2.960 1632.470 3.020 ;
        RECT 1629.390 2.820 1632.470 2.960 ;
        RECT 1629.390 2.760 1629.710 2.820 ;
        RECT 1632.150 2.760 1632.470 2.820 ;
      LAYER via ;
        RECT 1510.740 591.980 1511.000 592.240 ;
        RECT 1629.420 591.980 1629.680 592.240 ;
        RECT 1629.420 2.760 1629.680 3.020 ;
        RECT 1632.180 2.760 1632.440 3.020 ;
      LAYER met2 ;
        RECT 1510.050 600.170 1510.330 604.000 ;
        RECT 1510.050 600.030 1510.940 600.170 ;
        RECT 1510.050 600.000 1510.330 600.030 ;
        RECT 1510.800 592.270 1510.940 600.030 ;
        RECT 1510.740 591.950 1511.000 592.270 ;
        RECT 1629.420 591.950 1629.680 592.270 ;
        RECT 1629.480 3.050 1629.620 591.950 ;
        RECT 1629.420 2.730 1629.680 3.050 ;
        RECT 1632.180 2.730 1632.440 3.050 ;
        RECT 1632.240 2.400 1632.380 2.730 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1520.830 591.840 1521.150 591.900 ;
        RECT 1650.090 591.840 1650.410 591.900 ;
        RECT 1520.830 591.700 1650.410 591.840 ;
        RECT 1520.830 591.640 1521.150 591.700 ;
        RECT 1650.090 591.640 1650.410 591.700 ;
      LAYER via ;
        RECT 1520.860 591.640 1521.120 591.900 ;
        RECT 1650.120 591.640 1650.380 591.900 ;
      LAYER met2 ;
        RECT 1519.250 600.170 1519.530 604.000 ;
        RECT 1519.250 600.030 1521.060 600.170 ;
        RECT 1519.250 600.000 1519.530 600.030 ;
        RECT 1520.920 591.930 1521.060 600.030 ;
        RECT 1520.860 591.610 1521.120 591.930 ;
        RECT 1650.120 591.610 1650.380 591.930 ;
        RECT 1650.180 2.400 1650.320 591.610 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1530.030 591.500 1530.350 591.560 ;
        RECT 1664.350 591.500 1664.670 591.560 ;
        RECT 1530.030 591.360 1664.670 591.500 ;
        RECT 1530.030 591.300 1530.350 591.360 ;
        RECT 1664.350 591.300 1664.670 591.360 ;
        RECT 1664.350 2.960 1664.670 3.020 ;
        RECT 1668.030 2.960 1668.350 3.020 ;
        RECT 1664.350 2.820 1668.350 2.960 ;
        RECT 1664.350 2.760 1664.670 2.820 ;
        RECT 1668.030 2.760 1668.350 2.820 ;
      LAYER via ;
        RECT 1530.060 591.300 1530.320 591.560 ;
        RECT 1664.380 591.300 1664.640 591.560 ;
        RECT 1664.380 2.760 1664.640 3.020 ;
        RECT 1668.060 2.760 1668.320 3.020 ;
      LAYER met2 ;
        RECT 1528.450 600.170 1528.730 604.000 ;
        RECT 1528.450 600.030 1530.260 600.170 ;
        RECT 1528.450 600.000 1528.730 600.030 ;
        RECT 1530.120 591.590 1530.260 600.030 ;
        RECT 1530.060 591.270 1530.320 591.590 ;
        RECT 1664.380 591.270 1664.640 591.590 ;
        RECT 1664.440 3.050 1664.580 591.270 ;
        RECT 1664.380 2.730 1664.640 3.050 ;
        RECT 1668.060 2.730 1668.320 3.050 ;
        RECT 1668.120 2.400 1668.260 2.730 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1538.310 591.160 1538.630 591.220 ;
        RECT 1684.590 591.160 1684.910 591.220 ;
        RECT 1538.310 591.020 1684.910 591.160 ;
        RECT 1538.310 590.960 1538.630 591.020 ;
        RECT 1684.590 590.960 1684.910 591.020 ;
        RECT 1684.590 14.180 1684.910 14.240 ;
        RECT 1684.590 14.040 1685.280 14.180 ;
        RECT 1684.590 13.980 1684.910 14.040 ;
        RECT 1685.140 13.900 1685.280 14.040 ;
        RECT 1685.050 13.640 1685.370 13.900 ;
        RECT 1685.050 2.960 1685.370 3.020 ;
        RECT 1685.510 2.960 1685.830 3.020 ;
        RECT 1685.050 2.820 1685.830 2.960 ;
        RECT 1685.050 2.760 1685.370 2.820 ;
        RECT 1685.510 2.760 1685.830 2.820 ;
      LAYER via ;
        RECT 1538.340 590.960 1538.600 591.220 ;
        RECT 1684.620 590.960 1684.880 591.220 ;
        RECT 1684.620 13.980 1684.880 14.240 ;
        RECT 1685.080 13.640 1685.340 13.900 ;
        RECT 1685.080 2.760 1685.340 3.020 ;
        RECT 1685.540 2.760 1685.800 3.020 ;
      LAYER met2 ;
        RECT 1537.650 600.170 1537.930 604.000 ;
        RECT 1537.650 600.030 1538.540 600.170 ;
        RECT 1537.650 600.000 1537.930 600.030 ;
        RECT 1538.400 591.250 1538.540 600.030 ;
        RECT 1538.340 590.930 1538.600 591.250 ;
        RECT 1684.620 590.930 1684.880 591.250 ;
        RECT 1684.680 14.270 1684.820 590.930 ;
        RECT 1684.620 13.950 1684.880 14.270 ;
        RECT 1685.080 13.610 1685.340 13.930 ;
        RECT 1685.140 3.050 1685.280 13.610 ;
        RECT 1685.080 2.730 1685.340 3.050 ;
        RECT 1685.540 2.730 1685.800 3.050 ;
        RECT 1685.600 2.400 1685.740 2.730 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 722.270 38.320 722.590 38.380 ;
        RECT 1042.890 38.320 1043.210 38.380 ;
        RECT 722.270 38.180 1043.210 38.320 ;
        RECT 722.270 38.120 722.590 38.180 ;
        RECT 1042.890 38.120 1043.210 38.180 ;
      LAYER via ;
        RECT 722.300 38.120 722.560 38.380 ;
        RECT 1042.920 38.120 1043.180 38.380 ;
      LAYER met2 ;
        RECT 1041.770 600.170 1042.050 604.000 ;
        RECT 1041.770 600.030 1043.120 600.170 ;
        RECT 1041.770 600.000 1042.050 600.030 ;
        RECT 1042.980 38.410 1043.120 600.030 ;
        RECT 722.300 38.090 722.560 38.410 ;
        RECT 1042.920 38.090 1043.180 38.410 ;
        RECT 722.360 2.400 722.500 38.090 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1583.390 590.820 1583.710 590.880 ;
        RECT 1698.390 590.820 1698.710 590.880 ;
        RECT 1583.390 590.680 1698.710 590.820 ;
        RECT 1583.390 590.620 1583.710 590.680 ;
        RECT 1698.390 590.620 1698.710 590.680 ;
        RECT 1548.430 587.760 1548.750 587.820 ;
        RECT 1583.390 587.760 1583.710 587.820 ;
        RECT 1548.430 587.620 1583.710 587.760 ;
        RECT 1548.430 587.560 1548.750 587.620 ;
        RECT 1583.390 587.560 1583.710 587.620 ;
        RECT 1698.390 579.600 1698.710 579.660 ;
        RECT 1699.310 579.600 1699.630 579.660 ;
        RECT 1698.390 579.460 1699.630 579.600 ;
        RECT 1698.390 579.400 1698.710 579.460 ;
        RECT 1699.310 579.400 1699.630 579.460 ;
        RECT 1698.390 531.660 1698.710 531.720 ;
        RECT 1699.310 531.660 1699.630 531.720 ;
        RECT 1698.390 531.520 1699.630 531.660 ;
        RECT 1698.390 531.460 1698.710 531.520 ;
        RECT 1699.310 531.460 1699.630 531.520 ;
        RECT 1698.390 13.980 1698.710 14.240 ;
        RECT 1698.480 13.840 1698.620 13.980 ;
        RECT 1700.690 13.840 1701.010 13.900 ;
        RECT 1698.480 13.700 1701.010 13.840 ;
        RECT 1700.690 13.640 1701.010 13.700 ;
        RECT 1700.690 2.960 1701.010 3.020 ;
        RECT 1703.450 2.960 1703.770 3.020 ;
        RECT 1700.690 2.820 1703.770 2.960 ;
        RECT 1700.690 2.760 1701.010 2.820 ;
        RECT 1703.450 2.760 1703.770 2.820 ;
      LAYER via ;
        RECT 1583.420 590.620 1583.680 590.880 ;
        RECT 1698.420 590.620 1698.680 590.880 ;
        RECT 1548.460 587.560 1548.720 587.820 ;
        RECT 1583.420 587.560 1583.680 587.820 ;
        RECT 1698.420 579.400 1698.680 579.660 ;
        RECT 1699.340 579.400 1699.600 579.660 ;
        RECT 1698.420 531.460 1698.680 531.720 ;
        RECT 1699.340 531.460 1699.600 531.720 ;
        RECT 1698.420 13.980 1698.680 14.240 ;
        RECT 1700.720 13.640 1700.980 13.900 ;
        RECT 1700.720 2.760 1700.980 3.020 ;
        RECT 1703.480 2.760 1703.740 3.020 ;
      LAYER met2 ;
        RECT 1546.850 600.170 1547.130 604.000 ;
        RECT 1546.850 600.030 1548.660 600.170 ;
        RECT 1546.850 600.000 1547.130 600.030 ;
        RECT 1548.520 587.850 1548.660 600.030 ;
        RECT 1583.420 590.590 1583.680 590.910 ;
        RECT 1698.420 590.590 1698.680 590.910 ;
        RECT 1583.480 587.850 1583.620 590.590 ;
        RECT 1548.460 587.530 1548.720 587.850 ;
        RECT 1583.420 587.530 1583.680 587.850 ;
        RECT 1698.480 579.690 1698.620 590.590 ;
        RECT 1698.420 579.370 1698.680 579.690 ;
        RECT 1699.340 579.370 1699.600 579.690 ;
        RECT 1699.400 531.750 1699.540 579.370 ;
        RECT 1698.420 531.430 1698.680 531.750 ;
        RECT 1699.340 531.430 1699.600 531.750 ;
        RECT 1698.480 14.270 1698.620 531.430 ;
        RECT 1698.420 13.950 1698.680 14.270 ;
        RECT 1700.720 13.610 1700.980 13.930 ;
        RECT 1700.780 3.050 1700.920 13.610 ;
        RECT 1700.720 2.730 1700.980 3.050 ;
        RECT 1703.480 2.730 1703.740 3.050 ;
        RECT 1703.540 2.400 1703.680 2.730 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1582.930 590.480 1583.250 590.540 ;
        RECT 1719.550 590.480 1719.870 590.540 ;
        RECT 1582.930 590.340 1719.870 590.480 ;
        RECT 1582.930 590.280 1583.250 590.340 ;
        RECT 1719.550 590.280 1719.870 590.340 ;
        RECT 1557.630 588.100 1557.950 588.160 ;
        RECT 1582.930 588.100 1583.250 588.160 ;
        RECT 1557.630 587.960 1583.250 588.100 ;
        RECT 1557.630 587.900 1557.950 587.960 ;
        RECT 1582.930 587.900 1583.250 587.960 ;
        RECT 1719.550 579.600 1719.870 579.660 ;
        RECT 1720.470 579.600 1720.790 579.660 ;
        RECT 1719.550 579.460 1720.790 579.600 ;
        RECT 1719.550 579.400 1719.870 579.460 ;
        RECT 1720.470 579.400 1720.790 579.460 ;
        RECT 1719.550 531.660 1719.870 531.720 ;
        RECT 1720.470 531.660 1720.790 531.720 ;
        RECT 1719.550 531.520 1720.790 531.660 ;
        RECT 1719.550 531.460 1719.870 531.520 ;
        RECT 1720.470 531.460 1720.790 531.520 ;
        RECT 1719.550 483.040 1719.870 483.100 ;
        RECT 1720.470 483.040 1720.790 483.100 ;
        RECT 1719.550 482.900 1720.790 483.040 ;
        RECT 1719.550 482.840 1719.870 482.900 ;
        RECT 1720.470 482.840 1720.790 482.900 ;
        RECT 1719.550 435.100 1719.870 435.160 ;
        RECT 1720.470 435.100 1720.790 435.160 ;
        RECT 1719.550 434.960 1720.790 435.100 ;
        RECT 1719.550 434.900 1719.870 434.960 ;
        RECT 1720.470 434.900 1720.790 434.960 ;
        RECT 1719.550 13.980 1719.870 14.240 ;
        RECT 1719.640 13.840 1719.780 13.980 ;
        RECT 1720.010 13.840 1720.330 13.900 ;
        RECT 1719.640 13.700 1720.330 13.840 ;
        RECT 1720.010 13.640 1720.330 13.700 ;
        RECT 1720.010 2.960 1720.330 3.020 ;
        RECT 1721.390 2.960 1721.710 3.020 ;
        RECT 1720.010 2.820 1721.710 2.960 ;
        RECT 1720.010 2.760 1720.330 2.820 ;
        RECT 1721.390 2.760 1721.710 2.820 ;
      LAYER via ;
        RECT 1582.960 590.280 1583.220 590.540 ;
        RECT 1719.580 590.280 1719.840 590.540 ;
        RECT 1557.660 587.900 1557.920 588.160 ;
        RECT 1582.960 587.900 1583.220 588.160 ;
        RECT 1719.580 579.400 1719.840 579.660 ;
        RECT 1720.500 579.400 1720.760 579.660 ;
        RECT 1719.580 531.460 1719.840 531.720 ;
        RECT 1720.500 531.460 1720.760 531.720 ;
        RECT 1719.580 482.840 1719.840 483.100 ;
        RECT 1720.500 482.840 1720.760 483.100 ;
        RECT 1719.580 434.900 1719.840 435.160 ;
        RECT 1720.500 434.900 1720.760 435.160 ;
        RECT 1719.580 13.980 1719.840 14.240 ;
        RECT 1720.040 13.640 1720.300 13.900 ;
        RECT 1720.040 2.760 1720.300 3.020 ;
        RECT 1721.420 2.760 1721.680 3.020 ;
      LAYER met2 ;
        RECT 1556.050 600.170 1556.330 604.000 ;
        RECT 1556.050 600.030 1557.860 600.170 ;
        RECT 1556.050 600.000 1556.330 600.030 ;
        RECT 1557.720 588.190 1557.860 600.030 ;
        RECT 1582.960 590.250 1583.220 590.570 ;
        RECT 1719.580 590.250 1719.840 590.570 ;
        RECT 1583.020 588.190 1583.160 590.250 ;
        RECT 1557.660 587.870 1557.920 588.190 ;
        RECT 1582.960 587.870 1583.220 588.190 ;
        RECT 1719.640 579.690 1719.780 590.250 ;
        RECT 1719.580 579.370 1719.840 579.690 ;
        RECT 1720.500 579.370 1720.760 579.690 ;
        RECT 1720.560 531.750 1720.700 579.370 ;
        RECT 1719.580 531.430 1719.840 531.750 ;
        RECT 1720.500 531.430 1720.760 531.750 ;
        RECT 1719.640 483.130 1719.780 531.430 ;
        RECT 1719.580 482.810 1719.840 483.130 ;
        RECT 1720.500 482.810 1720.760 483.130 ;
        RECT 1720.560 435.190 1720.700 482.810 ;
        RECT 1719.580 434.870 1719.840 435.190 ;
        RECT 1720.500 434.870 1720.760 435.190 ;
        RECT 1719.640 14.270 1719.780 434.870 ;
        RECT 1719.580 13.950 1719.840 14.270 ;
        RECT 1720.040 13.610 1720.300 13.930 ;
        RECT 1720.100 3.050 1720.240 13.610 ;
        RECT 1720.040 2.730 1720.300 3.050 ;
        RECT 1721.420 2.730 1721.680 3.050 ;
        RECT 1721.480 2.400 1721.620 2.730 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1565.910 590.140 1566.230 590.200 ;
        RECT 1739.790 590.140 1740.110 590.200 ;
        RECT 1565.910 590.000 1740.110 590.140 ;
        RECT 1565.910 589.940 1566.230 590.000 ;
        RECT 1739.790 589.940 1740.110 590.000 ;
      LAYER via ;
        RECT 1565.940 589.940 1566.200 590.200 ;
        RECT 1739.820 589.940 1740.080 590.200 ;
      LAYER met2 ;
        RECT 1565.250 600.170 1565.530 604.000 ;
        RECT 1565.250 600.030 1566.140 600.170 ;
        RECT 1565.250 600.000 1565.530 600.030 ;
        RECT 1566.000 590.230 1566.140 600.030 ;
        RECT 1565.940 589.910 1566.200 590.230 ;
        RECT 1739.820 589.910 1740.080 590.230 ;
        RECT 1739.880 3.130 1740.020 589.910 ;
        RECT 1739.420 2.990 1740.020 3.130 ;
        RECT 1739.420 2.400 1739.560 2.990 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1576.030 588.780 1576.350 588.840 ;
        RECT 1579.710 588.780 1580.030 588.840 ;
        RECT 1576.030 588.640 1580.030 588.780 ;
        RECT 1576.030 588.580 1576.350 588.640 ;
        RECT 1579.710 588.580 1580.030 588.640 ;
        RECT 1579.710 32.880 1580.030 32.940 ;
        RECT 1755.430 32.880 1755.750 32.940 ;
        RECT 1579.710 32.740 1755.750 32.880 ;
        RECT 1579.710 32.680 1580.030 32.740 ;
        RECT 1755.430 32.680 1755.750 32.740 ;
      LAYER via ;
        RECT 1576.060 588.580 1576.320 588.840 ;
        RECT 1579.740 588.580 1580.000 588.840 ;
        RECT 1579.740 32.680 1580.000 32.940 ;
        RECT 1755.460 32.680 1755.720 32.940 ;
      LAYER met2 ;
        RECT 1574.450 600.170 1574.730 604.000 ;
        RECT 1574.450 600.030 1576.260 600.170 ;
        RECT 1574.450 600.000 1574.730 600.030 ;
        RECT 1576.120 588.870 1576.260 600.030 ;
        RECT 1576.060 588.550 1576.320 588.870 ;
        RECT 1579.740 588.550 1580.000 588.870 ;
        RECT 1579.800 32.970 1579.940 588.550 ;
        RECT 1579.740 32.650 1580.000 32.970 ;
        RECT 1755.460 32.650 1755.720 32.970 ;
        RECT 1755.520 32.370 1755.660 32.650 ;
        RECT 1755.520 32.230 1757.040 32.370 ;
        RECT 1756.900 2.400 1757.040 32.230 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1585.230 532.000 1585.550 532.060 ;
        RECT 1586.150 532.000 1586.470 532.060 ;
        RECT 1585.230 531.860 1586.470 532.000 ;
        RECT 1585.230 531.800 1585.550 531.860 ;
        RECT 1586.150 531.800 1586.470 531.860 ;
        RECT 1584.310 524.180 1584.630 524.240 ;
        RECT 1585.230 524.180 1585.550 524.240 ;
        RECT 1584.310 524.040 1585.550 524.180 ;
        RECT 1584.310 523.980 1584.630 524.040 ;
        RECT 1585.230 523.980 1585.550 524.040 ;
        RECT 1584.310 476.240 1584.630 476.300 ;
        RECT 1585.230 476.240 1585.550 476.300 ;
        RECT 1584.310 476.100 1585.550 476.240 ;
        RECT 1584.310 476.040 1584.630 476.100 ;
        RECT 1585.230 476.040 1585.550 476.100 ;
        RECT 1584.770 434.760 1585.090 434.820 ;
        RECT 1585.690 434.760 1586.010 434.820 ;
        RECT 1584.770 434.620 1586.010 434.760 ;
        RECT 1584.770 434.560 1585.090 434.620 ;
        RECT 1585.690 434.560 1586.010 434.620 ;
        RECT 1584.770 386.480 1585.090 386.540 ;
        RECT 1586.150 386.480 1586.470 386.540 ;
        RECT 1584.770 386.340 1586.470 386.480 ;
        RECT 1584.770 386.280 1585.090 386.340 ;
        RECT 1586.150 386.280 1586.470 386.340 ;
        RECT 1585.690 241.640 1586.010 241.700 ;
        RECT 1586.150 241.640 1586.470 241.700 ;
        RECT 1585.690 241.500 1586.470 241.640 ;
        RECT 1585.690 241.440 1586.010 241.500 ;
        RECT 1586.150 241.440 1586.470 241.500 ;
        RECT 1585.690 145.080 1586.010 145.140 ;
        RECT 1586.150 145.080 1586.470 145.140 ;
        RECT 1585.690 144.940 1586.470 145.080 ;
        RECT 1585.690 144.880 1586.010 144.940 ;
        RECT 1586.150 144.880 1586.470 144.940 ;
        RECT 1585.230 29.480 1585.550 29.540 ;
        RECT 1774.750 29.480 1775.070 29.540 ;
        RECT 1585.230 29.340 1775.070 29.480 ;
        RECT 1585.230 29.280 1585.550 29.340 ;
        RECT 1774.750 29.280 1775.070 29.340 ;
      LAYER via ;
        RECT 1585.260 531.800 1585.520 532.060 ;
        RECT 1586.180 531.800 1586.440 532.060 ;
        RECT 1584.340 523.980 1584.600 524.240 ;
        RECT 1585.260 523.980 1585.520 524.240 ;
        RECT 1584.340 476.040 1584.600 476.300 ;
        RECT 1585.260 476.040 1585.520 476.300 ;
        RECT 1584.800 434.560 1585.060 434.820 ;
        RECT 1585.720 434.560 1585.980 434.820 ;
        RECT 1584.800 386.280 1585.060 386.540 ;
        RECT 1586.180 386.280 1586.440 386.540 ;
        RECT 1585.720 241.440 1585.980 241.700 ;
        RECT 1586.180 241.440 1586.440 241.700 ;
        RECT 1585.720 144.880 1585.980 145.140 ;
        RECT 1586.180 144.880 1586.440 145.140 ;
        RECT 1585.260 29.280 1585.520 29.540 ;
        RECT 1774.780 29.280 1775.040 29.540 ;
      LAYER met2 ;
        RECT 1583.650 600.850 1583.930 604.000 ;
        RECT 1583.650 600.710 1585.460 600.850 ;
        RECT 1583.650 600.000 1583.930 600.710 ;
        RECT 1585.320 555.290 1585.460 600.710 ;
        RECT 1585.320 555.150 1586.380 555.290 ;
        RECT 1586.240 532.090 1586.380 555.150 ;
        RECT 1585.260 531.770 1585.520 532.090 ;
        RECT 1586.180 531.770 1586.440 532.090 ;
        RECT 1585.320 524.270 1585.460 531.770 ;
        RECT 1584.340 523.950 1584.600 524.270 ;
        RECT 1585.260 523.950 1585.520 524.270 ;
        RECT 1584.400 476.330 1584.540 523.950 ;
        RECT 1584.340 476.010 1584.600 476.330 ;
        RECT 1585.260 476.010 1585.520 476.330 ;
        RECT 1585.320 434.930 1585.460 476.010 ;
        RECT 1585.320 434.850 1585.920 434.930 ;
        RECT 1584.800 434.530 1585.060 434.850 ;
        RECT 1585.320 434.790 1585.980 434.850 ;
        RECT 1585.720 434.530 1585.980 434.790 ;
        RECT 1584.860 386.570 1585.000 434.530 ;
        RECT 1584.800 386.250 1585.060 386.570 ;
        RECT 1586.180 386.250 1586.440 386.570 ;
        RECT 1586.240 351.970 1586.380 386.250 ;
        RECT 1585.780 351.830 1586.380 351.970 ;
        RECT 1585.780 303.690 1585.920 351.830 ;
        RECT 1585.780 303.550 1586.380 303.690 ;
        RECT 1586.240 241.730 1586.380 303.550 ;
        RECT 1585.720 241.410 1585.980 241.730 ;
        RECT 1586.180 241.410 1586.440 241.730 ;
        RECT 1585.780 207.130 1585.920 241.410 ;
        RECT 1585.780 206.990 1586.380 207.130 ;
        RECT 1586.240 145.170 1586.380 206.990 ;
        RECT 1585.720 144.850 1585.980 145.170 ;
        RECT 1586.180 144.850 1586.440 145.170 ;
        RECT 1585.780 110.570 1585.920 144.850 ;
        RECT 1585.780 110.430 1586.380 110.570 ;
        RECT 1586.240 62.290 1586.380 110.430 ;
        RECT 1585.320 62.150 1586.380 62.290 ;
        RECT 1585.320 29.570 1585.460 62.150 ;
        RECT 1585.260 29.250 1585.520 29.570 ;
        RECT 1774.780 29.250 1775.040 29.570 ;
        RECT 1774.840 2.400 1774.980 29.250 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.050 30.500 1593.370 30.560 ;
        RECT 1792.690 30.500 1793.010 30.560 ;
        RECT 1593.050 30.360 1793.010 30.500 ;
        RECT 1593.050 30.300 1593.370 30.360 ;
        RECT 1792.690 30.300 1793.010 30.360 ;
      LAYER via ;
        RECT 1593.080 30.300 1593.340 30.560 ;
        RECT 1792.720 30.300 1792.980 30.560 ;
      LAYER met2 ;
        RECT 1592.850 600.000 1593.130 604.000 ;
        RECT 1592.910 598.810 1593.050 600.000 ;
        RECT 1592.910 598.670 1593.280 598.810 ;
        RECT 1593.140 30.590 1593.280 598.670 ;
        RECT 1593.080 30.270 1593.340 30.590 ;
        RECT 1792.720 30.270 1792.980 30.590 ;
        RECT 1792.780 2.400 1792.920 30.270 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1603.630 588.780 1603.950 588.840 ;
        RECT 1606.850 588.780 1607.170 588.840 ;
        RECT 1603.630 588.640 1607.170 588.780 ;
        RECT 1603.630 588.580 1603.950 588.640 ;
        RECT 1606.850 588.580 1607.170 588.640 ;
        RECT 1606.850 34.240 1607.170 34.300 ;
        RECT 1810.630 34.240 1810.950 34.300 ;
        RECT 1606.850 34.100 1810.950 34.240 ;
        RECT 1606.850 34.040 1607.170 34.100 ;
        RECT 1810.630 34.040 1810.950 34.100 ;
      LAYER via ;
        RECT 1603.660 588.580 1603.920 588.840 ;
        RECT 1606.880 588.580 1607.140 588.840 ;
        RECT 1606.880 34.040 1607.140 34.300 ;
        RECT 1810.660 34.040 1810.920 34.300 ;
      LAYER met2 ;
        RECT 1602.050 600.170 1602.330 604.000 ;
        RECT 1602.050 600.030 1603.860 600.170 ;
        RECT 1602.050 600.000 1602.330 600.030 ;
        RECT 1603.720 588.870 1603.860 600.030 ;
        RECT 1603.660 588.550 1603.920 588.870 ;
        RECT 1606.880 588.550 1607.140 588.870 ;
        RECT 1606.940 34.330 1607.080 588.550 ;
        RECT 1606.880 34.010 1607.140 34.330 ;
        RECT 1810.660 34.010 1810.920 34.330 ;
        RECT 1810.720 2.400 1810.860 34.010 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1612.830 586.740 1613.150 586.800 ;
        RECT 1614.210 586.740 1614.530 586.800 ;
        RECT 1612.830 586.600 1614.530 586.740 ;
        RECT 1612.830 586.540 1613.150 586.600 ;
        RECT 1614.210 586.540 1614.530 586.600 ;
        RECT 1614.210 21.320 1614.530 21.380 ;
        RECT 1828.570 21.320 1828.890 21.380 ;
        RECT 1614.210 21.180 1828.890 21.320 ;
        RECT 1614.210 21.120 1614.530 21.180 ;
        RECT 1828.570 21.120 1828.890 21.180 ;
      LAYER via ;
        RECT 1612.860 586.540 1613.120 586.800 ;
        RECT 1614.240 586.540 1614.500 586.800 ;
        RECT 1614.240 21.120 1614.500 21.380 ;
        RECT 1828.600 21.120 1828.860 21.380 ;
      LAYER met2 ;
        RECT 1611.250 600.170 1611.530 604.000 ;
        RECT 1611.250 600.030 1613.060 600.170 ;
        RECT 1611.250 600.000 1611.530 600.030 ;
        RECT 1612.920 586.830 1613.060 600.030 ;
        RECT 1612.860 586.510 1613.120 586.830 ;
        RECT 1614.240 586.510 1614.500 586.830 ;
        RECT 1614.300 21.410 1614.440 586.510 ;
        RECT 1614.240 21.090 1614.500 21.410 ;
        RECT 1828.600 21.090 1828.860 21.410 ;
        RECT 1828.660 2.400 1828.800 21.090 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1620.650 21.660 1620.970 21.720 ;
        RECT 1846.050 21.660 1846.370 21.720 ;
        RECT 1620.650 21.520 1846.370 21.660 ;
        RECT 1620.650 21.460 1620.970 21.520 ;
        RECT 1846.050 21.460 1846.370 21.520 ;
      LAYER via ;
        RECT 1620.680 21.460 1620.940 21.720 ;
        RECT 1846.080 21.460 1846.340 21.720 ;
      LAYER met2 ;
        RECT 1620.450 600.000 1620.730 604.000 ;
        RECT 1620.510 598.810 1620.650 600.000 ;
        RECT 1620.510 598.670 1620.880 598.810 ;
        RECT 1620.740 21.750 1620.880 598.670 ;
        RECT 1620.680 21.430 1620.940 21.750 ;
        RECT 1846.080 21.430 1846.340 21.750 ;
        RECT 1846.140 2.400 1846.280 21.430 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1631.230 586.740 1631.550 586.800 ;
        RECT 1634.910 586.740 1635.230 586.800 ;
        RECT 1631.230 586.600 1635.230 586.740 ;
        RECT 1631.230 586.540 1631.550 586.600 ;
        RECT 1634.910 586.540 1635.230 586.600 ;
        RECT 1634.910 22.000 1635.230 22.060 ;
        RECT 1863.990 22.000 1864.310 22.060 ;
        RECT 1634.910 21.860 1864.310 22.000 ;
        RECT 1634.910 21.800 1635.230 21.860 ;
        RECT 1863.990 21.800 1864.310 21.860 ;
      LAYER via ;
        RECT 1631.260 586.540 1631.520 586.800 ;
        RECT 1634.940 586.540 1635.200 586.800 ;
        RECT 1634.940 21.800 1635.200 22.060 ;
        RECT 1864.020 21.800 1864.280 22.060 ;
      LAYER met2 ;
        RECT 1629.650 600.170 1629.930 604.000 ;
        RECT 1629.650 600.030 1631.460 600.170 ;
        RECT 1629.650 600.000 1629.930 600.030 ;
        RECT 1631.320 586.830 1631.460 600.030 ;
        RECT 1631.260 586.510 1631.520 586.830 ;
        RECT 1634.940 586.510 1635.200 586.830 ;
        RECT 1635.000 22.090 1635.140 586.510 ;
        RECT 1634.940 21.770 1635.200 22.090 ;
        RECT 1864.020 21.770 1864.280 22.090 ;
        RECT 1864.080 2.400 1864.220 21.770 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1025.870 598.980 1026.190 599.040 ;
        RECT 1050.940 598.980 1051.260 599.040 ;
        RECT 1025.870 598.840 1051.260 598.980 ;
        RECT 1025.870 598.780 1026.190 598.840 ;
        RECT 1050.940 598.780 1051.260 598.840 ;
        RECT 955.490 588.780 955.810 588.840 ;
        RECT 1025.870 588.780 1026.190 588.840 ;
        RECT 955.490 588.640 1026.190 588.780 ;
        RECT 955.490 588.580 955.810 588.640 ;
        RECT 1025.870 588.580 1026.190 588.640 ;
        RECT 740.210 15.200 740.530 15.260 ;
        RECT 955.490 15.200 955.810 15.260 ;
        RECT 740.210 15.060 955.810 15.200 ;
        RECT 740.210 15.000 740.530 15.060 ;
        RECT 955.490 15.000 955.810 15.060 ;
      LAYER via ;
        RECT 1025.900 598.780 1026.160 599.040 ;
        RECT 1050.970 598.780 1051.230 599.040 ;
        RECT 955.520 588.580 955.780 588.840 ;
        RECT 1025.900 588.580 1026.160 588.840 ;
        RECT 740.240 15.000 740.500 15.260 ;
        RECT 955.520 15.000 955.780 15.260 ;
      LAYER met2 ;
        RECT 1050.970 600.000 1051.250 604.000 ;
        RECT 1051.030 599.070 1051.170 600.000 ;
        RECT 1025.900 598.750 1026.160 599.070 ;
        RECT 1050.970 598.750 1051.230 599.070 ;
        RECT 1025.960 588.870 1026.100 598.750 ;
        RECT 955.520 588.550 955.780 588.870 ;
        RECT 1025.900 588.550 1026.160 588.870 ;
        RECT 955.580 15.290 955.720 588.550 ;
        RECT 740.240 14.970 740.500 15.290 ;
        RECT 955.520 14.970 955.780 15.290 ;
        RECT 740.300 2.400 740.440 14.970 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1640.430 586.740 1640.750 586.800 ;
        RECT 1641.810 586.740 1642.130 586.800 ;
        RECT 1640.430 586.600 1642.130 586.740 ;
        RECT 1640.430 586.540 1640.750 586.600 ;
        RECT 1641.810 586.540 1642.130 586.600 ;
        RECT 1641.810 22.340 1642.130 22.400 ;
        RECT 1881.930 22.340 1882.250 22.400 ;
        RECT 1641.810 22.200 1882.250 22.340 ;
        RECT 1641.810 22.140 1642.130 22.200 ;
        RECT 1881.930 22.140 1882.250 22.200 ;
      LAYER via ;
        RECT 1640.460 586.540 1640.720 586.800 ;
        RECT 1641.840 586.540 1642.100 586.800 ;
        RECT 1641.840 22.140 1642.100 22.400 ;
        RECT 1881.960 22.140 1882.220 22.400 ;
      LAYER met2 ;
        RECT 1638.850 600.170 1639.130 604.000 ;
        RECT 1638.850 600.030 1640.660 600.170 ;
        RECT 1638.850 600.000 1639.130 600.030 ;
        RECT 1640.520 586.830 1640.660 600.030 ;
        RECT 1640.460 586.510 1640.720 586.830 ;
        RECT 1641.840 586.510 1642.100 586.830 ;
        RECT 1641.900 22.430 1642.040 586.510 ;
        RECT 1641.840 22.110 1642.100 22.430 ;
        RECT 1881.960 22.110 1882.220 22.430 ;
        RECT 1882.020 2.400 1882.160 22.110 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1648.250 23.020 1648.570 23.080 ;
        RECT 1899.870 23.020 1900.190 23.080 ;
        RECT 1648.250 22.880 1900.190 23.020 ;
        RECT 1648.250 22.820 1648.570 22.880 ;
        RECT 1899.870 22.820 1900.190 22.880 ;
      LAYER via ;
        RECT 1648.280 22.820 1648.540 23.080 ;
        RECT 1899.900 22.820 1900.160 23.080 ;
      LAYER met2 ;
        RECT 1647.590 600.170 1647.870 604.000 ;
        RECT 1647.590 600.030 1648.480 600.170 ;
        RECT 1647.590 600.000 1647.870 600.030 ;
        RECT 1648.340 23.110 1648.480 600.030 ;
        RECT 1648.280 22.790 1648.540 23.110 ;
        RECT 1899.900 22.790 1900.160 23.110 ;
        RECT 1899.960 2.400 1900.100 22.790 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1658.370 586.740 1658.690 586.800 ;
        RECT 1662.510 586.740 1662.830 586.800 ;
        RECT 1658.370 586.600 1662.830 586.740 ;
        RECT 1658.370 586.540 1658.690 586.600 ;
        RECT 1662.510 586.540 1662.830 586.600 ;
        RECT 1662.510 22.680 1662.830 22.740 ;
        RECT 1917.810 22.680 1918.130 22.740 ;
        RECT 1662.510 22.540 1918.130 22.680 ;
        RECT 1662.510 22.480 1662.830 22.540 ;
        RECT 1917.810 22.480 1918.130 22.540 ;
      LAYER via ;
        RECT 1658.400 586.540 1658.660 586.800 ;
        RECT 1662.540 586.540 1662.800 586.800 ;
        RECT 1662.540 22.480 1662.800 22.740 ;
        RECT 1917.840 22.480 1918.100 22.740 ;
      LAYER met2 ;
        RECT 1656.790 600.170 1657.070 604.000 ;
        RECT 1656.790 600.030 1658.600 600.170 ;
        RECT 1656.790 600.000 1657.070 600.030 ;
        RECT 1658.460 586.830 1658.600 600.030 ;
        RECT 1658.400 586.510 1658.660 586.830 ;
        RECT 1662.540 586.510 1662.800 586.830 ;
        RECT 1662.600 22.770 1662.740 586.510 ;
        RECT 1662.540 22.450 1662.800 22.770 ;
        RECT 1917.840 22.450 1918.100 22.770 ;
        RECT 1917.900 2.400 1918.040 22.450 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1667.570 586.740 1667.890 586.800 ;
        RECT 1668.950 586.740 1669.270 586.800 ;
        RECT 1667.570 586.600 1669.270 586.740 ;
        RECT 1667.570 586.540 1667.890 586.600 ;
        RECT 1668.950 586.540 1669.270 586.600 ;
        RECT 1668.950 23.360 1669.270 23.420 ;
        RECT 1935.290 23.360 1935.610 23.420 ;
        RECT 1668.950 23.220 1935.610 23.360 ;
        RECT 1668.950 23.160 1669.270 23.220 ;
        RECT 1935.290 23.160 1935.610 23.220 ;
      LAYER via ;
        RECT 1667.600 586.540 1667.860 586.800 ;
        RECT 1668.980 586.540 1669.240 586.800 ;
        RECT 1668.980 23.160 1669.240 23.420 ;
        RECT 1935.320 23.160 1935.580 23.420 ;
      LAYER met2 ;
        RECT 1665.990 600.170 1666.270 604.000 ;
        RECT 1665.990 600.030 1667.800 600.170 ;
        RECT 1665.990 600.000 1666.270 600.030 ;
        RECT 1667.660 586.830 1667.800 600.030 ;
        RECT 1667.600 586.510 1667.860 586.830 ;
        RECT 1668.980 586.510 1669.240 586.830 ;
        RECT 1669.040 23.450 1669.180 586.510 ;
        RECT 1668.980 23.130 1669.240 23.450 ;
        RECT 1935.320 23.130 1935.580 23.450 ;
        RECT 1935.380 2.400 1935.520 23.130 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1676.310 27.440 1676.630 27.500 ;
        RECT 1953.230 27.440 1953.550 27.500 ;
        RECT 1676.310 27.300 1953.550 27.440 ;
        RECT 1676.310 27.240 1676.630 27.300 ;
        RECT 1953.230 27.240 1953.550 27.300 ;
      LAYER via ;
        RECT 1676.340 27.240 1676.600 27.500 ;
        RECT 1953.260 27.240 1953.520 27.500 ;
      LAYER met2 ;
        RECT 1675.190 600.170 1675.470 604.000 ;
        RECT 1675.190 600.030 1676.540 600.170 ;
        RECT 1675.190 600.000 1675.470 600.030 ;
        RECT 1676.400 27.530 1676.540 600.030 ;
        RECT 1676.340 27.210 1676.600 27.530 ;
        RECT 1953.260 27.210 1953.520 27.530 ;
        RECT 1953.320 2.400 1953.460 27.210 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.970 586.740 1686.290 586.800 ;
        RECT 1690.110 586.740 1690.430 586.800 ;
        RECT 1685.970 586.600 1690.430 586.740 ;
        RECT 1685.970 586.540 1686.290 586.600 ;
        RECT 1690.110 586.540 1690.430 586.600 ;
        RECT 1690.110 23.700 1690.430 23.760 ;
        RECT 1971.170 23.700 1971.490 23.760 ;
        RECT 1690.110 23.560 1971.490 23.700 ;
        RECT 1690.110 23.500 1690.430 23.560 ;
        RECT 1971.170 23.500 1971.490 23.560 ;
      LAYER via ;
        RECT 1686.000 586.540 1686.260 586.800 ;
        RECT 1690.140 586.540 1690.400 586.800 ;
        RECT 1690.140 23.500 1690.400 23.760 ;
        RECT 1971.200 23.500 1971.460 23.760 ;
      LAYER met2 ;
        RECT 1684.390 600.170 1684.670 604.000 ;
        RECT 1684.390 600.030 1686.200 600.170 ;
        RECT 1684.390 600.000 1684.670 600.030 ;
        RECT 1686.060 586.830 1686.200 600.030 ;
        RECT 1686.000 586.510 1686.260 586.830 ;
        RECT 1690.140 586.510 1690.400 586.830 ;
        RECT 1690.200 23.790 1690.340 586.510 ;
        RECT 1690.140 23.470 1690.400 23.790 ;
        RECT 1971.200 23.470 1971.460 23.790 ;
        RECT 1971.260 2.400 1971.400 23.470 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1695.630 427.620 1695.950 427.680 ;
        RECT 1696.090 427.620 1696.410 427.680 ;
        RECT 1695.630 427.480 1696.410 427.620 ;
        RECT 1695.630 427.420 1695.950 427.480 ;
        RECT 1696.090 427.420 1696.410 427.480 ;
        RECT 1694.710 420.820 1695.030 420.880 ;
        RECT 1695.630 420.820 1695.950 420.880 ;
        RECT 1694.710 420.680 1695.950 420.820 ;
        RECT 1694.710 420.620 1695.030 420.680 ;
        RECT 1695.630 420.620 1695.950 420.680 ;
        RECT 1696.090 331.740 1696.410 331.800 ;
        RECT 1696.550 331.740 1696.870 331.800 ;
        RECT 1696.090 331.600 1696.870 331.740 ;
        RECT 1696.090 331.540 1696.410 331.600 ;
        RECT 1696.550 331.540 1696.870 331.600 ;
        RECT 1695.630 324.260 1695.950 324.320 ;
        RECT 1697.470 324.260 1697.790 324.320 ;
        RECT 1695.630 324.120 1697.790 324.260 ;
        RECT 1695.630 324.060 1695.950 324.120 ;
        RECT 1697.470 324.060 1697.790 324.120 ;
        RECT 1696.090 228.040 1696.410 228.100 ;
        RECT 1697.470 228.040 1697.790 228.100 ;
        RECT 1696.090 227.900 1697.790 228.040 ;
        RECT 1696.090 227.840 1696.410 227.900 ;
        RECT 1697.470 227.840 1697.790 227.900 ;
        RECT 1696.090 186.900 1696.410 186.960 ;
        RECT 1695.720 186.760 1696.410 186.900 ;
        RECT 1695.720 186.280 1695.860 186.760 ;
        RECT 1696.090 186.700 1696.410 186.760 ;
        RECT 1695.630 186.020 1695.950 186.280 ;
        RECT 1696.550 90.000 1696.870 90.060 ;
        RECT 1697.010 90.000 1697.330 90.060 ;
        RECT 1696.550 89.860 1697.330 90.000 ;
        RECT 1696.550 89.800 1696.870 89.860 ;
        RECT 1697.010 89.800 1697.330 89.860 ;
        RECT 1695.630 48.520 1695.950 48.580 ;
        RECT 1697.010 48.520 1697.330 48.580 ;
        RECT 1695.630 48.380 1697.330 48.520 ;
        RECT 1695.630 48.320 1695.950 48.380 ;
        RECT 1697.010 48.320 1697.330 48.380 ;
        RECT 1695.630 47.840 1695.950 47.900 ;
        RECT 1715.410 47.840 1715.730 47.900 ;
        RECT 1695.630 47.700 1715.730 47.840 ;
        RECT 1695.630 47.640 1695.950 47.700 ;
        RECT 1715.410 47.640 1715.730 47.700 ;
        RECT 1715.410 27.100 1715.730 27.160 ;
        RECT 1989.110 27.100 1989.430 27.160 ;
        RECT 1715.410 26.960 1989.430 27.100 ;
        RECT 1715.410 26.900 1715.730 26.960 ;
        RECT 1989.110 26.900 1989.430 26.960 ;
      LAYER via ;
        RECT 1695.660 427.420 1695.920 427.680 ;
        RECT 1696.120 427.420 1696.380 427.680 ;
        RECT 1694.740 420.620 1695.000 420.880 ;
        RECT 1695.660 420.620 1695.920 420.880 ;
        RECT 1696.120 331.540 1696.380 331.800 ;
        RECT 1696.580 331.540 1696.840 331.800 ;
        RECT 1695.660 324.060 1695.920 324.320 ;
        RECT 1697.500 324.060 1697.760 324.320 ;
        RECT 1696.120 227.840 1696.380 228.100 ;
        RECT 1697.500 227.840 1697.760 228.100 ;
        RECT 1696.120 186.700 1696.380 186.960 ;
        RECT 1695.660 186.020 1695.920 186.280 ;
        RECT 1696.580 89.800 1696.840 90.060 ;
        RECT 1697.040 89.800 1697.300 90.060 ;
        RECT 1695.660 48.320 1695.920 48.580 ;
        RECT 1697.040 48.320 1697.300 48.580 ;
        RECT 1695.660 47.640 1695.920 47.900 ;
        RECT 1715.440 47.640 1715.700 47.900 ;
        RECT 1715.440 26.900 1715.700 27.160 ;
        RECT 1989.140 26.900 1989.400 27.160 ;
      LAYER met2 ;
        RECT 1693.590 600.000 1693.870 604.000 ;
        RECT 1693.650 598.810 1693.790 600.000 ;
        RECT 1693.420 598.670 1693.790 598.810 ;
        RECT 1693.420 579.885 1693.560 598.670 ;
        RECT 1693.350 579.515 1693.630 579.885 ;
        RECT 1695.190 579.515 1695.470 579.885 ;
        RECT 1695.260 545.090 1695.400 579.515 ;
        RECT 1695.260 544.950 1696.780 545.090 ;
        RECT 1696.640 483.210 1696.780 544.950 ;
        RECT 1696.640 483.070 1697.240 483.210 ;
        RECT 1697.100 428.130 1697.240 483.070 ;
        RECT 1696.180 427.990 1697.240 428.130 ;
        RECT 1696.180 427.710 1696.320 427.990 ;
        RECT 1695.660 427.390 1695.920 427.710 ;
        RECT 1696.120 427.390 1696.380 427.710 ;
        RECT 1695.720 420.910 1695.860 427.390 ;
        RECT 1694.740 420.590 1695.000 420.910 ;
        RECT 1695.660 420.590 1695.920 420.910 ;
        RECT 1694.800 376.450 1694.940 420.590 ;
        RECT 1694.800 376.310 1695.860 376.450 ;
        RECT 1695.720 339.050 1695.860 376.310 ;
        RECT 1695.720 338.910 1696.780 339.050 ;
        RECT 1696.640 331.830 1696.780 338.910 ;
        RECT 1696.120 331.570 1696.380 331.830 ;
        RECT 1695.720 331.510 1696.380 331.570 ;
        RECT 1696.580 331.510 1696.840 331.830 ;
        RECT 1695.720 331.430 1696.320 331.510 ;
        RECT 1695.720 324.350 1695.860 331.430 ;
        RECT 1695.660 324.030 1695.920 324.350 ;
        RECT 1697.500 324.030 1697.760 324.350 ;
        RECT 1697.560 228.130 1697.700 324.030 ;
        RECT 1696.120 227.810 1696.380 228.130 ;
        RECT 1697.500 227.810 1697.760 228.130 ;
        RECT 1696.180 186.990 1696.320 227.810 ;
        RECT 1696.120 186.670 1696.380 186.990 ;
        RECT 1695.660 185.990 1695.920 186.310 ;
        RECT 1695.720 145.250 1695.860 185.990 ;
        RECT 1695.260 145.110 1695.860 145.250 ;
        RECT 1695.260 143.890 1695.400 145.110 ;
        RECT 1695.260 143.750 1696.320 143.890 ;
        RECT 1696.180 137.770 1696.320 143.750 ;
        RECT 1696.180 137.630 1696.780 137.770 ;
        RECT 1696.640 90.090 1696.780 137.630 ;
        RECT 1696.580 89.770 1696.840 90.090 ;
        RECT 1697.040 89.770 1697.300 90.090 ;
        RECT 1697.100 48.610 1697.240 89.770 ;
        RECT 1695.660 48.290 1695.920 48.610 ;
        RECT 1697.040 48.290 1697.300 48.610 ;
        RECT 1695.720 47.930 1695.860 48.290 ;
        RECT 1695.660 47.610 1695.920 47.930 ;
        RECT 1715.440 47.610 1715.700 47.930 ;
        RECT 1715.500 27.190 1715.640 47.610 ;
        RECT 1715.440 26.870 1715.700 27.190 ;
        RECT 1989.140 26.870 1989.400 27.190 ;
        RECT 1989.200 2.400 1989.340 26.870 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
      LAYER via2 ;
        RECT 1693.350 579.560 1693.630 579.840 ;
        RECT 1695.190 579.560 1695.470 579.840 ;
      LAYER met3 ;
        RECT 1693.325 579.850 1693.655 579.865 ;
        RECT 1695.165 579.850 1695.495 579.865 ;
        RECT 1693.325 579.550 1695.495 579.850 ;
        RECT 1693.325 579.535 1693.655 579.550 ;
        RECT 1695.165 579.535 1695.495 579.550 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.910 26.760 1704.230 26.820 ;
        RECT 2006.590 26.760 2006.910 26.820 ;
        RECT 1703.910 26.620 2006.910 26.760 ;
        RECT 1703.910 26.560 1704.230 26.620 ;
        RECT 2006.590 26.560 2006.910 26.620 ;
      LAYER via ;
        RECT 1703.940 26.560 1704.200 26.820 ;
        RECT 2006.620 26.560 2006.880 26.820 ;
      LAYER met2 ;
        RECT 1702.790 600.170 1703.070 604.000 ;
        RECT 1702.790 600.030 1704.140 600.170 ;
        RECT 1702.790 600.000 1703.070 600.030 ;
        RECT 1704.000 26.850 1704.140 600.030 ;
        RECT 1703.940 26.530 1704.200 26.850 ;
        RECT 2006.620 26.530 2006.880 26.850 ;
        RECT 2006.680 2.400 2006.820 26.530 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1713.570 586.740 1713.890 586.800 ;
        RECT 1717.710 586.740 1718.030 586.800 ;
        RECT 1713.570 586.600 1718.030 586.740 ;
        RECT 1713.570 586.540 1713.890 586.600 ;
        RECT 1717.710 586.540 1718.030 586.600 ;
        RECT 1717.710 26.420 1718.030 26.480 ;
        RECT 2024.530 26.420 2024.850 26.480 ;
        RECT 1717.710 26.280 2024.850 26.420 ;
        RECT 1717.710 26.220 1718.030 26.280 ;
        RECT 2024.530 26.220 2024.850 26.280 ;
      LAYER via ;
        RECT 1713.600 586.540 1713.860 586.800 ;
        RECT 1717.740 586.540 1718.000 586.800 ;
        RECT 1717.740 26.220 1718.000 26.480 ;
        RECT 2024.560 26.220 2024.820 26.480 ;
      LAYER met2 ;
        RECT 1711.990 600.170 1712.270 604.000 ;
        RECT 1711.990 600.030 1713.800 600.170 ;
        RECT 1711.990 600.000 1712.270 600.030 ;
        RECT 1713.660 586.830 1713.800 600.030 ;
        RECT 1713.600 586.510 1713.860 586.830 ;
        RECT 1717.740 586.510 1718.000 586.830 ;
        RECT 1717.800 26.510 1717.940 586.510 ;
        RECT 1717.740 26.190 1718.000 26.510 ;
        RECT 2024.560 26.190 2024.820 26.510 ;
        RECT 2024.620 2.400 2024.760 26.190 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1722.770 586.740 1723.090 586.800 ;
        RECT 1724.610 586.740 1724.930 586.800 ;
        RECT 1722.770 586.600 1724.930 586.740 ;
        RECT 1722.770 586.540 1723.090 586.600 ;
        RECT 1724.610 586.540 1724.930 586.600 ;
        RECT 1724.610 26.080 1724.930 26.140 ;
        RECT 2042.470 26.080 2042.790 26.140 ;
        RECT 1724.610 25.940 2042.790 26.080 ;
        RECT 1724.610 25.880 1724.930 25.940 ;
        RECT 2042.470 25.880 2042.790 25.940 ;
      LAYER via ;
        RECT 1722.800 586.540 1723.060 586.800 ;
        RECT 1724.640 586.540 1724.900 586.800 ;
        RECT 1724.640 25.880 1724.900 26.140 ;
        RECT 2042.500 25.880 2042.760 26.140 ;
      LAYER met2 ;
        RECT 1721.190 600.170 1721.470 604.000 ;
        RECT 1721.190 600.030 1723.000 600.170 ;
        RECT 1721.190 600.000 1721.470 600.030 ;
        RECT 1722.860 586.830 1723.000 600.030 ;
        RECT 1722.800 586.510 1723.060 586.830 ;
        RECT 1724.640 586.510 1724.900 586.830 ;
        RECT 1724.700 26.170 1724.840 586.510 ;
        RECT 1724.640 25.850 1724.900 26.170 ;
        RECT 2042.500 25.850 2042.760 26.170 ;
        RECT 2042.560 2.400 2042.700 25.850 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 983.090 588.100 983.410 588.160 ;
        RECT 1058.530 588.100 1058.850 588.160 ;
        RECT 983.090 587.960 1058.850 588.100 ;
        RECT 983.090 587.900 983.410 587.960 ;
        RECT 1058.530 587.900 1058.850 587.960 ;
        RECT 757.690 19.280 758.010 19.340 ;
        RECT 983.090 19.280 983.410 19.340 ;
        RECT 757.690 19.140 983.410 19.280 ;
        RECT 757.690 19.080 758.010 19.140 ;
        RECT 983.090 19.080 983.410 19.140 ;
      LAYER via ;
        RECT 983.120 587.900 983.380 588.160 ;
        RECT 1058.560 587.900 1058.820 588.160 ;
        RECT 757.720 19.080 757.980 19.340 ;
        RECT 983.120 19.080 983.380 19.340 ;
      LAYER met2 ;
        RECT 1060.170 600.170 1060.450 604.000 ;
        RECT 1058.620 600.030 1060.450 600.170 ;
        RECT 1058.620 588.190 1058.760 600.030 ;
        RECT 1060.170 600.000 1060.450 600.030 ;
        RECT 983.120 587.870 983.380 588.190 ;
        RECT 1058.560 587.870 1058.820 588.190 ;
        RECT 983.180 19.370 983.320 587.870 ;
        RECT 757.720 19.050 757.980 19.370 ;
        RECT 983.120 19.050 983.380 19.370 ;
        RECT 757.780 2.400 757.920 19.050 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1731.510 25.740 1731.830 25.800 ;
        RECT 2060.410 25.740 2060.730 25.800 ;
        RECT 1731.510 25.600 2060.730 25.740 ;
        RECT 1731.510 25.540 1731.830 25.600 ;
        RECT 2060.410 25.540 2060.730 25.600 ;
      LAYER via ;
        RECT 1731.540 25.540 1731.800 25.800 ;
        RECT 2060.440 25.540 2060.700 25.800 ;
      LAYER met2 ;
        RECT 1730.390 600.170 1730.670 604.000 ;
        RECT 1730.390 600.030 1731.740 600.170 ;
        RECT 1730.390 600.000 1730.670 600.030 ;
        RECT 1731.600 25.830 1731.740 600.030 ;
        RECT 1731.540 25.510 1731.800 25.830 ;
        RECT 2060.440 25.510 2060.700 25.830 ;
        RECT 2060.500 2.400 2060.640 25.510 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1741.170 586.740 1741.490 586.800 ;
        RECT 1745.310 586.740 1745.630 586.800 ;
        RECT 1741.170 586.600 1745.630 586.740 ;
        RECT 1741.170 586.540 1741.490 586.600 ;
        RECT 1745.310 586.540 1745.630 586.600 ;
        RECT 1745.310 25.400 1745.630 25.460 ;
        RECT 2078.350 25.400 2078.670 25.460 ;
        RECT 1745.310 25.260 2078.670 25.400 ;
        RECT 1745.310 25.200 1745.630 25.260 ;
        RECT 2078.350 25.200 2078.670 25.260 ;
      LAYER via ;
        RECT 1741.200 586.540 1741.460 586.800 ;
        RECT 1745.340 586.540 1745.600 586.800 ;
        RECT 1745.340 25.200 1745.600 25.460 ;
        RECT 2078.380 25.200 2078.640 25.460 ;
      LAYER met2 ;
        RECT 1739.590 600.170 1739.870 604.000 ;
        RECT 1739.590 600.030 1741.400 600.170 ;
        RECT 1739.590 600.000 1739.870 600.030 ;
        RECT 1741.260 586.830 1741.400 600.030 ;
        RECT 1741.200 586.510 1741.460 586.830 ;
        RECT 1745.340 586.510 1745.600 586.830 ;
        RECT 1745.400 25.490 1745.540 586.510 ;
        RECT 1745.340 25.170 1745.600 25.490 ;
        RECT 2078.380 25.170 2078.640 25.490 ;
        RECT 2078.440 2.400 2078.580 25.170 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1750.370 586.740 1750.690 586.800 ;
        RECT 1752.210 586.740 1752.530 586.800 ;
        RECT 1750.370 586.600 1752.530 586.740 ;
        RECT 1750.370 586.540 1750.690 586.600 ;
        RECT 1752.210 586.540 1752.530 586.600 ;
        RECT 1752.210 25.060 1752.530 25.120 ;
        RECT 2095.830 25.060 2096.150 25.120 ;
        RECT 1752.210 24.920 2096.150 25.060 ;
        RECT 1752.210 24.860 1752.530 24.920 ;
        RECT 2095.830 24.860 2096.150 24.920 ;
      LAYER via ;
        RECT 1750.400 586.540 1750.660 586.800 ;
        RECT 1752.240 586.540 1752.500 586.800 ;
        RECT 1752.240 24.860 1752.500 25.120 ;
        RECT 2095.860 24.860 2096.120 25.120 ;
      LAYER met2 ;
        RECT 1748.790 600.170 1749.070 604.000 ;
        RECT 1748.790 600.030 1750.600 600.170 ;
        RECT 1748.790 600.000 1749.070 600.030 ;
        RECT 1750.460 586.830 1750.600 600.030 ;
        RECT 1750.400 586.510 1750.660 586.830 ;
        RECT 1752.240 586.510 1752.500 586.830 ;
        RECT 1752.300 25.150 1752.440 586.510 ;
        RECT 1752.240 24.830 1752.500 25.150 ;
        RECT 2095.860 24.830 2096.120 25.150 ;
        RECT 2095.920 2.400 2096.060 24.830 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1759.110 24.720 1759.430 24.780 ;
        RECT 2113.770 24.720 2114.090 24.780 ;
        RECT 1759.110 24.580 2114.090 24.720 ;
        RECT 1759.110 24.520 1759.430 24.580 ;
        RECT 2113.770 24.520 2114.090 24.580 ;
      LAYER via ;
        RECT 1759.140 24.520 1759.400 24.780 ;
        RECT 2113.800 24.520 2114.060 24.780 ;
      LAYER met2 ;
        RECT 1757.990 600.170 1758.270 604.000 ;
        RECT 1757.990 600.030 1759.340 600.170 ;
        RECT 1757.990 600.000 1758.270 600.030 ;
        RECT 1759.200 24.810 1759.340 600.030 ;
        RECT 1759.140 24.490 1759.400 24.810 ;
        RECT 2113.800 24.490 2114.060 24.810 ;
        RECT 2113.860 2.400 2114.000 24.490 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.770 586.740 1769.090 586.800 ;
        RECT 1772.910 586.740 1773.230 586.800 ;
        RECT 1768.770 586.600 1773.230 586.740 ;
        RECT 1768.770 586.540 1769.090 586.600 ;
        RECT 1772.910 586.540 1773.230 586.600 ;
        RECT 1772.910 24.380 1773.230 24.440 ;
        RECT 2131.710 24.380 2132.030 24.440 ;
        RECT 1772.910 24.240 2132.030 24.380 ;
        RECT 1772.910 24.180 1773.230 24.240 ;
        RECT 2131.710 24.180 2132.030 24.240 ;
      LAYER via ;
        RECT 1768.800 586.540 1769.060 586.800 ;
        RECT 1772.940 586.540 1773.200 586.800 ;
        RECT 1772.940 24.180 1773.200 24.440 ;
        RECT 2131.740 24.180 2132.000 24.440 ;
      LAYER met2 ;
        RECT 1767.190 600.170 1767.470 604.000 ;
        RECT 1767.190 600.030 1769.000 600.170 ;
        RECT 1767.190 600.000 1767.470 600.030 ;
        RECT 1768.860 586.830 1769.000 600.030 ;
        RECT 1768.800 586.510 1769.060 586.830 ;
        RECT 1772.940 586.510 1773.200 586.830 ;
        RECT 1773.000 24.470 1773.140 586.510 ;
        RECT 1772.940 24.150 1773.200 24.470 ;
        RECT 2131.740 24.150 2132.000 24.470 ;
        RECT 2131.800 2.400 2131.940 24.150 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1777.970 586.740 1778.290 586.800 ;
        RECT 1779.810 586.740 1780.130 586.800 ;
        RECT 1777.970 586.600 1780.130 586.740 ;
        RECT 1777.970 586.540 1778.290 586.600 ;
        RECT 1779.810 586.540 1780.130 586.600 ;
        RECT 1779.810 24.040 1780.130 24.100 ;
        RECT 2149.650 24.040 2149.970 24.100 ;
        RECT 1779.810 23.900 2149.970 24.040 ;
        RECT 1779.810 23.840 1780.130 23.900 ;
        RECT 2149.650 23.840 2149.970 23.900 ;
      LAYER via ;
        RECT 1778.000 586.540 1778.260 586.800 ;
        RECT 1779.840 586.540 1780.100 586.800 ;
        RECT 1779.840 23.840 1780.100 24.100 ;
        RECT 2149.680 23.840 2149.940 24.100 ;
      LAYER met2 ;
        RECT 1776.390 600.170 1776.670 604.000 ;
        RECT 1776.390 600.030 1778.200 600.170 ;
        RECT 1776.390 600.000 1776.670 600.030 ;
        RECT 1778.060 586.830 1778.200 600.030 ;
        RECT 1778.000 586.510 1778.260 586.830 ;
        RECT 1779.840 586.510 1780.100 586.830 ;
        RECT 1779.900 24.130 1780.040 586.510 ;
        RECT 1779.840 23.810 1780.100 24.130 ;
        RECT 2149.680 23.810 2149.940 24.130 ;
        RECT 2149.740 2.400 2149.880 23.810 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.710 36.620 1787.030 36.680 ;
        RECT 2167.590 36.620 2167.910 36.680 ;
        RECT 1786.710 36.480 2167.910 36.620 ;
        RECT 1786.710 36.420 1787.030 36.480 ;
        RECT 2167.590 36.420 2167.910 36.480 ;
      LAYER via ;
        RECT 1786.740 36.420 1787.000 36.680 ;
        RECT 2167.620 36.420 2167.880 36.680 ;
      LAYER met2 ;
        RECT 1785.590 600.170 1785.870 604.000 ;
        RECT 1785.590 600.030 1786.940 600.170 ;
        RECT 1785.590 600.000 1785.870 600.030 ;
        RECT 1786.800 36.710 1786.940 600.030 ;
        RECT 1786.740 36.390 1787.000 36.710 ;
        RECT 2167.620 36.390 2167.880 36.710 ;
        RECT 2167.680 2.400 2167.820 36.390 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1796.370 590.820 1796.690 590.880 ;
        RECT 1800.510 590.820 1800.830 590.880 ;
        RECT 1796.370 590.680 1800.830 590.820 ;
        RECT 1796.370 590.620 1796.690 590.680 ;
        RECT 1800.510 590.620 1800.830 590.680 ;
        RECT 1800.510 43.080 1800.830 43.140 ;
        RECT 2185.070 43.080 2185.390 43.140 ;
        RECT 1800.510 42.940 2185.390 43.080 ;
        RECT 1800.510 42.880 1800.830 42.940 ;
        RECT 2185.070 42.880 2185.390 42.940 ;
      LAYER via ;
        RECT 1796.400 590.620 1796.660 590.880 ;
        RECT 1800.540 590.620 1800.800 590.880 ;
        RECT 1800.540 42.880 1800.800 43.140 ;
        RECT 2185.100 42.880 2185.360 43.140 ;
      LAYER met2 ;
        RECT 1794.790 600.170 1795.070 604.000 ;
        RECT 1794.790 600.030 1796.600 600.170 ;
        RECT 1794.790 600.000 1795.070 600.030 ;
        RECT 1796.460 590.910 1796.600 600.030 ;
        RECT 1796.400 590.590 1796.660 590.910 ;
        RECT 1800.540 590.590 1800.800 590.910 ;
        RECT 1800.600 43.170 1800.740 590.590 ;
        RECT 1800.540 42.850 1800.800 43.170 ;
        RECT 2185.100 42.850 2185.360 43.170 ;
        RECT 2185.160 2.400 2185.300 42.850 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1805.570 586.740 1805.890 586.800 ;
        RECT 1807.410 586.740 1807.730 586.800 ;
        RECT 1805.570 586.600 1807.730 586.740 ;
        RECT 1805.570 586.540 1805.890 586.600 ;
        RECT 1807.410 586.540 1807.730 586.600 ;
        RECT 1807.410 43.420 1807.730 43.480 ;
        RECT 2203.010 43.420 2203.330 43.480 ;
        RECT 1807.410 43.280 2203.330 43.420 ;
        RECT 1807.410 43.220 1807.730 43.280 ;
        RECT 2203.010 43.220 2203.330 43.280 ;
      LAYER via ;
        RECT 1805.600 586.540 1805.860 586.800 ;
        RECT 1807.440 586.540 1807.700 586.800 ;
        RECT 1807.440 43.220 1807.700 43.480 ;
        RECT 2203.040 43.220 2203.300 43.480 ;
      LAYER met2 ;
        RECT 1803.990 600.170 1804.270 604.000 ;
        RECT 1803.990 600.030 1805.800 600.170 ;
        RECT 1803.990 600.000 1804.270 600.030 ;
        RECT 1805.660 586.830 1805.800 600.030 ;
        RECT 1805.600 586.510 1805.860 586.830 ;
        RECT 1807.440 586.510 1807.700 586.830 ;
        RECT 1807.500 43.510 1807.640 586.510 ;
        RECT 1807.440 43.190 1807.700 43.510 ;
        RECT 2203.040 43.190 2203.300 43.510 ;
        RECT 2203.100 2.400 2203.240 43.190 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.310 43.760 1814.630 43.820 ;
        RECT 2220.950 43.760 2221.270 43.820 ;
        RECT 1814.310 43.620 2221.270 43.760 ;
        RECT 1814.310 43.560 1814.630 43.620 ;
        RECT 2220.950 43.560 2221.270 43.620 ;
      LAYER via ;
        RECT 1814.340 43.560 1814.600 43.820 ;
        RECT 2220.980 43.560 2221.240 43.820 ;
      LAYER met2 ;
        RECT 1813.190 600.170 1813.470 604.000 ;
        RECT 1813.190 600.030 1814.540 600.170 ;
        RECT 1813.190 600.000 1813.470 600.030 ;
        RECT 1814.400 43.850 1814.540 600.030 ;
        RECT 1814.340 43.530 1814.600 43.850 ;
        RECT 2220.980 43.530 2221.240 43.850 ;
        RECT 2221.040 2.400 2221.180 43.530 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.470 26.760 869.790 26.820 ;
        RECT 1069.570 26.760 1069.890 26.820 ;
        RECT 869.470 26.620 1069.890 26.760 ;
        RECT 869.470 26.560 869.790 26.620 ;
        RECT 1069.570 26.560 1069.890 26.620 ;
        RECT 775.630 18.600 775.950 18.660 ;
        RECT 869.470 18.600 869.790 18.660 ;
        RECT 775.630 18.460 869.790 18.600 ;
        RECT 775.630 18.400 775.950 18.460 ;
        RECT 869.470 18.400 869.790 18.460 ;
      LAYER via ;
        RECT 869.500 26.560 869.760 26.820 ;
        RECT 1069.600 26.560 1069.860 26.820 ;
        RECT 775.660 18.400 775.920 18.660 ;
        RECT 869.500 18.400 869.760 18.660 ;
      LAYER met2 ;
        RECT 1069.370 600.000 1069.650 604.000 ;
        RECT 1069.430 598.810 1069.570 600.000 ;
        RECT 1069.430 598.670 1069.800 598.810 ;
        RECT 1069.660 26.850 1069.800 598.670 ;
        RECT 869.500 26.530 869.760 26.850 ;
        RECT 1069.600 26.530 1069.860 26.850 ;
        RECT 869.560 18.690 869.700 26.530 ;
        RECT 775.660 18.370 775.920 18.690 ;
        RECT 869.500 18.370 869.760 18.690 ;
        RECT 775.720 2.400 775.860 18.370 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1823.970 586.740 1824.290 586.800 ;
        RECT 1828.110 586.740 1828.430 586.800 ;
        RECT 1823.970 586.600 1828.430 586.740 ;
        RECT 1823.970 586.540 1824.290 586.600 ;
        RECT 1828.110 586.540 1828.430 586.600 ;
        RECT 1828.110 44.100 1828.430 44.160 ;
        RECT 2238.890 44.100 2239.210 44.160 ;
        RECT 1828.110 43.960 2239.210 44.100 ;
        RECT 1828.110 43.900 1828.430 43.960 ;
        RECT 2238.890 43.900 2239.210 43.960 ;
      LAYER via ;
        RECT 1824.000 586.540 1824.260 586.800 ;
        RECT 1828.140 586.540 1828.400 586.800 ;
        RECT 1828.140 43.900 1828.400 44.160 ;
        RECT 2238.920 43.900 2239.180 44.160 ;
      LAYER met2 ;
        RECT 1822.390 600.170 1822.670 604.000 ;
        RECT 1822.390 600.030 1824.200 600.170 ;
        RECT 1822.390 600.000 1822.670 600.030 ;
        RECT 1824.060 586.830 1824.200 600.030 ;
        RECT 1824.000 586.510 1824.260 586.830 ;
        RECT 1828.140 586.510 1828.400 586.830 ;
        RECT 1828.200 44.190 1828.340 586.510 ;
        RECT 1828.140 43.870 1828.400 44.190 ;
        RECT 2238.920 43.870 2239.180 44.190 ;
        RECT 2238.980 2.400 2239.120 43.870 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1833.170 586.740 1833.490 586.800 ;
        RECT 1835.010 586.740 1835.330 586.800 ;
        RECT 1833.170 586.600 1835.330 586.740 ;
        RECT 1833.170 586.540 1833.490 586.600 ;
        RECT 1835.010 586.540 1835.330 586.600 ;
        RECT 1835.010 44.440 1835.330 44.500 ;
        RECT 2256.830 44.440 2257.150 44.500 ;
        RECT 1835.010 44.300 2257.150 44.440 ;
        RECT 1835.010 44.240 1835.330 44.300 ;
        RECT 2256.830 44.240 2257.150 44.300 ;
      LAYER via ;
        RECT 1833.200 586.540 1833.460 586.800 ;
        RECT 1835.040 586.540 1835.300 586.800 ;
        RECT 1835.040 44.240 1835.300 44.500 ;
        RECT 2256.860 44.240 2257.120 44.500 ;
      LAYER met2 ;
        RECT 1831.590 600.170 1831.870 604.000 ;
        RECT 1831.590 600.030 1833.400 600.170 ;
        RECT 1831.590 600.000 1831.870 600.030 ;
        RECT 1833.260 586.830 1833.400 600.030 ;
        RECT 1833.200 586.510 1833.460 586.830 ;
        RECT 1835.040 586.510 1835.300 586.830 ;
        RECT 1835.100 44.530 1835.240 586.510 ;
        RECT 1835.040 44.210 1835.300 44.530 ;
        RECT 2256.860 44.210 2257.120 44.530 ;
        RECT 2256.920 7.210 2257.060 44.210 ;
        RECT 2256.460 7.070 2257.060 7.210 ;
        RECT 2256.460 2.400 2256.600 7.070 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1841.910 48.180 1842.230 48.240 ;
        RECT 2274.310 48.180 2274.630 48.240 ;
        RECT 1841.910 48.040 2274.630 48.180 ;
        RECT 1841.910 47.980 1842.230 48.040 ;
        RECT 2274.310 47.980 2274.630 48.040 ;
      LAYER via ;
        RECT 1841.940 47.980 1842.200 48.240 ;
        RECT 2274.340 47.980 2274.600 48.240 ;
      LAYER met2 ;
        RECT 1840.790 600.170 1841.070 604.000 ;
        RECT 1840.790 600.030 1842.140 600.170 ;
        RECT 1840.790 600.000 1841.070 600.030 ;
        RECT 1842.000 48.270 1842.140 600.030 ;
        RECT 1841.940 47.950 1842.200 48.270 ;
        RECT 2274.340 47.950 2274.600 48.270 ;
        RECT 2274.400 2.400 2274.540 47.950 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1851.570 586.740 1851.890 586.800 ;
        RECT 1855.710 586.740 1856.030 586.800 ;
        RECT 1851.570 586.600 1856.030 586.740 ;
        RECT 1851.570 586.540 1851.890 586.600 ;
        RECT 1855.710 586.540 1856.030 586.600 ;
        RECT 1855.710 47.840 1856.030 47.900 ;
        RECT 2292.250 47.840 2292.570 47.900 ;
        RECT 1855.710 47.700 2292.570 47.840 ;
        RECT 1855.710 47.640 1856.030 47.700 ;
        RECT 2292.250 47.640 2292.570 47.700 ;
      LAYER via ;
        RECT 1851.600 586.540 1851.860 586.800 ;
        RECT 1855.740 586.540 1856.000 586.800 ;
        RECT 1855.740 47.640 1856.000 47.900 ;
        RECT 2292.280 47.640 2292.540 47.900 ;
      LAYER met2 ;
        RECT 1849.990 600.170 1850.270 604.000 ;
        RECT 1849.990 600.030 1851.800 600.170 ;
        RECT 1849.990 600.000 1850.270 600.030 ;
        RECT 1851.660 586.830 1851.800 600.030 ;
        RECT 1851.600 586.510 1851.860 586.830 ;
        RECT 1855.740 586.510 1856.000 586.830 ;
        RECT 1855.800 47.930 1855.940 586.510 ;
        RECT 1855.740 47.610 1856.000 47.930 ;
        RECT 2292.280 47.610 2292.540 47.930 ;
        RECT 2292.340 2.400 2292.480 47.610 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1860.770 586.740 1861.090 586.800 ;
        RECT 1862.610 586.740 1862.930 586.800 ;
        RECT 1860.770 586.600 1862.930 586.740 ;
        RECT 1860.770 586.540 1861.090 586.600 ;
        RECT 1862.610 586.540 1862.930 586.600 ;
        RECT 1862.610 47.500 1862.930 47.560 ;
        RECT 2310.190 47.500 2310.510 47.560 ;
        RECT 1862.610 47.360 2310.510 47.500 ;
        RECT 1862.610 47.300 1862.930 47.360 ;
        RECT 2310.190 47.300 2310.510 47.360 ;
      LAYER via ;
        RECT 1860.800 586.540 1861.060 586.800 ;
        RECT 1862.640 586.540 1862.900 586.800 ;
        RECT 1862.640 47.300 1862.900 47.560 ;
        RECT 2310.220 47.300 2310.480 47.560 ;
      LAYER met2 ;
        RECT 1859.190 600.170 1859.470 604.000 ;
        RECT 1859.190 600.030 1861.000 600.170 ;
        RECT 1859.190 600.000 1859.470 600.030 ;
        RECT 1860.860 586.830 1861.000 600.030 ;
        RECT 1860.800 586.510 1861.060 586.830 ;
        RECT 1862.640 586.510 1862.900 586.830 ;
        RECT 1862.700 47.590 1862.840 586.510 ;
        RECT 1862.640 47.270 1862.900 47.590 ;
        RECT 2310.220 47.270 2310.480 47.590 ;
        RECT 2310.280 2.400 2310.420 47.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1869.510 28.460 1869.830 28.520 ;
        RECT 2328.130 28.460 2328.450 28.520 ;
        RECT 1869.510 28.320 2328.450 28.460 ;
        RECT 1869.510 28.260 1869.830 28.320 ;
        RECT 2328.130 28.260 2328.450 28.320 ;
      LAYER via ;
        RECT 1869.540 28.260 1869.800 28.520 ;
        RECT 2328.160 28.260 2328.420 28.520 ;
      LAYER met2 ;
        RECT 1868.390 600.170 1868.670 604.000 ;
        RECT 1868.390 600.030 1869.740 600.170 ;
        RECT 1868.390 600.000 1868.670 600.030 ;
        RECT 1869.600 28.550 1869.740 600.030 ;
        RECT 1869.540 28.230 1869.800 28.550 ;
        RECT 2328.160 28.230 2328.420 28.550 ;
        RECT 2328.220 2.400 2328.360 28.230 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1879.170 586.740 1879.490 586.800 ;
        RECT 1883.310 586.740 1883.630 586.800 ;
        RECT 1879.170 586.600 1883.630 586.740 ;
        RECT 1879.170 586.540 1879.490 586.600 ;
        RECT 1883.310 586.540 1883.630 586.600 ;
        RECT 1881.930 37.640 1882.250 37.700 ;
        RECT 1883.310 37.640 1883.630 37.700 ;
        RECT 1881.930 37.500 1883.630 37.640 ;
        RECT 1881.930 37.440 1882.250 37.500 ;
        RECT 1883.310 37.440 1883.630 37.500 ;
        RECT 1881.930 28.120 1882.250 28.180 ;
        RECT 2345.610 28.120 2345.930 28.180 ;
        RECT 1881.930 27.980 2345.930 28.120 ;
        RECT 1881.930 27.920 1882.250 27.980 ;
        RECT 2345.610 27.920 2345.930 27.980 ;
      LAYER via ;
        RECT 1879.200 586.540 1879.460 586.800 ;
        RECT 1883.340 586.540 1883.600 586.800 ;
        RECT 1881.960 37.440 1882.220 37.700 ;
        RECT 1883.340 37.440 1883.600 37.700 ;
        RECT 1881.960 27.920 1882.220 28.180 ;
        RECT 2345.640 27.920 2345.900 28.180 ;
      LAYER met2 ;
        RECT 1877.590 600.170 1877.870 604.000 ;
        RECT 1877.590 600.030 1879.400 600.170 ;
        RECT 1877.590 600.000 1877.870 600.030 ;
        RECT 1879.260 586.830 1879.400 600.030 ;
        RECT 1879.200 586.510 1879.460 586.830 ;
        RECT 1883.340 586.510 1883.600 586.830 ;
        RECT 1883.400 37.730 1883.540 586.510 ;
        RECT 1881.960 37.410 1882.220 37.730 ;
        RECT 1883.340 37.410 1883.600 37.730 ;
        RECT 1882.020 28.210 1882.160 37.410 ;
        RECT 1881.960 27.890 1882.220 28.210 ;
        RECT 2345.640 27.890 2345.900 28.210 ;
        RECT 2345.700 2.400 2345.840 27.890 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1888.370 586.740 1888.690 586.800 ;
        RECT 1890.210 586.740 1890.530 586.800 ;
        RECT 1888.370 586.600 1890.530 586.740 ;
        RECT 1888.370 586.540 1888.690 586.600 ;
        RECT 1890.210 586.540 1890.530 586.600 ;
        RECT 1890.210 28.800 1890.530 28.860 ;
        RECT 2363.550 28.800 2363.870 28.860 ;
        RECT 1890.210 28.660 2363.870 28.800 ;
        RECT 1890.210 28.600 1890.530 28.660 ;
        RECT 2363.550 28.600 2363.870 28.660 ;
      LAYER via ;
        RECT 1888.400 586.540 1888.660 586.800 ;
        RECT 1890.240 586.540 1890.500 586.800 ;
        RECT 1890.240 28.600 1890.500 28.860 ;
        RECT 2363.580 28.600 2363.840 28.860 ;
      LAYER met2 ;
        RECT 1886.790 600.170 1887.070 604.000 ;
        RECT 1886.790 600.030 1888.600 600.170 ;
        RECT 1886.790 600.000 1887.070 600.030 ;
        RECT 1888.460 586.830 1888.600 600.030 ;
        RECT 1888.400 586.510 1888.660 586.830 ;
        RECT 1890.240 586.510 1890.500 586.830 ;
        RECT 1890.300 28.890 1890.440 586.510 ;
        RECT 1890.240 28.570 1890.500 28.890 ;
        RECT 2363.580 28.570 2363.840 28.890 ;
        RECT 2363.640 2.400 2363.780 28.570 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1896.650 29.480 1896.970 29.540 ;
        RECT 2381.490 29.480 2381.810 29.540 ;
        RECT 1896.650 29.340 2381.810 29.480 ;
        RECT 1896.650 29.280 1896.970 29.340 ;
        RECT 2381.490 29.280 2381.810 29.340 ;
      LAYER via ;
        RECT 1896.680 29.280 1896.940 29.540 ;
        RECT 2381.520 29.280 2381.780 29.540 ;
      LAYER met2 ;
        RECT 1895.990 600.170 1896.270 604.000 ;
        RECT 1895.990 600.030 1896.880 600.170 ;
        RECT 1895.990 600.000 1896.270 600.030 ;
        RECT 1896.740 29.570 1896.880 600.030 ;
        RECT 1896.680 29.250 1896.940 29.570 ;
        RECT 2381.520 29.250 2381.780 29.570 ;
        RECT 2381.580 2.400 2381.720 29.250 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1906.770 586.740 1907.090 586.800 ;
        RECT 1910.910 586.740 1911.230 586.800 ;
        RECT 1906.770 586.600 1911.230 586.740 ;
        RECT 1906.770 586.540 1907.090 586.600 ;
        RECT 1910.910 586.540 1911.230 586.600 ;
        RECT 1910.910 29.140 1911.230 29.200 ;
        RECT 2399.430 29.140 2399.750 29.200 ;
        RECT 1910.910 29.000 2399.750 29.140 ;
        RECT 1910.910 28.940 1911.230 29.000 ;
        RECT 2399.430 28.940 2399.750 29.000 ;
      LAYER via ;
        RECT 1906.800 586.540 1907.060 586.800 ;
        RECT 1910.940 586.540 1911.200 586.800 ;
        RECT 1910.940 28.940 1911.200 29.200 ;
        RECT 2399.460 28.940 2399.720 29.200 ;
      LAYER met2 ;
        RECT 1905.190 600.170 1905.470 604.000 ;
        RECT 1905.190 600.030 1907.000 600.170 ;
        RECT 1905.190 600.000 1905.470 600.030 ;
        RECT 1906.860 586.830 1907.000 600.030 ;
        RECT 1906.800 586.510 1907.060 586.830 ;
        RECT 1910.940 586.510 1911.200 586.830 ;
        RECT 1911.000 29.230 1911.140 586.510 ;
        RECT 1910.940 28.910 1911.200 29.230 ;
        RECT 2399.460 28.910 2399.720 29.230 ;
        RECT 2399.520 2.400 2399.660 28.910 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.570 24.720 793.890 24.780 ;
        RECT 1076.470 24.720 1076.790 24.780 ;
        RECT 793.570 24.580 1076.790 24.720 ;
        RECT 793.570 24.520 793.890 24.580 ;
        RECT 1076.470 24.520 1076.790 24.580 ;
      LAYER via ;
        RECT 793.600 24.520 793.860 24.780 ;
        RECT 1076.500 24.520 1076.760 24.780 ;
      LAYER met2 ;
        RECT 1078.570 600.170 1078.850 604.000 ;
        RECT 1076.560 600.030 1078.850 600.170 ;
        RECT 1076.560 24.810 1076.700 600.030 ;
        RECT 1078.570 600.000 1078.850 600.030 ;
        RECT 793.600 24.490 793.860 24.810 ;
        RECT 1076.500 24.490 1076.760 24.810 ;
        RECT 793.660 2.400 793.800 24.490 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 993.670 553.080 993.990 553.140 ;
        RECT 997.350 553.080 997.670 553.140 ;
        RECT 993.670 552.940 997.670 553.080 ;
        RECT 993.670 552.880 993.990 552.940 ;
        RECT 997.350 552.880 997.670 552.940 ;
        RECT 639.010 36.620 639.330 36.680 ;
        RECT 993.670 36.620 993.990 36.680 ;
        RECT 639.010 36.480 993.990 36.620 ;
        RECT 639.010 36.420 639.330 36.480 ;
        RECT 993.670 36.420 993.990 36.480 ;
      LAYER via ;
        RECT 993.700 552.880 993.960 553.140 ;
        RECT 997.380 552.880 997.640 553.140 ;
        RECT 639.040 36.420 639.300 36.680 ;
        RECT 993.700 36.420 993.960 36.680 ;
      LAYER met2 ;
        RECT 998.990 600.170 999.270 604.000 ;
        RECT 997.440 600.030 999.270 600.170 ;
        RECT 997.440 553.170 997.580 600.030 ;
        RECT 998.990 600.000 999.270 600.030 ;
        RECT 993.700 552.850 993.960 553.170 ;
        RECT 997.380 552.850 997.640 553.170 ;
        RECT 993.760 36.710 993.900 552.850 ;
        RECT 639.040 36.390 639.300 36.710 ;
        RECT 993.700 36.390 993.960 36.710 ;
        RECT 639.100 2.400 639.240 36.390 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1917.350 30.160 1917.670 30.220 ;
        RECT 2422.890 30.160 2423.210 30.220 ;
        RECT 1917.350 30.020 2423.210 30.160 ;
        RECT 1917.350 29.960 1917.670 30.020 ;
        RECT 2422.890 29.960 2423.210 30.020 ;
      LAYER via ;
        RECT 1917.380 29.960 1917.640 30.220 ;
        RECT 2422.920 29.960 2423.180 30.220 ;
      LAYER met2 ;
        RECT 1917.150 600.000 1917.430 604.000 ;
        RECT 1917.210 598.810 1917.350 600.000 ;
        RECT 1917.210 598.670 1917.580 598.810 ;
        RECT 1917.440 30.250 1917.580 598.670 ;
        RECT 1917.380 29.930 1917.640 30.250 ;
        RECT 2422.920 29.930 2423.180 30.250 ;
        RECT 2422.980 2.400 2423.120 29.930 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1927.930 586.740 1928.250 586.800 ;
        RECT 1931.610 586.740 1931.930 586.800 ;
        RECT 1927.930 586.600 1931.930 586.740 ;
        RECT 1927.930 586.540 1928.250 586.600 ;
        RECT 1931.610 586.540 1931.930 586.600 ;
        RECT 1931.610 29.820 1931.930 29.880 ;
        RECT 2440.830 29.820 2441.150 29.880 ;
        RECT 1931.610 29.680 2441.150 29.820 ;
        RECT 1931.610 29.620 1931.930 29.680 ;
        RECT 2440.830 29.620 2441.150 29.680 ;
      LAYER via ;
        RECT 1927.960 586.540 1928.220 586.800 ;
        RECT 1931.640 586.540 1931.900 586.800 ;
        RECT 1931.640 29.620 1931.900 29.880 ;
        RECT 2440.860 29.620 2441.120 29.880 ;
      LAYER met2 ;
        RECT 1926.350 600.170 1926.630 604.000 ;
        RECT 1926.350 600.030 1928.160 600.170 ;
        RECT 1926.350 600.000 1926.630 600.030 ;
        RECT 1928.020 586.830 1928.160 600.030 ;
        RECT 1927.960 586.510 1928.220 586.830 ;
        RECT 1931.640 586.510 1931.900 586.830 ;
        RECT 1931.700 29.910 1931.840 586.510 ;
        RECT 1931.640 29.590 1931.900 29.910 ;
        RECT 2440.860 29.590 2441.120 29.910 ;
        RECT 2440.920 2.400 2441.060 29.590 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1938.510 30.500 1938.830 30.560 ;
        RECT 2458.770 30.500 2459.090 30.560 ;
        RECT 1938.510 30.360 2459.090 30.500 ;
        RECT 1938.510 30.300 1938.830 30.360 ;
        RECT 2458.770 30.300 2459.090 30.360 ;
      LAYER via ;
        RECT 1938.540 30.300 1938.800 30.560 ;
        RECT 2458.800 30.300 2459.060 30.560 ;
      LAYER met2 ;
        RECT 1935.550 600.170 1935.830 604.000 ;
        RECT 1935.550 600.030 1938.280 600.170 ;
        RECT 1935.550 600.000 1935.830 600.030 ;
        RECT 1938.140 587.250 1938.280 600.030 ;
        RECT 1938.140 587.110 1938.740 587.250 ;
        RECT 1938.600 30.590 1938.740 587.110 ;
        RECT 1938.540 30.270 1938.800 30.590 ;
        RECT 2458.800 30.270 2459.060 30.590 ;
        RECT 2458.860 2.400 2459.000 30.270 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1945.410 34.240 1945.730 34.300 ;
        RECT 2476.710 34.240 2477.030 34.300 ;
        RECT 1945.410 34.100 2477.030 34.240 ;
        RECT 1945.410 34.040 1945.730 34.100 ;
        RECT 2476.710 34.040 2477.030 34.100 ;
      LAYER via ;
        RECT 1945.440 34.040 1945.700 34.300 ;
        RECT 2476.740 34.040 2477.000 34.300 ;
      LAYER met2 ;
        RECT 1944.750 600.170 1945.030 604.000 ;
        RECT 1944.750 600.030 1945.640 600.170 ;
        RECT 1944.750 600.000 1945.030 600.030 ;
        RECT 1945.500 34.330 1945.640 600.030 ;
        RECT 1945.440 34.010 1945.700 34.330 ;
        RECT 2476.740 34.010 2477.000 34.330 ;
        RECT 2476.800 2.400 2476.940 34.010 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1955.530 586.740 1955.850 586.800 ;
        RECT 1959.210 586.740 1959.530 586.800 ;
        RECT 1955.530 586.600 1959.530 586.740 ;
        RECT 1955.530 586.540 1955.850 586.600 ;
        RECT 1959.210 586.540 1959.530 586.600 ;
        RECT 2494.650 33.900 2494.970 33.960 ;
        RECT 1959.760 33.760 2494.970 33.900 ;
        RECT 1958.750 33.560 1959.070 33.620 ;
        RECT 1959.760 33.560 1959.900 33.760 ;
        RECT 2494.650 33.700 2494.970 33.760 ;
        RECT 1958.750 33.420 1959.900 33.560 ;
        RECT 1958.750 33.360 1959.070 33.420 ;
      LAYER via ;
        RECT 1955.560 586.540 1955.820 586.800 ;
        RECT 1959.240 586.540 1959.500 586.800 ;
        RECT 1958.780 33.360 1959.040 33.620 ;
        RECT 2494.680 33.700 2494.940 33.960 ;
      LAYER met2 ;
        RECT 1953.950 600.170 1954.230 604.000 ;
        RECT 1953.950 600.030 1955.760 600.170 ;
        RECT 1953.950 600.000 1954.230 600.030 ;
        RECT 1955.620 586.830 1955.760 600.030 ;
        RECT 1955.560 586.510 1955.820 586.830 ;
        RECT 1959.240 586.510 1959.500 586.830 ;
        RECT 1959.300 51.410 1959.440 586.510 ;
        RECT 1958.840 51.270 1959.440 51.410 ;
        RECT 1958.840 33.650 1958.980 51.270 ;
        RECT 2494.680 33.670 2494.940 33.990 ;
        RECT 1958.780 33.330 1959.040 33.650 ;
        RECT 2494.740 2.400 2494.880 33.670 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1966.110 33.560 1966.430 33.620 ;
        RECT 2512.130 33.560 2512.450 33.620 ;
        RECT 1966.110 33.420 2512.450 33.560 ;
        RECT 1966.110 33.360 1966.430 33.420 ;
        RECT 2512.130 33.360 2512.450 33.420 ;
      LAYER via ;
        RECT 1966.140 33.360 1966.400 33.620 ;
        RECT 2512.160 33.360 2512.420 33.620 ;
      LAYER met2 ;
        RECT 1963.150 600.170 1963.430 604.000 ;
        RECT 1963.150 600.030 1965.880 600.170 ;
        RECT 1963.150 600.000 1963.430 600.030 ;
        RECT 1965.740 587.250 1965.880 600.030 ;
        RECT 1965.740 587.110 1966.340 587.250 ;
        RECT 1966.200 33.650 1966.340 587.110 ;
        RECT 1966.140 33.330 1966.400 33.650 ;
        RECT 2512.160 33.330 2512.420 33.650 ;
        RECT 2512.220 2.400 2512.360 33.330 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1973.010 33.220 1973.330 33.280 ;
        RECT 2530.070 33.220 2530.390 33.280 ;
        RECT 1973.010 33.080 2530.390 33.220 ;
        RECT 1973.010 33.020 1973.330 33.080 ;
        RECT 2530.070 33.020 2530.390 33.080 ;
      LAYER via ;
        RECT 1973.040 33.020 1973.300 33.280 ;
        RECT 2530.100 33.020 2530.360 33.280 ;
      LAYER met2 ;
        RECT 1972.350 600.170 1972.630 604.000 ;
        RECT 1972.350 600.030 1973.240 600.170 ;
        RECT 1972.350 600.000 1972.630 600.030 ;
        RECT 1973.100 33.310 1973.240 600.030 ;
        RECT 1973.040 32.990 1973.300 33.310 ;
        RECT 2530.100 32.990 2530.360 33.310 ;
        RECT 2530.160 2.400 2530.300 32.990 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1983.130 586.740 1983.450 586.800 ;
        RECT 1986.810 586.740 1987.130 586.800 ;
        RECT 1983.130 586.600 1987.130 586.740 ;
        RECT 1983.130 586.540 1983.450 586.600 ;
        RECT 1986.810 586.540 1987.130 586.600 ;
        RECT 1986.810 32.880 1987.130 32.940 ;
        RECT 2548.010 32.880 2548.330 32.940 ;
        RECT 1986.810 32.740 2548.330 32.880 ;
        RECT 1986.810 32.680 1987.130 32.740 ;
        RECT 2548.010 32.680 2548.330 32.740 ;
      LAYER via ;
        RECT 1983.160 586.540 1983.420 586.800 ;
        RECT 1986.840 586.540 1987.100 586.800 ;
        RECT 1986.840 32.680 1987.100 32.940 ;
        RECT 2548.040 32.680 2548.300 32.940 ;
      LAYER met2 ;
        RECT 1981.550 600.170 1981.830 604.000 ;
        RECT 1981.550 600.030 1983.360 600.170 ;
        RECT 1981.550 600.000 1981.830 600.030 ;
        RECT 1983.220 586.830 1983.360 600.030 ;
        RECT 1983.160 586.510 1983.420 586.830 ;
        RECT 1986.840 586.510 1987.100 586.830 ;
        RECT 1986.900 32.970 1987.040 586.510 ;
        RECT 1986.840 32.650 1987.100 32.970 ;
        RECT 2548.040 32.650 2548.300 32.970 ;
        RECT 2548.100 2.400 2548.240 32.650 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1993.710 32.540 1994.030 32.600 ;
        RECT 2565.950 32.540 2566.270 32.600 ;
        RECT 1993.710 32.400 2566.270 32.540 ;
        RECT 1993.710 32.340 1994.030 32.400 ;
        RECT 2565.950 32.340 2566.270 32.400 ;
      LAYER via ;
        RECT 1993.740 32.340 1994.000 32.600 ;
        RECT 2565.980 32.340 2566.240 32.600 ;
      LAYER met2 ;
        RECT 1990.750 600.170 1991.030 604.000 ;
        RECT 1990.750 600.030 1993.480 600.170 ;
        RECT 1990.750 600.000 1991.030 600.030 ;
        RECT 1993.340 587.250 1993.480 600.030 ;
        RECT 1993.340 587.110 1993.940 587.250 ;
        RECT 1993.800 32.630 1993.940 587.110 ;
        RECT 1993.740 32.310 1994.000 32.630 ;
        RECT 2565.980 32.310 2566.240 32.630 ;
        RECT 2566.040 2.400 2566.180 32.310 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2000.150 32.200 2000.470 32.260 ;
        RECT 2583.890 32.200 2584.210 32.260 ;
        RECT 2000.150 32.060 2584.210 32.200 ;
        RECT 2000.150 32.000 2000.470 32.060 ;
        RECT 2583.890 32.000 2584.210 32.060 ;
      LAYER via ;
        RECT 2000.180 32.000 2000.440 32.260 ;
        RECT 2583.920 32.000 2584.180 32.260 ;
      LAYER met2 ;
        RECT 1999.950 600.000 2000.230 604.000 ;
        RECT 2000.010 598.810 2000.150 600.000 ;
        RECT 2000.010 598.670 2000.380 598.810 ;
        RECT 2000.240 32.290 2000.380 598.670 ;
        RECT 2000.180 31.970 2000.440 32.290 ;
        RECT 2583.920 31.970 2584.180 32.290 ;
        RECT 2583.980 2.400 2584.120 31.970 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.490 25.060 817.810 25.120 ;
        RECT 1090.270 25.060 1090.590 25.120 ;
        RECT 817.490 24.920 1090.590 25.060 ;
        RECT 817.490 24.860 817.810 24.920 ;
        RECT 1090.270 24.860 1090.590 24.920 ;
      LAYER via ;
        RECT 817.520 24.860 817.780 25.120 ;
        RECT 1090.300 24.860 1090.560 25.120 ;
      LAYER met2 ;
        RECT 1090.530 600.000 1090.810 604.000 ;
        RECT 1090.590 598.810 1090.730 600.000 ;
        RECT 1090.360 598.670 1090.730 598.810 ;
        RECT 1090.360 25.150 1090.500 598.670 ;
        RECT 817.520 24.830 817.780 25.150 ;
        RECT 1090.300 24.830 1090.560 25.150 ;
        RECT 817.580 2.400 817.720 24.830 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2010.730 586.740 2011.050 586.800 ;
        RECT 2013.950 586.740 2014.270 586.800 ;
        RECT 2010.730 586.600 2014.270 586.740 ;
        RECT 2010.730 586.540 2011.050 586.600 ;
        RECT 2013.950 586.540 2014.270 586.600 ;
        RECT 2013.950 31.860 2014.270 31.920 ;
        RECT 2601.370 31.860 2601.690 31.920 ;
        RECT 2013.950 31.720 2601.690 31.860 ;
        RECT 2013.950 31.660 2014.270 31.720 ;
        RECT 2601.370 31.660 2601.690 31.720 ;
      LAYER via ;
        RECT 2010.760 586.540 2011.020 586.800 ;
        RECT 2013.980 586.540 2014.240 586.800 ;
        RECT 2013.980 31.660 2014.240 31.920 ;
        RECT 2601.400 31.660 2601.660 31.920 ;
      LAYER met2 ;
        RECT 2009.150 600.170 2009.430 604.000 ;
        RECT 2009.150 600.030 2010.960 600.170 ;
        RECT 2009.150 600.000 2009.430 600.030 ;
        RECT 2010.820 586.830 2010.960 600.030 ;
        RECT 2010.760 586.510 2011.020 586.830 ;
        RECT 2013.980 586.510 2014.240 586.830 ;
        RECT 2014.040 31.950 2014.180 586.510 ;
        RECT 2013.980 31.630 2014.240 31.950 ;
        RECT 2601.400 31.630 2601.660 31.950 ;
        RECT 2601.460 2.400 2601.600 31.630 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2018.550 572.800 2018.870 572.860 ;
        RECT 2019.470 572.800 2019.790 572.860 ;
        RECT 2018.550 572.660 2019.790 572.800 ;
        RECT 2018.550 572.600 2018.870 572.660 ;
        RECT 2019.470 572.600 2019.790 572.660 ;
        RECT 2019.470 545.260 2019.790 545.320 ;
        RECT 2019.470 545.120 2020.160 545.260 ;
        RECT 2019.470 545.060 2019.790 545.120 ;
        RECT 2020.020 544.980 2020.160 545.120 ;
        RECT 2019.930 544.720 2020.250 544.980 ;
        RECT 2019.930 531.320 2020.250 531.380 ;
        RECT 2020.390 531.320 2020.710 531.380 ;
        RECT 2019.930 531.180 2020.710 531.320 ;
        RECT 2019.930 531.120 2020.250 531.180 ;
        RECT 2020.390 531.120 2020.710 531.180 ;
        RECT 2018.550 483.040 2018.870 483.100 ;
        RECT 2019.930 483.040 2020.250 483.100 ;
        RECT 2018.550 482.900 2020.250 483.040 ;
        RECT 2018.550 482.840 2018.870 482.900 ;
        RECT 2019.930 482.840 2020.250 482.900 ;
        RECT 2018.550 435.100 2018.870 435.160 ;
        RECT 2019.470 435.100 2019.790 435.160 ;
        RECT 2018.550 434.960 2019.790 435.100 ;
        RECT 2018.550 434.900 2018.870 434.960 ;
        RECT 2019.470 434.900 2019.790 434.960 ;
        RECT 2019.470 434.420 2019.790 434.480 ;
        RECT 2019.930 434.420 2020.250 434.480 ;
        RECT 2019.470 434.280 2020.250 434.420 ;
        RECT 2019.470 434.220 2019.790 434.280 ;
        RECT 2019.930 434.220 2020.250 434.280 ;
        RECT 2019.010 331.400 2019.330 331.460 ;
        RECT 2020.390 331.400 2020.710 331.460 ;
        RECT 2019.010 331.260 2020.710 331.400 ;
        RECT 2019.010 331.200 2019.330 331.260 ;
        RECT 2020.390 331.200 2020.710 331.260 ;
        RECT 2019.010 282.780 2019.330 282.840 ;
        RECT 2019.930 282.780 2020.250 282.840 ;
        RECT 2019.010 282.640 2020.250 282.780 ;
        RECT 2019.010 282.580 2019.330 282.640 ;
        RECT 2019.930 282.580 2020.250 282.640 ;
        RECT 2019.010 234.840 2019.330 234.900 ;
        RECT 2020.390 234.840 2020.710 234.900 ;
        RECT 2019.010 234.700 2020.710 234.840 ;
        RECT 2019.010 234.640 2019.330 234.700 ;
        RECT 2020.390 234.640 2020.710 234.700 ;
        RECT 2020.390 158.820 2020.710 159.080 ;
        RECT 2020.480 158.400 2020.620 158.820 ;
        RECT 2020.390 158.140 2020.710 158.400 ;
        RECT 2020.850 31.520 2021.170 31.580 ;
        RECT 2619.310 31.520 2619.630 31.580 ;
        RECT 2020.850 31.380 2619.630 31.520 ;
        RECT 2020.850 31.320 2021.170 31.380 ;
        RECT 2619.310 31.320 2619.630 31.380 ;
      LAYER via ;
        RECT 2018.580 572.600 2018.840 572.860 ;
        RECT 2019.500 572.600 2019.760 572.860 ;
        RECT 2019.500 545.060 2019.760 545.320 ;
        RECT 2019.960 544.720 2020.220 544.980 ;
        RECT 2019.960 531.120 2020.220 531.380 ;
        RECT 2020.420 531.120 2020.680 531.380 ;
        RECT 2018.580 482.840 2018.840 483.100 ;
        RECT 2019.960 482.840 2020.220 483.100 ;
        RECT 2018.580 434.900 2018.840 435.160 ;
        RECT 2019.500 434.900 2019.760 435.160 ;
        RECT 2019.500 434.220 2019.760 434.480 ;
        RECT 2019.960 434.220 2020.220 434.480 ;
        RECT 2019.040 331.200 2019.300 331.460 ;
        RECT 2020.420 331.200 2020.680 331.460 ;
        RECT 2019.040 282.580 2019.300 282.840 ;
        RECT 2019.960 282.580 2020.220 282.840 ;
        RECT 2019.040 234.640 2019.300 234.900 ;
        RECT 2020.420 234.640 2020.680 234.900 ;
        RECT 2020.420 158.820 2020.680 159.080 ;
        RECT 2020.420 158.140 2020.680 158.400 ;
        RECT 2020.880 31.320 2021.140 31.580 ;
        RECT 2619.340 31.320 2619.600 31.580 ;
      LAYER met2 ;
        RECT 2018.350 600.000 2018.630 604.000 ;
        RECT 2018.410 598.810 2018.550 600.000 ;
        RECT 2018.410 598.670 2018.780 598.810 ;
        RECT 2018.640 572.890 2018.780 598.670 ;
        RECT 2018.580 572.570 2018.840 572.890 ;
        RECT 2019.500 572.570 2019.760 572.890 ;
        RECT 2019.560 545.350 2019.700 572.570 ;
        RECT 2019.500 545.030 2019.760 545.350 ;
        RECT 2019.960 544.690 2020.220 545.010 ;
        RECT 2020.020 531.410 2020.160 544.690 ;
        RECT 2019.960 531.090 2020.220 531.410 ;
        RECT 2020.420 531.090 2020.680 531.410 ;
        RECT 2020.480 496.810 2020.620 531.090 ;
        RECT 2019.560 496.670 2020.620 496.810 ;
        RECT 2019.560 483.210 2019.700 496.670 ;
        RECT 2019.560 483.130 2020.160 483.210 ;
        RECT 2018.580 482.810 2018.840 483.130 ;
        RECT 2019.560 483.070 2020.220 483.130 ;
        RECT 2019.960 482.810 2020.220 483.070 ;
        RECT 2018.640 435.190 2018.780 482.810 ;
        RECT 2020.020 482.655 2020.160 482.810 ;
        RECT 2018.580 434.870 2018.840 435.190 ;
        RECT 2019.500 434.870 2019.760 435.190 ;
        RECT 2019.560 434.510 2019.700 434.870 ;
        RECT 2019.500 434.190 2019.760 434.510 ;
        RECT 2019.960 434.190 2020.220 434.510 ;
        RECT 2020.020 356.050 2020.160 434.190 ;
        RECT 2019.100 355.910 2020.160 356.050 ;
        RECT 2019.100 331.490 2019.240 355.910 ;
        RECT 2019.040 331.170 2019.300 331.490 ;
        RECT 2020.420 331.170 2020.680 331.490 ;
        RECT 2020.480 330.890 2020.620 331.170 ;
        RECT 2020.480 330.750 2021.080 330.890 ;
        RECT 2020.940 303.010 2021.080 330.750 ;
        RECT 2020.020 302.870 2021.080 303.010 ;
        RECT 2020.020 282.870 2020.160 302.870 ;
        RECT 2019.040 282.550 2019.300 282.870 ;
        RECT 2019.960 282.550 2020.220 282.870 ;
        RECT 2019.100 234.930 2019.240 282.550 ;
        RECT 2019.040 234.610 2019.300 234.930 ;
        RECT 2020.420 234.610 2020.680 234.930 ;
        RECT 2020.480 218.010 2020.620 234.610 ;
        RECT 2020.020 217.870 2020.620 218.010 ;
        RECT 2020.020 210.530 2020.160 217.870 ;
        RECT 2020.020 210.390 2020.620 210.530 ;
        RECT 2020.480 159.110 2020.620 210.390 ;
        RECT 2020.420 158.790 2020.680 159.110 ;
        RECT 2020.420 158.110 2020.680 158.430 ;
        RECT 2020.480 109.890 2020.620 158.110 ;
        RECT 2020.480 109.750 2021.080 109.890 ;
        RECT 2020.940 31.610 2021.080 109.750 ;
        RECT 2020.880 31.290 2021.140 31.610 ;
        RECT 2619.340 31.290 2619.600 31.610 ;
        RECT 2619.400 2.400 2619.540 31.290 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2027.750 30.840 2028.070 30.900 ;
        RECT 2637.250 30.840 2637.570 30.900 ;
        RECT 2027.750 30.700 2637.570 30.840 ;
        RECT 2027.750 30.640 2028.070 30.700 ;
        RECT 2637.250 30.640 2637.570 30.700 ;
      LAYER via ;
        RECT 2027.780 30.640 2028.040 30.900 ;
        RECT 2637.280 30.640 2637.540 30.900 ;
      LAYER met2 ;
        RECT 2027.550 600.000 2027.830 604.000 ;
        RECT 2027.610 598.810 2027.750 600.000 ;
        RECT 2027.610 598.670 2027.980 598.810 ;
        RECT 2027.840 30.930 2027.980 598.670 ;
        RECT 2027.780 30.610 2028.040 30.930 ;
        RECT 2637.280 30.610 2637.540 30.930 ;
        RECT 2637.340 2.400 2637.480 30.610 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2038.330 586.740 2038.650 586.800 ;
        RECT 2042.010 586.740 2042.330 586.800 ;
        RECT 2038.330 586.600 2042.330 586.740 ;
        RECT 2038.330 586.540 2038.650 586.600 ;
        RECT 2042.010 586.540 2042.330 586.600 ;
        RECT 2042.010 31.180 2042.330 31.240 ;
        RECT 2655.190 31.180 2655.510 31.240 ;
        RECT 2042.010 31.040 2655.510 31.180 ;
        RECT 2042.010 30.980 2042.330 31.040 ;
        RECT 2655.190 30.980 2655.510 31.040 ;
      LAYER via ;
        RECT 2038.360 586.540 2038.620 586.800 ;
        RECT 2042.040 586.540 2042.300 586.800 ;
        RECT 2042.040 30.980 2042.300 31.240 ;
        RECT 2655.220 30.980 2655.480 31.240 ;
      LAYER met2 ;
        RECT 2036.750 600.170 2037.030 604.000 ;
        RECT 2036.750 600.030 2038.560 600.170 ;
        RECT 2036.750 600.000 2037.030 600.030 ;
        RECT 2038.420 586.830 2038.560 600.030 ;
        RECT 2038.360 586.510 2038.620 586.830 ;
        RECT 2042.040 586.510 2042.300 586.830 ;
        RECT 2042.100 31.270 2042.240 586.510 ;
        RECT 2042.040 30.950 2042.300 31.270 ;
        RECT 2655.220 30.950 2655.480 31.270 ;
        RECT 2655.280 2.400 2655.420 30.950 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2046.610 573.140 2046.930 573.200 ;
        RECT 2047.990 573.140 2048.310 573.200 ;
        RECT 2046.610 573.000 2048.310 573.140 ;
        RECT 2046.610 572.940 2046.930 573.000 ;
        RECT 2047.990 572.940 2048.310 573.000 ;
        RECT 2047.070 572.460 2047.390 572.520 ;
        RECT 2047.990 572.460 2048.310 572.520 ;
        RECT 2047.070 572.320 2048.310 572.460 ;
        RECT 2047.070 572.260 2047.390 572.320 ;
        RECT 2047.990 572.260 2048.310 572.320 ;
        RECT 2046.610 524.520 2046.930 524.580 ;
        RECT 2047.070 524.520 2047.390 524.580 ;
        RECT 2046.610 524.380 2047.390 524.520 ;
        RECT 2046.610 524.320 2046.930 524.380 ;
        RECT 2047.070 524.320 2047.390 524.380 ;
        RECT 2046.610 476.240 2046.930 476.300 ;
        RECT 2047.990 476.240 2048.310 476.300 ;
        RECT 2046.610 476.100 2048.310 476.240 ;
        RECT 2046.610 476.040 2046.930 476.100 ;
        RECT 2047.990 476.040 2048.310 476.100 ;
        RECT 2047.530 448.700 2047.850 448.760 ;
        RECT 2047.530 448.560 2048.220 448.700 ;
        RECT 2047.530 448.500 2047.850 448.560 ;
        RECT 2048.080 448.420 2048.220 448.560 ;
        RECT 2047.990 448.160 2048.310 448.420 ;
        RECT 2047.530 338.200 2047.850 338.260 ;
        RECT 2047.990 338.200 2048.310 338.260 ;
        RECT 2047.530 338.060 2048.310 338.200 ;
        RECT 2047.530 338.000 2047.850 338.060 ;
        RECT 2047.990 338.000 2048.310 338.060 ;
        RECT 2047.070 331.060 2047.390 331.120 ;
        RECT 2047.530 331.060 2047.850 331.120 ;
        RECT 2047.070 330.920 2047.850 331.060 ;
        RECT 2047.070 330.860 2047.390 330.920 ;
        RECT 2047.530 330.860 2047.850 330.920 ;
        RECT 2046.610 283.120 2046.930 283.180 ;
        RECT 2047.070 283.120 2047.390 283.180 ;
        RECT 2046.610 282.980 2047.390 283.120 ;
        RECT 2046.610 282.920 2046.930 282.980 ;
        RECT 2047.070 282.920 2047.390 282.980 ;
        RECT 2046.610 255.240 2046.930 255.300 ;
        RECT 2047.530 255.240 2047.850 255.300 ;
        RECT 2046.610 255.100 2047.850 255.240 ;
        RECT 2046.610 255.040 2046.930 255.100 ;
        RECT 2047.530 255.040 2047.850 255.100 ;
        RECT 2046.610 193.020 2046.930 193.080 ;
        RECT 2047.990 193.020 2048.310 193.080 ;
        RECT 2046.610 192.880 2048.310 193.020 ;
        RECT 2046.610 192.820 2046.930 192.880 ;
        RECT 2047.990 192.820 2048.310 192.880 ;
        RECT 2046.610 145.080 2046.930 145.140 ;
        RECT 2047.070 145.080 2047.390 145.140 ;
        RECT 2046.610 144.940 2047.390 145.080 ;
        RECT 2046.610 144.880 2046.930 144.940 ;
        RECT 2047.070 144.880 2047.390 144.940 ;
        RECT 2047.070 96.800 2047.390 96.860 ;
        RECT 2047.990 96.800 2048.310 96.860 ;
        RECT 2047.070 96.660 2048.310 96.800 ;
        RECT 2047.070 96.600 2047.390 96.660 ;
        RECT 2047.990 96.600 2048.310 96.660 ;
        RECT 2047.990 40.700 2048.310 40.760 ;
        RECT 2672.670 40.700 2672.990 40.760 ;
        RECT 2047.990 40.560 2672.990 40.700 ;
        RECT 2047.990 40.500 2048.310 40.560 ;
        RECT 2672.670 40.500 2672.990 40.560 ;
      LAYER via ;
        RECT 2046.640 572.940 2046.900 573.200 ;
        RECT 2048.020 572.940 2048.280 573.200 ;
        RECT 2047.100 572.260 2047.360 572.520 ;
        RECT 2048.020 572.260 2048.280 572.520 ;
        RECT 2046.640 524.320 2046.900 524.580 ;
        RECT 2047.100 524.320 2047.360 524.580 ;
        RECT 2046.640 476.040 2046.900 476.300 ;
        RECT 2048.020 476.040 2048.280 476.300 ;
        RECT 2047.560 448.500 2047.820 448.760 ;
        RECT 2048.020 448.160 2048.280 448.420 ;
        RECT 2047.560 338.000 2047.820 338.260 ;
        RECT 2048.020 338.000 2048.280 338.260 ;
        RECT 2047.100 330.860 2047.360 331.120 ;
        RECT 2047.560 330.860 2047.820 331.120 ;
        RECT 2046.640 282.920 2046.900 283.180 ;
        RECT 2047.100 282.920 2047.360 283.180 ;
        RECT 2046.640 255.040 2046.900 255.300 ;
        RECT 2047.560 255.040 2047.820 255.300 ;
        RECT 2046.640 192.820 2046.900 193.080 ;
        RECT 2048.020 192.820 2048.280 193.080 ;
        RECT 2046.640 144.880 2046.900 145.140 ;
        RECT 2047.100 144.880 2047.360 145.140 ;
        RECT 2047.100 96.600 2047.360 96.860 ;
        RECT 2048.020 96.600 2048.280 96.860 ;
        RECT 2048.020 40.500 2048.280 40.760 ;
        RECT 2672.700 40.500 2672.960 40.760 ;
      LAYER met2 ;
        RECT 2045.950 600.170 2046.230 604.000 ;
        RECT 2045.950 600.030 2046.840 600.170 ;
        RECT 2045.950 600.000 2046.230 600.030 ;
        RECT 2046.700 573.230 2046.840 600.030 ;
        RECT 2046.640 572.910 2046.900 573.230 ;
        RECT 2048.020 572.910 2048.280 573.230 ;
        RECT 2048.080 572.550 2048.220 572.910 ;
        RECT 2047.100 572.230 2047.360 572.550 ;
        RECT 2048.020 572.230 2048.280 572.550 ;
        RECT 2047.160 524.610 2047.300 572.230 ;
        RECT 2046.640 524.290 2046.900 524.610 ;
        RECT 2047.100 524.290 2047.360 524.610 ;
        RECT 2046.700 476.330 2046.840 524.290 ;
        RECT 2046.640 476.010 2046.900 476.330 ;
        RECT 2048.020 476.010 2048.280 476.330 ;
        RECT 2048.080 475.730 2048.220 476.010 ;
        RECT 2047.620 475.590 2048.220 475.730 ;
        RECT 2047.620 448.790 2047.760 475.590 ;
        RECT 2047.560 448.470 2047.820 448.790 ;
        RECT 2048.020 448.130 2048.280 448.450 ;
        RECT 2048.080 338.290 2048.220 448.130 ;
        RECT 2047.560 337.970 2047.820 338.290 ;
        RECT 2048.020 337.970 2048.280 338.290 ;
        RECT 2047.620 331.150 2047.760 337.970 ;
        RECT 2047.100 330.830 2047.360 331.150 ;
        RECT 2047.560 330.830 2047.820 331.150 ;
        RECT 2047.160 283.210 2047.300 330.830 ;
        RECT 2046.640 282.890 2046.900 283.210 ;
        RECT 2047.100 282.890 2047.360 283.210 ;
        RECT 2046.700 255.330 2046.840 282.890 ;
        RECT 2046.640 255.010 2046.900 255.330 ;
        RECT 2047.560 255.010 2047.820 255.330 ;
        RECT 2047.620 206.450 2047.760 255.010 ;
        RECT 2047.620 206.310 2048.220 206.450 ;
        RECT 2048.080 193.110 2048.220 206.310 ;
        RECT 2046.640 192.790 2046.900 193.110 ;
        RECT 2048.020 192.790 2048.280 193.110 ;
        RECT 2046.700 145.170 2046.840 192.790 ;
        RECT 2046.640 144.850 2046.900 145.170 ;
        RECT 2047.100 144.850 2047.360 145.170 ;
        RECT 2047.160 96.890 2047.300 144.850 ;
        RECT 2047.100 96.570 2047.360 96.890 ;
        RECT 2048.020 96.570 2048.280 96.890 ;
        RECT 2048.080 40.790 2048.220 96.570 ;
        RECT 2048.020 40.470 2048.280 40.790 ;
        RECT 2672.700 40.470 2672.960 40.790 ;
        RECT 2672.760 2.400 2672.900 40.470 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2055.350 40.360 2055.670 40.420 ;
        RECT 2690.610 40.360 2690.930 40.420 ;
        RECT 2055.350 40.220 2690.930 40.360 ;
        RECT 2055.350 40.160 2055.670 40.220 ;
        RECT 2690.610 40.160 2690.930 40.220 ;
      LAYER via ;
        RECT 2055.380 40.160 2055.640 40.420 ;
        RECT 2690.640 40.160 2690.900 40.420 ;
      LAYER met2 ;
        RECT 2055.150 600.000 2055.430 604.000 ;
        RECT 2055.210 598.810 2055.350 600.000 ;
        RECT 2055.210 598.670 2055.580 598.810 ;
        RECT 2055.440 40.450 2055.580 598.670 ;
        RECT 2055.380 40.130 2055.640 40.450 ;
        RECT 2690.640 40.130 2690.900 40.450 ;
        RECT 2690.700 2.400 2690.840 40.130 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2065.930 586.740 2066.250 586.800 ;
        RECT 2069.610 586.740 2069.930 586.800 ;
        RECT 2065.930 586.600 2069.930 586.740 ;
        RECT 2065.930 586.540 2066.250 586.600 ;
        RECT 2069.610 586.540 2069.930 586.600 ;
        RECT 2069.610 40.020 2069.930 40.080 ;
        RECT 2708.550 40.020 2708.870 40.080 ;
        RECT 2069.610 39.880 2708.870 40.020 ;
        RECT 2069.610 39.820 2069.930 39.880 ;
        RECT 2708.550 39.820 2708.870 39.880 ;
      LAYER via ;
        RECT 2065.960 586.540 2066.220 586.800 ;
        RECT 2069.640 586.540 2069.900 586.800 ;
        RECT 2069.640 39.820 2069.900 40.080 ;
        RECT 2708.580 39.820 2708.840 40.080 ;
      LAYER met2 ;
        RECT 2064.350 600.170 2064.630 604.000 ;
        RECT 2064.350 600.030 2066.160 600.170 ;
        RECT 2064.350 600.000 2064.630 600.030 ;
        RECT 2066.020 586.830 2066.160 600.030 ;
        RECT 2065.960 586.510 2066.220 586.830 ;
        RECT 2069.640 586.510 2069.900 586.830 ;
        RECT 2069.700 40.110 2069.840 586.510 ;
        RECT 2069.640 39.790 2069.900 40.110 ;
        RECT 2708.580 39.790 2708.840 40.110 ;
        RECT 2708.640 2.400 2708.780 39.790 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2073.750 566.000 2074.070 566.060 ;
        RECT 2076.050 566.000 2076.370 566.060 ;
        RECT 2073.750 565.860 2076.370 566.000 ;
        RECT 2073.750 565.800 2074.070 565.860 ;
        RECT 2076.050 565.800 2076.370 565.860 ;
        RECT 2076.050 531.460 2076.370 531.720 ;
        RECT 2076.140 531.040 2076.280 531.460 ;
        RECT 2076.050 530.780 2076.370 531.040 ;
        RECT 2074.670 517.380 2074.990 517.440 ;
        RECT 2075.590 517.380 2075.910 517.440 ;
        RECT 2074.670 517.240 2075.910 517.380 ;
        RECT 2074.670 517.180 2074.990 517.240 ;
        RECT 2075.590 517.180 2075.910 517.240 ;
        RECT 2075.590 448.500 2075.910 448.760 ;
        RECT 2075.680 448.080 2075.820 448.500 ;
        RECT 2075.590 447.820 2075.910 448.080 ;
        RECT 2075.130 420.820 2075.450 420.880 ;
        RECT 2075.590 420.820 2075.910 420.880 ;
        RECT 2075.130 420.680 2075.910 420.820 ;
        RECT 2075.130 420.620 2075.450 420.680 ;
        RECT 2075.590 420.620 2075.910 420.680 ;
        RECT 2074.670 372.880 2074.990 372.940 ;
        RECT 2075.130 372.880 2075.450 372.940 ;
        RECT 2074.670 372.740 2075.450 372.880 ;
        RECT 2074.670 372.680 2074.990 372.740 ;
        RECT 2075.130 372.680 2075.450 372.740 ;
        RECT 2073.750 331.060 2074.070 331.120 ;
        RECT 2074.670 331.060 2074.990 331.120 ;
        RECT 2073.750 330.920 2074.990 331.060 ;
        RECT 2073.750 330.860 2074.070 330.920 ;
        RECT 2074.670 330.860 2074.990 330.920 ;
        RECT 2073.750 283.120 2074.070 283.180 ;
        RECT 2076.050 283.120 2076.370 283.180 ;
        RECT 2073.750 282.980 2076.370 283.120 ;
        RECT 2073.750 282.920 2074.070 282.980 ;
        RECT 2076.050 282.920 2076.370 282.980 ;
        RECT 2074.670 241.640 2074.990 241.700 ;
        RECT 2076.050 241.640 2076.370 241.700 ;
        RECT 2074.670 241.500 2076.370 241.640 ;
        RECT 2074.670 241.440 2074.990 241.500 ;
        RECT 2076.050 241.440 2076.370 241.500 ;
        RECT 2075.590 158.820 2075.910 159.080 ;
        RECT 2075.130 158.680 2075.450 158.740 ;
        RECT 2075.680 158.680 2075.820 158.820 ;
        RECT 2075.130 158.540 2075.820 158.680 ;
        RECT 2075.130 158.480 2075.450 158.540 ;
        RECT 2075.130 145.080 2075.450 145.140 ;
        RECT 2076.050 145.080 2076.370 145.140 ;
        RECT 2075.130 144.940 2076.370 145.080 ;
        RECT 2075.130 144.880 2075.450 144.940 ;
        RECT 2076.050 144.880 2076.370 144.940 ;
        RECT 2075.590 39.680 2075.910 39.740 ;
        RECT 2726.490 39.680 2726.810 39.740 ;
        RECT 2075.590 39.540 2726.810 39.680 ;
        RECT 2075.590 39.480 2075.910 39.540 ;
        RECT 2726.490 39.480 2726.810 39.540 ;
      LAYER via ;
        RECT 2073.780 565.800 2074.040 566.060 ;
        RECT 2076.080 565.800 2076.340 566.060 ;
        RECT 2076.080 531.460 2076.340 531.720 ;
        RECT 2076.080 530.780 2076.340 531.040 ;
        RECT 2074.700 517.180 2074.960 517.440 ;
        RECT 2075.620 517.180 2075.880 517.440 ;
        RECT 2075.620 448.500 2075.880 448.760 ;
        RECT 2075.620 447.820 2075.880 448.080 ;
        RECT 2075.160 420.620 2075.420 420.880 ;
        RECT 2075.620 420.620 2075.880 420.880 ;
        RECT 2074.700 372.680 2074.960 372.940 ;
        RECT 2075.160 372.680 2075.420 372.940 ;
        RECT 2073.780 330.860 2074.040 331.120 ;
        RECT 2074.700 330.860 2074.960 331.120 ;
        RECT 2073.780 282.920 2074.040 283.180 ;
        RECT 2076.080 282.920 2076.340 283.180 ;
        RECT 2074.700 241.440 2074.960 241.700 ;
        RECT 2076.080 241.440 2076.340 241.700 ;
        RECT 2075.620 158.820 2075.880 159.080 ;
        RECT 2075.160 158.480 2075.420 158.740 ;
        RECT 2075.160 144.880 2075.420 145.140 ;
        RECT 2076.080 144.880 2076.340 145.140 ;
        RECT 2075.620 39.480 2075.880 39.740 ;
        RECT 2726.520 39.480 2726.780 39.740 ;
      LAYER met2 ;
        RECT 2073.550 600.000 2073.830 604.000 ;
        RECT 2073.610 598.810 2073.750 600.000 ;
        RECT 2073.610 598.670 2073.980 598.810 ;
        RECT 2073.840 566.090 2073.980 598.670 ;
        RECT 2073.780 565.770 2074.040 566.090 ;
        RECT 2076.080 565.770 2076.340 566.090 ;
        RECT 2076.140 531.750 2076.280 565.770 ;
        RECT 2076.080 531.430 2076.340 531.750 ;
        RECT 2076.080 530.750 2076.340 531.070 ;
        RECT 2076.140 524.010 2076.280 530.750 ;
        RECT 2075.680 523.870 2076.280 524.010 ;
        RECT 2075.680 517.470 2075.820 523.870 ;
        RECT 2074.700 517.150 2074.960 517.470 ;
        RECT 2075.620 517.150 2075.880 517.470 ;
        RECT 2074.760 473.010 2074.900 517.150 ;
        RECT 2074.760 472.870 2075.820 473.010 ;
        RECT 2075.680 448.790 2075.820 472.870 ;
        RECT 2075.620 448.470 2075.880 448.790 ;
        RECT 2075.620 447.790 2075.880 448.110 ;
        RECT 2075.680 420.910 2075.820 447.790 ;
        RECT 2075.160 420.590 2075.420 420.910 ;
        RECT 2075.620 420.590 2075.880 420.910 ;
        RECT 2075.220 372.970 2075.360 420.590 ;
        RECT 2074.700 372.650 2074.960 372.970 ;
        RECT 2075.160 372.650 2075.420 372.970 ;
        RECT 2074.760 331.150 2074.900 372.650 ;
        RECT 2073.780 330.830 2074.040 331.150 ;
        RECT 2074.700 330.830 2074.960 331.150 ;
        RECT 2073.840 283.210 2073.980 330.830 ;
        RECT 2073.780 282.890 2074.040 283.210 ;
        RECT 2076.080 282.890 2076.340 283.210 ;
        RECT 2076.140 241.730 2076.280 282.890 ;
        RECT 2074.700 241.410 2074.960 241.730 ;
        RECT 2076.080 241.410 2076.340 241.730 ;
        RECT 2074.760 217.330 2074.900 241.410 ;
        RECT 2074.760 217.190 2075.820 217.330 ;
        RECT 2075.680 159.110 2075.820 217.190 ;
        RECT 2075.620 158.790 2075.880 159.110 ;
        RECT 2075.160 158.450 2075.420 158.770 ;
        RECT 2075.220 145.170 2075.360 158.450 ;
        RECT 2075.160 144.850 2075.420 145.170 ;
        RECT 2076.080 144.850 2076.340 145.170 ;
        RECT 2076.140 62.290 2076.280 144.850 ;
        RECT 2075.680 62.150 2076.280 62.290 ;
        RECT 2075.680 39.770 2075.820 62.150 ;
        RECT 2075.620 39.450 2075.880 39.770 ;
        RECT 2726.520 39.450 2726.780 39.770 ;
        RECT 2726.580 2.400 2726.720 39.450 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2082.950 39.340 2083.270 39.400 ;
        RECT 2744.430 39.340 2744.750 39.400 ;
        RECT 2082.950 39.200 2744.750 39.340 ;
        RECT 2082.950 39.140 2083.270 39.200 ;
        RECT 2744.430 39.140 2744.750 39.200 ;
      LAYER via ;
        RECT 2082.980 39.140 2083.240 39.400 ;
        RECT 2744.460 39.140 2744.720 39.400 ;
      LAYER met2 ;
        RECT 2082.750 600.000 2083.030 604.000 ;
        RECT 2082.810 598.810 2082.950 600.000 ;
        RECT 2082.810 598.670 2083.180 598.810 ;
        RECT 2083.040 39.430 2083.180 598.670 ;
        RECT 2082.980 39.110 2083.240 39.430 ;
        RECT 2744.460 39.110 2744.720 39.430 ;
        RECT 2744.520 2.400 2744.660 39.110 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2093.070 586.740 2093.390 586.800 ;
        RECT 2097.210 586.740 2097.530 586.800 ;
        RECT 2093.070 586.600 2097.530 586.740 ;
        RECT 2093.070 586.540 2093.390 586.600 ;
        RECT 2097.210 586.540 2097.530 586.600 ;
        RECT 2097.210 39.000 2097.530 39.060 ;
        RECT 2761.910 39.000 2762.230 39.060 ;
        RECT 2097.210 38.860 2762.230 39.000 ;
        RECT 2097.210 38.800 2097.530 38.860 ;
        RECT 2761.910 38.800 2762.230 38.860 ;
      LAYER via ;
        RECT 2093.100 586.540 2093.360 586.800 ;
        RECT 2097.240 586.540 2097.500 586.800 ;
        RECT 2097.240 38.800 2097.500 39.060 ;
        RECT 2761.940 38.800 2762.200 39.060 ;
      LAYER met2 ;
        RECT 2091.490 600.170 2091.770 604.000 ;
        RECT 2091.490 600.030 2093.300 600.170 ;
        RECT 2091.490 600.000 2091.770 600.030 ;
        RECT 2093.160 586.830 2093.300 600.030 ;
        RECT 2093.100 586.510 2093.360 586.830 ;
        RECT 2097.240 586.510 2097.500 586.830 ;
        RECT 2097.300 39.090 2097.440 586.510 ;
        RECT 2097.240 38.770 2097.500 39.090 ;
        RECT 2761.940 38.770 2762.200 39.090 ;
        RECT 2762.000 2.400 2762.140 38.770 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 835.430 25.400 835.750 25.460 ;
        RECT 1097.630 25.400 1097.950 25.460 ;
        RECT 835.430 25.260 1097.950 25.400 ;
        RECT 835.430 25.200 835.750 25.260 ;
        RECT 1097.630 25.200 1097.950 25.260 ;
      LAYER via ;
        RECT 835.460 25.200 835.720 25.460 ;
        RECT 1097.660 25.200 1097.920 25.460 ;
      LAYER met2 ;
        RECT 1099.730 600.170 1100.010 604.000 ;
        RECT 1097.720 600.030 1100.010 600.170 ;
        RECT 1097.720 25.490 1097.860 600.030 ;
        RECT 1099.730 600.000 1100.010 600.030 ;
        RECT 835.460 25.170 835.720 25.490 ;
        RECT 1097.660 25.170 1097.920 25.490 ;
        RECT 835.520 2.400 835.660 25.170 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2101.350 579.940 2101.670 580.000 ;
        RECT 2102.270 579.940 2102.590 580.000 ;
        RECT 2101.350 579.800 2102.590 579.940 ;
        RECT 2101.350 579.740 2101.670 579.800 ;
        RECT 2102.270 579.740 2102.590 579.800 ;
        RECT 2102.730 524.180 2103.050 524.240 ;
        RECT 2103.190 524.180 2103.510 524.240 ;
        RECT 2102.730 524.040 2103.510 524.180 ;
        RECT 2102.730 523.980 2103.050 524.040 ;
        RECT 2103.190 523.980 2103.510 524.040 ;
        RECT 2102.730 476.240 2103.050 476.300 ;
        RECT 2103.650 476.240 2103.970 476.300 ;
        RECT 2102.730 476.100 2103.970 476.240 ;
        RECT 2102.730 476.040 2103.050 476.100 ;
        RECT 2103.650 476.040 2103.970 476.100 ;
        RECT 2102.730 434.760 2103.050 434.820 ;
        RECT 2103.190 434.760 2103.510 434.820 ;
        RECT 2102.730 434.620 2103.510 434.760 ;
        RECT 2102.730 434.560 2103.050 434.620 ;
        RECT 2103.190 434.560 2103.510 434.620 ;
        RECT 2102.730 386.820 2103.050 386.880 ;
        RECT 2103.650 386.820 2103.970 386.880 ;
        RECT 2102.730 386.680 2103.970 386.820 ;
        RECT 2102.730 386.620 2103.050 386.680 ;
        RECT 2103.650 386.620 2103.970 386.680 ;
        RECT 2103.190 338.200 2103.510 338.260 ;
        RECT 2105.030 338.200 2105.350 338.260 ;
        RECT 2103.190 338.060 2105.350 338.200 ;
        RECT 2103.190 338.000 2103.510 338.060 ;
        RECT 2105.030 338.000 2105.350 338.060 ;
        RECT 2103.650 303.860 2103.970 303.920 ;
        RECT 2103.280 303.720 2103.970 303.860 ;
        RECT 2103.280 303.580 2103.420 303.720 ;
        RECT 2103.650 303.660 2103.970 303.720 ;
        RECT 2103.190 303.320 2103.510 303.580 ;
        RECT 2102.270 289.580 2102.590 289.640 ;
        RECT 2103.650 289.580 2103.970 289.640 ;
        RECT 2102.270 289.440 2103.970 289.580 ;
        RECT 2102.270 289.380 2102.590 289.440 ;
        RECT 2103.650 289.380 2103.970 289.440 ;
        RECT 2102.730 241.300 2103.050 241.360 ;
        RECT 2103.190 241.300 2103.510 241.360 ;
        RECT 2102.730 241.160 2103.510 241.300 ;
        RECT 2102.730 241.100 2103.050 241.160 ;
        RECT 2103.190 241.100 2103.510 241.160 ;
        RECT 2102.270 169.220 2102.590 169.280 ;
        RECT 2103.190 169.220 2103.510 169.280 ;
        RECT 2102.270 169.080 2103.510 169.220 ;
        RECT 2102.270 169.020 2102.590 169.080 ;
        RECT 2103.190 169.020 2103.510 169.080 ;
        RECT 2102.730 144.740 2103.050 144.800 ;
        RECT 2103.190 144.740 2103.510 144.800 ;
        RECT 2102.730 144.600 2103.510 144.740 ;
        RECT 2102.730 144.540 2103.050 144.600 ;
        RECT 2103.190 144.540 2103.510 144.600 ;
        RECT 2102.270 72.660 2102.590 72.720 ;
        RECT 2103.190 72.660 2103.510 72.720 ;
        RECT 2102.270 72.520 2103.510 72.660 ;
        RECT 2102.270 72.460 2102.590 72.520 ;
        RECT 2103.190 72.460 2103.510 72.520 ;
        RECT 2102.270 48.520 2102.590 48.580 ;
        RECT 2103.190 48.520 2103.510 48.580 ;
        RECT 2102.270 48.380 2103.510 48.520 ;
        RECT 2102.270 48.320 2102.590 48.380 ;
        RECT 2103.190 48.320 2103.510 48.380 ;
        RECT 2103.190 38.660 2103.510 38.720 ;
        RECT 2779.850 38.660 2780.170 38.720 ;
        RECT 2103.190 38.520 2780.170 38.660 ;
        RECT 2103.190 38.460 2103.510 38.520 ;
        RECT 2779.850 38.460 2780.170 38.520 ;
      LAYER via ;
        RECT 2101.380 579.740 2101.640 580.000 ;
        RECT 2102.300 579.740 2102.560 580.000 ;
        RECT 2102.760 523.980 2103.020 524.240 ;
        RECT 2103.220 523.980 2103.480 524.240 ;
        RECT 2102.760 476.040 2103.020 476.300 ;
        RECT 2103.680 476.040 2103.940 476.300 ;
        RECT 2102.760 434.560 2103.020 434.820 ;
        RECT 2103.220 434.560 2103.480 434.820 ;
        RECT 2102.760 386.620 2103.020 386.880 ;
        RECT 2103.680 386.620 2103.940 386.880 ;
        RECT 2103.220 338.000 2103.480 338.260 ;
        RECT 2105.060 338.000 2105.320 338.260 ;
        RECT 2103.680 303.660 2103.940 303.920 ;
        RECT 2103.220 303.320 2103.480 303.580 ;
        RECT 2102.300 289.380 2102.560 289.640 ;
        RECT 2103.680 289.380 2103.940 289.640 ;
        RECT 2102.760 241.100 2103.020 241.360 ;
        RECT 2103.220 241.100 2103.480 241.360 ;
        RECT 2102.300 169.020 2102.560 169.280 ;
        RECT 2103.220 169.020 2103.480 169.280 ;
        RECT 2102.760 144.540 2103.020 144.800 ;
        RECT 2103.220 144.540 2103.480 144.800 ;
        RECT 2102.300 72.460 2102.560 72.720 ;
        RECT 2103.220 72.460 2103.480 72.720 ;
        RECT 2102.300 48.320 2102.560 48.580 ;
        RECT 2103.220 48.320 2103.480 48.580 ;
        RECT 2103.220 38.460 2103.480 38.720 ;
        RECT 2779.880 38.460 2780.140 38.720 ;
      LAYER met2 ;
        RECT 2100.690 600.170 2100.970 604.000 ;
        RECT 2100.690 600.030 2101.580 600.170 ;
        RECT 2100.690 600.000 2100.970 600.030 ;
        RECT 2101.440 580.030 2101.580 600.030 ;
        RECT 2101.380 579.710 2101.640 580.030 ;
        RECT 2102.300 579.710 2102.560 580.030 ;
        RECT 2102.360 545.090 2102.500 579.710 ;
        RECT 2102.360 544.950 2103.420 545.090 ;
        RECT 2103.280 524.270 2103.420 544.950 ;
        RECT 2102.760 523.950 2103.020 524.270 ;
        RECT 2103.220 523.950 2103.480 524.270 ;
        RECT 2102.820 476.330 2102.960 523.950 ;
        RECT 2102.760 476.010 2103.020 476.330 ;
        RECT 2103.680 476.010 2103.940 476.330 ;
        RECT 2103.740 434.930 2103.880 476.010 ;
        RECT 2103.280 434.850 2103.880 434.930 ;
        RECT 2102.760 434.530 2103.020 434.850 ;
        RECT 2103.220 434.790 2103.880 434.850 ;
        RECT 2103.220 434.530 2103.480 434.790 ;
        RECT 2102.820 386.910 2102.960 434.530 ;
        RECT 2102.760 386.590 2103.020 386.910 ;
        RECT 2103.680 386.590 2103.940 386.910 ;
        RECT 2103.740 386.085 2103.880 386.590 ;
        RECT 2103.670 385.715 2103.950 386.085 ;
        RECT 2105.050 385.715 2105.330 386.085 ;
        RECT 2105.120 338.290 2105.260 385.715 ;
        RECT 2103.220 337.970 2103.480 338.290 ;
        RECT 2105.060 337.970 2105.320 338.290 ;
        RECT 2103.280 337.690 2103.420 337.970 ;
        RECT 2103.280 337.550 2103.880 337.690 ;
        RECT 2103.740 303.950 2103.880 337.550 ;
        RECT 2103.680 303.630 2103.940 303.950 ;
        RECT 2103.220 303.290 2103.480 303.610 ;
        RECT 2103.280 290.090 2103.420 303.290 ;
        RECT 2103.280 289.950 2103.880 290.090 ;
        RECT 2103.740 289.670 2103.880 289.950 ;
        RECT 2102.300 289.350 2102.560 289.670 ;
        RECT 2103.680 289.350 2103.940 289.670 ;
        RECT 2102.360 241.925 2102.500 289.350 ;
        RECT 2102.290 241.555 2102.570 241.925 ;
        RECT 2103.210 241.555 2103.490 241.925 ;
        RECT 2103.280 241.390 2103.420 241.555 ;
        RECT 2102.760 241.070 2103.020 241.390 ;
        RECT 2103.220 241.070 2103.480 241.390 ;
        RECT 2102.820 206.450 2102.960 241.070 ;
        RECT 2102.820 206.310 2103.420 206.450 ;
        RECT 2103.280 169.310 2103.420 206.310 ;
        RECT 2102.300 168.990 2102.560 169.310 ;
        RECT 2103.220 168.990 2103.480 169.310 ;
        RECT 2102.360 145.365 2102.500 168.990 ;
        RECT 2102.290 144.995 2102.570 145.365 ;
        RECT 2102.760 144.510 2103.020 144.830 ;
        RECT 2103.210 144.825 2103.490 145.195 ;
        RECT 2103.220 144.510 2103.480 144.825 ;
        RECT 2102.820 109.890 2102.960 144.510 ;
        RECT 2102.820 109.750 2103.420 109.890 ;
        RECT 2103.280 72.750 2103.420 109.750 ;
        RECT 2102.300 72.430 2102.560 72.750 ;
        RECT 2103.220 72.430 2103.480 72.750 ;
        RECT 2102.360 48.610 2102.500 72.430 ;
        RECT 2102.300 48.290 2102.560 48.610 ;
        RECT 2103.220 48.290 2103.480 48.610 ;
        RECT 2103.280 38.750 2103.420 48.290 ;
        RECT 2103.220 38.430 2103.480 38.750 ;
        RECT 2779.880 38.430 2780.140 38.750 ;
        RECT 2779.940 2.400 2780.080 38.430 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
      LAYER via2 ;
        RECT 2103.670 385.760 2103.950 386.040 ;
        RECT 2105.050 385.760 2105.330 386.040 ;
        RECT 2102.290 241.600 2102.570 241.880 ;
        RECT 2103.210 241.600 2103.490 241.880 ;
        RECT 2102.290 145.040 2102.570 145.320 ;
        RECT 2103.210 144.870 2103.490 145.150 ;
      LAYER met3 ;
        RECT 2103.645 386.050 2103.975 386.065 ;
        RECT 2105.025 386.050 2105.355 386.065 ;
        RECT 2103.645 385.750 2105.355 386.050 ;
        RECT 2103.645 385.735 2103.975 385.750 ;
        RECT 2105.025 385.735 2105.355 385.750 ;
        RECT 2102.265 241.890 2102.595 241.905 ;
        RECT 2103.185 241.890 2103.515 241.905 ;
        RECT 2102.265 241.590 2103.515 241.890 ;
        RECT 2102.265 241.575 2102.595 241.590 ;
        RECT 2103.185 241.575 2103.515 241.590 ;
        RECT 2102.265 145.330 2102.595 145.345 ;
        RECT 2102.265 145.160 2102.810 145.330 ;
        RECT 2103.185 145.160 2103.515 145.175 ;
        RECT 2102.265 145.015 2103.515 145.160 ;
        RECT 2102.510 144.860 2103.515 145.015 ;
        RECT 2103.185 144.845 2103.515 144.860 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2110.550 38.320 2110.870 38.380 ;
        RECT 2797.790 38.320 2798.110 38.380 ;
        RECT 2110.550 38.180 2798.110 38.320 ;
        RECT 2110.550 38.120 2110.870 38.180 ;
        RECT 2797.790 38.120 2798.110 38.180 ;
      LAYER via ;
        RECT 2110.580 38.120 2110.840 38.380 ;
        RECT 2797.820 38.120 2798.080 38.380 ;
      LAYER met2 ;
        RECT 2109.890 600.170 2110.170 604.000 ;
        RECT 2109.890 600.030 2110.780 600.170 ;
        RECT 2109.890 600.000 2110.170 600.030 ;
        RECT 2110.640 38.410 2110.780 600.030 ;
        RECT 2110.580 38.090 2110.840 38.410 ;
        RECT 2797.820 38.090 2798.080 38.410 ;
        RECT 2797.880 2.400 2798.020 38.090 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2120.670 586.740 2120.990 586.800 ;
        RECT 2124.810 586.740 2125.130 586.800 ;
        RECT 2120.670 586.600 2125.130 586.740 ;
        RECT 2120.670 586.540 2120.990 586.600 ;
        RECT 2124.810 586.540 2125.130 586.600 ;
        RECT 2124.810 37.980 2125.130 38.040 ;
        RECT 2815.730 37.980 2816.050 38.040 ;
        RECT 2124.810 37.840 2816.050 37.980 ;
        RECT 2124.810 37.780 2125.130 37.840 ;
        RECT 2815.730 37.780 2816.050 37.840 ;
      LAYER via ;
        RECT 2120.700 586.540 2120.960 586.800 ;
        RECT 2124.840 586.540 2125.100 586.800 ;
        RECT 2124.840 37.780 2125.100 38.040 ;
        RECT 2815.760 37.780 2816.020 38.040 ;
      LAYER met2 ;
        RECT 2119.090 600.170 2119.370 604.000 ;
        RECT 2119.090 600.030 2120.900 600.170 ;
        RECT 2119.090 600.000 2119.370 600.030 ;
        RECT 2120.760 586.830 2120.900 600.030 ;
        RECT 2120.700 586.510 2120.960 586.830 ;
        RECT 2124.840 586.510 2125.100 586.830 ;
        RECT 2124.900 38.070 2125.040 586.510 ;
        RECT 2124.840 37.750 2125.100 38.070 ;
        RECT 2815.760 37.750 2816.020 38.070 ;
        RECT 2815.820 2.400 2815.960 37.750 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2129.870 572.260 2130.190 572.520 ;
        RECT 2129.960 572.120 2130.100 572.260 ;
        RECT 2130.790 572.120 2131.110 572.180 ;
        RECT 2129.960 571.980 2131.110 572.120 ;
        RECT 2130.790 571.920 2131.110 571.980 ;
        RECT 2129.870 524.180 2130.190 524.240 ;
        RECT 2130.790 524.180 2131.110 524.240 ;
        RECT 2129.870 524.040 2131.110 524.180 ;
        RECT 2129.870 523.980 2130.190 524.040 ;
        RECT 2130.790 523.980 2131.110 524.040 ;
        RECT 2130.330 403.480 2130.650 403.540 ;
        RECT 2130.790 403.480 2131.110 403.540 ;
        RECT 2130.330 403.340 2131.110 403.480 ;
        RECT 2130.330 403.280 2130.650 403.340 ;
        RECT 2130.790 403.280 2131.110 403.340 ;
        RECT 2130.330 372.540 2130.650 372.600 ;
        RECT 2132.170 372.540 2132.490 372.600 ;
        RECT 2130.330 372.400 2132.490 372.540 ;
        RECT 2130.330 372.340 2130.650 372.400 ;
        RECT 2132.170 372.340 2132.490 372.400 ;
        RECT 2129.870 324.260 2130.190 324.320 ;
        RECT 2130.330 324.260 2130.650 324.320 ;
        RECT 2129.870 324.120 2130.650 324.260 ;
        RECT 2129.870 324.060 2130.190 324.120 ;
        RECT 2130.330 324.060 2130.650 324.120 ;
        RECT 2129.870 276.660 2130.190 276.720 ;
        RECT 2130.330 276.660 2130.650 276.720 ;
        RECT 2129.870 276.520 2130.650 276.660 ;
        RECT 2129.870 276.460 2130.190 276.520 ;
        RECT 2130.330 276.460 2130.650 276.520 ;
        RECT 2128.950 275.980 2129.270 276.040 ;
        RECT 2130.330 275.980 2130.650 276.040 ;
        RECT 2128.950 275.840 2130.650 275.980 ;
        RECT 2128.950 275.780 2129.270 275.840 ;
        RECT 2130.330 275.780 2130.650 275.840 ;
        RECT 2128.950 228.040 2129.270 228.100 ;
        RECT 2129.870 228.040 2130.190 228.100 ;
        RECT 2128.950 227.900 2130.190 228.040 ;
        RECT 2128.950 227.840 2129.270 227.900 ;
        RECT 2129.870 227.840 2130.190 227.900 ;
        RECT 2128.950 227.360 2129.270 227.420 ;
        RECT 2129.870 227.360 2130.190 227.420 ;
        RECT 2128.950 227.220 2130.190 227.360 ;
        RECT 2128.950 227.160 2129.270 227.220 ;
        RECT 2129.870 227.160 2130.190 227.220 ;
        RECT 2129.870 172.620 2130.190 172.680 ;
        RECT 2130.330 172.620 2130.650 172.680 ;
        RECT 2129.870 172.480 2130.650 172.620 ;
        RECT 2129.870 172.420 2130.190 172.480 ;
        RECT 2130.330 172.420 2130.650 172.480 ;
        RECT 2130.330 124.000 2130.650 124.060 ;
        RECT 2130.790 124.000 2131.110 124.060 ;
        RECT 2130.330 123.860 2131.110 124.000 ;
        RECT 2130.330 123.800 2130.650 123.860 ;
        RECT 2130.790 123.800 2131.110 123.860 ;
        RECT 2130.790 45.800 2131.110 45.860 ;
        RECT 2833.670 45.800 2833.990 45.860 ;
        RECT 2130.790 45.660 2833.990 45.800 ;
        RECT 2130.790 45.600 2131.110 45.660 ;
        RECT 2833.670 45.600 2833.990 45.660 ;
      LAYER via ;
        RECT 2129.900 572.260 2130.160 572.520 ;
        RECT 2130.820 571.920 2131.080 572.180 ;
        RECT 2129.900 523.980 2130.160 524.240 ;
        RECT 2130.820 523.980 2131.080 524.240 ;
        RECT 2130.360 403.280 2130.620 403.540 ;
        RECT 2130.820 403.280 2131.080 403.540 ;
        RECT 2130.360 372.340 2130.620 372.600 ;
        RECT 2132.200 372.340 2132.460 372.600 ;
        RECT 2129.900 324.060 2130.160 324.320 ;
        RECT 2130.360 324.060 2130.620 324.320 ;
        RECT 2129.900 276.460 2130.160 276.720 ;
        RECT 2130.360 276.460 2130.620 276.720 ;
        RECT 2128.980 275.780 2129.240 276.040 ;
        RECT 2130.360 275.780 2130.620 276.040 ;
        RECT 2128.980 227.840 2129.240 228.100 ;
        RECT 2129.900 227.840 2130.160 228.100 ;
        RECT 2128.980 227.160 2129.240 227.420 ;
        RECT 2129.900 227.160 2130.160 227.420 ;
        RECT 2129.900 172.420 2130.160 172.680 ;
        RECT 2130.360 172.420 2130.620 172.680 ;
        RECT 2130.360 123.800 2130.620 124.060 ;
        RECT 2130.820 123.800 2131.080 124.060 ;
        RECT 2130.820 45.600 2131.080 45.860 ;
        RECT 2833.700 45.600 2833.960 45.860 ;
      LAYER met2 ;
        RECT 2128.290 600.170 2128.570 604.000 ;
        RECT 2128.290 600.030 2130.100 600.170 ;
        RECT 2128.290 600.000 2128.570 600.030 ;
        RECT 2129.960 572.550 2130.100 600.030 ;
        RECT 2129.900 572.230 2130.160 572.550 ;
        RECT 2130.820 571.890 2131.080 572.210 ;
        RECT 2130.880 524.270 2131.020 571.890 ;
        RECT 2129.900 523.950 2130.160 524.270 ;
        RECT 2130.820 523.950 2131.080 524.270 ;
        RECT 2129.960 435.045 2130.100 523.950 ;
        RECT 2129.890 434.675 2130.170 435.045 ;
        RECT 2130.810 434.675 2131.090 435.045 ;
        RECT 2130.880 403.570 2131.020 434.675 ;
        RECT 2130.360 403.250 2130.620 403.570 ;
        RECT 2130.820 403.250 2131.080 403.570 ;
        RECT 2130.420 372.630 2130.560 403.250 ;
        RECT 2130.360 372.310 2130.620 372.630 ;
        RECT 2132.200 372.310 2132.460 372.630 ;
        RECT 2132.260 324.885 2132.400 372.310 ;
        RECT 2130.350 324.515 2130.630 324.885 ;
        RECT 2132.190 324.515 2132.470 324.885 ;
        RECT 2130.420 324.350 2130.560 324.515 ;
        RECT 2129.900 324.030 2130.160 324.350 ;
        RECT 2130.360 324.030 2130.620 324.350 ;
        RECT 2129.960 276.750 2130.100 324.030 ;
        RECT 2129.900 276.430 2130.160 276.750 ;
        RECT 2130.360 276.430 2130.620 276.750 ;
        RECT 2130.420 276.070 2130.560 276.430 ;
        RECT 2128.980 275.750 2129.240 276.070 ;
        RECT 2130.360 275.750 2130.620 276.070 ;
        RECT 2129.040 228.130 2129.180 275.750 ;
        RECT 2128.980 227.810 2129.240 228.130 ;
        RECT 2129.900 227.810 2130.160 228.130 ;
        RECT 2129.960 227.450 2130.100 227.810 ;
        RECT 2128.980 227.130 2129.240 227.450 ;
        RECT 2129.900 227.130 2130.160 227.450 ;
        RECT 2129.040 220.845 2129.180 227.130 ;
        RECT 2128.970 220.475 2129.250 220.845 ;
        RECT 2129.890 220.475 2130.170 220.845 ;
        RECT 2129.960 172.710 2130.100 220.475 ;
        RECT 2129.900 172.390 2130.160 172.710 ;
        RECT 2130.360 172.390 2130.620 172.710 ;
        RECT 2130.420 124.090 2130.560 172.390 ;
        RECT 2130.360 123.770 2130.620 124.090 ;
        RECT 2130.820 123.770 2131.080 124.090 ;
        RECT 2130.880 45.890 2131.020 123.770 ;
        RECT 2130.820 45.570 2131.080 45.890 ;
        RECT 2833.700 45.570 2833.960 45.890 ;
        RECT 2833.760 2.400 2833.900 45.570 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
      LAYER via2 ;
        RECT 2129.890 434.720 2130.170 435.000 ;
        RECT 2130.810 434.720 2131.090 435.000 ;
        RECT 2130.350 324.560 2130.630 324.840 ;
        RECT 2132.190 324.560 2132.470 324.840 ;
        RECT 2128.970 220.520 2129.250 220.800 ;
        RECT 2129.890 220.520 2130.170 220.800 ;
      LAYER met3 ;
        RECT 2129.865 435.010 2130.195 435.025 ;
        RECT 2130.785 435.010 2131.115 435.025 ;
        RECT 2129.865 434.710 2131.115 435.010 ;
        RECT 2129.865 434.695 2130.195 434.710 ;
        RECT 2130.785 434.695 2131.115 434.710 ;
        RECT 2130.325 324.850 2130.655 324.865 ;
        RECT 2132.165 324.850 2132.495 324.865 ;
        RECT 2130.325 324.550 2132.495 324.850 ;
        RECT 2130.325 324.535 2130.655 324.550 ;
        RECT 2132.165 324.535 2132.495 324.550 ;
        RECT 2128.945 220.810 2129.275 220.825 ;
        RECT 2129.865 220.810 2130.195 220.825 ;
        RECT 2128.945 220.510 2130.195 220.810 ;
        RECT 2128.945 220.495 2129.275 220.510 ;
        RECT 2129.865 220.495 2130.195 220.510 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2138.150 45.120 2138.470 45.180 ;
        RECT 2851.150 45.120 2851.470 45.180 ;
        RECT 2138.150 44.980 2851.470 45.120 ;
        RECT 2138.150 44.920 2138.470 44.980 ;
        RECT 2851.150 44.920 2851.470 44.980 ;
      LAYER via ;
        RECT 2138.180 44.920 2138.440 45.180 ;
        RECT 2851.180 44.920 2851.440 45.180 ;
      LAYER met2 ;
        RECT 2137.490 600.170 2137.770 604.000 ;
        RECT 2137.490 600.030 2138.380 600.170 ;
        RECT 2137.490 600.000 2137.770 600.030 ;
        RECT 2138.240 45.210 2138.380 600.030 ;
        RECT 2138.180 44.890 2138.440 45.210 ;
        RECT 2851.180 44.890 2851.440 45.210 ;
        RECT 2851.240 2.400 2851.380 44.890 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2148.270 586.740 2148.590 586.800 ;
        RECT 2152.410 586.740 2152.730 586.800 ;
        RECT 2148.270 586.600 2152.730 586.740 ;
        RECT 2148.270 586.540 2148.590 586.600 ;
        RECT 2152.410 586.540 2152.730 586.600 ;
        RECT 2152.410 45.460 2152.730 45.520 ;
        RECT 2869.090 45.460 2869.410 45.520 ;
        RECT 2152.410 45.320 2869.410 45.460 ;
        RECT 2152.410 45.260 2152.730 45.320 ;
        RECT 2869.090 45.260 2869.410 45.320 ;
      LAYER via ;
        RECT 2148.300 586.540 2148.560 586.800 ;
        RECT 2152.440 586.540 2152.700 586.800 ;
        RECT 2152.440 45.260 2152.700 45.520 ;
        RECT 2869.120 45.260 2869.380 45.520 ;
      LAYER met2 ;
        RECT 2146.690 600.170 2146.970 604.000 ;
        RECT 2146.690 600.030 2148.500 600.170 ;
        RECT 2146.690 600.000 2146.970 600.030 ;
        RECT 2148.360 586.830 2148.500 600.030 ;
        RECT 2148.300 586.510 2148.560 586.830 ;
        RECT 2152.440 586.510 2152.700 586.830 ;
        RECT 2152.500 45.550 2152.640 586.510 ;
        RECT 2152.440 45.230 2152.700 45.550 ;
        RECT 2869.120 45.230 2869.380 45.550 ;
        RECT 2869.180 2.400 2869.320 45.230 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2157.930 572.460 2158.250 572.520 ;
        RECT 2158.390 572.460 2158.710 572.520 ;
        RECT 2157.930 572.320 2158.710 572.460 ;
        RECT 2157.930 572.260 2158.250 572.320 ;
        RECT 2158.390 572.260 2158.710 572.320 ;
        RECT 2158.390 531.460 2158.710 531.720 ;
        RECT 2157.930 531.320 2158.250 531.380 ;
        RECT 2158.480 531.320 2158.620 531.460 ;
        RECT 2157.930 531.180 2158.620 531.320 ;
        RECT 2157.930 531.120 2158.250 531.180 ;
        RECT 2157.010 524.180 2157.330 524.240 ;
        RECT 2158.390 524.180 2158.710 524.240 ;
        RECT 2157.010 524.040 2158.710 524.180 ;
        RECT 2157.010 523.980 2157.330 524.040 ;
        RECT 2158.390 523.980 2158.710 524.040 ;
        RECT 2157.010 475.900 2157.330 475.960 ;
        RECT 2157.470 475.900 2157.790 475.960 ;
        RECT 2157.010 475.760 2157.790 475.900 ;
        RECT 2157.010 475.700 2157.330 475.760 ;
        RECT 2157.470 475.700 2157.790 475.760 ;
        RECT 2157.470 427.960 2157.790 428.020 ;
        RECT 2157.930 427.960 2158.250 428.020 ;
        RECT 2157.470 427.820 2158.250 427.960 ;
        RECT 2157.470 427.760 2157.790 427.820 ;
        RECT 2157.930 427.760 2158.250 427.820 ;
        RECT 2157.930 400.420 2158.250 400.480 ;
        RECT 2158.850 400.420 2159.170 400.480 ;
        RECT 2157.930 400.280 2159.170 400.420 ;
        RECT 2157.930 400.220 2158.250 400.280 ;
        RECT 2158.850 400.220 2159.170 400.280 ;
        RECT 2157.930 379.340 2158.250 379.400 ;
        RECT 2158.850 379.340 2159.170 379.400 ;
        RECT 2157.930 379.200 2159.170 379.340 ;
        RECT 2157.930 379.140 2158.250 379.200 ;
        RECT 2158.850 379.140 2159.170 379.200 ;
        RECT 2157.010 324.260 2157.330 324.320 ;
        RECT 2157.930 324.260 2158.250 324.320 ;
        RECT 2157.010 324.120 2158.250 324.260 ;
        RECT 2157.010 324.060 2157.330 324.120 ;
        RECT 2157.930 324.060 2158.250 324.120 ;
        RECT 2157.010 276.320 2157.330 276.380 ;
        RECT 2157.930 276.320 2158.250 276.380 ;
        RECT 2157.010 276.180 2158.250 276.320 ;
        RECT 2157.010 276.120 2157.330 276.180 ;
        RECT 2157.930 276.120 2158.250 276.180 ;
        RECT 2157.470 227.700 2157.790 227.760 ;
        RECT 2157.930 227.700 2158.250 227.760 ;
        RECT 2157.470 227.560 2158.250 227.700 ;
        RECT 2157.470 227.500 2157.790 227.560 ;
        RECT 2157.930 227.500 2158.250 227.560 ;
        RECT 2157.010 179.760 2157.330 179.820 ;
        RECT 2157.470 179.760 2157.790 179.820 ;
        RECT 2157.010 179.620 2157.790 179.760 ;
        RECT 2157.010 179.560 2157.330 179.620 ;
        RECT 2157.470 179.560 2157.790 179.620 ;
        RECT 2157.010 138.280 2157.330 138.340 ;
        RECT 2158.390 138.280 2158.710 138.340 ;
        RECT 2157.010 138.140 2158.710 138.280 ;
        RECT 2157.010 138.080 2157.330 138.140 ;
        RECT 2158.390 138.080 2158.710 138.140 ;
        RECT 2158.390 44.780 2158.710 44.840 ;
        RECT 2887.030 44.780 2887.350 44.840 ;
        RECT 2158.390 44.640 2887.350 44.780 ;
        RECT 2158.390 44.580 2158.710 44.640 ;
        RECT 2887.030 44.580 2887.350 44.640 ;
      LAYER via ;
        RECT 2157.960 572.260 2158.220 572.520 ;
        RECT 2158.420 572.260 2158.680 572.520 ;
        RECT 2158.420 531.460 2158.680 531.720 ;
        RECT 2157.960 531.120 2158.220 531.380 ;
        RECT 2157.040 523.980 2157.300 524.240 ;
        RECT 2158.420 523.980 2158.680 524.240 ;
        RECT 2157.040 475.700 2157.300 475.960 ;
        RECT 2157.500 475.700 2157.760 475.960 ;
        RECT 2157.500 427.760 2157.760 428.020 ;
        RECT 2157.960 427.760 2158.220 428.020 ;
        RECT 2157.960 400.220 2158.220 400.480 ;
        RECT 2158.880 400.220 2159.140 400.480 ;
        RECT 2157.960 379.140 2158.220 379.400 ;
        RECT 2158.880 379.140 2159.140 379.400 ;
        RECT 2157.040 324.060 2157.300 324.320 ;
        RECT 2157.960 324.060 2158.220 324.320 ;
        RECT 2157.040 276.120 2157.300 276.380 ;
        RECT 2157.960 276.120 2158.220 276.380 ;
        RECT 2157.500 227.500 2157.760 227.760 ;
        RECT 2157.960 227.500 2158.220 227.760 ;
        RECT 2157.040 179.560 2157.300 179.820 ;
        RECT 2157.500 179.560 2157.760 179.820 ;
        RECT 2157.040 138.080 2157.300 138.340 ;
        RECT 2158.420 138.080 2158.680 138.340 ;
        RECT 2158.420 44.580 2158.680 44.840 ;
        RECT 2887.060 44.580 2887.320 44.840 ;
      LAYER met2 ;
        RECT 2155.890 600.170 2156.170 604.000 ;
        RECT 2155.890 600.030 2156.780 600.170 ;
        RECT 2155.890 600.000 2156.170 600.030 ;
        RECT 2156.640 573.765 2156.780 600.030 ;
        RECT 2156.570 573.395 2156.850 573.765 ;
        RECT 2157.950 572.715 2158.230 573.085 ;
        RECT 2158.020 572.550 2158.160 572.715 ;
        RECT 2157.960 572.230 2158.220 572.550 ;
        RECT 2158.420 572.230 2158.680 572.550 ;
        RECT 2158.480 531.750 2158.620 572.230 ;
        RECT 2158.420 531.430 2158.680 531.750 ;
        RECT 2157.960 531.090 2158.220 531.410 ;
        RECT 2158.020 524.690 2158.160 531.090 ;
        RECT 2158.020 524.550 2158.620 524.690 ;
        RECT 2158.480 524.270 2158.620 524.550 ;
        RECT 2157.040 523.950 2157.300 524.270 ;
        RECT 2158.420 523.950 2158.680 524.270 ;
        RECT 2157.100 475.990 2157.240 523.950 ;
        RECT 2157.040 475.670 2157.300 475.990 ;
        RECT 2157.500 475.670 2157.760 475.990 ;
        RECT 2157.560 428.050 2157.700 475.670 ;
        RECT 2157.500 427.730 2157.760 428.050 ;
        RECT 2157.960 427.730 2158.220 428.050 ;
        RECT 2158.020 400.510 2158.160 427.730 ;
        RECT 2158.940 400.510 2159.080 400.665 ;
        RECT 2157.960 400.250 2158.220 400.510 ;
        RECT 2158.880 400.250 2159.140 400.510 ;
        RECT 2157.960 400.190 2159.140 400.250 ;
        RECT 2158.020 400.110 2159.080 400.190 ;
        RECT 2158.020 379.430 2158.160 400.110 ;
        RECT 2157.960 379.110 2158.220 379.430 ;
        RECT 2158.880 379.110 2159.140 379.430 ;
        RECT 2158.940 331.685 2159.080 379.110 ;
        RECT 2157.950 331.315 2158.230 331.685 ;
        RECT 2158.870 331.315 2159.150 331.685 ;
        RECT 2158.020 324.350 2158.160 331.315 ;
        RECT 2157.040 324.030 2157.300 324.350 ;
        RECT 2157.960 324.030 2158.220 324.350 ;
        RECT 2157.100 276.410 2157.240 324.030 ;
        RECT 2157.040 276.090 2157.300 276.410 ;
        RECT 2157.960 276.090 2158.220 276.410 ;
        RECT 2158.020 227.790 2158.160 276.090 ;
        RECT 2157.500 227.470 2157.760 227.790 ;
        RECT 2157.960 227.470 2158.220 227.790 ;
        RECT 2157.560 179.850 2157.700 227.470 ;
        RECT 2157.040 179.530 2157.300 179.850 ;
        RECT 2157.500 179.530 2157.760 179.850 ;
        RECT 2157.100 138.370 2157.240 179.530 ;
        RECT 2157.040 138.050 2157.300 138.370 ;
        RECT 2158.420 138.050 2158.680 138.370 ;
        RECT 2158.480 110.570 2158.620 138.050 ;
        RECT 2158.480 110.430 2159.080 110.570 ;
        RECT 2158.940 62.290 2159.080 110.430 ;
        RECT 2158.480 62.150 2159.080 62.290 ;
        RECT 2158.480 44.870 2158.620 62.150 ;
        RECT 2158.420 44.550 2158.680 44.870 ;
        RECT 2887.060 44.550 2887.320 44.870 ;
        RECT 2887.120 2.400 2887.260 44.550 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
      LAYER via2 ;
        RECT 2156.570 573.440 2156.850 573.720 ;
        RECT 2157.950 572.760 2158.230 573.040 ;
        RECT 2157.950 331.360 2158.230 331.640 ;
        RECT 2158.870 331.360 2159.150 331.640 ;
      LAYER met3 ;
        RECT 2156.545 573.730 2156.875 573.745 ;
        RECT 2156.545 573.430 2158.930 573.730 ;
        RECT 2156.545 573.415 2156.875 573.430 ;
        RECT 2157.925 573.050 2158.255 573.065 ;
        RECT 2158.630 573.050 2158.930 573.430 ;
        RECT 2157.925 572.750 2158.930 573.050 ;
        RECT 2157.925 572.735 2158.255 572.750 ;
        RECT 2157.925 331.650 2158.255 331.665 ;
        RECT 2158.845 331.650 2159.175 331.665 ;
        RECT 2157.925 331.350 2159.175 331.650 ;
        RECT 2157.925 331.335 2158.255 331.350 ;
        RECT 2158.845 331.335 2159.175 331.350 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2165.750 51.580 2166.070 51.640 ;
        RECT 2905.430 51.580 2905.750 51.640 ;
        RECT 2165.750 51.440 2905.750 51.580 ;
        RECT 2165.750 51.380 2166.070 51.440 ;
        RECT 2905.430 51.380 2905.750 51.440 ;
      LAYER via ;
        RECT 2165.780 51.380 2166.040 51.640 ;
        RECT 2905.460 51.380 2905.720 51.640 ;
      LAYER met2 ;
        RECT 2165.090 600.170 2165.370 604.000 ;
        RECT 2165.090 600.030 2165.980 600.170 ;
        RECT 2165.090 600.000 2165.370 600.030 ;
        RECT 2165.840 51.670 2165.980 600.030 ;
        RECT 2165.780 51.350 2166.040 51.670 ;
        RECT 2905.460 51.350 2905.720 51.670 ;
        RECT 2905.520 3.130 2905.660 51.350 ;
        RECT 2905.060 2.990 2905.660 3.130 ;
        RECT 2905.060 2.400 2905.200 2.990 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1106.370 524.180 1106.690 524.240 ;
        RECT 1107.290 524.180 1107.610 524.240 ;
        RECT 1106.370 524.040 1107.610 524.180 ;
        RECT 1106.370 523.980 1106.690 524.040 ;
        RECT 1107.290 523.980 1107.610 524.040 ;
        RECT 1104.990 379.340 1105.310 379.400 ;
        RECT 1106.370 379.340 1106.690 379.400 ;
        RECT 1104.990 379.200 1106.690 379.340 ;
        RECT 1104.990 379.140 1105.310 379.200 ;
        RECT 1106.370 379.140 1106.690 379.200 ;
        RECT 1104.990 331.060 1105.310 331.120 ;
        RECT 1105.450 331.060 1105.770 331.120 ;
        RECT 1104.990 330.920 1105.770 331.060 ;
        RECT 1104.990 330.860 1105.310 330.920 ;
        RECT 1105.450 330.860 1105.770 330.920 ;
        RECT 1104.990 324.260 1105.310 324.320 ;
        RECT 1105.910 324.260 1106.230 324.320 ;
        RECT 1104.990 324.120 1106.230 324.260 ;
        RECT 1104.990 324.060 1105.310 324.120 ;
        RECT 1105.910 324.060 1106.230 324.120 ;
        RECT 1104.990 276.320 1105.310 276.380 ;
        RECT 1105.910 276.320 1106.230 276.380 ;
        RECT 1104.990 276.180 1106.230 276.320 ;
        RECT 1104.990 276.120 1105.310 276.180 ;
        RECT 1105.910 276.120 1106.230 276.180 ;
        RECT 1104.990 227.700 1105.310 227.760 ;
        RECT 1106.370 227.700 1106.690 227.760 ;
        RECT 1104.990 227.560 1106.690 227.700 ;
        RECT 1104.990 227.500 1105.310 227.560 ;
        RECT 1106.370 227.500 1106.690 227.560 ;
        RECT 1105.450 138.280 1105.770 138.340 ;
        RECT 1106.370 138.280 1106.690 138.340 ;
        RECT 1105.450 138.140 1106.690 138.280 ;
        RECT 1105.450 138.080 1105.770 138.140 ;
        RECT 1106.370 138.080 1106.690 138.140 ;
        RECT 1104.990 90.000 1105.310 90.060 ;
        RECT 1105.450 90.000 1105.770 90.060 ;
        RECT 1104.990 89.860 1105.770 90.000 ;
        RECT 1104.990 89.800 1105.310 89.860 ;
        RECT 1105.450 89.800 1105.770 89.860 ;
        RECT 852.910 26.080 853.230 26.140 ;
        RECT 1104.990 26.080 1105.310 26.140 ;
        RECT 852.910 25.940 1105.310 26.080 ;
        RECT 852.910 25.880 853.230 25.940 ;
        RECT 1104.990 25.880 1105.310 25.940 ;
      LAYER via ;
        RECT 1106.400 523.980 1106.660 524.240 ;
        RECT 1107.320 523.980 1107.580 524.240 ;
        RECT 1105.020 379.140 1105.280 379.400 ;
        RECT 1106.400 379.140 1106.660 379.400 ;
        RECT 1105.020 330.860 1105.280 331.120 ;
        RECT 1105.480 330.860 1105.740 331.120 ;
        RECT 1105.020 324.060 1105.280 324.320 ;
        RECT 1105.940 324.060 1106.200 324.320 ;
        RECT 1105.020 276.120 1105.280 276.380 ;
        RECT 1105.940 276.120 1106.200 276.380 ;
        RECT 1105.020 227.500 1105.280 227.760 ;
        RECT 1106.400 227.500 1106.660 227.760 ;
        RECT 1105.480 138.080 1105.740 138.340 ;
        RECT 1106.400 138.080 1106.660 138.340 ;
        RECT 1105.020 89.800 1105.280 90.060 ;
        RECT 1105.480 89.800 1105.740 90.060 ;
        RECT 852.940 25.880 853.200 26.140 ;
        RECT 1105.020 25.880 1105.280 26.140 ;
      LAYER met2 ;
        RECT 1108.930 600.170 1109.210 604.000 ;
        RECT 1108.300 600.030 1109.210 600.170 ;
        RECT 1108.300 579.885 1108.440 600.030 ;
        RECT 1108.930 600.000 1109.210 600.030 ;
        RECT 1107.310 579.515 1107.590 579.885 ;
        RECT 1108.230 579.515 1108.510 579.885 ;
        RECT 1107.380 524.270 1107.520 579.515 ;
        RECT 1106.400 523.950 1106.660 524.270 ;
        RECT 1107.320 523.950 1107.580 524.270 ;
        RECT 1106.460 495.450 1106.600 523.950 ;
        RECT 1105.540 495.310 1106.600 495.450 ;
        RECT 1105.540 400.250 1105.680 495.310 ;
        RECT 1105.080 400.110 1105.680 400.250 ;
        RECT 1105.080 379.430 1105.220 400.110 ;
        RECT 1105.020 379.110 1105.280 379.430 ;
        RECT 1106.400 379.110 1106.660 379.430 ;
        RECT 1106.460 331.685 1106.600 379.110 ;
        RECT 1105.470 331.315 1105.750 331.685 ;
        RECT 1106.390 331.315 1106.670 331.685 ;
        RECT 1105.540 331.150 1105.680 331.315 ;
        RECT 1105.020 330.830 1105.280 331.150 ;
        RECT 1105.480 330.830 1105.740 331.150 ;
        RECT 1105.080 324.350 1105.220 330.830 ;
        RECT 1105.020 324.030 1105.280 324.350 ;
        RECT 1105.940 324.030 1106.200 324.350 ;
        RECT 1106.000 276.410 1106.140 324.030 ;
        RECT 1105.020 276.090 1105.280 276.410 ;
        RECT 1105.940 276.090 1106.200 276.410 ;
        RECT 1105.080 227.790 1105.220 276.090 ;
        RECT 1105.020 227.470 1105.280 227.790 ;
        RECT 1106.400 227.470 1106.660 227.790 ;
        RECT 1106.460 138.370 1106.600 227.470 ;
        RECT 1105.480 138.050 1105.740 138.370 ;
        RECT 1106.400 138.050 1106.660 138.370 ;
        RECT 1105.540 90.090 1105.680 138.050 ;
        RECT 1105.020 89.770 1105.280 90.090 ;
        RECT 1105.480 89.770 1105.740 90.090 ;
        RECT 1105.080 26.170 1105.220 89.770 ;
        RECT 852.940 25.850 853.200 26.170 ;
        RECT 1105.020 25.850 1105.280 26.170 ;
        RECT 853.000 2.400 853.140 25.850 ;
        RECT 852.790 -4.800 853.350 2.400 ;
      LAYER via2 ;
        RECT 1107.310 579.560 1107.590 579.840 ;
        RECT 1108.230 579.560 1108.510 579.840 ;
        RECT 1105.470 331.360 1105.750 331.640 ;
        RECT 1106.390 331.360 1106.670 331.640 ;
      LAYER met3 ;
        RECT 1107.285 579.850 1107.615 579.865 ;
        RECT 1108.205 579.850 1108.535 579.865 ;
        RECT 1107.285 579.550 1108.535 579.850 ;
        RECT 1107.285 579.535 1107.615 579.550 ;
        RECT 1108.205 579.535 1108.535 579.550 ;
        RECT 1105.445 331.650 1105.775 331.665 ;
        RECT 1106.365 331.650 1106.695 331.665 ;
        RECT 1105.445 331.350 1106.695 331.650 ;
        RECT 1105.445 331.335 1105.775 331.350 ;
        RECT 1106.365 331.335 1106.695 331.350 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 26.420 871.170 26.480 ;
        RECT 1118.330 26.420 1118.650 26.480 ;
        RECT 870.850 26.280 1118.650 26.420 ;
        RECT 870.850 26.220 871.170 26.280 ;
        RECT 1118.330 26.220 1118.650 26.280 ;
      LAYER via ;
        RECT 870.880 26.220 871.140 26.480 ;
        RECT 1118.360 26.220 1118.620 26.480 ;
      LAYER met2 ;
        RECT 1118.130 600.000 1118.410 604.000 ;
        RECT 1118.190 598.810 1118.330 600.000 ;
        RECT 1118.190 598.670 1118.560 598.810 ;
        RECT 1118.420 26.510 1118.560 598.670 ;
        RECT 870.880 26.190 871.140 26.510 ;
        RECT 1118.360 26.190 1118.620 26.510 ;
        RECT 870.940 2.400 871.080 26.190 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 889.710 589.800 890.030 589.860 ;
        RECT 1125.690 589.800 1126.010 589.860 ;
        RECT 889.710 589.660 1126.010 589.800 ;
        RECT 889.710 589.600 890.030 589.660 ;
        RECT 1125.690 589.600 1126.010 589.660 ;
      LAYER via ;
        RECT 889.740 589.600 890.000 589.860 ;
        RECT 1125.720 589.600 1125.980 589.860 ;
      LAYER met2 ;
        RECT 1127.330 600.170 1127.610 604.000 ;
        RECT 1125.780 600.030 1127.610 600.170 ;
        RECT 1125.780 589.890 1125.920 600.030 ;
        RECT 1127.330 600.000 1127.610 600.030 ;
        RECT 889.740 589.570 890.000 589.890 ;
        RECT 1125.720 589.570 1125.980 589.890 ;
        RECT 889.800 3.130 889.940 589.570 ;
        RECT 888.880 2.990 889.940 3.130 ;
        RECT 888.880 2.400 889.020 2.990 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 910.410 590.140 910.730 590.200 ;
        RECT 1134.890 590.140 1135.210 590.200 ;
        RECT 910.410 590.000 1135.210 590.140 ;
        RECT 910.410 589.940 910.730 590.000 ;
        RECT 1134.890 589.940 1135.210 590.000 ;
        RECT 906.730 20.640 907.050 20.700 ;
        RECT 910.410 20.640 910.730 20.700 ;
        RECT 906.730 20.500 910.730 20.640 ;
        RECT 906.730 20.440 907.050 20.500 ;
        RECT 910.410 20.440 910.730 20.500 ;
      LAYER via ;
        RECT 910.440 589.940 910.700 590.200 ;
        RECT 1134.920 589.940 1135.180 590.200 ;
        RECT 906.760 20.440 907.020 20.700 ;
        RECT 910.440 20.440 910.700 20.700 ;
      LAYER met2 ;
        RECT 1136.530 600.170 1136.810 604.000 ;
        RECT 1134.980 600.030 1136.810 600.170 ;
        RECT 1134.980 590.230 1135.120 600.030 ;
        RECT 1136.530 600.000 1136.810 600.030 ;
        RECT 910.440 589.910 910.700 590.230 ;
        RECT 1134.920 589.910 1135.180 590.230 ;
        RECT 910.500 20.730 910.640 589.910 ;
        RECT 906.760 20.410 907.020 20.730 ;
        RECT 910.440 20.410 910.700 20.730 ;
        RECT 906.820 2.400 906.960 20.410 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 591.160 924.530 591.220 ;
        RECT 1145.930 591.160 1146.250 591.220 ;
        RECT 924.210 591.020 1146.250 591.160 ;
        RECT 924.210 590.960 924.530 591.020 ;
        RECT 1145.930 590.960 1146.250 591.020 ;
      LAYER via ;
        RECT 924.240 590.960 924.500 591.220 ;
        RECT 1145.960 590.960 1146.220 591.220 ;
      LAYER met2 ;
        RECT 1145.730 600.000 1146.010 604.000 ;
        RECT 1145.790 598.810 1145.930 600.000 ;
        RECT 1145.790 598.670 1146.160 598.810 ;
        RECT 1146.020 591.250 1146.160 598.670 ;
        RECT 924.240 590.930 924.500 591.250 ;
        RECT 1145.960 590.930 1146.220 591.250 ;
        RECT 924.300 2.400 924.440 590.930 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 944.910 592.520 945.230 592.580 ;
        RECT 1153.290 592.520 1153.610 592.580 ;
        RECT 944.910 592.380 1153.610 592.520 ;
        RECT 944.910 592.320 945.230 592.380 ;
        RECT 1153.290 592.320 1153.610 592.380 ;
        RECT 942.150 20.640 942.470 20.700 ;
        RECT 944.910 20.640 945.230 20.700 ;
        RECT 942.150 20.500 945.230 20.640 ;
        RECT 942.150 20.440 942.470 20.500 ;
        RECT 944.910 20.440 945.230 20.500 ;
      LAYER via ;
        RECT 944.940 592.320 945.200 592.580 ;
        RECT 1153.320 592.320 1153.580 592.580 ;
        RECT 942.180 20.440 942.440 20.700 ;
        RECT 944.940 20.440 945.200 20.700 ;
      LAYER met2 ;
        RECT 1154.930 600.170 1155.210 604.000 ;
        RECT 1153.380 600.030 1155.210 600.170 ;
        RECT 1153.380 592.610 1153.520 600.030 ;
        RECT 1154.930 600.000 1155.210 600.030 ;
        RECT 944.940 592.290 945.200 592.610 ;
        RECT 1153.320 592.290 1153.580 592.610 ;
        RECT 945.000 20.730 945.140 592.290 ;
        RECT 942.180 20.410 942.440 20.730 ;
        RECT 944.940 20.410 945.200 20.730 ;
        RECT 942.240 2.400 942.380 20.410 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1065.890 588.440 1066.210 588.500 ;
        RECT 1162.490 588.440 1162.810 588.500 ;
        RECT 1065.890 588.300 1162.810 588.440 ;
        RECT 1065.890 588.240 1066.210 588.300 ;
        RECT 1162.490 588.240 1162.810 588.300 ;
        RECT 960.090 15.880 960.410 15.940 ;
        RECT 1065.890 15.880 1066.210 15.940 ;
        RECT 960.090 15.740 1066.210 15.880 ;
        RECT 960.090 15.680 960.410 15.740 ;
        RECT 1065.890 15.680 1066.210 15.740 ;
      LAYER via ;
        RECT 1065.920 588.240 1066.180 588.500 ;
        RECT 1162.520 588.240 1162.780 588.500 ;
        RECT 960.120 15.680 960.380 15.940 ;
        RECT 1065.920 15.680 1066.180 15.940 ;
      LAYER met2 ;
        RECT 1164.130 600.170 1164.410 604.000 ;
        RECT 1162.580 600.030 1164.410 600.170 ;
        RECT 1162.580 588.530 1162.720 600.030 ;
        RECT 1164.130 600.000 1164.410 600.030 ;
        RECT 1065.920 588.210 1066.180 588.530 ;
        RECT 1162.520 588.210 1162.780 588.530 ;
        RECT 1065.980 15.970 1066.120 588.210 ;
        RECT 960.120 15.650 960.380 15.970 ;
        RECT 1065.920 15.650 1066.180 15.970 ;
        RECT 960.180 2.400 960.320 15.650 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 979.410 592.860 979.730 592.920 ;
        RECT 1173.530 592.860 1173.850 592.920 ;
        RECT 979.410 592.720 1173.850 592.860 ;
        RECT 979.410 592.660 979.730 592.720 ;
        RECT 1173.530 592.660 1173.850 592.720 ;
      LAYER via ;
        RECT 979.440 592.660 979.700 592.920 ;
        RECT 1173.560 592.660 1173.820 592.920 ;
      LAYER met2 ;
        RECT 1173.330 600.000 1173.610 604.000 ;
        RECT 1173.390 598.810 1173.530 600.000 ;
        RECT 1173.390 598.670 1173.760 598.810 ;
        RECT 1173.620 592.950 1173.760 598.670 ;
        RECT 979.440 592.630 979.700 592.950 ;
        RECT 1173.560 592.630 1173.820 592.950 ;
        RECT 979.500 3.130 979.640 592.630 ;
        RECT 978.120 2.990 979.640 3.130 ;
        RECT 978.120 2.400 978.260 2.990 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 43.760 657.270 43.820 ;
        RECT 1007.930 43.760 1008.250 43.820 ;
        RECT 656.950 43.620 1008.250 43.760 ;
        RECT 656.950 43.560 657.270 43.620 ;
        RECT 1007.930 43.560 1008.250 43.620 ;
      LAYER via ;
        RECT 656.980 43.560 657.240 43.820 ;
        RECT 1007.960 43.560 1008.220 43.820 ;
      LAYER met2 ;
        RECT 1008.190 600.000 1008.470 604.000 ;
        RECT 1008.250 598.810 1008.390 600.000 ;
        RECT 1008.020 598.670 1008.390 598.810 ;
        RECT 1008.020 43.850 1008.160 598.670 ;
        RECT 656.980 43.530 657.240 43.850 ;
        RECT 1007.960 43.530 1008.220 43.850 ;
        RECT 657.040 2.400 657.180 43.530 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1000.110 593.200 1000.430 593.260 ;
        RECT 1180.890 593.200 1181.210 593.260 ;
        RECT 1000.110 593.060 1181.210 593.200 ;
        RECT 1000.110 593.000 1000.430 593.060 ;
        RECT 1180.890 593.000 1181.210 593.060 ;
        RECT 995.970 20.640 996.290 20.700 ;
        RECT 1000.110 20.640 1000.430 20.700 ;
        RECT 995.970 20.500 1000.430 20.640 ;
        RECT 995.970 20.440 996.290 20.500 ;
        RECT 1000.110 20.440 1000.430 20.500 ;
      LAYER via ;
        RECT 1000.140 593.000 1000.400 593.260 ;
        RECT 1180.920 593.000 1181.180 593.260 ;
        RECT 996.000 20.440 996.260 20.700 ;
        RECT 1000.140 20.440 1000.400 20.700 ;
      LAYER met2 ;
        RECT 1182.530 600.170 1182.810 604.000 ;
        RECT 1180.980 600.030 1182.810 600.170 ;
        RECT 1180.980 593.290 1181.120 600.030 ;
        RECT 1182.530 600.000 1182.810 600.030 ;
        RECT 1000.140 592.970 1000.400 593.290 ;
        RECT 1180.920 592.970 1181.180 593.290 ;
        RECT 1000.200 20.730 1000.340 592.970 ;
        RECT 996.000 20.410 996.260 20.730 ;
        RECT 1000.140 20.410 1000.400 20.730 ;
        RECT 996.060 2.400 996.200 20.410 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1190.550 591.840 1190.870 591.900 ;
        RECT 1166.720 591.700 1190.870 591.840 ;
        RECT 1155.590 591.500 1155.910 591.560 ;
        RECT 1166.720 591.500 1166.860 591.700 ;
        RECT 1190.550 591.640 1190.870 591.700 ;
        RECT 1155.590 591.360 1166.860 591.500 ;
        RECT 1155.590 591.300 1155.910 591.360 ;
        RECT 1013.450 19.620 1013.770 19.680 ;
        RECT 1155.590 19.620 1155.910 19.680 ;
        RECT 1013.450 19.480 1155.910 19.620 ;
        RECT 1013.450 19.420 1013.770 19.480 ;
        RECT 1155.590 19.420 1155.910 19.480 ;
      LAYER via ;
        RECT 1155.620 591.300 1155.880 591.560 ;
        RECT 1190.580 591.640 1190.840 591.900 ;
        RECT 1013.480 19.420 1013.740 19.680 ;
        RECT 1155.620 19.420 1155.880 19.680 ;
      LAYER met2 ;
        RECT 1191.730 600.170 1192.010 604.000 ;
        RECT 1190.640 600.030 1192.010 600.170 ;
        RECT 1190.640 591.930 1190.780 600.030 ;
        RECT 1191.730 600.000 1192.010 600.030 ;
        RECT 1190.580 591.610 1190.840 591.930 ;
        RECT 1155.620 591.270 1155.880 591.590 ;
        RECT 1155.680 19.710 1155.820 591.270 ;
        RECT 1013.480 19.390 1013.740 19.710 ;
        RECT 1155.620 19.390 1155.880 19.710 ;
        RECT 1013.540 2.400 1013.680 19.390 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1201.130 587.420 1201.450 587.480 ;
        RECT 1194.780 587.280 1201.450 587.420 ;
        RECT 1162.490 587.080 1162.810 587.140 ;
        RECT 1162.490 586.940 1187.100 587.080 ;
        RECT 1162.490 586.880 1162.810 586.940 ;
        RECT 1186.960 586.740 1187.100 586.940 ;
        RECT 1194.780 586.740 1194.920 587.280 ;
        RECT 1201.130 587.220 1201.450 587.280 ;
        RECT 1186.960 586.600 1194.920 586.740 ;
        RECT 1031.390 16.900 1031.710 16.960 ;
        RECT 1161.570 16.900 1161.890 16.960 ;
        RECT 1031.390 16.760 1161.890 16.900 ;
        RECT 1031.390 16.700 1031.710 16.760 ;
        RECT 1161.570 16.700 1161.890 16.760 ;
      LAYER via ;
        RECT 1162.520 586.880 1162.780 587.140 ;
        RECT 1201.160 587.220 1201.420 587.480 ;
        RECT 1031.420 16.700 1031.680 16.960 ;
        RECT 1161.600 16.700 1161.860 16.960 ;
      LAYER met2 ;
        RECT 1200.930 600.000 1201.210 604.000 ;
        RECT 1200.990 598.810 1201.130 600.000 ;
        RECT 1200.990 598.670 1201.360 598.810 ;
        RECT 1201.220 587.510 1201.360 598.670 ;
        RECT 1201.160 587.190 1201.420 587.510 ;
        RECT 1162.520 586.850 1162.780 587.170 ;
        RECT 1162.580 21.490 1162.720 586.850 ;
        RECT 1161.660 21.350 1162.720 21.490 ;
        RECT 1161.660 16.990 1161.800 21.350 ;
        RECT 1031.420 16.670 1031.680 16.990 ;
        RECT 1161.600 16.670 1161.860 16.990 ;
        RECT 1031.480 2.400 1031.620 16.670 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1208.490 589.800 1208.810 589.860 ;
        RECT 1197.540 589.660 1208.810 589.800 ;
        RECT 1190.550 589.460 1190.870 589.520 ;
        RECT 1197.540 589.460 1197.680 589.660 ;
        RECT 1208.490 589.600 1208.810 589.660 ;
        RECT 1190.550 589.320 1197.680 589.460 ;
        RECT 1190.550 589.260 1190.870 589.320 ;
        RECT 1190.090 110.200 1190.410 110.460 ;
        RECT 1190.180 110.060 1190.320 110.200 ;
        RECT 1190.550 110.060 1190.870 110.120 ;
        RECT 1190.180 109.920 1190.870 110.060 ;
        RECT 1190.550 109.860 1190.870 109.920 ;
        RECT 1049.330 19.960 1049.650 20.020 ;
        RECT 1190.550 19.960 1190.870 20.020 ;
        RECT 1049.330 19.820 1190.870 19.960 ;
        RECT 1049.330 19.760 1049.650 19.820 ;
        RECT 1190.550 19.760 1190.870 19.820 ;
      LAYER via ;
        RECT 1190.580 589.260 1190.840 589.520 ;
        RECT 1208.520 589.600 1208.780 589.860 ;
        RECT 1190.120 110.200 1190.380 110.460 ;
        RECT 1190.580 109.860 1190.840 110.120 ;
        RECT 1049.360 19.760 1049.620 20.020 ;
        RECT 1190.580 19.760 1190.840 20.020 ;
      LAYER met2 ;
        RECT 1210.130 600.170 1210.410 604.000 ;
        RECT 1208.580 600.030 1210.410 600.170 ;
        RECT 1208.580 589.890 1208.720 600.030 ;
        RECT 1210.130 600.000 1210.410 600.030 ;
        RECT 1208.520 589.570 1208.780 589.890 ;
        RECT 1190.580 589.230 1190.840 589.550 ;
        RECT 1190.640 483.210 1190.780 589.230 ;
        RECT 1190.180 483.070 1190.780 483.210 ;
        RECT 1190.180 351.970 1190.320 483.070 ;
        RECT 1189.720 351.830 1190.320 351.970 ;
        RECT 1189.720 351.290 1189.860 351.830 ;
        RECT 1189.720 351.150 1190.320 351.290 ;
        RECT 1190.180 255.410 1190.320 351.150 ;
        RECT 1189.720 255.270 1190.320 255.410 ;
        RECT 1189.720 254.730 1189.860 255.270 ;
        RECT 1189.720 254.590 1190.320 254.730 ;
        RECT 1190.180 158.850 1190.320 254.590 ;
        RECT 1189.720 158.710 1190.320 158.850 ;
        RECT 1189.720 158.170 1189.860 158.710 ;
        RECT 1189.720 158.030 1190.320 158.170 ;
        RECT 1190.180 110.490 1190.320 158.030 ;
        RECT 1190.120 110.170 1190.380 110.490 ;
        RECT 1190.580 109.830 1190.840 110.150 ;
        RECT 1190.640 20.050 1190.780 109.830 ;
        RECT 1049.360 19.730 1049.620 20.050 ;
        RECT 1190.580 19.730 1190.840 20.050 ;
        RECT 1049.420 2.400 1049.560 19.730 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 589.120 1069.430 589.180 ;
        RECT 1218.150 589.120 1218.470 589.180 ;
        RECT 1069.110 588.980 1218.470 589.120 ;
        RECT 1069.110 588.920 1069.430 588.980 ;
        RECT 1218.150 588.920 1218.470 588.980 ;
      LAYER via ;
        RECT 1069.140 588.920 1069.400 589.180 ;
        RECT 1218.180 588.920 1218.440 589.180 ;
      LAYER met2 ;
        RECT 1219.330 600.170 1219.610 604.000 ;
        RECT 1218.240 600.030 1219.610 600.170 ;
        RECT 1218.240 589.210 1218.380 600.030 ;
        RECT 1219.330 600.000 1219.610 600.030 ;
        RECT 1069.140 588.890 1069.400 589.210 ;
        RECT 1218.180 588.890 1218.440 589.210 ;
        RECT 1069.200 3.130 1069.340 588.890 ;
        RECT 1067.360 2.990 1069.340 3.130 ;
        RECT 1067.360 2.400 1067.500 2.990 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 588.780 1090.130 588.840 ;
        RECT 1228.270 588.780 1228.590 588.840 ;
        RECT 1089.810 588.640 1228.590 588.780 ;
        RECT 1089.810 588.580 1090.130 588.640 ;
        RECT 1228.270 588.580 1228.590 588.640 ;
        RECT 1085.210 15.200 1085.530 15.260 ;
        RECT 1089.810 15.200 1090.130 15.260 ;
        RECT 1085.210 15.060 1090.130 15.200 ;
        RECT 1085.210 15.000 1085.530 15.060 ;
        RECT 1089.810 15.000 1090.130 15.060 ;
      LAYER via ;
        RECT 1089.840 588.580 1090.100 588.840 ;
        RECT 1228.300 588.580 1228.560 588.840 ;
        RECT 1085.240 15.000 1085.500 15.260 ;
        RECT 1089.840 15.000 1090.100 15.260 ;
      LAYER met2 ;
        RECT 1228.530 600.000 1228.810 604.000 ;
        RECT 1228.590 598.810 1228.730 600.000 ;
        RECT 1228.360 598.670 1228.730 598.810 ;
        RECT 1228.360 588.870 1228.500 598.670 ;
        RECT 1089.840 588.550 1090.100 588.870 ;
        RECT 1228.300 588.550 1228.560 588.870 ;
        RECT 1089.900 15.290 1090.040 588.550 ;
        RECT 1085.240 14.970 1085.500 15.290 ;
        RECT 1089.840 14.970 1090.100 15.290 ;
        RECT 1085.300 2.400 1085.440 14.970 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1210.790 587.080 1211.110 587.140 ;
        RECT 1236.090 587.080 1236.410 587.140 ;
        RECT 1210.790 586.940 1236.410 587.080 ;
        RECT 1210.790 586.880 1211.110 586.940 ;
        RECT 1236.090 586.880 1236.410 586.940 ;
        RECT 1102.690 15.880 1103.010 15.940 ;
        RECT 1102.690 15.740 1173.300 15.880 ;
        RECT 1102.690 15.680 1103.010 15.740 ;
        RECT 1173.160 15.540 1173.300 15.740 ;
        RECT 1210.790 15.540 1211.110 15.600 ;
        RECT 1173.160 15.400 1211.110 15.540 ;
        RECT 1210.790 15.340 1211.110 15.400 ;
      LAYER via ;
        RECT 1210.820 586.880 1211.080 587.140 ;
        RECT 1236.120 586.880 1236.380 587.140 ;
        RECT 1102.720 15.680 1102.980 15.940 ;
        RECT 1210.820 15.340 1211.080 15.600 ;
      LAYER met2 ;
        RECT 1237.730 600.170 1238.010 604.000 ;
        RECT 1236.180 600.030 1238.010 600.170 ;
        RECT 1236.180 587.170 1236.320 600.030 ;
        RECT 1237.730 600.000 1238.010 600.030 ;
        RECT 1210.820 586.850 1211.080 587.170 ;
        RECT 1236.120 586.850 1236.380 587.170 ;
        RECT 1102.720 15.650 1102.980 15.970 ;
        RECT 1102.780 2.400 1102.920 15.650 ;
        RECT 1210.880 15.630 1211.020 586.850 ;
        RECT 1210.820 15.310 1211.080 15.630 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1217.690 587.420 1218.010 587.480 ;
        RECT 1245.290 587.420 1245.610 587.480 ;
        RECT 1217.690 587.280 1245.610 587.420 ;
        RECT 1217.690 587.220 1218.010 587.280 ;
        RECT 1245.290 587.220 1245.610 587.280 ;
        RECT 1120.630 15.200 1120.950 15.260 ;
        RECT 1217.690 15.200 1218.010 15.260 ;
        RECT 1120.630 15.060 1218.010 15.200 ;
        RECT 1120.630 15.000 1120.950 15.060 ;
        RECT 1217.690 15.000 1218.010 15.060 ;
      LAYER via ;
        RECT 1217.720 587.220 1217.980 587.480 ;
        RECT 1245.320 587.220 1245.580 587.480 ;
        RECT 1120.660 15.000 1120.920 15.260 ;
        RECT 1217.720 15.000 1217.980 15.260 ;
      LAYER met2 ;
        RECT 1246.930 600.170 1247.210 604.000 ;
        RECT 1245.380 600.030 1247.210 600.170 ;
        RECT 1245.380 587.510 1245.520 600.030 ;
        RECT 1246.930 600.000 1247.210 600.030 ;
        RECT 1217.720 587.190 1217.980 587.510 ;
        RECT 1245.320 587.190 1245.580 587.510 ;
        RECT 1217.780 15.290 1217.920 587.190 ;
        RECT 1120.660 14.970 1120.920 15.290 ;
        RECT 1217.720 14.970 1217.980 15.290 ;
        RECT 1120.720 2.400 1120.860 14.970 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 590.140 1145.330 590.200 ;
        RECT 1256.330 590.140 1256.650 590.200 ;
        RECT 1145.010 590.000 1256.650 590.140 ;
        RECT 1145.010 589.940 1145.330 590.000 ;
        RECT 1256.330 589.940 1256.650 590.000 ;
        RECT 1138.570 18.260 1138.890 18.320 ;
        RECT 1145.010 18.260 1145.330 18.320 ;
        RECT 1138.570 18.120 1145.330 18.260 ;
        RECT 1138.570 18.060 1138.890 18.120 ;
        RECT 1145.010 18.060 1145.330 18.120 ;
      LAYER via ;
        RECT 1145.040 589.940 1145.300 590.200 ;
        RECT 1256.360 589.940 1256.620 590.200 ;
        RECT 1138.600 18.060 1138.860 18.320 ;
        RECT 1145.040 18.060 1145.300 18.320 ;
      LAYER met2 ;
        RECT 1256.130 600.000 1256.410 604.000 ;
        RECT 1256.190 598.810 1256.330 600.000 ;
        RECT 1256.190 598.670 1256.560 598.810 ;
        RECT 1256.420 590.230 1256.560 598.670 ;
        RECT 1145.040 589.910 1145.300 590.230 ;
        RECT 1256.360 589.910 1256.620 590.230 ;
        RECT 1145.100 18.350 1145.240 589.910 ;
        RECT 1138.600 18.030 1138.860 18.350 ;
        RECT 1145.040 18.030 1145.300 18.350 ;
        RECT 1138.660 2.400 1138.800 18.030 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.810 590.480 1159.130 590.540 ;
        RECT 1263.690 590.480 1264.010 590.540 ;
        RECT 1158.810 590.340 1264.010 590.480 ;
        RECT 1158.810 590.280 1159.130 590.340 ;
        RECT 1263.690 590.280 1264.010 590.340 ;
        RECT 1156.510 20.640 1156.830 20.700 ;
        RECT 1158.810 20.640 1159.130 20.700 ;
        RECT 1156.510 20.500 1159.130 20.640 ;
        RECT 1156.510 20.440 1156.830 20.500 ;
        RECT 1158.810 20.440 1159.130 20.500 ;
      LAYER via ;
        RECT 1158.840 590.280 1159.100 590.540 ;
        RECT 1263.720 590.280 1263.980 590.540 ;
        RECT 1156.540 20.440 1156.800 20.700 ;
        RECT 1158.840 20.440 1159.100 20.700 ;
      LAYER met2 ;
        RECT 1265.330 600.170 1265.610 604.000 ;
        RECT 1263.780 600.030 1265.610 600.170 ;
        RECT 1263.780 590.570 1263.920 600.030 ;
        RECT 1265.330 600.000 1265.610 600.030 ;
        RECT 1158.840 590.250 1159.100 590.570 ;
        RECT 1263.720 590.250 1263.980 590.570 ;
        RECT 1158.900 20.730 1159.040 590.250 ;
        RECT 1156.540 20.410 1156.800 20.730 ;
        RECT 1158.840 20.410 1159.100 20.730 ;
        RECT 1156.600 2.400 1156.740 20.410 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 674.430 45.460 674.750 45.520 ;
        RECT 1014.830 45.460 1015.150 45.520 ;
        RECT 674.430 45.320 1015.150 45.460 ;
        RECT 674.430 45.260 674.750 45.320 ;
        RECT 1014.830 45.260 1015.150 45.320 ;
      LAYER via ;
        RECT 674.460 45.260 674.720 45.520 ;
        RECT 1014.860 45.260 1015.120 45.520 ;
      LAYER met2 ;
        RECT 1017.390 600.170 1017.670 604.000 ;
        RECT 1014.920 600.030 1017.670 600.170 ;
        RECT 1014.920 45.550 1015.060 600.030 ;
        RECT 1017.390 600.000 1017.670 600.030 ;
        RECT 674.460 45.230 674.720 45.550 ;
        RECT 1014.860 45.230 1015.120 45.550 ;
        RECT 674.520 2.400 674.660 45.230 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1179.510 592.180 1179.830 592.240 ;
        RECT 1272.890 592.180 1273.210 592.240 ;
        RECT 1179.510 592.040 1273.210 592.180 ;
        RECT 1179.510 591.980 1179.830 592.040 ;
        RECT 1272.890 591.980 1273.210 592.040 ;
        RECT 1173.990 20.640 1174.310 20.700 ;
        RECT 1179.510 20.640 1179.830 20.700 ;
        RECT 1173.990 20.500 1179.830 20.640 ;
        RECT 1173.990 20.440 1174.310 20.500 ;
        RECT 1179.510 20.440 1179.830 20.500 ;
      LAYER via ;
        RECT 1179.540 591.980 1179.800 592.240 ;
        RECT 1272.920 591.980 1273.180 592.240 ;
        RECT 1174.020 20.440 1174.280 20.700 ;
        RECT 1179.540 20.440 1179.800 20.700 ;
      LAYER met2 ;
        RECT 1274.530 600.170 1274.810 604.000 ;
        RECT 1272.980 600.030 1274.810 600.170 ;
        RECT 1272.980 592.270 1273.120 600.030 ;
        RECT 1274.530 600.000 1274.810 600.030 ;
        RECT 1179.540 591.950 1179.800 592.270 ;
        RECT 1272.920 591.950 1273.180 592.270 ;
        RECT 1179.600 20.730 1179.740 591.950 ;
        RECT 1174.020 20.410 1174.280 20.730 ;
        RECT 1179.540 20.410 1179.800 20.730 ;
        RECT 1174.080 2.400 1174.220 20.410 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1193.310 591.840 1193.630 591.900 ;
        RECT 1283.470 591.840 1283.790 591.900 ;
        RECT 1193.310 591.700 1283.790 591.840 ;
        RECT 1193.310 591.640 1193.630 591.700 ;
        RECT 1283.470 591.640 1283.790 591.700 ;
        RECT 1191.930 2.960 1192.250 3.020 ;
        RECT 1193.310 2.960 1193.630 3.020 ;
        RECT 1191.930 2.820 1193.630 2.960 ;
        RECT 1191.930 2.760 1192.250 2.820 ;
        RECT 1193.310 2.760 1193.630 2.820 ;
      LAYER via ;
        RECT 1193.340 591.640 1193.600 591.900 ;
        RECT 1283.500 591.640 1283.760 591.900 ;
        RECT 1191.960 2.760 1192.220 3.020 ;
        RECT 1193.340 2.760 1193.600 3.020 ;
      LAYER met2 ;
        RECT 1283.730 600.000 1284.010 604.000 ;
        RECT 1283.790 598.810 1283.930 600.000 ;
        RECT 1283.560 598.670 1283.930 598.810 ;
        RECT 1283.560 591.930 1283.700 598.670 ;
        RECT 1193.340 591.610 1193.600 591.930 ;
        RECT 1283.500 591.610 1283.760 591.930 ;
        RECT 1193.400 3.050 1193.540 591.610 ;
        RECT 1191.960 2.730 1192.220 3.050 ;
        RECT 1193.340 2.730 1193.600 3.050 ;
        RECT 1192.020 2.400 1192.160 2.730 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1249.430 593.200 1249.750 593.260 ;
        RECT 1291.290 593.200 1291.610 593.260 ;
        RECT 1249.430 593.060 1291.610 593.200 ;
        RECT 1249.430 593.000 1249.750 593.060 ;
        RECT 1291.290 593.000 1291.610 593.060 ;
        RECT 1214.010 586.740 1214.330 586.800 ;
        RECT 1249.430 586.740 1249.750 586.800 ;
        RECT 1214.010 586.600 1249.750 586.740 ;
        RECT 1214.010 586.540 1214.330 586.600 ;
        RECT 1249.430 586.540 1249.750 586.600 ;
        RECT 1209.870 15.880 1210.190 15.940 ;
        RECT 1214.010 15.880 1214.330 15.940 ;
        RECT 1209.870 15.740 1214.330 15.880 ;
        RECT 1209.870 15.680 1210.190 15.740 ;
        RECT 1214.010 15.680 1214.330 15.740 ;
      LAYER via ;
        RECT 1249.460 593.000 1249.720 593.260 ;
        RECT 1291.320 593.000 1291.580 593.260 ;
        RECT 1214.040 586.540 1214.300 586.800 ;
        RECT 1249.460 586.540 1249.720 586.800 ;
        RECT 1209.900 15.680 1210.160 15.940 ;
        RECT 1214.040 15.680 1214.300 15.940 ;
      LAYER met2 ;
        RECT 1292.470 600.170 1292.750 604.000 ;
        RECT 1291.380 600.030 1292.750 600.170 ;
        RECT 1291.380 593.290 1291.520 600.030 ;
        RECT 1292.470 600.000 1292.750 600.030 ;
        RECT 1249.460 592.970 1249.720 593.290 ;
        RECT 1291.320 592.970 1291.580 593.290 ;
        RECT 1249.520 586.830 1249.660 592.970 ;
        RECT 1214.040 586.510 1214.300 586.830 ;
        RECT 1249.460 586.510 1249.720 586.830 ;
        RECT 1214.100 15.970 1214.240 586.510 ;
        RECT 1209.900 15.650 1210.160 15.970 ;
        RECT 1214.040 15.650 1214.300 15.970 ;
        RECT 1209.960 2.400 1210.100 15.650 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1228.730 589.120 1229.050 589.180 ;
        RECT 1300.030 589.120 1300.350 589.180 ;
        RECT 1228.730 588.980 1300.350 589.120 ;
        RECT 1228.730 588.920 1229.050 588.980 ;
        RECT 1300.030 588.920 1300.350 588.980 ;
        RECT 1226.890 572.800 1227.210 572.860 ;
        RECT 1228.730 572.800 1229.050 572.860 ;
        RECT 1226.890 572.660 1229.050 572.800 ;
        RECT 1226.890 572.600 1227.210 572.660 ;
        RECT 1228.730 572.600 1229.050 572.660 ;
        RECT 1226.890 531.660 1227.210 531.720 ;
        RECT 1227.350 531.660 1227.670 531.720 ;
        RECT 1226.890 531.520 1227.670 531.660 ;
        RECT 1226.890 531.460 1227.210 531.520 ;
        RECT 1227.350 531.460 1227.670 531.520 ;
        RECT 1226.890 47.980 1227.210 48.240 ;
        RECT 1226.980 47.840 1227.120 47.980 ;
        RECT 1227.350 47.840 1227.670 47.900 ;
        RECT 1226.980 47.700 1227.670 47.840 ;
        RECT 1227.350 47.640 1227.670 47.700 ;
      LAYER via ;
        RECT 1228.760 588.920 1229.020 589.180 ;
        RECT 1300.060 588.920 1300.320 589.180 ;
        RECT 1226.920 572.600 1227.180 572.860 ;
        RECT 1228.760 572.600 1229.020 572.860 ;
        RECT 1226.920 531.460 1227.180 531.720 ;
        RECT 1227.380 531.460 1227.640 531.720 ;
        RECT 1226.920 47.980 1227.180 48.240 ;
        RECT 1227.380 47.640 1227.640 47.900 ;
      LAYER met2 ;
        RECT 1301.670 600.170 1301.950 604.000 ;
        RECT 1300.120 600.030 1301.950 600.170 ;
        RECT 1300.120 589.210 1300.260 600.030 ;
        RECT 1301.670 600.000 1301.950 600.030 ;
        RECT 1228.760 588.890 1229.020 589.210 ;
        RECT 1300.060 588.890 1300.320 589.210 ;
        RECT 1228.820 572.890 1228.960 588.890 ;
        RECT 1226.920 572.570 1227.180 572.890 ;
        RECT 1228.760 572.570 1229.020 572.890 ;
        RECT 1226.980 531.750 1227.120 572.570 ;
        RECT 1226.920 531.430 1227.180 531.750 ;
        RECT 1227.380 531.430 1227.640 531.750 ;
        RECT 1227.440 62.290 1227.580 531.430 ;
        RECT 1226.520 62.150 1227.580 62.290 ;
        RECT 1226.520 48.690 1226.660 62.150 ;
        RECT 1226.520 48.550 1227.120 48.690 ;
        RECT 1226.980 48.270 1227.120 48.550 ;
        RECT 1226.920 47.950 1227.180 48.270 ;
        RECT 1227.380 47.610 1227.640 47.930 ;
        RECT 1227.440 20.130 1227.580 47.610 ;
        RECT 1227.440 19.990 1228.040 20.130 ;
        RECT 1227.900 2.400 1228.040 19.990 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 587.420 1248.830 587.480 ;
        RECT 1311.070 587.420 1311.390 587.480 ;
        RECT 1248.510 587.280 1311.390 587.420 ;
        RECT 1248.510 587.220 1248.830 587.280 ;
        RECT 1311.070 587.220 1311.390 587.280 ;
        RECT 1245.750 20.640 1246.070 20.700 ;
        RECT 1248.510 20.640 1248.830 20.700 ;
        RECT 1245.750 20.500 1248.830 20.640 ;
        RECT 1245.750 20.440 1246.070 20.500 ;
        RECT 1248.510 20.440 1248.830 20.500 ;
      LAYER via ;
        RECT 1248.540 587.220 1248.800 587.480 ;
        RECT 1311.100 587.220 1311.360 587.480 ;
        RECT 1245.780 20.440 1246.040 20.700 ;
        RECT 1248.540 20.440 1248.800 20.700 ;
      LAYER met2 ;
        RECT 1310.870 600.000 1311.150 604.000 ;
        RECT 1310.930 598.810 1311.070 600.000 ;
        RECT 1310.930 598.670 1311.300 598.810 ;
        RECT 1311.160 587.510 1311.300 598.670 ;
        RECT 1248.540 587.190 1248.800 587.510 ;
        RECT 1311.100 587.190 1311.360 587.510 ;
        RECT 1248.600 20.730 1248.740 587.190 ;
        RECT 1245.780 20.410 1246.040 20.730 ;
        RECT 1248.540 20.410 1248.800 20.730 ;
        RECT 1245.840 2.400 1245.980 20.410 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1269.210 591.160 1269.530 591.220 ;
        RECT 1318.430 591.160 1318.750 591.220 ;
        RECT 1269.210 591.020 1318.750 591.160 ;
        RECT 1269.210 590.960 1269.530 591.020 ;
        RECT 1318.430 590.960 1318.750 591.020 ;
        RECT 1263.230 20.640 1263.550 20.700 ;
        RECT 1269.210 20.640 1269.530 20.700 ;
        RECT 1263.230 20.500 1269.530 20.640 ;
        RECT 1263.230 20.440 1263.550 20.500 ;
        RECT 1269.210 20.440 1269.530 20.500 ;
      LAYER via ;
        RECT 1269.240 590.960 1269.500 591.220 ;
        RECT 1318.460 590.960 1318.720 591.220 ;
        RECT 1263.260 20.440 1263.520 20.700 ;
        RECT 1269.240 20.440 1269.500 20.700 ;
      LAYER met2 ;
        RECT 1320.070 600.170 1320.350 604.000 ;
        RECT 1318.520 600.030 1320.350 600.170 ;
        RECT 1318.520 591.250 1318.660 600.030 ;
        RECT 1320.070 600.000 1320.350 600.030 ;
        RECT 1269.240 590.930 1269.500 591.250 ;
        RECT 1318.460 590.930 1318.720 591.250 ;
        RECT 1269.300 20.730 1269.440 590.930 ;
        RECT 1263.260 20.410 1263.520 20.730 ;
        RECT 1269.240 20.410 1269.500 20.730 ;
        RECT 1263.320 2.400 1263.460 20.410 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 591.500 1283.330 591.560 ;
        RECT 1327.630 591.500 1327.950 591.560 ;
        RECT 1283.010 591.360 1327.950 591.500 ;
        RECT 1283.010 591.300 1283.330 591.360 ;
        RECT 1327.630 591.300 1327.950 591.360 ;
      LAYER via ;
        RECT 1283.040 591.300 1283.300 591.560 ;
        RECT 1327.660 591.300 1327.920 591.560 ;
      LAYER met2 ;
        RECT 1329.270 600.170 1329.550 604.000 ;
        RECT 1327.720 600.030 1329.550 600.170 ;
        RECT 1327.720 591.590 1327.860 600.030 ;
        RECT 1329.270 600.000 1329.550 600.030 ;
        RECT 1283.040 591.270 1283.300 591.590 ;
        RECT 1327.660 591.270 1327.920 591.590 ;
        RECT 1283.100 16.730 1283.240 591.270 ;
        RECT 1281.260 16.590 1283.240 16.730 ;
        RECT 1281.260 2.400 1281.400 16.590 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.710 591.840 1304.030 591.900 ;
        RECT 1338.670 591.840 1338.990 591.900 ;
        RECT 1303.710 591.700 1338.990 591.840 ;
        RECT 1303.710 591.640 1304.030 591.700 ;
        RECT 1338.670 591.640 1338.990 591.700 ;
        RECT 1299.110 17.580 1299.430 17.640 ;
        RECT 1303.710 17.580 1304.030 17.640 ;
        RECT 1299.110 17.440 1304.030 17.580 ;
        RECT 1299.110 17.380 1299.430 17.440 ;
        RECT 1303.710 17.380 1304.030 17.440 ;
      LAYER via ;
        RECT 1303.740 591.640 1304.000 591.900 ;
        RECT 1338.700 591.640 1338.960 591.900 ;
        RECT 1299.140 17.380 1299.400 17.640 ;
        RECT 1303.740 17.380 1304.000 17.640 ;
      LAYER met2 ;
        RECT 1338.470 600.000 1338.750 604.000 ;
        RECT 1338.530 598.810 1338.670 600.000 ;
        RECT 1338.530 598.670 1338.900 598.810 ;
        RECT 1338.760 591.930 1338.900 598.670 ;
        RECT 1303.740 591.610 1304.000 591.930 ;
        RECT 1338.700 591.610 1338.960 591.930 ;
        RECT 1303.800 17.670 1303.940 591.610 ;
        RECT 1299.140 17.350 1299.400 17.670 ;
        RECT 1303.740 17.350 1304.000 17.670 ;
        RECT 1299.200 2.400 1299.340 17.350 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.050 589.120 1317.370 589.180 ;
        RECT 1346.030 589.120 1346.350 589.180 ;
        RECT 1317.050 588.980 1346.350 589.120 ;
        RECT 1317.050 588.920 1317.370 588.980 ;
        RECT 1346.030 588.920 1346.350 588.980 ;
      LAYER via ;
        RECT 1317.080 588.920 1317.340 589.180 ;
        RECT 1346.060 588.920 1346.320 589.180 ;
      LAYER met2 ;
        RECT 1347.670 600.170 1347.950 604.000 ;
        RECT 1346.120 600.030 1347.950 600.170 ;
        RECT 1346.120 589.210 1346.260 600.030 ;
        RECT 1347.670 600.000 1347.950 600.030 ;
        RECT 1317.080 588.890 1317.340 589.210 ;
        RECT 1346.060 588.890 1346.320 589.210 ;
        RECT 1317.140 2.400 1317.280 588.890 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 590.820 1338.530 590.880 ;
        RECT 1355.230 590.820 1355.550 590.880 ;
        RECT 1338.210 590.680 1355.550 590.820 ;
        RECT 1338.210 590.620 1338.530 590.680 ;
        RECT 1355.230 590.620 1355.550 590.680 ;
        RECT 1334.990 17.240 1335.310 17.300 ;
        RECT 1338.210 17.240 1338.530 17.300 ;
        RECT 1334.990 17.100 1338.530 17.240 ;
        RECT 1334.990 17.040 1335.310 17.100 ;
        RECT 1338.210 17.040 1338.530 17.100 ;
      LAYER via ;
        RECT 1338.240 590.620 1338.500 590.880 ;
        RECT 1355.260 590.620 1355.520 590.880 ;
        RECT 1335.020 17.040 1335.280 17.300 ;
        RECT 1338.240 17.040 1338.500 17.300 ;
      LAYER met2 ;
        RECT 1356.870 600.170 1357.150 604.000 ;
        RECT 1355.320 600.030 1357.150 600.170 ;
        RECT 1355.320 590.910 1355.460 600.030 ;
        RECT 1356.870 600.000 1357.150 600.030 ;
        RECT 1338.240 590.590 1338.500 590.910 ;
        RECT 1355.260 590.590 1355.520 590.910 ;
        RECT 1338.300 17.330 1338.440 590.590 ;
        RECT 1335.020 17.010 1335.280 17.330 ;
        RECT 1338.240 17.010 1338.500 17.330 ;
        RECT 1335.080 2.400 1335.220 17.010 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1023.110 483.040 1023.430 483.100 ;
        RECT 1024.030 483.040 1024.350 483.100 ;
        RECT 1023.110 482.900 1024.350 483.040 ;
        RECT 1023.110 482.840 1023.430 482.900 ;
        RECT 1024.030 482.840 1024.350 482.900 ;
        RECT 1021.730 386.480 1022.050 386.540 ;
        RECT 1023.110 386.480 1023.430 386.540 ;
        RECT 1021.730 386.340 1023.430 386.480 ;
        RECT 1021.730 386.280 1022.050 386.340 ;
        RECT 1023.110 386.280 1023.430 386.340 ;
        RECT 1021.730 144.740 1022.050 144.800 ;
        RECT 1022.650 144.740 1022.970 144.800 ;
        RECT 1021.730 144.600 1022.970 144.740 ;
        RECT 1021.730 144.540 1022.050 144.600 ;
        RECT 1022.650 144.540 1022.970 144.600 ;
        RECT 1021.730 96.800 1022.050 96.860 ;
        RECT 1022.190 96.800 1022.510 96.860 ;
        RECT 1021.730 96.660 1022.510 96.800 ;
        RECT 1021.730 96.600 1022.050 96.660 ;
        RECT 1022.190 96.600 1022.510 96.660 ;
        RECT 1022.190 62.460 1022.510 62.520 ;
        RECT 1021.820 62.320 1022.510 62.460 ;
        RECT 1021.820 62.180 1021.960 62.320 ;
        RECT 1022.190 62.260 1022.510 62.320 ;
        RECT 1021.730 61.920 1022.050 62.180 ;
        RECT 692.370 44.780 692.690 44.840 ;
        RECT 1021.730 44.780 1022.050 44.840 ;
        RECT 692.370 44.640 1022.050 44.780 ;
        RECT 692.370 44.580 692.690 44.640 ;
        RECT 1021.730 44.580 1022.050 44.640 ;
      LAYER via ;
        RECT 1023.140 482.840 1023.400 483.100 ;
        RECT 1024.060 482.840 1024.320 483.100 ;
        RECT 1021.760 386.280 1022.020 386.540 ;
        RECT 1023.140 386.280 1023.400 386.540 ;
        RECT 1021.760 144.540 1022.020 144.800 ;
        RECT 1022.680 144.540 1022.940 144.800 ;
        RECT 1021.760 96.600 1022.020 96.860 ;
        RECT 1022.220 96.600 1022.480 96.860 ;
        RECT 1022.220 62.260 1022.480 62.520 ;
        RECT 1021.760 61.920 1022.020 62.180 ;
        RECT 692.400 44.580 692.660 44.840 ;
        RECT 1021.760 44.580 1022.020 44.840 ;
      LAYER met2 ;
        RECT 1026.130 600.170 1026.410 604.000 ;
        RECT 1024.580 600.030 1026.410 600.170 ;
        RECT 1024.580 579.885 1024.720 600.030 ;
        RECT 1026.130 600.000 1026.410 600.030 ;
        RECT 1022.670 579.515 1022.950 579.885 ;
        RECT 1024.510 579.515 1024.790 579.885 ;
        RECT 1022.740 497.490 1022.880 579.515 ;
        RECT 1022.280 497.350 1022.880 497.490 ;
        RECT 1022.280 496.810 1022.420 497.350 ;
        RECT 1022.280 496.670 1023.340 496.810 ;
        RECT 1023.200 483.130 1023.340 496.670 ;
        RECT 1023.140 482.810 1023.400 483.130 ;
        RECT 1024.060 482.810 1024.320 483.130 ;
        RECT 1024.120 435.045 1024.260 482.810 ;
        RECT 1023.130 434.675 1023.410 435.045 ;
        RECT 1024.050 434.675 1024.330 435.045 ;
        RECT 1023.200 386.570 1023.340 434.675 ;
        RECT 1021.760 386.250 1022.020 386.570 ;
        RECT 1023.140 386.250 1023.400 386.570 ;
        RECT 1021.820 351.970 1021.960 386.250 ;
        RECT 1021.820 351.830 1022.880 351.970 ;
        RECT 1022.740 317.290 1022.880 351.830 ;
        RECT 1022.280 317.150 1022.880 317.290 ;
        RECT 1022.280 303.010 1022.420 317.150 ;
        RECT 1022.280 302.870 1022.880 303.010 ;
        RECT 1022.740 207.130 1022.880 302.870 ;
        RECT 1022.280 206.990 1022.880 207.130 ;
        RECT 1022.280 206.450 1022.420 206.990 ;
        RECT 1022.280 206.310 1022.880 206.450 ;
        RECT 1022.740 144.830 1022.880 206.310 ;
        RECT 1021.760 144.510 1022.020 144.830 ;
        RECT 1022.680 144.510 1022.940 144.830 ;
        RECT 1021.820 96.890 1021.960 144.510 ;
        RECT 1021.760 96.570 1022.020 96.890 ;
        RECT 1022.220 96.570 1022.480 96.890 ;
        RECT 1022.280 62.550 1022.420 96.570 ;
        RECT 1022.220 62.230 1022.480 62.550 ;
        RECT 1021.760 61.890 1022.020 62.210 ;
        RECT 1021.820 44.870 1021.960 61.890 ;
        RECT 692.400 44.550 692.660 44.870 ;
        RECT 1021.760 44.550 1022.020 44.870 ;
        RECT 692.460 2.400 692.600 44.550 ;
        RECT 692.250 -4.800 692.810 2.400 ;
      LAYER via2 ;
        RECT 1022.670 579.560 1022.950 579.840 ;
        RECT 1024.510 579.560 1024.790 579.840 ;
        RECT 1023.130 434.720 1023.410 435.000 ;
        RECT 1024.050 434.720 1024.330 435.000 ;
      LAYER met3 ;
        RECT 1022.645 579.850 1022.975 579.865 ;
        RECT 1024.485 579.850 1024.815 579.865 ;
        RECT 1022.645 579.550 1024.815 579.850 ;
        RECT 1022.645 579.535 1022.975 579.550 ;
        RECT 1024.485 579.535 1024.815 579.550 ;
        RECT 1023.105 435.010 1023.435 435.025 ;
        RECT 1024.025 435.010 1024.355 435.025 ;
        RECT 1023.105 434.710 1024.355 435.010 ;
        RECT 1023.105 434.695 1023.435 434.710 ;
        RECT 1024.025 434.695 1024.355 434.710 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1358.910 587.420 1359.230 587.480 ;
        RECT 1366.270 587.420 1366.590 587.480 ;
        RECT 1358.910 587.280 1366.590 587.420 ;
        RECT 1358.910 587.220 1359.230 587.280 ;
        RECT 1366.270 587.220 1366.590 587.280 ;
        RECT 1352.470 17.240 1352.790 17.300 ;
        RECT 1358.910 17.240 1359.230 17.300 ;
        RECT 1352.470 17.100 1359.230 17.240 ;
        RECT 1352.470 17.040 1352.790 17.100 ;
        RECT 1358.910 17.040 1359.230 17.100 ;
      LAYER via ;
        RECT 1358.940 587.220 1359.200 587.480 ;
        RECT 1366.300 587.220 1366.560 587.480 ;
        RECT 1352.500 17.040 1352.760 17.300 ;
        RECT 1358.940 17.040 1359.200 17.300 ;
      LAYER met2 ;
        RECT 1366.070 600.000 1366.350 604.000 ;
        RECT 1366.130 598.810 1366.270 600.000 ;
        RECT 1366.130 598.670 1366.500 598.810 ;
        RECT 1366.360 587.510 1366.500 598.670 ;
        RECT 1358.940 587.190 1359.200 587.510 ;
        RECT 1366.300 587.190 1366.560 587.510 ;
        RECT 1359.000 17.330 1359.140 587.190 ;
        RECT 1352.500 17.010 1352.760 17.330 ;
        RECT 1358.940 17.010 1359.200 17.330 ;
        RECT 1352.560 2.400 1352.700 17.010 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.410 20.640 1370.730 20.700 ;
        RECT 1372.710 20.640 1373.030 20.700 ;
        RECT 1370.410 20.500 1373.030 20.640 ;
        RECT 1370.410 20.440 1370.730 20.500 ;
        RECT 1372.710 20.440 1373.030 20.500 ;
      LAYER via ;
        RECT 1370.440 20.440 1370.700 20.700 ;
        RECT 1372.740 20.440 1373.000 20.700 ;
      LAYER met2 ;
        RECT 1375.270 600.170 1375.550 604.000 ;
        RECT 1373.260 600.030 1375.550 600.170 ;
        RECT 1373.260 586.570 1373.400 600.030 ;
        RECT 1375.270 600.000 1375.550 600.030 ;
        RECT 1372.800 586.430 1373.400 586.570 ;
        RECT 1372.800 20.730 1372.940 586.430 ;
        RECT 1370.440 20.410 1370.700 20.730 ;
        RECT 1372.740 20.410 1373.000 20.730 ;
        RECT 1370.500 2.400 1370.640 20.410 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1386.510 20.640 1386.830 20.700 ;
        RECT 1388.350 20.640 1388.670 20.700 ;
        RECT 1386.510 20.500 1388.670 20.640 ;
        RECT 1386.510 20.440 1386.830 20.500 ;
        RECT 1388.350 20.440 1388.670 20.500 ;
      LAYER via ;
        RECT 1386.540 20.440 1386.800 20.700 ;
        RECT 1388.380 20.440 1388.640 20.700 ;
      LAYER met2 ;
        RECT 1384.470 600.170 1384.750 604.000 ;
        RECT 1384.470 600.030 1386.740 600.170 ;
        RECT 1384.470 600.000 1384.750 600.030 ;
        RECT 1386.600 20.730 1386.740 600.030 ;
        RECT 1386.540 20.410 1386.800 20.730 ;
        RECT 1388.380 20.410 1388.640 20.730 ;
        RECT 1388.440 2.400 1388.580 20.410 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1395.250 589.800 1395.570 589.860 ;
        RECT 1401.690 589.800 1402.010 589.860 ;
        RECT 1395.250 589.660 1402.010 589.800 ;
        RECT 1395.250 589.600 1395.570 589.660 ;
        RECT 1401.690 589.600 1402.010 589.660 ;
        RECT 1401.690 2.960 1402.010 3.020 ;
        RECT 1406.290 2.960 1406.610 3.020 ;
        RECT 1401.690 2.820 1406.610 2.960 ;
        RECT 1401.690 2.760 1402.010 2.820 ;
        RECT 1406.290 2.760 1406.610 2.820 ;
      LAYER via ;
        RECT 1395.280 589.600 1395.540 589.860 ;
        RECT 1401.720 589.600 1401.980 589.860 ;
        RECT 1401.720 2.760 1401.980 3.020 ;
        RECT 1406.320 2.760 1406.580 3.020 ;
      LAYER met2 ;
        RECT 1393.670 600.170 1393.950 604.000 ;
        RECT 1393.670 600.030 1395.480 600.170 ;
        RECT 1393.670 600.000 1393.950 600.030 ;
        RECT 1395.340 589.890 1395.480 600.030 ;
        RECT 1395.280 589.570 1395.540 589.890 ;
        RECT 1401.720 589.570 1401.980 589.890 ;
        RECT 1401.780 3.050 1401.920 589.570 ;
        RECT 1401.720 2.730 1401.980 3.050 ;
        RECT 1406.320 2.730 1406.580 3.050 ;
        RECT 1406.380 2.400 1406.520 2.730 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1404.450 589.800 1404.770 589.860 ;
        RECT 1407.210 589.800 1407.530 589.860 ;
        RECT 1404.450 589.660 1407.530 589.800 ;
        RECT 1404.450 589.600 1404.770 589.660 ;
        RECT 1407.210 589.600 1407.530 589.660 ;
        RECT 1407.210 17.580 1407.530 17.640 ;
        RECT 1423.770 17.580 1424.090 17.640 ;
        RECT 1407.210 17.440 1424.090 17.580 ;
        RECT 1407.210 17.380 1407.530 17.440 ;
        RECT 1423.770 17.380 1424.090 17.440 ;
      LAYER via ;
        RECT 1404.480 589.600 1404.740 589.860 ;
        RECT 1407.240 589.600 1407.500 589.860 ;
        RECT 1407.240 17.380 1407.500 17.640 ;
        RECT 1423.800 17.380 1424.060 17.640 ;
      LAYER met2 ;
        RECT 1402.870 600.170 1403.150 604.000 ;
        RECT 1402.870 600.030 1404.680 600.170 ;
        RECT 1402.870 600.000 1403.150 600.030 ;
        RECT 1404.540 589.890 1404.680 600.030 ;
        RECT 1404.480 589.570 1404.740 589.890 ;
        RECT 1407.240 589.570 1407.500 589.890 ;
        RECT 1407.300 17.670 1407.440 589.570 ;
        RECT 1407.240 17.350 1407.500 17.670 ;
        RECT 1423.800 17.350 1424.060 17.670 ;
        RECT 1423.860 2.400 1424.000 17.350 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1413.650 16.560 1413.970 16.620 ;
        RECT 1413.650 16.420 1430.440 16.560 ;
        RECT 1413.650 16.360 1413.970 16.420 ;
        RECT 1430.300 15.880 1430.440 16.420 ;
        RECT 1441.710 15.880 1442.030 15.940 ;
        RECT 1430.300 15.740 1442.030 15.880 ;
        RECT 1441.710 15.680 1442.030 15.740 ;
      LAYER via ;
        RECT 1413.680 16.360 1413.940 16.620 ;
        RECT 1441.740 15.680 1442.000 15.940 ;
      LAYER met2 ;
        RECT 1412.070 600.170 1412.350 604.000 ;
        RECT 1412.070 600.030 1413.880 600.170 ;
        RECT 1412.070 600.000 1412.350 600.030 ;
        RECT 1413.740 16.650 1413.880 600.030 ;
        RECT 1413.680 16.330 1413.940 16.650 ;
        RECT 1441.740 15.650 1442.000 15.970 ;
        RECT 1441.800 2.400 1441.940 15.650 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1422.850 587.080 1423.170 587.140 ;
        RECT 1427.450 587.080 1427.770 587.140 ;
        RECT 1422.850 586.940 1427.770 587.080 ;
        RECT 1422.850 586.880 1423.170 586.940 ;
        RECT 1427.450 586.880 1427.770 586.940 ;
        RECT 1427.450 17.240 1427.770 17.300 ;
        RECT 1459.650 17.240 1459.970 17.300 ;
        RECT 1427.450 17.100 1459.970 17.240 ;
        RECT 1427.450 17.040 1427.770 17.100 ;
        RECT 1459.650 17.040 1459.970 17.100 ;
      LAYER via ;
        RECT 1422.880 586.880 1423.140 587.140 ;
        RECT 1427.480 586.880 1427.740 587.140 ;
        RECT 1427.480 17.040 1427.740 17.300 ;
        RECT 1459.680 17.040 1459.940 17.300 ;
      LAYER met2 ;
        RECT 1421.270 600.170 1421.550 604.000 ;
        RECT 1421.270 600.030 1423.080 600.170 ;
        RECT 1421.270 600.000 1421.550 600.030 ;
        RECT 1422.940 587.170 1423.080 600.030 ;
        RECT 1422.880 586.850 1423.140 587.170 ;
        RECT 1427.480 586.850 1427.740 587.170 ;
        RECT 1427.540 17.330 1427.680 586.850 ;
        RECT 1427.480 17.010 1427.740 17.330 ;
        RECT 1459.680 17.010 1459.940 17.330 ;
        RECT 1459.740 2.400 1459.880 17.010 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1432.050 586.740 1432.370 586.800 ;
        RECT 1434.810 586.740 1435.130 586.800 ;
        RECT 1432.050 586.600 1435.130 586.740 ;
        RECT 1432.050 586.540 1432.370 586.600 ;
        RECT 1434.810 586.540 1435.130 586.600 ;
        RECT 1434.810 19.960 1435.130 20.020 ;
        RECT 1477.590 19.960 1477.910 20.020 ;
        RECT 1434.810 19.820 1477.910 19.960 ;
        RECT 1434.810 19.760 1435.130 19.820 ;
        RECT 1477.590 19.760 1477.910 19.820 ;
      LAYER via ;
        RECT 1432.080 586.540 1432.340 586.800 ;
        RECT 1434.840 586.540 1435.100 586.800 ;
        RECT 1434.840 19.760 1435.100 20.020 ;
        RECT 1477.620 19.760 1477.880 20.020 ;
      LAYER met2 ;
        RECT 1430.470 600.170 1430.750 604.000 ;
        RECT 1430.470 600.030 1432.280 600.170 ;
        RECT 1430.470 600.000 1430.750 600.030 ;
        RECT 1432.140 586.830 1432.280 600.030 ;
        RECT 1432.080 586.510 1432.340 586.830 ;
        RECT 1434.840 586.510 1435.100 586.830 ;
        RECT 1434.900 20.050 1435.040 586.510 ;
        RECT 1434.840 19.730 1435.100 20.050 ;
        RECT 1477.620 19.730 1477.880 20.050 ;
        RECT 1477.680 2.400 1477.820 19.730 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.250 18.940 1441.570 19.000 ;
        RECT 1495.530 18.940 1495.850 19.000 ;
        RECT 1441.250 18.800 1495.850 18.940 ;
        RECT 1441.250 18.740 1441.570 18.800 ;
        RECT 1495.530 18.740 1495.850 18.800 ;
      LAYER via ;
        RECT 1441.280 18.740 1441.540 19.000 ;
        RECT 1495.560 18.740 1495.820 19.000 ;
      LAYER met2 ;
        RECT 1439.670 600.170 1439.950 604.000 ;
        RECT 1439.670 600.030 1441.480 600.170 ;
        RECT 1439.670 600.000 1439.950 600.030 ;
        RECT 1441.340 19.030 1441.480 600.030 ;
        RECT 1441.280 18.710 1441.540 19.030 ;
        RECT 1495.560 18.710 1495.820 19.030 ;
        RECT 1495.620 2.400 1495.760 18.710 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1450.450 586.740 1450.770 586.800 ;
        RECT 1453.670 586.740 1453.990 586.800 ;
        RECT 1450.450 586.600 1453.990 586.740 ;
        RECT 1450.450 586.540 1450.770 586.600 ;
        RECT 1453.670 586.540 1453.990 586.600 ;
        RECT 1455.050 18.600 1455.370 18.660 ;
        RECT 1513.010 18.600 1513.330 18.660 ;
        RECT 1455.050 18.460 1513.330 18.600 ;
        RECT 1455.050 18.400 1455.370 18.460 ;
        RECT 1513.010 18.400 1513.330 18.460 ;
      LAYER via ;
        RECT 1450.480 586.540 1450.740 586.800 ;
        RECT 1453.700 586.540 1453.960 586.800 ;
        RECT 1455.080 18.400 1455.340 18.660 ;
        RECT 1513.040 18.400 1513.300 18.660 ;
      LAYER met2 ;
        RECT 1448.870 600.170 1449.150 604.000 ;
        RECT 1448.870 600.030 1450.680 600.170 ;
        RECT 1448.870 600.000 1449.150 600.030 ;
        RECT 1450.540 586.830 1450.680 600.030 ;
        RECT 1450.480 586.510 1450.740 586.830 ;
        RECT 1453.700 586.510 1453.960 586.830 ;
        RECT 1453.760 582.490 1453.900 586.510 ;
        RECT 1453.760 582.350 1455.280 582.490 ;
        RECT 1455.140 18.690 1455.280 582.350 ;
        RECT 1455.080 18.370 1455.340 18.690 ;
        RECT 1513.040 18.370 1513.300 18.690 ;
        RECT 1513.100 2.400 1513.240 18.370 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 710.310 24.040 710.630 24.100 ;
        RECT 1035.070 24.040 1035.390 24.100 ;
        RECT 710.310 23.900 1035.390 24.040 ;
        RECT 710.310 23.840 710.630 23.900 ;
        RECT 1035.070 23.840 1035.390 23.900 ;
      LAYER via ;
        RECT 710.340 23.840 710.600 24.100 ;
        RECT 1035.100 23.840 1035.360 24.100 ;
      LAYER met2 ;
        RECT 1035.330 600.000 1035.610 604.000 ;
        RECT 1035.390 598.810 1035.530 600.000 ;
        RECT 1035.160 598.670 1035.530 598.810 ;
        RECT 1035.160 24.130 1035.300 598.670 ;
        RECT 710.340 23.810 710.600 24.130 ;
        RECT 1035.100 23.810 1035.360 24.130 ;
        RECT 710.400 2.400 710.540 23.810 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1459.650 586.740 1459.970 586.800 ;
        RECT 1461.950 586.740 1462.270 586.800 ;
        RECT 1459.650 586.600 1462.270 586.740 ;
        RECT 1459.650 586.540 1459.970 586.600 ;
        RECT 1461.950 586.540 1462.270 586.600 ;
        RECT 1530.950 18.600 1531.270 18.660 ;
        RECT 1513.560 18.460 1531.270 18.600 ;
        RECT 1461.950 18.260 1462.270 18.320 ;
        RECT 1513.560 18.260 1513.700 18.460 ;
        RECT 1530.950 18.400 1531.270 18.460 ;
        RECT 1461.950 18.120 1513.700 18.260 ;
        RECT 1461.950 18.060 1462.270 18.120 ;
      LAYER via ;
        RECT 1459.680 586.540 1459.940 586.800 ;
        RECT 1461.980 586.540 1462.240 586.800 ;
        RECT 1461.980 18.060 1462.240 18.320 ;
        RECT 1530.980 18.400 1531.240 18.660 ;
      LAYER met2 ;
        RECT 1458.070 600.170 1458.350 604.000 ;
        RECT 1458.070 600.030 1459.880 600.170 ;
        RECT 1458.070 600.000 1458.350 600.030 ;
        RECT 1459.740 586.830 1459.880 600.030 ;
        RECT 1459.680 586.510 1459.940 586.830 ;
        RECT 1461.980 586.510 1462.240 586.830 ;
        RECT 1462.040 18.350 1462.180 586.510 ;
        RECT 1530.980 18.370 1531.240 18.690 ;
        RECT 1461.980 18.030 1462.240 18.350 ;
        RECT 1531.040 2.400 1531.180 18.370 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1469.310 19.620 1469.630 19.680 ;
        RECT 1548.890 19.620 1549.210 19.680 ;
        RECT 1469.310 19.480 1549.210 19.620 ;
        RECT 1469.310 19.420 1469.630 19.480 ;
        RECT 1548.890 19.420 1549.210 19.480 ;
      LAYER via ;
        RECT 1469.340 19.420 1469.600 19.680 ;
        RECT 1548.920 19.420 1549.180 19.680 ;
      LAYER met2 ;
        RECT 1467.270 600.170 1467.550 604.000 ;
        RECT 1467.270 600.030 1469.540 600.170 ;
        RECT 1467.270 600.000 1467.550 600.030 ;
        RECT 1469.400 19.710 1469.540 600.030 ;
        RECT 1469.340 19.390 1469.600 19.710 ;
        RECT 1548.920 19.390 1549.180 19.710 ;
        RECT 1548.980 2.400 1549.120 19.390 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1478.050 586.740 1478.370 586.800 ;
        RECT 1483.110 586.740 1483.430 586.800 ;
        RECT 1478.050 586.600 1483.430 586.740 ;
        RECT 1478.050 586.540 1478.370 586.600 ;
        RECT 1483.110 586.540 1483.430 586.600 ;
        RECT 1483.110 17.580 1483.430 17.640 ;
        RECT 1483.110 17.440 1543.140 17.580 ;
        RECT 1483.110 17.380 1483.430 17.440 ;
        RECT 1543.000 17.240 1543.140 17.440 ;
        RECT 1566.830 17.240 1567.150 17.300 ;
        RECT 1543.000 17.100 1567.150 17.240 ;
        RECT 1566.830 17.040 1567.150 17.100 ;
      LAYER via ;
        RECT 1478.080 586.540 1478.340 586.800 ;
        RECT 1483.140 586.540 1483.400 586.800 ;
        RECT 1483.140 17.380 1483.400 17.640 ;
        RECT 1566.860 17.040 1567.120 17.300 ;
      LAYER met2 ;
        RECT 1476.470 600.170 1476.750 604.000 ;
        RECT 1476.470 600.030 1478.280 600.170 ;
        RECT 1476.470 600.000 1476.750 600.030 ;
        RECT 1478.140 586.830 1478.280 600.030 ;
        RECT 1478.080 586.510 1478.340 586.830 ;
        RECT 1483.140 586.510 1483.400 586.830 ;
        RECT 1483.200 17.670 1483.340 586.510 ;
        RECT 1483.140 17.350 1483.400 17.670 ;
        RECT 1566.860 17.010 1567.120 17.330 ;
        RECT 1566.920 2.400 1567.060 17.010 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1487.250 586.740 1487.570 586.800 ;
        RECT 1489.550 586.740 1489.870 586.800 ;
        RECT 1487.250 586.600 1489.870 586.740 ;
        RECT 1487.250 586.540 1487.570 586.600 ;
        RECT 1489.550 586.540 1489.870 586.600 ;
        RECT 1489.550 19.960 1489.870 20.020 ;
        RECT 1584.770 19.960 1585.090 20.020 ;
        RECT 1489.550 19.820 1585.090 19.960 ;
        RECT 1489.550 19.760 1489.870 19.820 ;
        RECT 1584.770 19.760 1585.090 19.820 ;
      LAYER via ;
        RECT 1487.280 586.540 1487.540 586.800 ;
        RECT 1489.580 586.540 1489.840 586.800 ;
        RECT 1489.580 19.760 1489.840 20.020 ;
        RECT 1584.800 19.760 1585.060 20.020 ;
      LAYER met2 ;
        RECT 1485.670 600.170 1485.950 604.000 ;
        RECT 1485.670 600.030 1487.480 600.170 ;
        RECT 1485.670 600.000 1485.950 600.030 ;
        RECT 1487.340 586.830 1487.480 600.030 ;
        RECT 1487.280 586.510 1487.540 586.830 ;
        RECT 1489.580 586.510 1489.840 586.830 ;
        RECT 1489.640 20.050 1489.780 586.510 ;
        RECT 1489.580 19.730 1489.840 20.050 ;
        RECT 1584.800 19.730 1585.060 20.050 ;
        RECT 1584.860 2.400 1585.000 19.730 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1496.450 592.520 1496.770 592.580 ;
        RECT 1601.790 592.520 1602.110 592.580 ;
        RECT 1496.450 592.380 1602.110 592.520 ;
        RECT 1496.450 592.320 1496.770 592.380 ;
        RECT 1601.790 592.320 1602.110 592.380 ;
      LAYER via ;
        RECT 1496.480 592.320 1496.740 592.580 ;
        RECT 1601.820 592.320 1602.080 592.580 ;
      LAYER met2 ;
        RECT 1494.870 600.170 1495.150 604.000 ;
        RECT 1494.870 600.030 1496.680 600.170 ;
        RECT 1494.870 600.000 1495.150 600.030 ;
        RECT 1496.540 592.610 1496.680 600.030 ;
        RECT 1496.480 592.290 1496.740 592.610 ;
        RECT 1601.820 592.290 1602.080 592.610 ;
        RECT 1601.880 2.960 1602.020 592.290 ;
        RECT 1601.880 2.820 1602.480 2.960 ;
        RECT 1602.340 2.400 1602.480 2.820 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1505.650 592.860 1505.970 592.920 ;
        RECT 1615.590 592.860 1615.910 592.920 ;
        RECT 1505.650 592.720 1615.910 592.860 ;
        RECT 1505.650 592.660 1505.970 592.720 ;
        RECT 1615.590 592.660 1615.910 592.720 ;
        RECT 1615.590 2.960 1615.910 3.020 ;
        RECT 1620.190 2.960 1620.510 3.020 ;
        RECT 1615.590 2.820 1620.510 2.960 ;
        RECT 1615.590 2.760 1615.910 2.820 ;
        RECT 1620.190 2.760 1620.510 2.820 ;
      LAYER via ;
        RECT 1505.680 592.660 1505.940 592.920 ;
        RECT 1615.620 592.660 1615.880 592.920 ;
        RECT 1615.620 2.760 1615.880 3.020 ;
        RECT 1620.220 2.760 1620.480 3.020 ;
      LAYER met2 ;
        RECT 1504.070 600.170 1504.350 604.000 ;
        RECT 1504.070 600.030 1505.880 600.170 ;
        RECT 1504.070 600.000 1504.350 600.030 ;
        RECT 1505.740 592.950 1505.880 600.030 ;
        RECT 1505.680 592.630 1505.940 592.950 ;
        RECT 1615.620 592.630 1615.880 592.950 ;
        RECT 1615.680 3.050 1615.820 592.630 ;
        RECT 1615.620 2.730 1615.880 3.050 ;
        RECT 1620.220 2.730 1620.480 3.050 ;
        RECT 1620.280 2.400 1620.420 2.730 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1514.850 586.740 1515.170 586.800 ;
        RECT 1517.610 586.740 1517.930 586.800 ;
        RECT 1514.850 586.600 1517.930 586.740 ;
        RECT 1514.850 586.540 1515.170 586.600 ;
        RECT 1517.610 586.540 1517.930 586.600 ;
        RECT 1517.610 26.080 1517.930 26.140 ;
        RECT 1638.130 26.080 1638.450 26.140 ;
        RECT 1517.610 25.940 1638.450 26.080 ;
        RECT 1517.610 25.880 1517.930 25.940 ;
        RECT 1638.130 25.880 1638.450 25.940 ;
      LAYER via ;
        RECT 1514.880 586.540 1515.140 586.800 ;
        RECT 1517.640 586.540 1517.900 586.800 ;
        RECT 1517.640 25.880 1517.900 26.140 ;
        RECT 1638.160 25.880 1638.420 26.140 ;
      LAYER met2 ;
        RECT 1513.270 600.170 1513.550 604.000 ;
        RECT 1513.270 600.030 1515.080 600.170 ;
        RECT 1513.270 600.000 1513.550 600.030 ;
        RECT 1514.940 586.830 1515.080 600.030 ;
        RECT 1514.880 586.510 1515.140 586.830 ;
        RECT 1517.640 586.510 1517.900 586.830 ;
        RECT 1517.700 26.170 1517.840 586.510 ;
        RECT 1517.640 25.850 1517.900 26.170 ;
        RECT 1638.160 25.850 1638.420 26.170 ;
        RECT 1638.220 2.400 1638.360 25.850 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1524.510 25.400 1524.830 25.460 ;
        RECT 1656.070 25.400 1656.390 25.460 ;
        RECT 1524.510 25.260 1656.390 25.400 ;
        RECT 1524.510 25.200 1524.830 25.260 ;
        RECT 1656.070 25.200 1656.390 25.260 ;
      LAYER via ;
        RECT 1524.540 25.200 1524.800 25.460 ;
        RECT 1656.100 25.200 1656.360 25.460 ;
      LAYER met2 ;
        RECT 1522.470 600.170 1522.750 604.000 ;
        RECT 1522.470 600.030 1524.740 600.170 ;
        RECT 1522.470 600.000 1522.750 600.030 ;
        RECT 1524.600 25.490 1524.740 600.030 ;
        RECT 1524.540 25.170 1524.800 25.490 ;
        RECT 1656.100 25.170 1656.360 25.490 ;
        RECT 1656.160 2.400 1656.300 25.170 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1533.250 586.740 1533.570 586.800 ;
        RECT 1538.310 586.740 1538.630 586.800 ;
        RECT 1533.250 586.600 1538.630 586.740 ;
        RECT 1533.250 586.540 1533.570 586.600 ;
        RECT 1538.310 586.540 1538.630 586.600 ;
        RECT 1538.310 25.740 1538.630 25.800 ;
        RECT 1673.550 25.740 1673.870 25.800 ;
        RECT 1538.310 25.600 1673.870 25.740 ;
        RECT 1538.310 25.540 1538.630 25.600 ;
        RECT 1673.550 25.540 1673.870 25.600 ;
      LAYER via ;
        RECT 1533.280 586.540 1533.540 586.800 ;
        RECT 1538.340 586.540 1538.600 586.800 ;
        RECT 1538.340 25.540 1538.600 25.800 ;
        RECT 1673.580 25.540 1673.840 25.800 ;
      LAYER met2 ;
        RECT 1531.670 600.170 1531.950 604.000 ;
        RECT 1531.670 600.030 1533.480 600.170 ;
        RECT 1531.670 600.000 1531.950 600.030 ;
        RECT 1533.340 586.830 1533.480 600.030 ;
        RECT 1533.280 586.510 1533.540 586.830 ;
        RECT 1538.340 586.510 1538.600 586.830 ;
        RECT 1538.400 25.830 1538.540 586.510 ;
        RECT 1538.340 25.510 1538.600 25.830 ;
        RECT 1673.580 25.510 1673.840 25.830 ;
        RECT 1673.640 2.400 1673.780 25.510 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1542.450 588.100 1542.770 588.160 ;
        RECT 1544.750 588.100 1545.070 588.160 ;
        RECT 1542.450 587.960 1545.070 588.100 ;
        RECT 1542.450 587.900 1542.770 587.960 ;
        RECT 1544.750 587.900 1545.070 587.960 ;
        RECT 1544.750 25.060 1545.070 25.120 ;
        RECT 1691.490 25.060 1691.810 25.120 ;
        RECT 1544.750 24.920 1691.810 25.060 ;
        RECT 1544.750 24.860 1545.070 24.920 ;
        RECT 1691.490 24.860 1691.810 24.920 ;
      LAYER via ;
        RECT 1542.480 587.900 1542.740 588.160 ;
        RECT 1544.780 587.900 1545.040 588.160 ;
        RECT 1544.780 24.860 1545.040 25.120 ;
        RECT 1691.520 24.860 1691.780 25.120 ;
      LAYER met2 ;
        RECT 1540.870 600.170 1541.150 604.000 ;
        RECT 1540.870 600.030 1542.680 600.170 ;
        RECT 1540.870 600.000 1541.150 600.030 ;
        RECT 1542.540 588.190 1542.680 600.030 ;
        RECT 1542.480 587.870 1542.740 588.190 ;
        RECT 1544.780 587.870 1545.040 588.190 ;
        RECT 1544.840 25.150 1544.980 587.870 ;
        RECT 1544.780 24.830 1545.040 25.150 ;
        RECT 1691.520 24.830 1691.780 25.150 ;
        RECT 1691.580 2.400 1691.720 24.830 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1041.970 583.000 1042.290 583.060 ;
        RECT 1043.350 583.000 1043.670 583.060 ;
        RECT 1041.970 582.860 1043.670 583.000 ;
        RECT 1041.970 582.800 1042.290 582.860 ;
        RECT 1043.350 582.800 1043.670 582.860 ;
        RECT 728.250 24.380 728.570 24.440 ;
        RECT 1041.970 24.380 1042.290 24.440 ;
        RECT 728.250 24.240 1042.290 24.380 ;
        RECT 728.250 24.180 728.570 24.240 ;
        RECT 1041.970 24.180 1042.290 24.240 ;
      LAYER via ;
        RECT 1042.000 582.800 1042.260 583.060 ;
        RECT 1043.380 582.800 1043.640 583.060 ;
        RECT 728.280 24.180 728.540 24.440 ;
        RECT 1042.000 24.180 1042.260 24.440 ;
      LAYER met2 ;
        RECT 1044.530 600.170 1044.810 604.000 ;
        RECT 1043.440 600.030 1044.810 600.170 ;
        RECT 1043.440 583.090 1043.580 600.030 ;
        RECT 1044.530 600.000 1044.810 600.030 ;
        RECT 1042.000 582.770 1042.260 583.090 ;
        RECT 1043.380 582.770 1043.640 583.090 ;
        RECT 1042.060 24.470 1042.200 582.770 ;
        RECT 728.280 24.150 728.540 24.470 ;
        RECT 1042.000 24.150 1042.260 24.470 ;
        RECT 728.340 2.400 728.480 24.150 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1552.110 24.720 1552.430 24.780 ;
        RECT 1709.430 24.720 1709.750 24.780 ;
        RECT 1552.110 24.580 1709.750 24.720 ;
        RECT 1552.110 24.520 1552.430 24.580 ;
        RECT 1709.430 24.520 1709.750 24.580 ;
      LAYER via ;
        RECT 1552.140 24.520 1552.400 24.780 ;
        RECT 1709.460 24.520 1709.720 24.780 ;
      LAYER met2 ;
        RECT 1550.070 600.170 1550.350 604.000 ;
        RECT 1550.070 600.030 1552.340 600.170 ;
        RECT 1550.070 600.000 1550.350 600.030 ;
        RECT 1552.200 24.810 1552.340 600.030 ;
        RECT 1552.140 24.490 1552.400 24.810 ;
        RECT 1709.460 24.490 1709.720 24.810 ;
        RECT 1709.520 2.400 1709.660 24.490 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1559.010 24.380 1559.330 24.440 ;
        RECT 1727.370 24.380 1727.690 24.440 ;
        RECT 1559.010 24.240 1727.690 24.380 ;
        RECT 1559.010 24.180 1559.330 24.240 ;
        RECT 1727.370 24.180 1727.690 24.240 ;
      LAYER via ;
        RECT 1559.040 24.180 1559.300 24.440 ;
        RECT 1727.400 24.180 1727.660 24.440 ;
      LAYER met2 ;
        RECT 1558.810 600.000 1559.090 604.000 ;
        RECT 1558.870 598.810 1559.010 600.000 ;
        RECT 1558.870 598.670 1559.240 598.810 ;
        RECT 1559.100 24.470 1559.240 598.670 ;
        RECT 1559.040 24.150 1559.300 24.470 ;
        RECT 1727.400 24.150 1727.660 24.470 ;
        RECT 1727.460 2.400 1727.600 24.150 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1569.590 586.740 1569.910 586.800 ;
        RECT 1572.810 586.740 1573.130 586.800 ;
        RECT 1569.590 586.600 1573.130 586.740 ;
        RECT 1569.590 586.540 1569.910 586.600 ;
        RECT 1572.810 586.540 1573.130 586.600 ;
        RECT 1572.810 24.040 1573.130 24.100 ;
        RECT 1745.310 24.040 1745.630 24.100 ;
        RECT 1572.810 23.900 1745.630 24.040 ;
        RECT 1572.810 23.840 1573.130 23.900 ;
        RECT 1745.310 23.840 1745.630 23.900 ;
      LAYER via ;
        RECT 1569.620 586.540 1569.880 586.800 ;
        RECT 1572.840 586.540 1573.100 586.800 ;
        RECT 1572.840 23.840 1573.100 24.100 ;
        RECT 1745.340 23.840 1745.600 24.100 ;
      LAYER met2 ;
        RECT 1568.010 600.170 1568.290 604.000 ;
        RECT 1568.010 600.030 1569.820 600.170 ;
        RECT 1568.010 600.000 1568.290 600.030 ;
        RECT 1569.680 586.830 1569.820 600.030 ;
        RECT 1569.620 586.510 1569.880 586.830 ;
        RECT 1572.840 586.510 1573.100 586.830 ;
        RECT 1572.900 24.130 1573.040 586.510 ;
        RECT 1572.840 23.810 1573.100 24.130 ;
        RECT 1745.340 23.810 1745.600 24.130 ;
        RECT 1745.400 2.400 1745.540 23.810 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1579.250 29.140 1579.570 29.200 ;
        RECT 1762.790 29.140 1763.110 29.200 ;
        RECT 1579.250 29.000 1763.110 29.140 ;
        RECT 1579.250 28.940 1579.570 29.000 ;
        RECT 1762.790 28.940 1763.110 29.000 ;
      LAYER via ;
        RECT 1579.280 28.940 1579.540 29.200 ;
        RECT 1762.820 28.940 1763.080 29.200 ;
      LAYER met2 ;
        RECT 1577.210 600.170 1577.490 604.000 ;
        RECT 1577.210 600.030 1579.480 600.170 ;
        RECT 1577.210 600.000 1577.490 600.030 ;
        RECT 1579.340 29.230 1579.480 600.030 ;
        RECT 1579.280 28.910 1579.540 29.230 ;
        RECT 1762.820 28.910 1763.080 29.230 ;
        RECT 1762.880 2.400 1763.020 28.910 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1586.610 30.160 1586.930 30.220 ;
        RECT 1780.730 30.160 1781.050 30.220 ;
        RECT 1586.610 30.020 1781.050 30.160 ;
        RECT 1586.610 29.960 1586.930 30.020 ;
        RECT 1780.730 29.960 1781.050 30.020 ;
      LAYER via ;
        RECT 1586.640 29.960 1586.900 30.220 ;
        RECT 1780.760 29.960 1781.020 30.220 ;
      LAYER met2 ;
        RECT 1586.410 600.000 1586.690 604.000 ;
        RECT 1586.470 598.810 1586.610 600.000 ;
        RECT 1586.470 598.670 1586.840 598.810 ;
        RECT 1586.700 30.250 1586.840 598.670 ;
        RECT 1586.640 29.930 1586.900 30.250 ;
        RECT 1780.760 29.930 1781.020 30.250 ;
        RECT 1780.820 2.400 1780.960 29.930 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1597.190 586.740 1597.510 586.800 ;
        RECT 1600.410 586.740 1600.730 586.800 ;
        RECT 1597.190 586.600 1600.730 586.740 ;
        RECT 1597.190 586.540 1597.510 586.600 ;
        RECT 1600.410 586.540 1600.730 586.600 ;
        RECT 1600.410 29.820 1600.730 29.880 ;
        RECT 1798.670 29.820 1798.990 29.880 ;
        RECT 1600.410 29.680 1798.990 29.820 ;
        RECT 1600.410 29.620 1600.730 29.680 ;
        RECT 1798.670 29.620 1798.990 29.680 ;
      LAYER via ;
        RECT 1597.220 586.540 1597.480 586.800 ;
        RECT 1600.440 586.540 1600.700 586.800 ;
        RECT 1600.440 29.620 1600.700 29.880 ;
        RECT 1798.700 29.620 1798.960 29.880 ;
      LAYER met2 ;
        RECT 1595.610 600.170 1595.890 604.000 ;
        RECT 1595.610 600.030 1597.420 600.170 ;
        RECT 1595.610 600.000 1595.890 600.030 ;
        RECT 1597.280 586.830 1597.420 600.030 ;
        RECT 1597.220 586.510 1597.480 586.830 ;
        RECT 1600.440 586.510 1600.700 586.830 ;
        RECT 1600.500 29.910 1600.640 586.510 ;
        RECT 1600.440 29.590 1600.700 29.910 ;
        RECT 1798.700 29.590 1798.960 29.910 ;
        RECT 1798.760 2.400 1798.900 29.590 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 33.900 1607.630 33.960 ;
        RECT 1816.610 33.900 1816.930 33.960 ;
        RECT 1607.310 33.760 1816.930 33.900 ;
        RECT 1607.310 33.700 1607.630 33.760 ;
        RECT 1816.610 33.700 1816.930 33.760 ;
      LAYER via ;
        RECT 1607.340 33.700 1607.600 33.960 ;
        RECT 1816.640 33.700 1816.900 33.960 ;
      LAYER met2 ;
        RECT 1604.810 600.170 1605.090 604.000 ;
        RECT 1604.810 600.030 1607.540 600.170 ;
        RECT 1604.810 600.000 1605.090 600.030 ;
        RECT 1607.400 33.990 1607.540 600.030 ;
        RECT 1607.340 33.670 1607.600 33.990 ;
        RECT 1816.640 33.670 1816.900 33.990 ;
        RECT 1816.700 2.400 1816.840 33.670 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1613.750 33.220 1614.070 33.280 ;
        RECT 1834.550 33.220 1834.870 33.280 ;
        RECT 1613.750 33.080 1834.870 33.220 ;
        RECT 1613.750 33.020 1614.070 33.080 ;
        RECT 1834.550 33.020 1834.870 33.080 ;
      LAYER via ;
        RECT 1613.780 33.020 1614.040 33.280 ;
        RECT 1834.580 33.020 1834.840 33.280 ;
      LAYER met2 ;
        RECT 1614.010 600.000 1614.290 604.000 ;
        RECT 1614.070 598.810 1614.210 600.000 ;
        RECT 1613.840 598.670 1614.210 598.810 ;
        RECT 1613.840 33.310 1613.980 598.670 ;
        RECT 1613.780 32.990 1614.040 33.310 ;
        RECT 1834.580 32.990 1834.840 33.310 ;
        RECT 1834.640 2.400 1834.780 32.990 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1624.790 586.740 1625.110 586.800 ;
        RECT 1627.550 586.740 1627.870 586.800 ;
        RECT 1624.790 586.600 1627.870 586.740 ;
        RECT 1624.790 586.540 1625.110 586.600 ;
        RECT 1627.550 586.540 1627.870 586.600 ;
        RECT 1627.550 32.540 1627.870 32.600 ;
        RECT 1852.030 32.540 1852.350 32.600 ;
        RECT 1627.550 32.400 1852.350 32.540 ;
        RECT 1627.550 32.340 1627.870 32.400 ;
        RECT 1852.030 32.340 1852.350 32.400 ;
      LAYER via ;
        RECT 1624.820 586.540 1625.080 586.800 ;
        RECT 1627.580 586.540 1627.840 586.800 ;
        RECT 1627.580 32.340 1627.840 32.600 ;
        RECT 1852.060 32.340 1852.320 32.600 ;
      LAYER met2 ;
        RECT 1623.210 600.170 1623.490 604.000 ;
        RECT 1623.210 600.030 1625.020 600.170 ;
        RECT 1623.210 600.000 1623.490 600.030 ;
        RECT 1624.880 586.830 1625.020 600.030 ;
        RECT 1624.820 586.510 1625.080 586.830 ;
        RECT 1627.580 586.510 1627.840 586.830 ;
        RECT 1627.640 32.630 1627.780 586.510 ;
        RECT 1627.580 32.310 1627.840 32.630 ;
        RECT 1852.060 32.310 1852.320 32.630 ;
        RECT 1852.120 2.400 1852.260 32.310 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1634.450 32.200 1634.770 32.260 ;
        RECT 1869.970 32.200 1870.290 32.260 ;
        RECT 1634.450 32.060 1870.290 32.200 ;
        RECT 1634.450 32.000 1634.770 32.060 ;
        RECT 1869.970 32.000 1870.290 32.060 ;
      LAYER via ;
        RECT 1634.480 32.000 1634.740 32.260 ;
        RECT 1870.000 32.000 1870.260 32.260 ;
      LAYER met2 ;
        RECT 1632.410 600.170 1632.690 604.000 ;
        RECT 1632.410 600.030 1634.680 600.170 ;
        RECT 1632.410 600.000 1632.690 600.030 ;
        RECT 1634.540 32.290 1634.680 600.030 ;
        RECT 1634.480 31.970 1634.740 32.290 ;
        RECT 1870.000 31.970 1870.260 32.290 ;
        RECT 1870.060 2.400 1870.200 31.970 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1049.790 483.040 1050.110 483.100 ;
        RECT 1050.710 483.040 1051.030 483.100 ;
        RECT 1049.790 482.900 1051.030 483.040 ;
        RECT 1049.790 482.840 1050.110 482.900 ;
        RECT 1050.710 482.840 1051.030 482.900 ;
        RECT 1049.330 338.200 1049.650 338.260 ;
        RECT 1049.790 338.200 1050.110 338.260 ;
        RECT 1049.330 338.060 1050.110 338.200 ;
        RECT 1049.330 338.000 1049.650 338.060 ;
        RECT 1049.790 338.000 1050.110 338.060 ;
        RECT 1048.410 289.580 1048.730 289.640 ;
        RECT 1049.790 289.580 1050.110 289.640 ;
        RECT 1048.410 289.440 1050.110 289.580 ;
        RECT 1048.410 289.380 1048.730 289.440 ;
        RECT 1049.790 289.380 1050.110 289.440 ;
        RECT 1047.950 145.080 1048.270 145.140 ;
        RECT 1049.790 145.080 1050.110 145.140 ;
        RECT 1047.950 144.940 1050.110 145.080 ;
        RECT 1047.950 144.880 1048.270 144.940 ;
        RECT 1049.790 144.880 1050.110 144.940 ;
        RECT 1047.950 96.800 1048.270 96.860 ;
        RECT 1048.870 96.800 1049.190 96.860 ;
        RECT 1047.950 96.660 1049.190 96.800 ;
        RECT 1047.950 96.600 1048.270 96.660 ;
        RECT 1048.870 96.600 1049.190 96.660 ;
        RECT 800.010 25.740 800.330 25.800 ;
        RECT 1049.330 25.740 1049.650 25.800 ;
        RECT 800.010 25.600 1049.650 25.740 ;
        RECT 800.010 25.540 800.330 25.600 ;
        RECT 1049.330 25.540 1049.650 25.600 ;
        RECT 746.190 17.240 746.510 17.300 ;
        RECT 800.010 17.240 800.330 17.300 ;
        RECT 746.190 17.100 800.330 17.240 ;
        RECT 746.190 17.040 746.510 17.100 ;
        RECT 800.010 17.040 800.330 17.100 ;
      LAYER via ;
        RECT 1049.820 482.840 1050.080 483.100 ;
        RECT 1050.740 482.840 1051.000 483.100 ;
        RECT 1049.360 338.000 1049.620 338.260 ;
        RECT 1049.820 338.000 1050.080 338.260 ;
        RECT 1048.440 289.380 1048.700 289.640 ;
        RECT 1049.820 289.380 1050.080 289.640 ;
        RECT 1047.980 144.880 1048.240 145.140 ;
        RECT 1049.820 144.880 1050.080 145.140 ;
        RECT 1047.980 96.600 1048.240 96.860 ;
        RECT 1048.900 96.600 1049.160 96.860 ;
        RECT 800.040 25.540 800.300 25.800 ;
        RECT 1049.360 25.540 1049.620 25.800 ;
        RECT 746.220 17.040 746.480 17.300 ;
        RECT 800.040 17.040 800.300 17.300 ;
      LAYER met2 ;
        RECT 1053.730 600.170 1054.010 604.000 ;
        RECT 1052.180 600.030 1054.010 600.170 ;
        RECT 1052.180 583.170 1052.320 600.030 ;
        RECT 1053.730 600.000 1054.010 600.030 ;
        RECT 1049.420 583.030 1052.320 583.170 ;
        RECT 1049.420 497.490 1049.560 583.030 ;
        RECT 1048.960 497.350 1049.560 497.490 ;
        RECT 1048.960 496.810 1049.100 497.350 ;
        RECT 1048.960 496.670 1050.020 496.810 ;
        RECT 1049.880 483.130 1050.020 496.670 ;
        RECT 1049.820 482.810 1050.080 483.130 ;
        RECT 1050.740 482.810 1051.000 483.130 ;
        RECT 1050.800 435.045 1050.940 482.810 ;
        RECT 1049.810 434.675 1050.090 435.045 ;
        RECT 1050.730 434.675 1051.010 435.045 ;
        RECT 1049.880 338.290 1050.020 434.675 ;
        RECT 1049.360 337.970 1049.620 338.290 ;
        RECT 1049.820 337.970 1050.080 338.290 ;
        RECT 1049.420 303.690 1049.560 337.970 ;
        RECT 1049.420 303.550 1050.020 303.690 ;
        RECT 1049.880 289.670 1050.020 303.550 ;
        RECT 1048.440 289.350 1048.700 289.670 ;
        RECT 1049.820 289.350 1050.080 289.670 ;
        RECT 1048.500 254.730 1048.640 289.350 ;
        RECT 1048.500 254.590 1049.560 254.730 ;
        RECT 1049.420 207.130 1049.560 254.590 ;
        RECT 1049.420 206.990 1050.020 207.130 ;
        RECT 1049.880 145.170 1050.020 206.990 ;
        RECT 1047.980 144.850 1048.240 145.170 ;
        RECT 1049.820 144.850 1050.080 145.170 ;
        RECT 1048.040 96.890 1048.180 144.850 ;
        RECT 1047.980 96.570 1048.240 96.890 ;
        RECT 1048.900 96.570 1049.160 96.890 ;
        RECT 1048.960 96.290 1049.100 96.570 ;
        RECT 1048.960 96.150 1049.560 96.290 ;
        RECT 1049.420 25.830 1049.560 96.150 ;
        RECT 800.040 25.510 800.300 25.830 ;
        RECT 1049.360 25.510 1049.620 25.830 ;
        RECT 800.100 17.330 800.240 25.510 ;
        RECT 746.220 17.010 746.480 17.330 ;
        RECT 800.040 17.010 800.300 17.330 ;
        RECT 746.280 2.400 746.420 17.010 ;
        RECT 746.070 -4.800 746.630 2.400 ;
      LAYER via2 ;
        RECT 1049.810 434.720 1050.090 435.000 ;
        RECT 1050.730 434.720 1051.010 435.000 ;
      LAYER met3 ;
        RECT 1049.785 435.010 1050.115 435.025 ;
        RECT 1050.705 435.010 1051.035 435.025 ;
        RECT 1049.785 434.710 1051.035 435.010 ;
        RECT 1049.785 434.695 1050.115 434.710 ;
        RECT 1050.705 434.695 1051.035 434.710 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1641.350 31.860 1641.670 31.920 ;
        RECT 1887.910 31.860 1888.230 31.920 ;
        RECT 1641.350 31.720 1888.230 31.860 ;
        RECT 1641.350 31.660 1641.670 31.720 ;
        RECT 1887.910 31.660 1888.230 31.720 ;
      LAYER via ;
        RECT 1641.380 31.660 1641.640 31.920 ;
        RECT 1887.940 31.660 1888.200 31.920 ;
      LAYER met2 ;
        RECT 1641.610 600.000 1641.890 604.000 ;
        RECT 1641.670 598.810 1641.810 600.000 ;
        RECT 1641.440 598.670 1641.810 598.810 ;
        RECT 1641.440 31.950 1641.580 598.670 ;
        RECT 1641.380 31.630 1641.640 31.950 ;
        RECT 1887.940 31.630 1888.200 31.950 ;
        RECT 1888.000 2.400 1888.140 31.630 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1652.390 586.740 1652.710 586.800 ;
        RECT 1655.610 586.740 1655.930 586.800 ;
        RECT 1652.390 586.600 1655.930 586.740 ;
        RECT 1652.390 586.540 1652.710 586.600 ;
        RECT 1655.610 586.540 1655.930 586.600 ;
        RECT 1655.610 31.520 1655.930 31.580 ;
        RECT 1905.850 31.520 1906.170 31.580 ;
        RECT 1655.610 31.380 1906.170 31.520 ;
        RECT 1655.610 31.320 1655.930 31.380 ;
        RECT 1905.850 31.320 1906.170 31.380 ;
      LAYER via ;
        RECT 1652.420 586.540 1652.680 586.800 ;
        RECT 1655.640 586.540 1655.900 586.800 ;
        RECT 1655.640 31.320 1655.900 31.580 ;
        RECT 1905.880 31.320 1906.140 31.580 ;
      LAYER met2 ;
        RECT 1650.810 600.170 1651.090 604.000 ;
        RECT 1650.810 600.030 1652.620 600.170 ;
        RECT 1650.810 600.000 1651.090 600.030 ;
        RECT 1652.480 586.830 1652.620 600.030 ;
        RECT 1652.420 586.510 1652.680 586.830 ;
        RECT 1655.640 586.510 1655.900 586.830 ;
        RECT 1655.700 31.610 1655.840 586.510 ;
        RECT 1655.640 31.290 1655.900 31.610 ;
        RECT 1905.880 31.290 1906.140 31.610 ;
        RECT 1905.940 2.400 1906.080 31.290 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.050 31.180 1662.370 31.240 ;
        RECT 1923.330 31.180 1923.650 31.240 ;
        RECT 1662.050 31.040 1923.650 31.180 ;
        RECT 1662.050 30.980 1662.370 31.040 ;
        RECT 1923.330 30.980 1923.650 31.040 ;
      LAYER via ;
        RECT 1662.080 30.980 1662.340 31.240 ;
        RECT 1923.360 30.980 1923.620 31.240 ;
      LAYER met2 ;
        RECT 1660.010 600.170 1660.290 604.000 ;
        RECT 1660.010 600.030 1662.280 600.170 ;
        RECT 1660.010 600.000 1660.290 600.030 ;
        RECT 1662.140 31.270 1662.280 600.030 ;
        RECT 1662.080 30.950 1662.340 31.270 ;
        RECT 1923.360 30.950 1923.620 31.270 ;
        RECT 1923.420 2.400 1923.560 30.950 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1668.490 30.840 1668.810 30.900 ;
        RECT 1941.270 30.840 1941.590 30.900 ;
        RECT 1668.490 30.700 1941.590 30.840 ;
        RECT 1668.490 30.640 1668.810 30.700 ;
        RECT 1941.270 30.640 1941.590 30.700 ;
      LAYER via ;
        RECT 1668.520 30.640 1668.780 30.900 ;
        RECT 1941.300 30.640 1941.560 30.900 ;
      LAYER met2 ;
        RECT 1669.210 600.170 1669.490 604.000 ;
        RECT 1668.580 600.030 1669.490 600.170 ;
        RECT 1668.580 30.930 1668.720 600.030 ;
        RECT 1669.210 600.000 1669.490 600.030 ;
        RECT 1668.520 30.610 1668.780 30.930 ;
        RECT 1941.300 30.610 1941.560 30.930 ;
        RECT 1941.360 2.400 1941.500 30.610 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1679.990 592.180 1680.310 592.240 ;
        RECT 1742.090 592.180 1742.410 592.240 ;
        RECT 1679.990 592.040 1742.410 592.180 ;
        RECT 1679.990 591.980 1680.310 592.040 ;
        RECT 1742.090 591.980 1742.410 592.040 ;
        RECT 1800.970 34.580 1801.290 34.640 ;
        RECT 1800.970 34.440 1811.320 34.580 ;
        RECT 1800.970 34.380 1801.290 34.440 ;
        RECT 1811.180 34.240 1811.320 34.440 ;
        RECT 1859.480 34.440 1883.540 34.580 ;
        RECT 1859.480 34.240 1859.620 34.440 ;
        RECT 1811.180 34.100 1859.620 34.240 ;
        RECT 1883.400 34.240 1883.540 34.440 ;
        RECT 1883.770 34.380 1884.090 34.640 ;
        RECT 1883.860 34.240 1884.000 34.380 ;
        RECT 1883.400 34.100 1884.000 34.240 ;
        RECT 1898.030 33.900 1898.350 33.960 ;
        RECT 1936.210 33.900 1936.530 33.960 ;
        RECT 1898.030 33.760 1936.530 33.900 ;
        RECT 1898.030 33.700 1898.350 33.760 ;
        RECT 1936.210 33.700 1936.530 33.760 ;
        RECT 1772.450 33.560 1772.770 33.620 ;
        RECT 1800.970 33.560 1801.290 33.620 ;
        RECT 1772.450 33.420 1801.290 33.560 ;
        RECT 1772.450 33.360 1772.770 33.420 ;
        RECT 1800.970 33.360 1801.290 33.420 ;
        RECT 1936.210 32.540 1936.530 32.600 ;
        RECT 1959.210 32.540 1959.530 32.600 ;
        RECT 1936.210 32.400 1959.530 32.540 ;
        RECT 1936.210 32.340 1936.530 32.400 ;
        RECT 1959.210 32.340 1959.530 32.400 ;
        RECT 1742.090 28.800 1742.410 28.860 ;
        RECT 1772.450 28.800 1772.770 28.860 ;
        RECT 1742.090 28.660 1772.770 28.800 ;
        RECT 1742.090 28.600 1742.410 28.660 ;
        RECT 1772.450 28.600 1772.770 28.660 ;
      LAYER via ;
        RECT 1680.020 591.980 1680.280 592.240 ;
        RECT 1742.120 591.980 1742.380 592.240 ;
        RECT 1801.000 34.380 1801.260 34.640 ;
        RECT 1883.800 34.380 1884.060 34.640 ;
        RECT 1898.060 33.700 1898.320 33.960 ;
        RECT 1936.240 33.700 1936.500 33.960 ;
        RECT 1772.480 33.360 1772.740 33.620 ;
        RECT 1801.000 33.360 1801.260 33.620 ;
        RECT 1936.240 32.340 1936.500 32.600 ;
        RECT 1959.240 32.340 1959.500 32.600 ;
        RECT 1742.120 28.600 1742.380 28.860 ;
        RECT 1772.480 28.600 1772.740 28.860 ;
      LAYER met2 ;
        RECT 1678.410 600.170 1678.690 604.000 ;
        RECT 1678.410 600.030 1680.220 600.170 ;
        RECT 1678.410 600.000 1678.690 600.030 ;
        RECT 1680.080 592.270 1680.220 600.030 ;
        RECT 1680.020 591.950 1680.280 592.270 ;
        RECT 1742.120 591.950 1742.380 592.270 ;
        RECT 1742.180 28.890 1742.320 591.950 ;
        RECT 1801.000 34.350 1801.260 34.670 ;
        RECT 1883.800 34.525 1884.060 34.670 ;
        RECT 1801.060 33.650 1801.200 34.350 ;
        RECT 1883.790 34.155 1884.070 34.525 ;
        RECT 1898.050 34.155 1898.330 34.525 ;
        RECT 1898.120 33.990 1898.260 34.155 ;
        RECT 1898.060 33.670 1898.320 33.990 ;
        RECT 1936.240 33.670 1936.500 33.990 ;
        RECT 1772.480 33.330 1772.740 33.650 ;
        RECT 1801.000 33.330 1801.260 33.650 ;
        RECT 1772.540 28.890 1772.680 33.330 ;
        RECT 1936.300 32.630 1936.440 33.670 ;
        RECT 1936.240 32.310 1936.500 32.630 ;
        RECT 1959.240 32.310 1959.500 32.630 ;
        RECT 1742.120 28.570 1742.380 28.890 ;
        RECT 1772.480 28.570 1772.740 28.890 ;
        RECT 1959.300 2.400 1959.440 32.310 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
      LAYER via2 ;
        RECT 1883.790 34.200 1884.070 34.480 ;
        RECT 1898.050 34.200 1898.330 34.480 ;
      LAYER met3 ;
        RECT 1883.765 34.490 1884.095 34.505 ;
        RECT 1898.025 34.490 1898.355 34.505 ;
        RECT 1883.765 34.190 1898.355 34.490 ;
        RECT 1883.765 34.175 1884.095 34.190 ;
        RECT 1898.025 34.175 1898.355 34.190 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1689.190 591.500 1689.510 591.560 ;
        RECT 1755.890 591.500 1756.210 591.560 ;
        RECT 1689.190 591.360 1756.210 591.500 ;
        RECT 1689.190 591.300 1689.510 591.360 ;
        RECT 1755.890 591.300 1756.210 591.360 ;
        RECT 1755.890 32.880 1756.210 32.940 ;
        RECT 1977.150 32.880 1977.470 32.940 ;
        RECT 1755.890 32.740 1977.470 32.880 ;
        RECT 1755.890 32.680 1756.210 32.740 ;
        RECT 1977.150 32.680 1977.470 32.740 ;
      LAYER via ;
        RECT 1689.220 591.300 1689.480 591.560 ;
        RECT 1755.920 591.300 1756.180 591.560 ;
        RECT 1755.920 32.680 1756.180 32.940 ;
        RECT 1977.180 32.680 1977.440 32.940 ;
      LAYER met2 ;
        RECT 1687.610 600.170 1687.890 604.000 ;
        RECT 1687.610 600.030 1689.420 600.170 ;
        RECT 1687.610 600.000 1687.890 600.030 ;
        RECT 1689.280 591.590 1689.420 600.030 ;
        RECT 1689.220 591.270 1689.480 591.590 ;
        RECT 1755.920 591.270 1756.180 591.590 ;
        RECT 1755.980 32.970 1756.120 591.270 ;
        RECT 1755.920 32.650 1756.180 32.970 ;
        RECT 1977.180 32.650 1977.440 32.970 ;
        RECT 1977.240 2.400 1977.380 32.650 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1697.010 591.160 1697.330 591.220 ;
        RECT 1769.690 591.160 1770.010 591.220 ;
        RECT 1697.010 591.020 1770.010 591.160 ;
        RECT 1697.010 590.960 1697.330 591.020 ;
        RECT 1769.690 590.960 1770.010 591.020 ;
        RECT 1769.690 27.780 1770.010 27.840 ;
        RECT 1995.090 27.780 1995.410 27.840 ;
        RECT 1769.690 27.640 1995.410 27.780 ;
        RECT 1769.690 27.580 1770.010 27.640 ;
        RECT 1995.090 27.580 1995.410 27.640 ;
      LAYER via ;
        RECT 1697.040 590.960 1697.300 591.220 ;
        RECT 1769.720 590.960 1769.980 591.220 ;
        RECT 1769.720 27.580 1769.980 27.840 ;
        RECT 1995.120 27.580 1995.380 27.840 ;
      LAYER met2 ;
        RECT 1696.810 600.000 1697.090 604.000 ;
        RECT 1696.870 598.810 1697.010 600.000 ;
        RECT 1696.870 598.670 1697.240 598.810 ;
        RECT 1697.100 591.250 1697.240 598.670 ;
        RECT 1697.040 590.930 1697.300 591.250 ;
        RECT 1769.720 590.930 1769.980 591.250 ;
        RECT 1769.780 27.870 1769.920 590.930 ;
        RECT 1769.720 27.550 1769.980 27.870 ;
        RECT 1995.120 27.550 1995.380 27.870 ;
        RECT 1995.180 2.400 1995.320 27.550 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1707.590 586.740 1707.910 586.800 ;
        RECT 1710.810 586.740 1711.130 586.800 ;
        RECT 1707.590 586.600 1711.130 586.740 ;
        RECT 1707.590 586.540 1707.910 586.600 ;
        RECT 1710.810 586.540 1711.130 586.600 ;
        RECT 1710.810 40.020 1711.130 40.080 ;
        RECT 2012.570 40.020 2012.890 40.080 ;
        RECT 1710.810 39.880 2012.890 40.020 ;
        RECT 1710.810 39.820 1711.130 39.880 ;
        RECT 2012.570 39.820 2012.890 39.880 ;
      LAYER via ;
        RECT 1707.620 586.540 1707.880 586.800 ;
        RECT 1710.840 586.540 1711.100 586.800 ;
        RECT 1710.840 39.820 1711.100 40.080 ;
        RECT 2012.600 39.820 2012.860 40.080 ;
      LAYER met2 ;
        RECT 1706.010 600.170 1706.290 604.000 ;
        RECT 1706.010 600.030 1707.820 600.170 ;
        RECT 1706.010 600.000 1706.290 600.030 ;
        RECT 1707.680 586.830 1707.820 600.030 ;
        RECT 1707.620 586.510 1707.880 586.830 ;
        RECT 1710.840 586.510 1711.100 586.830 ;
        RECT 1710.900 40.110 1711.040 586.510 ;
        RECT 1710.840 39.790 1711.100 40.110 ;
        RECT 2012.600 39.790 2012.860 40.110 ;
        RECT 2012.660 2.400 2012.800 39.790 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1717.250 39.680 1717.570 39.740 ;
        RECT 2030.510 39.680 2030.830 39.740 ;
        RECT 1717.250 39.540 2030.830 39.680 ;
        RECT 1717.250 39.480 1717.570 39.540 ;
        RECT 2030.510 39.480 2030.830 39.540 ;
      LAYER via ;
        RECT 1717.280 39.480 1717.540 39.740 ;
        RECT 2030.540 39.480 2030.800 39.740 ;
      LAYER met2 ;
        RECT 1715.210 600.170 1715.490 604.000 ;
        RECT 1715.210 600.030 1717.480 600.170 ;
        RECT 1715.210 600.000 1715.490 600.030 ;
        RECT 1717.340 39.770 1717.480 600.030 ;
        RECT 1717.280 39.450 1717.540 39.770 ;
        RECT 2030.540 39.450 2030.800 39.770 ;
        RECT 2030.600 2.400 2030.740 39.450 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1724.150 39.340 1724.470 39.400 ;
        RECT 2048.450 39.340 2048.770 39.400 ;
        RECT 1724.150 39.200 2048.770 39.340 ;
        RECT 1724.150 39.140 1724.470 39.200 ;
        RECT 2048.450 39.140 2048.770 39.200 ;
      LAYER via ;
        RECT 1724.180 39.140 1724.440 39.400 ;
        RECT 2048.480 39.140 2048.740 39.400 ;
      LAYER met2 ;
        RECT 1724.410 600.000 1724.690 604.000 ;
        RECT 1724.470 598.810 1724.610 600.000 ;
        RECT 1724.240 598.670 1724.610 598.810 ;
        RECT 1724.240 39.430 1724.380 598.670 ;
        RECT 1724.180 39.110 1724.440 39.430 ;
        RECT 2048.480 39.110 2048.740 39.430 ;
        RECT 2048.540 2.400 2048.680 39.110 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 985.850 33.560 986.170 33.620 ;
        RECT 1063.130 33.560 1063.450 33.620 ;
        RECT 985.850 33.420 1063.450 33.560 ;
        RECT 985.850 33.360 986.170 33.420 ;
        RECT 1063.130 33.360 1063.450 33.420 ;
        RECT 763.670 19.620 763.990 19.680 ;
        RECT 985.850 19.620 986.170 19.680 ;
        RECT 763.670 19.480 986.170 19.620 ;
        RECT 763.670 19.420 763.990 19.480 ;
        RECT 985.850 19.420 986.170 19.480 ;
      LAYER via ;
        RECT 985.880 33.360 986.140 33.620 ;
        RECT 1063.160 33.360 1063.420 33.620 ;
        RECT 763.700 19.420 763.960 19.680 ;
        RECT 985.880 19.420 986.140 19.680 ;
      LAYER met2 ;
        RECT 1062.930 600.000 1063.210 604.000 ;
        RECT 1062.990 598.810 1063.130 600.000 ;
        RECT 1062.990 598.670 1063.360 598.810 ;
        RECT 1063.220 33.650 1063.360 598.670 ;
        RECT 985.880 33.330 986.140 33.650 ;
        RECT 1063.160 33.330 1063.420 33.650 ;
        RECT 985.940 19.710 986.080 33.330 ;
        RECT 763.700 19.390 763.960 19.710 ;
        RECT 985.880 19.390 986.140 19.710 ;
        RECT 763.760 2.400 763.900 19.390 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1735.190 586.740 1735.510 586.800 ;
        RECT 1738.410 586.740 1738.730 586.800 ;
        RECT 1735.190 586.600 1738.730 586.740 ;
        RECT 1735.190 586.540 1735.510 586.600 ;
        RECT 1738.410 586.540 1738.730 586.600 ;
        RECT 1738.410 39.000 1738.730 39.060 ;
        RECT 2066.390 39.000 2066.710 39.060 ;
        RECT 1738.410 38.860 2066.710 39.000 ;
        RECT 1738.410 38.800 1738.730 38.860 ;
        RECT 2066.390 38.800 2066.710 38.860 ;
      LAYER via ;
        RECT 1735.220 586.540 1735.480 586.800 ;
        RECT 1738.440 586.540 1738.700 586.800 ;
        RECT 1738.440 38.800 1738.700 39.060 ;
        RECT 2066.420 38.800 2066.680 39.060 ;
      LAYER met2 ;
        RECT 1733.610 600.170 1733.890 604.000 ;
        RECT 1733.610 600.030 1735.420 600.170 ;
        RECT 1733.610 600.000 1733.890 600.030 ;
        RECT 1735.280 586.830 1735.420 600.030 ;
        RECT 1735.220 586.510 1735.480 586.830 ;
        RECT 1738.440 586.510 1738.700 586.830 ;
        RECT 1738.500 39.090 1738.640 586.510 ;
        RECT 1738.440 38.770 1738.700 39.090 ;
        RECT 2066.420 38.770 2066.680 39.090 ;
        RECT 2066.480 2.400 2066.620 38.770 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1744.850 38.660 1745.170 38.720 ;
        RECT 2084.330 38.660 2084.650 38.720 ;
        RECT 1744.850 38.520 2084.650 38.660 ;
        RECT 1744.850 38.460 1745.170 38.520 ;
        RECT 2084.330 38.460 2084.650 38.520 ;
      LAYER via ;
        RECT 1744.880 38.460 1745.140 38.720 ;
        RECT 2084.360 38.460 2084.620 38.720 ;
      LAYER met2 ;
        RECT 1742.810 600.170 1743.090 604.000 ;
        RECT 1742.810 600.030 1745.080 600.170 ;
        RECT 1742.810 600.000 1743.090 600.030 ;
        RECT 1744.940 38.750 1745.080 600.030 ;
        RECT 1744.880 38.430 1745.140 38.750 ;
        RECT 2084.360 38.430 2084.620 38.750 ;
        RECT 2084.420 2.400 2084.560 38.430 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1751.750 38.320 1752.070 38.380 ;
        RECT 2101.810 38.320 2102.130 38.380 ;
        RECT 1751.750 38.180 2102.130 38.320 ;
        RECT 1751.750 38.120 1752.070 38.180 ;
        RECT 2101.810 38.120 2102.130 38.180 ;
      LAYER via ;
        RECT 1751.780 38.120 1752.040 38.380 ;
        RECT 2101.840 38.120 2102.100 38.380 ;
      LAYER met2 ;
        RECT 1752.010 600.000 1752.290 604.000 ;
        RECT 1752.070 598.810 1752.210 600.000 ;
        RECT 1751.840 598.670 1752.210 598.810 ;
        RECT 1751.840 38.410 1751.980 598.670 ;
        RECT 1751.780 38.090 1752.040 38.410 ;
        RECT 2101.840 38.090 2102.100 38.410 ;
        RECT 2101.900 2.400 2102.040 38.090 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1762.790 586.740 1763.110 586.800 ;
        RECT 1766.010 586.740 1766.330 586.800 ;
        RECT 1762.790 586.600 1766.330 586.740 ;
        RECT 1762.790 586.540 1763.110 586.600 ;
        RECT 1766.010 586.540 1766.330 586.600 ;
        RECT 1766.010 37.980 1766.330 38.040 ;
        RECT 2119.750 37.980 2120.070 38.040 ;
        RECT 1766.010 37.840 2120.070 37.980 ;
        RECT 1766.010 37.780 1766.330 37.840 ;
        RECT 2119.750 37.780 2120.070 37.840 ;
      LAYER via ;
        RECT 1762.820 586.540 1763.080 586.800 ;
        RECT 1766.040 586.540 1766.300 586.800 ;
        RECT 1766.040 37.780 1766.300 38.040 ;
        RECT 2119.780 37.780 2120.040 38.040 ;
      LAYER met2 ;
        RECT 1761.210 600.170 1761.490 604.000 ;
        RECT 1761.210 600.030 1763.020 600.170 ;
        RECT 1761.210 600.000 1761.490 600.030 ;
        RECT 1762.880 586.830 1763.020 600.030 ;
        RECT 1762.820 586.510 1763.080 586.830 ;
        RECT 1766.040 586.510 1766.300 586.830 ;
        RECT 1766.100 38.070 1766.240 586.510 ;
        RECT 1766.040 37.750 1766.300 38.070 ;
        RECT 2119.780 37.750 2120.040 38.070 ;
        RECT 2119.840 2.400 2119.980 37.750 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.450 45.120 1772.770 45.180 ;
        RECT 2137.690 45.120 2138.010 45.180 ;
        RECT 1772.450 44.980 2138.010 45.120 ;
        RECT 1772.450 44.920 1772.770 44.980 ;
        RECT 2137.690 44.920 2138.010 44.980 ;
      LAYER via ;
        RECT 1772.480 44.920 1772.740 45.180 ;
        RECT 2137.720 44.920 2137.980 45.180 ;
      LAYER met2 ;
        RECT 1770.410 600.170 1770.690 604.000 ;
        RECT 1770.410 600.030 1772.680 600.170 ;
        RECT 1770.410 600.000 1770.690 600.030 ;
        RECT 1772.540 45.210 1772.680 600.030 ;
        RECT 1772.480 44.890 1772.740 45.210 ;
        RECT 2137.720 44.890 2137.980 45.210 ;
        RECT 2137.780 2.400 2137.920 44.890 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.350 44.780 1779.670 44.840 ;
        RECT 2155.630 44.780 2155.950 44.840 ;
        RECT 1779.350 44.640 2155.950 44.780 ;
        RECT 1779.350 44.580 1779.670 44.640 ;
        RECT 2155.630 44.580 2155.950 44.640 ;
      LAYER via ;
        RECT 1779.380 44.580 1779.640 44.840 ;
        RECT 2155.660 44.580 2155.920 44.840 ;
      LAYER met2 ;
        RECT 1779.610 600.000 1779.890 604.000 ;
        RECT 1779.670 598.810 1779.810 600.000 ;
        RECT 1779.440 598.670 1779.810 598.810 ;
        RECT 1779.440 44.870 1779.580 598.670 ;
        RECT 1779.380 44.550 1779.640 44.870 ;
        RECT 2155.660 44.550 2155.920 44.870 ;
        RECT 2155.720 2.400 2155.860 44.550 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1790.390 586.740 1790.710 586.800 ;
        RECT 1793.150 586.740 1793.470 586.800 ;
        RECT 1790.390 586.600 1793.470 586.740 ;
        RECT 1790.390 586.540 1790.710 586.600 ;
        RECT 1793.150 586.540 1793.470 586.600 ;
        RECT 1793.150 49.880 1793.470 49.940 ;
        RECT 2173.110 49.880 2173.430 49.940 ;
        RECT 1793.150 49.740 2173.430 49.880 ;
        RECT 1793.150 49.680 1793.470 49.740 ;
        RECT 2173.110 49.680 2173.430 49.740 ;
      LAYER via ;
        RECT 1790.420 586.540 1790.680 586.800 ;
        RECT 1793.180 586.540 1793.440 586.800 ;
        RECT 1793.180 49.680 1793.440 49.940 ;
        RECT 2173.140 49.680 2173.400 49.940 ;
      LAYER met2 ;
        RECT 1788.810 600.170 1789.090 604.000 ;
        RECT 1788.810 600.030 1790.620 600.170 ;
        RECT 1788.810 600.000 1789.090 600.030 ;
        RECT 1790.480 586.830 1790.620 600.030 ;
        RECT 1790.420 586.510 1790.680 586.830 ;
        RECT 1793.180 586.510 1793.440 586.830 ;
        RECT 1793.240 49.970 1793.380 586.510 ;
        RECT 1793.180 49.650 1793.440 49.970 ;
        RECT 2173.140 49.650 2173.400 49.970 ;
        RECT 2173.200 2.400 2173.340 49.650 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.050 50.220 1800.370 50.280 ;
        RECT 2187.370 50.220 2187.690 50.280 ;
        RECT 1800.050 50.080 2187.690 50.220 ;
        RECT 1800.050 50.020 1800.370 50.080 ;
        RECT 2187.370 50.020 2187.690 50.080 ;
      LAYER via ;
        RECT 1800.080 50.020 1800.340 50.280 ;
        RECT 2187.400 50.020 2187.660 50.280 ;
      LAYER met2 ;
        RECT 1798.010 600.170 1798.290 604.000 ;
        RECT 1798.010 600.030 1800.280 600.170 ;
        RECT 1798.010 600.000 1798.290 600.030 ;
        RECT 1800.140 50.310 1800.280 600.030 ;
        RECT 1800.080 49.990 1800.340 50.310 ;
        RECT 2187.400 49.990 2187.660 50.310 ;
        RECT 2187.460 3.130 2187.600 49.990 ;
        RECT 2187.460 2.990 2190.820 3.130 ;
        RECT 2190.680 2.960 2190.820 2.990 ;
        RECT 2190.680 2.820 2191.280 2.960 ;
        RECT 2191.140 2.400 2191.280 2.820 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1806.950 50.900 1807.270 50.960 ;
        RECT 2208.070 50.900 2208.390 50.960 ;
        RECT 1806.950 50.760 2208.390 50.900 ;
        RECT 1806.950 50.700 1807.270 50.760 ;
        RECT 2208.070 50.700 2208.390 50.760 ;
        RECT 2208.070 2.960 2208.390 3.020 ;
        RECT 2208.990 2.960 2209.310 3.020 ;
        RECT 2208.070 2.820 2209.310 2.960 ;
        RECT 2208.070 2.760 2208.390 2.820 ;
        RECT 2208.990 2.760 2209.310 2.820 ;
      LAYER via ;
        RECT 1806.980 50.700 1807.240 50.960 ;
        RECT 2208.100 50.700 2208.360 50.960 ;
        RECT 2208.100 2.760 2208.360 3.020 ;
        RECT 2209.020 2.760 2209.280 3.020 ;
      LAYER met2 ;
        RECT 1807.210 600.000 1807.490 604.000 ;
        RECT 1807.270 598.810 1807.410 600.000 ;
        RECT 1807.040 598.670 1807.410 598.810 ;
        RECT 1807.040 50.990 1807.180 598.670 ;
        RECT 1806.980 50.670 1807.240 50.990 ;
        RECT 2208.100 50.670 2208.360 50.990 ;
        RECT 2208.160 3.050 2208.300 50.670 ;
        RECT 2208.100 2.730 2208.360 3.050 ;
        RECT 2209.020 2.730 2209.280 3.050 ;
        RECT 2209.080 2.400 2209.220 2.730 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1817.990 586.740 1818.310 586.800 ;
        RECT 1821.210 586.740 1821.530 586.800 ;
        RECT 1817.990 586.600 1821.530 586.740 ;
        RECT 1817.990 586.540 1818.310 586.600 ;
        RECT 1821.210 586.540 1821.530 586.600 ;
        RECT 1821.210 50.560 1821.530 50.620 ;
        RECT 2221.870 50.560 2222.190 50.620 ;
        RECT 1821.210 50.420 2222.190 50.560 ;
        RECT 1821.210 50.360 1821.530 50.420 ;
        RECT 2221.870 50.360 2222.190 50.420 ;
        RECT 2221.870 2.960 2222.190 3.020 ;
        RECT 2226.930 2.960 2227.250 3.020 ;
        RECT 2221.870 2.820 2227.250 2.960 ;
        RECT 2221.870 2.760 2222.190 2.820 ;
        RECT 2226.930 2.760 2227.250 2.820 ;
      LAYER via ;
        RECT 1818.020 586.540 1818.280 586.800 ;
        RECT 1821.240 586.540 1821.500 586.800 ;
        RECT 1821.240 50.360 1821.500 50.620 ;
        RECT 2221.900 50.360 2222.160 50.620 ;
        RECT 2221.900 2.760 2222.160 3.020 ;
        RECT 2226.960 2.760 2227.220 3.020 ;
      LAYER met2 ;
        RECT 1816.410 600.170 1816.690 604.000 ;
        RECT 1816.410 600.030 1818.220 600.170 ;
        RECT 1816.410 600.000 1816.690 600.030 ;
        RECT 1818.080 586.830 1818.220 600.030 ;
        RECT 1818.020 586.510 1818.280 586.830 ;
        RECT 1821.240 586.510 1821.500 586.830 ;
        RECT 1821.300 50.650 1821.440 586.510 ;
        RECT 1821.240 50.330 1821.500 50.650 ;
        RECT 2221.900 50.330 2222.160 50.650 ;
        RECT 2221.960 3.050 2222.100 50.330 ;
        RECT 2221.900 2.730 2222.160 3.050 ;
        RECT 2226.960 2.730 2227.220 3.050 ;
        RECT 2227.020 2.400 2227.160 2.730 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 972.970 33.220 973.290 33.280 ;
        RECT 1070.490 33.220 1070.810 33.280 ;
        RECT 972.970 33.080 1070.810 33.220 ;
        RECT 972.970 33.020 973.290 33.080 ;
        RECT 1070.490 33.020 1070.810 33.080 ;
        RECT 781.610 19.960 781.930 20.020 ;
        RECT 972.970 19.960 973.290 20.020 ;
        RECT 781.610 19.820 973.290 19.960 ;
        RECT 781.610 19.760 781.930 19.820 ;
        RECT 972.970 19.760 973.290 19.820 ;
      LAYER via ;
        RECT 973.000 33.020 973.260 33.280 ;
        RECT 1070.520 33.020 1070.780 33.280 ;
        RECT 781.640 19.760 781.900 20.020 ;
        RECT 973.000 19.760 973.260 20.020 ;
      LAYER met2 ;
        RECT 1072.130 600.170 1072.410 604.000 ;
        RECT 1070.580 600.030 1072.410 600.170 ;
        RECT 1070.580 33.310 1070.720 600.030 ;
        RECT 1072.130 600.000 1072.410 600.030 ;
        RECT 973.000 32.990 973.260 33.310 ;
        RECT 1070.520 32.990 1070.780 33.310 ;
        RECT 973.060 20.050 973.200 32.990 ;
        RECT 781.640 19.730 781.900 20.050 ;
        RECT 973.000 19.730 973.260 20.050 ;
        RECT 781.700 2.400 781.840 19.730 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1827.650 51.240 1827.970 51.300 ;
        RECT 2242.570 51.240 2242.890 51.300 ;
        RECT 1827.650 51.100 2242.890 51.240 ;
        RECT 1827.650 51.040 1827.970 51.100 ;
        RECT 2242.570 51.040 2242.890 51.100 ;
        RECT 2242.570 2.960 2242.890 3.020 ;
        RECT 2244.870 2.960 2245.190 3.020 ;
        RECT 2242.570 2.820 2245.190 2.960 ;
        RECT 2242.570 2.760 2242.890 2.820 ;
        RECT 2244.870 2.760 2245.190 2.820 ;
      LAYER via ;
        RECT 1827.680 51.040 1827.940 51.300 ;
        RECT 2242.600 51.040 2242.860 51.300 ;
        RECT 2242.600 2.760 2242.860 3.020 ;
        RECT 2244.900 2.760 2245.160 3.020 ;
      LAYER met2 ;
        RECT 1825.150 600.170 1825.430 604.000 ;
        RECT 1825.150 600.030 1827.880 600.170 ;
        RECT 1825.150 600.000 1825.430 600.030 ;
        RECT 1827.740 51.330 1827.880 600.030 ;
        RECT 1827.680 51.010 1827.940 51.330 ;
        RECT 2242.600 51.010 2242.860 51.330 ;
        RECT 2242.660 3.050 2242.800 51.010 ;
        RECT 2242.600 2.730 2242.860 3.050 ;
        RECT 2244.900 2.730 2245.160 3.050 ;
        RECT 2244.960 2.400 2245.100 2.730 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1834.550 54.980 1834.870 55.040 ;
        RECT 2256.370 54.980 2256.690 55.040 ;
        RECT 1834.550 54.840 2256.690 54.980 ;
        RECT 1834.550 54.780 1834.870 54.840 ;
        RECT 2256.370 54.780 2256.690 54.840 ;
        RECT 2256.370 15.880 2256.690 15.940 ;
        RECT 2262.350 15.880 2262.670 15.940 ;
        RECT 2256.370 15.740 2262.670 15.880 ;
        RECT 2256.370 15.680 2256.690 15.740 ;
        RECT 2262.350 15.680 2262.670 15.740 ;
      LAYER via ;
        RECT 1834.580 54.780 1834.840 55.040 ;
        RECT 2256.400 54.780 2256.660 55.040 ;
        RECT 2256.400 15.680 2256.660 15.940 ;
        RECT 2262.380 15.680 2262.640 15.940 ;
      LAYER met2 ;
        RECT 1834.350 600.000 1834.630 604.000 ;
        RECT 1834.410 598.810 1834.550 600.000 ;
        RECT 1834.410 598.670 1834.780 598.810 ;
        RECT 1834.640 55.070 1834.780 598.670 ;
        RECT 1834.580 54.750 1834.840 55.070 ;
        RECT 2256.400 54.750 2256.660 55.070 ;
        RECT 2256.460 15.970 2256.600 54.750 ;
        RECT 2256.400 15.650 2256.660 15.970 ;
        RECT 2262.380 15.650 2262.640 15.970 ;
        RECT 2262.440 2.400 2262.580 15.650 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1845.130 586.740 1845.450 586.800 ;
        RECT 1848.810 586.740 1849.130 586.800 ;
        RECT 1845.130 586.600 1849.130 586.740 ;
        RECT 1845.130 586.540 1845.450 586.600 ;
        RECT 1848.810 586.540 1849.130 586.600 ;
        RECT 1848.810 54.640 1849.130 54.700 ;
        RECT 2277.070 54.640 2277.390 54.700 ;
        RECT 1848.810 54.500 2277.390 54.640 ;
        RECT 1848.810 54.440 1849.130 54.500 ;
        RECT 2277.070 54.440 2277.390 54.500 ;
        RECT 2277.070 2.960 2277.390 3.020 ;
        RECT 2280.290 2.960 2280.610 3.020 ;
        RECT 2277.070 2.820 2280.610 2.960 ;
        RECT 2277.070 2.760 2277.390 2.820 ;
        RECT 2280.290 2.760 2280.610 2.820 ;
      LAYER via ;
        RECT 1845.160 586.540 1845.420 586.800 ;
        RECT 1848.840 586.540 1849.100 586.800 ;
        RECT 1848.840 54.440 1849.100 54.700 ;
        RECT 2277.100 54.440 2277.360 54.700 ;
        RECT 2277.100 2.760 2277.360 3.020 ;
        RECT 2280.320 2.760 2280.580 3.020 ;
      LAYER met2 ;
        RECT 1843.550 600.170 1843.830 604.000 ;
        RECT 1843.550 600.030 1845.360 600.170 ;
        RECT 1843.550 600.000 1843.830 600.030 ;
        RECT 1845.220 586.830 1845.360 600.030 ;
        RECT 1845.160 586.510 1845.420 586.830 ;
        RECT 1848.840 586.510 1849.100 586.830 ;
        RECT 1848.900 54.730 1849.040 586.510 ;
        RECT 1848.840 54.410 1849.100 54.730 ;
        RECT 2277.100 54.410 2277.360 54.730 ;
        RECT 2277.160 3.050 2277.300 54.410 ;
        RECT 2277.100 2.730 2277.360 3.050 ;
        RECT 2280.320 2.730 2280.580 3.050 ;
        RECT 2280.380 2.400 2280.520 2.730 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.250 54.300 1855.570 54.360 ;
        RECT 2298.230 54.300 2298.550 54.360 ;
        RECT 1855.250 54.160 2298.550 54.300 ;
        RECT 1855.250 54.100 1855.570 54.160 ;
        RECT 2298.230 54.100 2298.550 54.160 ;
      LAYER via ;
        RECT 1855.280 54.100 1855.540 54.360 ;
        RECT 2298.260 54.100 2298.520 54.360 ;
      LAYER met2 ;
        RECT 1852.750 600.170 1853.030 604.000 ;
        RECT 1852.750 600.030 1855.480 600.170 ;
        RECT 1852.750 600.000 1853.030 600.030 ;
        RECT 1855.340 54.390 1855.480 600.030 ;
        RECT 1855.280 54.070 1855.540 54.390 ;
        RECT 2298.260 54.070 2298.520 54.390 ;
        RECT 2298.320 2.400 2298.460 54.070 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1862.150 53.960 1862.470 54.020 ;
        RECT 2311.570 53.960 2311.890 54.020 ;
        RECT 1862.150 53.820 2311.890 53.960 ;
        RECT 1862.150 53.760 1862.470 53.820 ;
        RECT 2311.570 53.760 2311.890 53.820 ;
      LAYER via ;
        RECT 1862.180 53.760 1862.440 54.020 ;
        RECT 2311.600 53.760 2311.860 54.020 ;
      LAYER met2 ;
        RECT 1861.950 600.000 1862.230 604.000 ;
        RECT 1862.010 598.810 1862.150 600.000 ;
        RECT 1862.010 598.670 1862.380 598.810 ;
        RECT 1862.240 54.050 1862.380 598.670 ;
        RECT 1862.180 53.730 1862.440 54.050 ;
        RECT 2311.600 53.730 2311.860 54.050 ;
        RECT 2311.660 17.410 2311.800 53.730 ;
        RECT 2311.660 17.270 2316.400 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1872.730 586.740 1873.050 586.800 ;
        RECT 1875.950 586.740 1876.270 586.800 ;
        RECT 1872.730 586.600 1876.270 586.740 ;
        RECT 1872.730 586.540 1873.050 586.600 ;
        RECT 1875.950 586.540 1876.270 586.600 ;
        RECT 1875.950 53.620 1876.270 53.680 ;
        RECT 2332.270 53.620 2332.590 53.680 ;
        RECT 1875.950 53.480 2332.590 53.620 ;
        RECT 1875.950 53.420 1876.270 53.480 ;
        RECT 2332.270 53.420 2332.590 53.480 ;
      LAYER via ;
        RECT 1872.760 586.540 1873.020 586.800 ;
        RECT 1875.980 586.540 1876.240 586.800 ;
        RECT 1875.980 53.420 1876.240 53.680 ;
        RECT 2332.300 53.420 2332.560 53.680 ;
      LAYER met2 ;
        RECT 1871.150 600.170 1871.430 604.000 ;
        RECT 1871.150 600.030 1872.960 600.170 ;
        RECT 1871.150 600.000 1871.430 600.030 ;
        RECT 1872.820 586.830 1872.960 600.030 ;
        RECT 1872.760 586.510 1873.020 586.830 ;
        RECT 1875.980 586.510 1876.240 586.830 ;
        RECT 1876.040 53.710 1876.180 586.510 ;
        RECT 1875.980 53.390 1876.240 53.710 ;
        RECT 2332.300 53.390 2332.560 53.710 ;
        RECT 2332.360 17.410 2332.500 53.390 ;
        RECT 2332.360 17.270 2334.340 17.410 ;
        RECT 2334.200 2.400 2334.340 17.270 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1882.850 53.280 1883.170 53.340 ;
        RECT 2346.070 53.280 2346.390 53.340 ;
        RECT 1882.850 53.140 2346.390 53.280 ;
        RECT 1882.850 53.080 1883.170 53.140 ;
        RECT 2346.070 53.080 2346.390 53.140 ;
      LAYER via ;
        RECT 1882.880 53.080 1883.140 53.340 ;
        RECT 2346.100 53.080 2346.360 53.340 ;
      LAYER met2 ;
        RECT 1880.350 600.170 1880.630 604.000 ;
        RECT 1880.350 600.030 1883.080 600.170 ;
        RECT 1880.350 600.000 1880.630 600.030 ;
        RECT 1882.940 53.370 1883.080 600.030 ;
        RECT 1882.880 53.050 1883.140 53.370 ;
        RECT 2346.100 53.050 2346.360 53.370 ;
        RECT 2346.160 17.410 2346.300 53.050 ;
        RECT 2346.160 17.270 2351.820 17.410 ;
        RECT 2351.680 2.400 2351.820 17.270 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1889.750 52.940 1890.070 53.000 ;
        RECT 2366.770 52.940 2367.090 53.000 ;
        RECT 1889.750 52.800 2367.090 52.940 ;
        RECT 1889.750 52.740 1890.070 52.800 ;
        RECT 2366.770 52.740 2367.090 52.800 ;
      LAYER via ;
        RECT 1889.780 52.740 1890.040 53.000 ;
        RECT 2366.800 52.740 2367.060 53.000 ;
      LAYER met2 ;
        RECT 1889.550 600.000 1889.830 604.000 ;
        RECT 1889.610 598.810 1889.750 600.000 ;
        RECT 1889.610 598.670 1889.980 598.810 ;
        RECT 1889.840 53.030 1889.980 598.670 ;
        RECT 1889.780 52.710 1890.040 53.030 ;
        RECT 2366.800 52.710 2367.060 53.030 ;
        RECT 2366.860 16.730 2367.000 52.710 ;
        RECT 2366.860 16.590 2369.760 16.730 ;
        RECT 2369.620 2.400 2369.760 16.590 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1900.330 586.740 1900.650 586.800 ;
        RECT 1904.010 586.740 1904.330 586.800 ;
        RECT 1900.330 586.600 1904.330 586.740 ;
        RECT 1900.330 586.540 1900.650 586.600 ;
        RECT 1904.010 586.540 1904.330 586.600 ;
        RECT 1904.010 52.600 1904.330 52.660 ;
        RECT 2387.930 52.600 2388.250 52.660 ;
        RECT 1904.010 52.460 2388.250 52.600 ;
        RECT 1904.010 52.400 1904.330 52.460 ;
        RECT 2387.930 52.400 2388.250 52.460 ;
      LAYER via ;
        RECT 1900.360 586.540 1900.620 586.800 ;
        RECT 1904.040 586.540 1904.300 586.800 ;
        RECT 1904.040 52.400 1904.300 52.660 ;
        RECT 2387.960 52.400 2388.220 52.660 ;
      LAYER met2 ;
        RECT 1898.750 600.170 1899.030 604.000 ;
        RECT 1898.750 600.030 1900.560 600.170 ;
        RECT 1898.750 600.000 1899.030 600.030 ;
        RECT 1900.420 586.830 1900.560 600.030 ;
        RECT 1900.360 586.510 1900.620 586.830 ;
        RECT 1904.040 586.510 1904.300 586.830 ;
        RECT 1904.100 52.690 1904.240 586.510 ;
        RECT 1904.040 52.370 1904.300 52.690 ;
        RECT 2387.960 52.370 2388.220 52.690 ;
        RECT 2388.020 17.410 2388.160 52.370 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1910.450 52.260 1910.770 52.320 ;
        RECT 2401.270 52.260 2401.590 52.320 ;
        RECT 1910.450 52.120 2401.590 52.260 ;
        RECT 1910.450 52.060 1910.770 52.120 ;
        RECT 2401.270 52.060 2401.590 52.120 ;
      LAYER via ;
        RECT 1910.480 52.060 1910.740 52.320 ;
        RECT 2401.300 52.060 2401.560 52.320 ;
      LAYER met2 ;
        RECT 1907.950 600.170 1908.230 604.000 ;
        RECT 1907.950 600.030 1910.680 600.170 ;
        RECT 1907.950 600.000 1908.230 600.030 ;
        RECT 1910.540 52.350 1910.680 600.030 ;
        RECT 1910.480 52.030 1910.740 52.350 ;
        RECT 2401.300 52.030 2401.560 52.350 ;
        RECT 2401.360 18.090 2401.500 52.030 ;
        RECT 2401.360 17.950 2405.640 18.090 ;
        RECT 2405.500 2.400 2405.640 17.950 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1077.850 476.240 1078.170 476.300 ;
        RECT 1079.690 476.240 1080.010 476.300 ;
        RECT 1077.850 476.100 1080.010 476.240 ;
        RECT 1077.850 476.040 1078.170 476.100 ;
        RECT 1079.690 476.040 1080.010 476.100 ;
        RECT 1077.390 434.760 1077.710 434.820 ;
        RECT 1077.850 434.760 1078.170 434.820 ;
        RECT 1077.390 434.620 1078.170 434.760 ;
        RECT 1077.390 434.560 1077.710 434.620 ;
        RECT 1077.850 434.560 1078.170 434.620 ;
        RECT 966.530 32.880 966.850 32.940 ;
        RECT 1077.390 32.880 1077.710 32.940 ;
        RECT 966.530 32.740 1077.710 32.880 ;
        RECT 966.530 32.680 966.850 32.740 ;
        RECT 1077.390 32.680 1077.710 32.740 ;
        RECT 799.550 14.860 799.870 14.920 ;
        RECT 966.530 14.860 966.850 14.920 ;
        RECT 799.550 14.720 966.850 14.860 ;
        RECT 799.550 14.660 799.870 14.720 ;
        RECT 966.530 14.660 966.850 14.720 ;
      LAYER via ;
        RECT 1077.880 476.040 1078.140 476.300 ;
        RECT 1079.720 476.040 1079.980 476.300 ;
        RECT 1077.420 434.560 1077.680 434.820 ;
        RECT 1077.880 434.560 1078.140 434.820 ;
        RECT 966.560 32.680 966.820 32.940 ;
        RECT 1077.420 32.680 1077.680 32.940 ;
        RECT 799.580 14.660 799.840 14.920 ;
        RECT 966.560 14.660 966.820 14.920 ;
      LAYER met2 ;
        RECT 1081.330 600.170 1081.610 604.000 ;
        RECT 1080.700 600.030 1081.610 600.170 ;
        RECT 1080.700 579.885 1080.840 600.030 ;
        RECT 1081.330 600.000 1081.610 600.030 ;
        RECT 1079.710 579.515 1079.990 579.885 ;
        RECT 1080.630 579.515 1080.910 579.885 ;
        RECT 1079.780 476.330 1079.920 579.515 ;
        RECT 1077.880 476.010 1078.140 476.330 ;
        RECT 1079.720 476.010 1079.980 476.330 ;
        RECT 1077.940 434.850 1078.080 476.010 ;
        RECT 1077.420 434.530 1077.680 434.850 ;
        RECT 1077.880 434.530 1078.140 434.850 ;
        RECT 1077.480 32.970 1077.620 434.530 ;
        RECT 966.560 32.650 966.820 32.970 ;
        RECT 1077.420 32.650 1077.680 32.970 ;
        RECT 966.620 14.950 966.760 32.650 ;
        RECT 799.580 14.630 799.840 14.950 ;
        RECT 966.560 14.630 966.820 14.950 ;
        RECT 799.640 2.400 799.780 14.630 ;
        RECT 799.430 -4.800 799.990 2.400 ;
      LAYER via2 ;
        RECT 1079.710 579.560 1079.990 579.840 ;
        RECT 1080.630 579.560 1080.910 579.840 ;
      LAYER met3 ;
        RECT 1079.685 579.850 1080.015 579.865 ;
        RECT 1080.605 579.850 1080.935 579.865 ;
        RECT 1079.685 579.550 1080.935 579.850 ;
        RECT 1079.685 579.535 1080.015 579.550 ;
        RECT 1080.605 579.535 1080.935 579.550 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 44.100 645.310 44.160 ;
        RECT 1001.030 44.100 1001.350 44.160 ;
        RECT 644.990 43.960 1001.350 44.100 ;
        RECT 644.990 43.900 645.310 43.960 ;
        RECT 1001.030 43.900 1001.350 43.960 ;
      LAYER via ;
        RECT 645.020 43.900 645.280 44.160 ;
        RECT 1001.060 43.900 1001.320 44.160 ;
      LAYER met2 ;
        RECT 1001.750 600.170 1002.030 604.000 ;
        RECT 1001.120 600.030 1002.030 600.170 ;
        RECT 1001.120 44.190 1001.260 600.030 ;
        RECT 1001.750 600.000 1002.030 600.030 ;
        RECT 645.020 43.870 645.280 44.190 ;
        RECT 1001.060 43.870 1001.320 44.190 ;
        RECT 645.080 2.400 645.220 43.870 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1921.950 586.740 1922.270 586.800 ;
        RECT 1924.250 586.740 1924.570 586.800 ;
        RECT 1921.950 586.600 1924.570 586.740 ;
        RECT 1921.950 586.540 1922.270 586.600 ;
        RECT 1924.250 586.540 1924.570 586.600 ;
        RECT 1924.250 51.920 1924.570 51.980 ;
        RECT 2428.870 51.920 2429.190 51.980 ;
        RECT 1924.250 51.780 2429.190 51.920 ;
        RECT 1924.250 51.720 1924.570 51.780 ;
        RECT 2428.870 51.720 2429.190 51.780 ;
      LAYER via ;
        RECT 1921.980 586.540 1922.240 586.800 ;
        RECT 1924.280 586.540 1924.540 586.800 ;
        RECT 1924.280 51.720 1924.540 51.980 ;
        RECT 2428.900 51.720 2429.160 51.980 ;
      LAYER met2 ;
        RECT 1920.370 600.170 1920.650 604.000 ;
        RECT 1920.370 600.030 1922.180 600.170 ;
        RECT 1920.370 600.000 1920.650 600.030 ;
        RECT 1922.040 586.830 1922.180 600.030 ;
        RECT 1921.980 586.510 1922.240 586.830 ;
        RECT 1924.280 586.510 1924.540 586.830 ;
        RECT 1924.340 52.010 1924.480 586.510 ;
        RECT 1924.280 51.690 1924.540 52.010 ;
        RECT 2428.900 51.690 2429.160 52.010 ;
        RECT 2428.960 2.400 2429.100 51.690 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1931.150 61.100 1931.470 61.160 ;
        RECT 2442.670 61.100 2442.990 61.160 ;
        RECT 1931.150 60.960 2442.990 61.100 ;
        RECT 1931.150 60.900 1931.470 60.960 ;
        RECT 2442.670 60.900 2442.990 60.960 ;
      LAYER via ;
        RECT 1931.180 60.900 1931.440 61.160 ;
        RECT 2442.700 60.900 2442.960 61.160 ;
      LAYER met2 ;
        RECT 1929.570 600.170 1929.850 604.000 ;
        RECT 1929.570 600.030 1931.380 600.170 ;
        RECT 1929.570 600.000 1929.850 600.030 ;
        RECT 1931.240 61.190 1931.380 600.030 ;
        RECT 1931.180 60.870 1931.440 61.190 ;
        RECT 2442.700 60.870 2442.960 61.190 ;
        RECT 2442.760 18.090 2442.900 60.870 ;
        RECT 2442.760 17.950 2447.040 18.090 ;
        RECT 2446.900 2.400 2447.040 17.950 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1940.350 586.740 1940.670 586.800 ;
        RECT 1944.490 586.740 1944.810 586.800 ;
        RECT 1940.350 586.600 1944.810 586.740 ;
        RECT 1940.350 586.540 1940.670 586.600 ;
        RECT 1944.490 586.540 1944.810 586.600 ;
        RECT 1944.490 60.760 1944.810 60.820 ;
        RECT 2463.370 60.760 2463.690 60.820 ;
        RECT 1944.490 60.620 2463.690 60.760 ;
        RECT 1944.490 60.560 1944.810 60.620 ;
        RECT 2463.370 60.560 2463.690 60.620 ;
      LAYER via ;
        RECT 1940.380 586.540 1940.640 586.800 ;
        RECT 1944.520 586.540 1944.780 586.800 ;
        RECT 1944.520 60.560 1944.780 60.820 ;
        RECT 2463.400 60.560 2463.660 60.820 ;
      LAYER met2 ;
        RECT 1938.770 600.170 1939.050 604.000 ;
        RECT 1938.770 600.030 1940.580 600.170 ;
        RECT 1938.770 600.000 1939.050 600.030 ;
        RECT 1940.440 586.830 1940.580 600.030 ;
        RECT 1940.380 586.510 1940.640 586.830 ;
        RECT 1944.520 586.510 1944.780 586.830 ;
        RECT 1944.580 60.850 1944.720 586.510 ;
        RECT 1944.520 60.530 1944.780 60.850 ;
        RECT 2463.400 60.530 2463.660 60.850 ;
        RECT 2463.460 17.410 2463.600 60.530 ;
        RECT 2463.460 17.270 2464.980 17.410 ;
        RECT 2464.840 2.400 2464.980 17.270 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1949.550 586.740 1949.870 586.800 ;
        RECT 1951.850 586.740 1952.170 586.800 ;
        RECT 1949.550 586.600 1952.170 586.740 ;
        RECT 1949.550 586.540 1949.870 586.600 ;
        RECT 1951.850 586.540 1952.170 586.600 ;
        RECT 1951.850 60.420 1952.170 60.480 ;
        RECT 2477.170 60.420 2477.490 60.480 ;
        RECT 1951.850 60.280 2477.490 60.420 ;
        RECT 1951.850 60.220 1952.170 60.280 ;
        RECT 2477.170 60.220 2477.490 60.280 ;
      LAYER via ;
        RECT 1949.580 586.540 1949.840 586.800 ;
        RECT 1951.880 586.540 1952.140 586.800 ;
        RECT 1951.880 60.220 1952.140 60.480 ;
        RECT 2477.200 60.220 2477.460 60.480 ;
      LAYER met2 ;
        RECT 1947.970 600.170 1948.250 604.000 ;
        RECT 1947.970 600.030 1949.780 600.170 ;
        RECT 1947.970 600.000 1948.250 600.030 ;
        RECT 1949.640 586.830 1949.780 600.030 ;
        RECT 1949.580 586.510 1949.840 586.830 ;
        RECT 1951.880 586.510 1952.140 586.830 ;
        RECT 1951.940 60.510 1952.080 586.510 ;
        RECT 1951.880 60.190 1952.140 60.510 ;
        RECT 2477.200 60.190 2477.460 60.510 ;
        RECT 2477.260 18.090 2477.400 60.190 ;
        RECT 2477.260 17.950 2482.920 18.090 ;
        RECT 2482.780 2.400 2482.920 17.950 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1958.750 60.080 1959.070 60.140 ;
        RECT 2497.870 60.080 2498.190 60.140 ;
        RECT 1958.750 59.940 2498.190 60.080 ;
        RECT 1958.750 59.880 1959.070 59.940 ;
        RECT 2497.870 59.880 2498.190 59.940 ;
        RECT 2497.870 2.960 2498.190 3.020 ;
        RECT 2500.630 2.960 2500.950 3.020 ;
        RECT 2497.870 2.820 2500.950 2.960 ;
        RECT 2497.870 2.760 2498.190 2.820 ;
        RECT 2500.630 2.760 2500.950 2.820 ;
      LAYER via ;
        RECT 1958.780 59.880 1959.040 60.140 ;
        RECT 2497.900 59.880 2498.160 60.140 ;
        RECT 2497.900 2.760 2498.160 3.020 ;
        RECT 2500.660 2.760 2500.920 3.020 ;
      LAYER met2 ;
        RECT 1957.170 600.170 1957.450 604.000 ;
        RECT 1957.170 600.030 1958.980 600.170 ;
        RECT 1957.170 600.000 1957.450 600.030 ;
        RECT 1958.840 60.170 1958.980 600.030 ;
        RECT 1958.780 59.850 1959.040 60.170 ;
        RECT 2497.900 59.850 2498.160 60.170 ;
        RECT 2497.960 3.050 2498.100 59.850 ;
        RECT 2497.900 2.730 2498.160 3.050 ;
        RECT 2500.660 2.730 2500.920 3.050 ;
        RECT 2500.720 2.400 2500.860 2.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1967.950 586.740 1968.270 586.800 ;
        RECT 1972.090 586.740 1972.410 586.800 ;
        RECT 1967.950 586.600 1972.410 586.740 ;
        RECT 1967.950 586.540 1968.270 586.600 ;
        RECT 1972.090 586.540 1972.410 586.600 ;
        RECT 1972.090 59.740 1972.410 59.800 ;
        RECT 2511.670 59.740 2511.990 59.800 ;
        RECT 1972.090 59.600 2511.990 59.740 ;
        RECT 1972.090 59.540 1972.410 59.600 ;
        RECT 2511.670 59.540 2511.990 59.600 ;
        RECT 2511.670 14.180 2511.990 14.240 ;
        RECT 2518.110 14.180 2518.430 14.240 ;
        RECT 2511.670 14.040 2518.430 14.180 ;
        RECT 2511.670 13.980 2511.990 14.040 ;
        RECT 2518.110 13.980 2518.430 14.040 ;
      LAYER via ;
        RECT 1967.980 586.540 1968.240 586.800 ;
        RECT 1972.120 586.540 1972.380 586.800 ;
        RECT 1972.120 59.540 1972.380 59.800 ;
        RECT 2511.700 59.540 2511.960 59.800 ;
        RECT 2511.700 13.980 2511.960 14.240 ;
        RECT 2518.140 13.980 2518.400 14.240 ;
      LAYER met2 ;
        RECT 1966.370 600.170 1966.650 604.000 ;
        RECT 1966.370 600.030 1968.180 600.170 ;
        RECT 1966.370 600.000 1966.650 600.030 ;
        RECT 1968.040 586.830 1968.180 600.030 ;
        RECT 1967.980 586.510 1968.240 586.830 ;
        RECT 1972.120 586.510 1972.380 586.830 ;
        RECT 1972.180 59.830 1972.320 586.510 ;
        RECT 1972.120 59.510 1972.380 59.830 ;
        RECT 2511.700 59.510 2511.960 59.830 ;
        RECT 2511.760 14.270 2511.900 59.510 ;
        RECT 2511.700 13.950 2511.960 14.270 ;
        RECT 2518.140 13.950 2518.400 14.270 ;
        RECT 2518.200 2.400 2518.340 13.950 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1977.150 586.740 1977.470 586.800 ;
        RECT 1979.450 586.740 1979.770 586.800 ;
        RECT 1977.150 586.600 1979.770 586.740 ;
        RECT 1977.150 586.540 1977.470 586.600 ;
        RECT 1979.450 586.540 1979.770 586.600 ;
        RECT 1979.450 59.400 1979.770 59.460 ;
        RECT 2532.370 59.400 2532.690 59.460 ;
        RECT 1979.450 59.260 2532.690 59.400 ;
        RECT 1979.450 59.200 1979.770 59.260 ;
        RECT 2532.370 59.200 2532.690 59.260 ;
        RECT 2532.370 2.960 2532.690 3.020 ;
        RECT 2536.050 2.960 2536.370 3.020 ;
        RECT 2532.370 2.820 2536.370 2.960 ;
        RECT 2532.370 2.760 2532.690 2.820 ;
        RECT 2536.050 2.760 2536.370 2.820 ;
      LAYER via ;
        RECT 1977.180 586.540 1977.440 586.800 ;
        RECT 1979.480 586.540 1979.740 586.800 ;
        RECT 1979.480 59.200 1979.740 59.460 ;
        RECT 2532.400 59.200 2532.660 59.460 ;
        RECT 2532.400 2.760 2532.660 3.020 ;
        RECT 2536.080 2.760 2536.340 3.020 ;
      LAYER met2 ;
        RECT 1975.570 600.170 1975.850 604.000 ;
        RECT 1975.570 600.030 1977.380 600.170 ;
        RECT 1975.570 600.000 1975.850 600.030 ;
        RECT 1977.240 586.830 1977.380 600.030 ;
        RECT 1977.180 586.510 1977.440 586.830 ;
        RECT 1979.480 586.510 1979.740 586.830 ;
        RECT 1979.540 59.490 1979.680 586.510 ;
        RECT 1979.480 59.170 1979.740 59.490 ;
        RECT 2532.400 59.170 2532.660 59.490 ;
        RECT 2532.460 3.050 2532.600 59.170 ;
        RECT 2532.400 2.730 2532.660 3.050 ;
        RECT 2536.080 2.730 2536.340 3.050 ;
        RECT 2536.140 2.400 2536.280 2.730 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1986.350 59.060 1986.670 59.120 ;
        RECT 2553.070 59.060 2553.390 59.120 ;
        RECT 1986.350 58.920 2553.390 59.060 ;
        RECT 1986.350 58.860 1986.670 58.920 ;
        RECT 2553.070 58.860 2553.390 58.920 ;
        RECT 2553.070 2.960 2553.390 3.020 ;
        RECT 2553.990 2.960 2554.310 3.020 ;
        RECT 2553.070 2.820 2554.310 2.960 ;
        RECT 2553.070 2.760 2553.390 2.820 ;
        RECT 2553.990 2.760 2554.310 2.820 ;
      LAYER via ;
        RECT 1986.380 58.860 1986.640 59.120 ;
        RECT 2553.100 58.860 2553.360 59.120 ;
        RECT 2553.100 2.760 2553.360 3.020 ;
        RECT 2554.020 2.760 2554.280 3.020 ;
      LAYER met2 ;
        RECT 1984.770 600.170 1985.050 604.000 ;
        RECT 1984.770 600.030 1986.580 600.170 ;
        RECT 1984.770 600.000 1985.050 600.030 ;
        RECT 1986.440 59.150 1986.580 600.030 ;
        RECT 1986.380 58.830 1986.640 59.150 ;
        RECT 2553.100 58.830 2553.360 59.150 ;
        RECT 2553.160 3.050 2553.300 58.830 ;
        RECT 2553.100 2.730 2553.360 3.050 ;
        RECT 2554.020 2.730 2554.280 3.050 ;
        RECT 2554.080 2.400 2554.220 2.730 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1995.550 586.740 1995.870 586.800 ;
        RECT 1999.690 586.740 2000.010 586.800 ;
        RECT 1995.550 586.600 2000.010 586.740 ;
        RECT 1995.550 586.540 1995.870 586.600 ;
        RECT 1999.690 586.540 2000.010 586.600 ;
        RECT 1999.690 58.720 2000.010 58.780 ;
        RECT 2566.870 58.720 2567.190 58.780 ;
        RECT 1999.690 58.580 2567.190 58.720 ;
        RECT 1999.690 58.520 2000.010 58.580 ;
        RECT 2566.870 58.520 2567.190 58.580 ;
        RECT 2566.870 2.960 2567.190 3.020 ;
        RECT 2571.930 2.960 2572.250 3.020 ;
        RECT 2566.870 2.820 2572.250 2.960 ;
        RECT 2566.870 2.760 2567.190 2.820 ;
        RECT 2571.930 2.760 2572.250 2.820 ;
      LAYER via ;
        RECT 1995.580 586.540 1995.840 586.800 ;
        RECT 1999.720 586.540 1999.980 586.800 ;
        RECT 1999.720 58.520 1999.980 58.780 ;
        RECT 2566.900 58.520 2567.160 58.780 ;
        RECT 2566.900 2.760 2567.160 3.020 ;
        RECT 2571.960 2.760 2572.220 3.020 ;
      LAYER met2 ;
        RECT 1993.970 600.170 1994.250 604.000 ;
        RECT 1993.970 600.030 1995.780 600.170 ;
        RECT 1993.970 600.000 1994.250 600.030 ;
        RECT 1995.640 586.830 1995.780 600.030 ;
        RECT 1995.580 586.510 1995.840 586.830 ;
        RECT 1999.720 586.510 1999.980 586.830 ;
        RECT 1999.780 58.810 1999.920 586.510 ;
        RECT 1999.720 58.490 1999.980 58.810 ;
        RECT 2566.900 58.490 2567.160 58.810 ;
        RECT 2566.960 3.050 2567.100 58.490 ;
        RECT 2566.900 2.730 2567.160 3.050 ;
        RECT 2571.960 2.730 2572.220 3.050 ;
        RECT 2572.020 2.400 2572.160 2.730 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2004.290 591.840 2004.610 591.900 ;
        RECT 2369.990 591.840 2370.310 591.900 ;
        RECT 2004.290 591.700 2370.310 591.840 ;
        RECT 2004.290 591.640 2004.610 591.700 ;
        RECT 2369.990 591.640 2370.310 591.700 ;
        RECT 2369.990 14.520 2370.310 14.580 ;
        RECT 2589.410 14.520 2589.730 14.580 ;
        RECT 2369.990 14.380 2589.730 14.520 ;
        RECT 2369.990 14.320 2370.310 14.380 ;
        RECT 2589.410 14.320 2589.730 14.380 ;
      LAYER via ;
        RECT 2004.320 591.640 2004.580 591.900 ;
        RECT 2370.020 591.640 2370.280 591.900 ;
        RECT 2370.020 14.320 2370.280 14.580 ;
        RECT 2589.440 14.320 2589.700 14.580 ;
      LAYER met2 ;
        RECT 2002.710 600.170 2002.990 604.000 ;
        RECT 2002.710 600.030 2004.520 600.170 ;
        RECT 2002.710 600.000 2002.990 600.030 ;
        RECT 2004.380 591.930 2004.520 600.030 ;
        RECT 2004.320 591.610 2004.580 591.930 ;
        RECT 2370.020 591.610 2370.280 591.930 ;
        RECT 2370.080 14.610 2370.220 591.610 ;
        RECT 2370.020 14.290 2370.280 14.610 ;
        RECT 2589.440 14.290 2589.700 14.610 ;
        RECT 2589.500 2.400 2589.640 14.290 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1091.190 524.520 1091.510 524.580 ;
        RECT 1091.650 524.520 1091.970 524.580 ;
        RECT 1091.190 524.380 1091.970 524.520 ;
        RECT 1091.190 524.320 1091.510 524.380 ;
        RECT 1091.650 524.320 1091.970 524.380 ;
        RECT 1091.650 476.240 1091.970 476.300 ;
        RECT 1092.110 476.240 1092.430 476.300 ;
        RECT 1091.650 476.100 1092.430 476.240 ;
        RECT 1091.650 476.040 1091.970 476.100 ;
        RECT 1092.110 476.040 1092.430 476.100 ;
        RECT 1091.190 434.760 1091.510 434.820 ;
        RECT 1091.650 434.760 1091.970 434.820 ;
        RECT 1091.190 434.620 1091.970 434.760 ;
        RECT 1091.190 434.560 1091.510 434.620 ;
        RECT 1091.650 434.560 1091.970 434.620 ;
        RECT 1091.190 427.620 1091.510 427.680 ;
        RECT 1092.110 427.620 1092.430 427.680 ;
        RECT 1091.190 427.480 1092.430 427.620 ;
        RECT 1091.190 427.420 1091.510 427.480 ;
        RECT 1092.110 427.420 1092.430 427.480 ;
        RECT 1091.190 379.680 1091.510 379.740 ;
        RECT 1092.110 379.680 1092.430 379.740 ;
        RECT 1091.190 379.540 1092.430 379.680 ;
        RECT 1091.190 379.480 1091.510 379.540 ;
        RECT 1092.110 379.480 1092.430 379.540 ;
        RECT 1090.730 282.780 1091.050 282.840 ;
        RECT 1091.190 282.780 1091.510 282.840 ;
        RECT 1090.730 282.640 1091.510 282.780 ;
        RECT 1090.730 282.580 1091.050 282.640 ;
        RECT 1091.190 282.580 1091.510 282.640 ;
        RECT 1090.730 234.840 1091.050 234.900 ;
        RECT 1092.110 234.840 1092.430 234.900 ;
        RECT 1090.730 234.700 1092.430 234.840 ;
        RECT 1090.730 234.640 1091.050 234.700 ;
        RECT 1092.110 234.640 1092.430 234.700 ;
        RECT 1091.190 145.080 1091.510 145.140 ;
        RECT 1092.110 145.080 1092.430 145.140 ;
        RECT 1091.190 144.940 1092.430 145.080 ;
        RECT 1091.190 144.880 1091.510 144.940 ;
        RECT 1092.110 144.880 1092.430 144.940 ;
        RECT 943.070 32.540 943.390 32.600 ;
        RECT 1091.190 32.540 1091.510 32.600 ;
        RECT 943.070 32.400 1091.510 32.540 ;
        RECT 943.070 32.340 943.390 32.400 ;
        RECT 1091.190 32.340 1091.510 32.400 ;
        RECT 823.470 20.300 823.790 20.360 ;
        RECT 943.070 20.300 943.390 20.360 ;
        RECT 823.470 20.160 943.390 20.300 ;
        RECT 823.470 20.100 823.790 20.160 ;
        RECT 943.070 20.100 943.390 20.160 ;
      LAYER via ;
        RECT 1091.220 524.320 1091.480 524.580 ;
        RECT 1091.680 524.320 1091.940 524.580 ;
        RECT 1091.680 476.040 1091.940 476.300 ;
        RECT 1092.140 476.040 1092.400 476.300 ;
        RECT 1091.220 434.560 1091.480 434.820 ;
        RECT 1091.680 434.560 1091.940 434.820 ;
        RECT 1091.220 427.420 1091.480 427.680 ;
        RECT 1092.140 427.420 1092.400 427.680 ;
        RECT 1091.220 379.480 1091.480 379.740 ;
        RECT 1092.140 379.480 1092.400 379.740 ;
        RECT 1090.760 282.580 1091.020 282.840 ;
        RECT 1091.220 282.580 1091.480 282.840 ;
        RECT 1090.760 234.640 1091.020 234.900 ;
        RECT 1092.140 234.640 1092.400 234.900 ;
        RECT 1091.220 144.880 1091.480 145.140 ;
        RECT 1092.140 144.880 1092.400 145.140 ;
        RECT 943.100 32.340 943.360 32.600 ;
        RECT 1091.220 32.340 1091.480 32.600 ;
        RECT 823.500 20.100 823.760 20.360 ;
        RECT 943.100 20.100 943.360 20.360 ;
      LAYER met2 ;
        RECT 1093.750 600.850 1094.030 604.000 ;
        RECT 1091.280 600.710 1094.030 600.850 ;
        RECT 1091.280 579.770 1091.420 600.710 ;
        RECT 1093.750 600.000 1094.030 600.710 ;
        RECT 1091.280 579.630 1091.880 579.770 ;
        RECT 1091.740 524.610 1091.880 579.630 ;
        RECT 1091.220 524.290 1091.480 524.610 ;
        RECT 1091.680 524.290 1091.940 524.610 ;
        RECT 1091.280 524.125 1091.420 524.290 ;
        RECT 1091.210 523.755 1091.490 524.125 ;
        RECT 1092.130 523.075 1092.410 523.445 ;
        RECT 1092.200 476.330 1092.340 523.075 ;
        RECT 1091.680 476.010 1091.940 476.330 ;
        RECT 1092.140 476.010 1092.400 476.330 ;
        RECT 1091.740 434.850 1091.880 476.010 ;
        RECT 1091.220 434.530 1091.480 434.850 ;
        RECT 1091.680 434.530 1091.940 434.850 ;
        RECT 1091.280 427.710 1091.420 434.530 ;
        RECT 1091.220 427.390 1091.480 427.710 ;
        RECT 1092.140 427.390 1092.400 427.710 ;
        RECT 1092.200 379.770 1092.340 427.390 ;
        RECT 1091.220 379.450 1091.480 379.770 ;
        RECT 1092.140 379.450 1092.400 379.770 ;
        RECT 1091.280 282.870 1091.420 379.450 ;
        RECT 1090.760 282.550 1091.020 282.870 ;
        RECT 1091.220 282.550 1091.480 282.870 ;
        RECT 1090.820 234.930 1090.960 282.550 ;
        RECT 1090.760 234.610 1091.020 234.930 ;
        RECT 1092.140 234.610 1092.400 234.930 ;
        RECT 1092.200 145.170 1092.340 234.610 ;
        RECT 1091.220 144.850 1091.480 145.170 ;
        RECT 1092.140 144.850 1092.400 145.170 ;
        RECT 1091.280 32.630 1091.420 144.850 ;
        RECT 943.100 32.310 943.360 32.630 ;
        RECT 1091.220 32.310 1091.480 32.630 ;
        RECT 943.160 20.390 943.300 32.310 ;
        RECT 823.500 20.070 823.760 20.390 ;
        RECT 943.100 20.070 943.360 20.390 ;
        RECT 823.560 2.400 823.700 20.070 ;
        RECT 823.350 -4.800 823.910 2.400 ;
      LAYER via2 ;
        RECT 1091.210 523.800 1091.490 524.080 ;
        RECT 1092.130 523.120 1092.410 523.400 ;
      LAYER met3 ;
        RECT 1091.185 524.090 1091.515 524.105 ;
        RECT 1090.510 523.790 1091.515 524.090 ;
        RECT 1090.510 523.410 1090.810 523.790 ;
        RECT 1091.185 523.775 1091.515 523.790 ;
        RECT 1092.105 523.410 1092.435 523.425 ;
        RECT 1090.510 523.110 1092.435 523.410 ;
        RECT 1092.105 523.095 1092.435 523.110 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2607.350 19.960 2607.670 20.020 ;
        RECT 2019.560 19.820 2607.670 19.960 ;
        RECT 2014.410 19.620 2014.730 19.680 ;
        RECT 2019.560 19.620 2019.700 19.820 ;
        RECT 2607.350 19.760 2607.670 19.820 ;
        RECT 2014.410 19.480 2019.700 19.620 ;
        RECT 2014.410 19.420 2014.730 19.480 ;
      LAYER via ;
        RECT 2014.440 19.420 2014.700 19.680 ;
        RECT 2607.380 19.760 2607.640 20.020 ;
      LAYER met2 ;
        RECT 2011.910 600.170 2012.190 604.000 ;
        RECT 2011.910 600.030 2014.640 600.170 ;
        RECT 2011.910 600.000 2012.190 600.030 ;
        RECT 2014.500 19.710 2014.640 600.030 ;
        RECT 2607.380 19.730 2607.640 20.050 ;
        RECT 2014.440 19.390 2014.700 19.710 ;
        RECT 2607.440 2.400 2607.580 19.730 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2021.310 592.520 2021.630 592.580 ;
        RECT 2376.890 592.520 2377.210 592.580 ;
        RECT 2021.310 592.380 2377.210 592.520 ;
        RECT 2021.310 592.320 2021.630 592.380 ;
        RECT 2376.890 592.320 2377.210 592.380 ;
        RECT 2376.890 14.860 2377.210 14.920 ;
        RECT 2625.290 14.860 2625.610 14.920 ;
        RECT 2376.890 14.720 2625.610 14.860 ;
        RECT 2376.890 14.660 2377.210 14.720 ;
        RECT 2625.290 14.660 2625.610 14.720 ;
      LAYER via ;
        RECT 2021.340 592.320 2021.600 592.580 ;
        RECT 2376.920 592.320 2377.180 592.580 ;
        RECT 2376.920 14.660 2377.180 14.920 ;
        RECT 2625.320 14.660 2625.580 14.920 ;
      LAYER met2 ;
        RECT 2021.110 600.000 2021.390 604.000 ;
        RECT 2021.170 598.810 2021.310 600.000 ;
        RECT 2021.170 598.670 2021.540 598.810 ;
        RECT 2021.400 592.610 2021.540 598.670 ;
        RECT 2021.340 592.290 2021.600 592.610 ;
        RECT 2376.920 592.290 2377.180 592.610 ;
        RECT 2376.980 14.950 2377.120 592.290 ;
        RECT 2376.920 14.630 2377.180 14.950 ;
        RECT 2625.320 14.630 2625.580 14.950 ;
        RECT 2625.380 2.400 2625.520 14.630 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2031.890 586.740 2032.210 586.800 ;
        RECT 2035.110 586.740 2035.430 586.800 ;
        RECT 2031.890 586.600 2035.430 586.740 ;
        RECT 2031.890 586.540 2032.210 586.600 ;
        RECT 2035.110 586.540 2035.430 586.600 ;
        RECT 2035.110 19.620 2035.430 19.680 ;
        RECT 2643.230 19.620 2643.550 19.680 ;
        RECT 2035.110 19.480 2643.550 19.620 ;
        RECT 2035.110 19.420 2035.430 19.480 ;
        RECT 2643.230 19.420 2643.550 19.480 ;
      LAYER via ;
        RECT 2031.920 586.540 2032.180 586.800 ;
        RECT 2035.140 586.540 2035.400 586.800 ;
        RECT 2035.140 19.420 2035.400 19.680 ;
        RECT 2643.260 19.420 2643.520 19.680 ;
      LAYER met2 ;
        RECT 2030.310 600.170 2030.590 604.000 ;
        RECT 2030.310 600.030 2032.120 600.170 ;
        RECT 2030.310 600.000 2030.590 600.030 ;
        RECT 2031.980 586.830 2032.120 600.030 ;
        RECT 2031.920 586.510 2032.180 586.830 ;
        RECT 2035.140 586.510 2035.400 586.830 ;
        RECT 2035.200 19.710 2035.340 586.510 ;
        RECT 2035.140 19.390 2035.400 19.710 ;
        RECT 2643.260 19.390 2643.520 19.710 ;
        RECT 2643.320 2.400 2643.460 19.390 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2041.090 592.860 2041.410 592.920 ;
        RECT 2390.690 592.860 2391.010 592.920 ;
        RECT 2041.090 592.720 2391.010 592.860 ;
        RECT 2041.090 592.660 2041.410 592.720 ;
        RECT 2390.690 592.660 2391.010 592.720 ;
        RECT 2390.690 15.200 2391.010 15.260 ;
        RECT 2661.170 15.200 2661.490 15.260 ;
        RECT 2390.690 15.060 2661.490 15.200 ;
        RECT 2390.690 15.000 2391.010 15.060 ;
        RECT 2661.170 15.000 2661.490 15.060 ;
      LAYER via ;
        RECT 2041.120 592.660 2041.380 592.920 ;
        RECT 2390.720 592.660 2390.980 592.920 ;
        RECT 2390.720 15.000 2390.980 15.260 ;
        RECT 2661.200 15.000 2661.460 15.260 ;
      LAYER met2 ;
        RECT 2039.510 600.170 2039.790 604.000 ;
        RECT 2039.510 600.030 2041.320 600.170 ;
        RECT 2039.510 600.000 2039.790 600.030 ;
        RECT 2041.180 592.950 2041.320 600.030 ;
        RECT 2041.120 592.630 2041.380 592.950 ;
        RECT 2390.720 592.630 2390.980 592.950 ;
        RECT 2390.780 15.290 2390.920 592.630 ;
        RECT 2390.720 14.970 2390.980 15.290 ;
        RECT 2661.200 14.970 2661.460 15.290 ;
        RECT 2661.260 2.400 2661.400 14.970 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2047.530 45.460 2047.850 45.520 ;
        RECT 2048.910 45.460 2049.230 45.520 ;
        RECT 2047.530 45.320 2049.230 45.460 ;
        RECT 2047.530 45.260 2047.850 45.320 ;
        RECT 2048.910 45.260 2049.230 45.320 ;
        RECT 2047.530 19.280 2047.850 19.340 ;
        RECT 2678.650 19.280 2678.970 19.340 ;
        RECT 2047.530 19.140 2678.970 19.280 ;
        RECT 2047.530 19.080 2047.850 19.140 ;
        RECT 2678.650 19.080 2678.970 19.140 ;
      LAYER via ;
        RECT 2047.560 45.260 2047.820 45.520 ;
        RECT 2048.940 45.260 2049.200 45.520 ;
        RECT 2047.560 19.080 2047.820 19.340 ;
        RECT 2678.680 19.080 2678.940 19.340 ;
      LAYER met2 ;
        RECT 2048.710 600.000 2048.990 604.000 ;
        RECT 2048.770 598.810 2048.910 600.000 ;
        RECT 2048.770 598.670 2049.140 598.810 ;
        RECT 2049.000 45.550 2049.140 598.670 ;
        RECT 2047.560 45.230 2047.820 45.550 ;
        RECT 2048.940 45.230 2049.200 45.550 ;
        RECT 2047.620 19.370 2047.760 45.230 ;
        RECT 2047.560 19.050 2047.820 19.370 ;
        RECT 2678.680 19.050 2678.940 19.370 ;
        RECT 2678.740 2.400 2678.880 19.050 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2059.490 588.780 2059.810 588.840 ;
        RECT 2404.490 588.780 2404.810 588.840 ;
        RECT 2059.490 588.640 2404.810 588.780 ;
        RECT 2059.490 588.580 2059.810 588.640 ;
        RECT 2404.490 588.580 2404.810 588.640 ;
        RECT 2404.490 20.640 2404.810 20.700 ;
        RECT 2406.330 20.640 2406.650 20.700 ;
        RECT 2404.490 20.500 2406.650 20.640 ;
        RECT 2404.490 20.440 2404.810 20.500 ;
        RECT 2406.330 20.440 2406.650 20.500 ;
        RECT 2406.330 15.540 2406.650 15.600 ;
        RECT 2696.590 15.540 2696.910 15.600 ;
        RECT 2406.330 15.400 2696.910 15.540 ;
        RECT 2406.330 15.340 2406.650 15.400 ;
        RECT 2696.590 15.340 2696.910 15.400 ;
      LAYER via ;
        RECT 2059.520 588.580 2059.780 588.840 ;
        RECT 2404.520 588.580 2404.780 588.840 ;
        RECT 2404.520 20.440 2404.780 20.700 ;
        RECT 2406.360 20.440 2406.620 20.700 ;
        RECT 2406.360 15.340 2406.620 15.600 ;
        RECT 2696.620 15.340 2696.880 15.600 ;
      LAYER met2 ;
        RECT 2057.910 600.170 2058.190 604.000 ;
        RECT 2057.910 600.030 2059.720 600.170 ;
        RECT 2057.910 600.000 2058.190 600.030 ;
        RECT 2059.580 588.870 2059.720 600.030 ;
        RECT 2059.520 588.550 2059.780 588.870 ;
        RECT 2404.520 588.550 2404.780 588.870 ;
        RECT 2404.580 20.730 2404.720 588.550 ;
        RECT 2404.520 20.410 2404.780 20.730 ;
        RECT 2406.360 20.410 2406.620 20.730 ;
        RECT 2406.420 15.630 2406.560 20.410 ;
        RECT 2406.360 15.310 2406.620 15.630 ;
        RECT 2696.620 15.310 2696.880 15.630 ;
        RECT 2696.680 2.400 2696.820 15.310 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2068.690 587.420 2069.010 587.480 ;
        RECT 2073.290 587.420 2073.610 587.480 ;
        RECT 2068.690 587.280 2073.610 587.420 ;
        RECT 2068.690 587.220 2069.010 587.280 ;
        RECT 2073.290 587.220 2073.610 587.280 ;
        RECT 2073.290 18.940 2073.610 19.000 ;
        RECT 2714.530 18.940 2714.850 19.000 ;
        RECT 2073.290 18.800 2714.850 18.940 ;
        RECT 2073.290 18.740 2073.610 18.800 ;
        RECT 2714.530 18.740 2714.850 18.800 ;
      LAYER via ;
        RECT 2068.720 587.220 2068.980 587.480 ;
        RECT 2073.320 587.220 2073.580 587.480 ;
        RECT 2073.320 18.740 2073.580 19.000 ;
        RECT 2714.560 18.740 2714.820 19.000 ;
      LAYER met2 ;
        RECT 2067.110 600.170 2067.390 604.000 ;
        RECT 2067.110 600.030 2068.920 600.170 ;
        RECT 2067.110 600.000 2067.390 600.030 ;
        RECT 2068.780 587.510 2068.920 600.030 ;
        RECT 2068.720 587.190 2068.980 587.510 ;
        RECT 2073.320 587.190 2073.580 587.510 ;
        RECT 2073.380 19.030 2073.520 587.190 ;
        RECT 2073.320 18.710 2073.580 19.030 ;
        RECT 2714.560 18.710 2714.820 19.030 ;
        RECT 2714.620 2.400 2714.760 18.710 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2076.510 588.440 2076.830 588.500 ;
        RECT 2411.390 588.440 2411.710 588.500 ;
        RECT 2076.510 588.300 2411.710 588.440 ;
        RECT 2076.510 588.240 2076.830 588.300 ;
        RECT 2411.390 588.240 2411.710 588.300 ;
        RECT 2410.930 16.220 2411.250 16.280 ;
        RECT 2732.470 16.220 2732.790 16.280 ;
        RECT 2410.930 16.080 2732.790 16.220 ;
        RECT 2410.930 16.020 2411.250 16.080 ;
        RECT 2732.470 16.020 2732.790 16.080 ;
      LAYER via ;
        RECT 2076.540 588.240 2076.800 588.500 ;
        RECT 2411.420 588.240 2411.680 588.500 ;
        RECT 2410.960 16.020 2411.220 16.280 ;
        RECT 2732.500 16.020 2732.760 16.280 ;
      LAYER met2 ;
        RECT 2076.310 600.000 2076.590 604.000 ;
        RECT 2076.370 598.810 2076.510 600.000 ;
        RECT 2076.370 598.670 2076.740 598.810 ;
        RECT 2076.600 588.530 2076.740 598.670 ;
        RECT 2076.540 588.210 2076.800 588.530 ;
        RECT 2411.420 588.210 2411.680 588.530 ;
        RECT 2411.480 34.410 2411.620 588.210 ;
        RECT 2411.020 34.270 2411.620 34.410 ;
        RECT 2411.020 16.310 2411.160 34.270 ;
        RECT 2410.960 15.990 2411.220 16.310 ;
        RECT 2732.500 15.990 2732.760 16.310 ;
        RECT 2732.560 2.400 2732.700 15.990 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2087.090 592.180 2087.410 592.240 ;
        RECT 2114.230 592.180 2114.550 592.240 ;
        RECT 2087.090 592.040 2114.550 592.180 ;
        RECT 2087.090 591.980 2087.410 592.040 ;
        RECT 2114.230 591.980 2114.550 592.040 ;
        RECT 2114.230 589.120 2114.550 589.180 ;
        RECT 2432.090 589.120 2432.410 589.180 ;
        RECT 2114.230 588.980 2432.410 589.120 ;
        RECT 2114.230 588.920 2114.550 588.980 ;
        RECT 2432.090 588.920 2432.410 588.980 ;
        RECT 2432.090 15.880 2432.410 15.940 ;
        RECT 2750.410 15.880 2750.730 15.940 ;
        RECT 2432.090 15.740 2750.730 15.880 ;
        RECT 2432.090 15.680 2432.410 15.740 ;
        RECT 2750.410 15.680 2750.730 15.740 ;
      LAYER via ;
        RECT 2087.120 591.980 2087.380 592.240 ;
        RECT 2114.260 591.980 2114.520 592.240 ;
        RECT 2114.260 588.920 2114.520 589.180 ;
        RECT 2432.120 588.920 2432.380 589.180 ;
        RECT 2432.120 15.680 2432.380 15.940 ;
        RECT 2750.440 15.680 2750.700 15.940 ;
      LAYER met2 ;
        RECT 2085.510 600.170 2085.790 604.000 ;
        RECT 2085.510 600.030 2087.320 600.170 ;
        RECT 2085.510 600.000 2085.790 600.030 ;
        RECT 2087.180 592.270 2087.320 600.030 ;
        RECT 2087.120 591.950 2087.380 592.270 ;
        RECT 2114.260 591.950 2114.520 592.270 ;
        RECT 2114.320 589.210 2114.460 591.950 ;
        RECT 2114.260 588.890 2114.520 589.210 ;
        RECT 2432.120 588.890 2432.380 589.210 ;
        RECT 2432.180 15.970 2432.320 588.890 ;
        RECT 2432.120 15.650 2432.380 15.970 ;
        RECT 2750.440 15.650 2750.700 15.970 ;
        RECT 2750.500 2.400 2750.640 15.650 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2096.290 587.760 2096.610 587.820 ;
        RECT 2100.890 587.760 2101.210 587.820 ;
        RECT 2096.290 587.620 2101.210 587.760 ;
        RECT 2096.290 587.560 2096.610 587.620 ;
        RECT 2100.890 587.560 2101.210 587.620 ;
        RECT 2100.890 18.600 2101.210 18.660 ;
        RECT 2767.890 18.600 2768.210 18.660 ;
        RECT 2100.890 18.460 2768.210 18.600 ;
        RECT 2100.890 18.400 2101.210 18.460 ;
        RECT 2767.890 18.400 2768.210 18.460 ;
      LAYER via ;
        RECT 2096.320 587.560 2096.580 587.820 ;
        RECT 2100.920 587.560 2101.180 587.820 ;
        RECT 2100.920 18.400 2101.180 18.660 ;
        RECT 2767.920 18.400 2768.180 18.660 ;
      LAYER met2 ;
        RECT 2094.710 600.170 2094.990 604.000 ;
        RECT 2094.710 600.030 2096.520 600.170 ;
        RECT 2094.710 600.000 2094.990 600.030 ;
        RECT 2096.380 587.850 2096.520 600.030 ;
        RECT 2096.320 587.530 2096.580 587.850 ;
        RECT 2100.920 587.530 2101.180 587.850 ;
        RECT 2100.980 18.690 2101.120 587.530 ;
        RECT 2100.920 18.370 2101.180 18.690 ;
        RECT 2767.920 18.370 2768.180 18.690 ;
        RECT 2767.980 2.400 2768.120 18.370 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1098.550 434.760 1098.870 434.820 ;
        RECT 1099.010 434.760 1099.330 434.820 ;
        RECT 1098.550 434.620 1099.330 434.760 ;
        RECT 1098.550 434.560 1098.870 434.620 ;
        RECT 1099.010 434.560 1099.330 434.620 ;
        RECT 1098.090 331.400 1098.410 331.460 ;
        RECT 1098.550 331.400 1098.870 331.460 ;
        RECT 1098.090 331.260 1098.870 331.400 ;
        RECT 1098.090 331.200 1098.410 331.260 ;
        RECT 1098.550 331.200 1098.870 331.260 ;
        RECT 1098.090 283.460 1098.410 283.520 ;
        RECT 1099.010 283.460 1099.330 283.520 ;
        RECT 1098.090 283.320 1099.330 283.460 ;
        RECT 1098.090 283.260 1098.410 283.320 ;
        RECT 1099.010 283.260 1099.330 283.320 ;
        RECT 1098.550 227.700 1098.870 227.760 ;
        RECT 1099.470 227.700 1099.790 227.760 ;
        RECT 1098.550 227.560 1099.790 227.700 ;
        RECT 1098.550 227.500 1098.870 227.560 ;
        RECT 1099.470 227.500 1099.790 227.560 ;
        RECT 1098.550 179.760 1098.870 179.820 ;
        RECT 1099.930 179.760 1100.250 179.820 ;
        RECT 1098.550 179.620 1100.250 179.760 ;
        RECT 1098.550 179.560 1098.870 179.620 ;
        RECT 1099.930 179.560 1100.250 179.620 ;
        RECT 1099.930 145.420 1100.250 145.480 ;
        RECT 1099.100 145.280 1100.250 145.420 ;
        RECT 1099.100 144.800 1099.240 145.280 ;
        RECT 1099.930 145.220 1100.250 145.280 ;
        RECT 1099.010 144.540 1099.330 144.800 ;
        RECT 1098.550 90.000 1098.870 90.060 ;
        RECT 1099.010 90.000 1099.330 90.060 ;
        RECT 1098.550 89.860 1099.330 90.000 ;
        RECT 1098.550 89.800 1098.870 89.860 ;
        RECT 1099.010 89.800 1099.330 89.860 ;
        RECT 940.310 32.200 940.630 32.260 ;
        RECT 1098.550 32.200 1098.870 32.260 ;
        RECT 940.310 32.060 1098.870 32.200 ;
        RECT 940.310 32.000 940.630 32.060 ;
        RECT 1098.550 32.000 1098.870 32.060 ;
        RECT 840.950 14.520 841.270 14.580 ;
        RECT 940.310 14.520 940.630 14.580 ;
        RECT 840.950 14.380 940.630 14.520 ;
        RECT 840.950 14.320 841.270 14.380 ;
        RECT 940.310 14.320 940.630 14.380 ;
      LAYER via ;
        RECT 1098.580 434.560 1098.840 434.820 ;
        RECT 1099.040 434.560 1099.300 434.820 ;
        RECT 1098.120 331.200 1098.380 331.460 ;
        RECT 1098.580 331.200 1098.840 331.460 ;
        RECT 1098.120 283.260 1098.380 283.520 ;
        RECT 1099.040 283.260 1099.300 283.520 ;
        RECT 1098.580 227.500 1098.840 227.760 ;
        RECT 1099.500 227.500 1099.760 227.760 ;
        RECT 1098.580 179.560 1098.840 179.820 ;
        RECT 1099.960 179.560 1100.220 179.820 ;
        RECT 1099.960 145.220 1100.220 145.480 ;
        RECT 1099.040 144.540 1099.300 144.800 ;
        RECT 1098.580 89.800 1098.840 90.060 ;
        RECT 1099.040 89.800 1099.300 90.060 ;
        RECT 940.340 32.000 940.600 32.260 ;
        RECT 1098.580 32.000 1098.840 32.260 ;
        RECT 840.980 14.320 841.240 14.580 ;
        RECT 940.340 14.320 940.600 14.580 ;
      LAYER met2 ;
        RECT 1102.950 600.170 1103.230 604.000 ;
        RECT 1101.860 600.030 1103.230 600.170 ;
        RECT 1101.860 579.885 1102.000 600.030 ;
        RECT 1102.950 600.000 1103.230 600.030 ;
        RECT 1100.870 579.515 1101.150 579.885 ;
        RECT 1101.790 579.515 1102.070 579.885 ;
        RECT 1100.940 495.450 1101.080 579.515 ;
        RECT 1099.100 495.310 1101.080 495.450 ;
        RECT 1099.100 434.850 1099.240 495.310 ;
        RECT 1098.580 434.530 1098.840 434.850 ;
        RECT 1099.040 434.530 1099.300 434.850 ;
        RECT 1098.640 331.490 1098.780 434.530 ;
        RECT 1098.120 331.170 1098.380 331.490 ;
        RECT 1098.580 331.170 1098.840 331.490 ;
        RECT 1098.180 283.550 1098.320 331.170 ;
        RECT 1098.120 283.230 1098.380 283.550 ;
        RECT 1099.040 283.230 1099.300 283.550 ;
        RECT 1099.100 266.290 1099.240 283.230 ;
        RECT 1099.100 266.150 1100.160 266.290 ;
        RECT 1100.020 235.010 1100.160 266.150 ;
        RECT 1099.560 234.870 1100.160 235.010 ;
        RECT 1099.560 227.790 1099.700 234.870 ;
        RECT 1098.580 227.470 1098.840 227.790 ;
        RECT 1099.500 227.470 1099.760 227.790 ;
        RECT 1098.640 179.850 1098.780 227.470 ;
        RECT 1098.580 179.530 1098.840 179.850 ;
        RECT 1099.960 179.530 1100.220 179.850 ;
        RECT 1100.020 145.510 1100.160 179.530 ;
        RECT 1099.960 145.190 1100.220 145.510 ;
        RECT 1099.040 144.510 1099.300 144.830 ;
        RECT 1099.100 90.090 1099.240 144.510 ;
        RECT 1098.580 89.770 1098.840 90.090 ;
        RECT 1099.040 89.770 1099.300 90.090 ;
        RECT 1098.640 32.290 1098.780 89.770 ;
        RECT 940.340 31.970 940.600 32.290 ;
        RECT 1098.580 31.970 1098.840 32.290 ;
        RECT 940.400 14.610 940.540 31.970 ;
        RECT 840.980 14.290 841.240 14.610 ;
        RECT 940.340 14.290 940.600 14.610 ;
        RECT 841.040 2.400 841.180 14.290 ;
        RECT 840.830 -4.800 841.390 2.400 ;
      LAYER via2 ;
        RECT 1100.870 579.560 1101.150 579.840 ;
        RECT 1101.790 579.560 1102.070 579.840 ;
      LAYER met3 ;
        RECT 1100.845 579.850 1101.175 579.865 ;
        RECT 1101.765 579.850 1102.095 579.865 ;
        RECT 1100.845 579.550 1102.095 579.850 ;
        RECT 1100.845 579.535 1101.175 579.550 ;
        RECT 1101.765 579.535 1102.095 579.550 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2104.110 589.460 2104.430 589.520 ;
        RECT 2445.890 589.460 2446.210 589.520 ;
        RECT 2104.110 589.320 2446.210 589.460 ;
        RECT 2104.110 589.260 2104.430 589.320 ;
        RECT 2445.890 589.260 2446.210 589.320 ;
        RECT 2445.890 20.640 2446.210 20.700 ;
        RECT 2447.730 20.640 2448.050 20.700 ;
        RECT 2445.890 20.500 2448.050 20.640 ;
        RECT 2445.890 20.440 2446.210 20.500 ;
        RECT 2447.730 20.440 2448.050 20.500 ;
        RECT 2447.730 16.560 2448.050 16.620 ;
        RECT 2785.830 16.560 2786.150 16.620 ;
        RECT 2447.730 16.420 2786.150 16.560 ;
        RECT 2447.730 16.360 2448.050 16.420 ;
        RECT 2785.830 16.360 2786.150 16.420 ;
      LAYER via ;
        RECT 2104.140 589.260 2104.400 589.520 ;
        RECT 2445.920 589.260 2446.180 589.520 ;
        RECT 2445.920 20.440 2446.180 20.700 ;
        RECT 2447.760 20.440 2448.020 20.700 ;
        RECT 2447.760 16.360 2448.020 16.620 ;
        RECT 2785.860 16.360 2786.120 16.620 ;
      LAYER met2 ;
        RECT 2103.910 600.000 2104.190 604.000 ;
        RECT 2103.970 598.810 2104.110 600.000 ;
        RECT 2103.970 598.670 2104.340 598.810 ;
        RECT 2104.200 589.550 2104.340 598.670 ;
        RECT 2104.140 589.230 2104.400 589.550 ;
        RECT 2445.920 589.230 2446.180 589.550 ;
        RECT 2445.980 20.730 2446.120 589.230 ;
        RECT 2445.920 20.410 2446.180 20.730 ;
        RECT 2447.760 20.410 2448.020 20.730 ;
        RECT 2447.820 16.650 2447.960 20.410 ;
        RECT 2447.760 16.330 2448.020 16.650 ;
        RECT 2785.860 16.330 2786.120 16.650 ;
        RECT 2785.920 2.400 2786.060 16.330 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2114.690 586.740 2115.010 586.800 ;
        RECT 2117.910 586.740 2118.230 586.800 ;
        RECT 2114.690 586.600 2118.230 586.740 ;
        RECT 2114.690 586.540 2115.010 586.600 ;
        RECT 2117.910 586.540 2118.230 586.600 ;
        RECT 2117.910 18.260 2118.230 18.320 ;
        RECT 2803.770 18.260 2804.090 18.320 ;
        RECT 2117.910 18.120 2804.090 18.260 ;
        RECT 2117.910 18.060 2118.230 18.120 ;
        RECT 2803.770 18.060 2804.090 18.120 ;
      LAYER via ;
        RECT 2114.720 586.540 2114.980 586.800 ;
        RECT 2117.940 586.540 2118.200 586.800 ;
        RECT 2117.940 18.060 2118.200 18.320 ;
        RECT 2803.800 18.060 2804.060 18.320 ;
      LAYER met2 ;
        RECT 2113.110 600.170 2113.390 604.000 ;
        RECT 2113.110 600.030 2114.920 600.170 ;
        RECT 2113.110 600.000 2113.390 600.030 ;
        RECT 2114.780 586.830 2114.920 600.030 ;
        RECT 2114.720 586.510 2114.980 586.830 ;
        RECT 2117.940 586.510 2118.200 586.830 ;
        RECT 2118.000 18.350 2118.140 586.510 ;
        RECT 2117.940 18.030 2118.200 18.350 ;
        RECT 2803.800 18.030 2804.060 18.350 ;
        RECT 2803.860 2.400 2804.000 18.030 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2123.890 593.200 2124.210 593.260 ;
        RECT 2466.590 593.200 2466.910 593.260 ;
        RECT 2123.890 593.060 2466.910 593.200 ;
        RECT 2123.890 593.000 2124.210 593.060 ;
        RECT 2466.590 593.000 2466.910 593.060 ;
        RECT 2466.590 16.900 2466.910 16.960 ;
        RECT 2821.710 16.900 2822.030 16.960 ;
        RECT 2466.590 16.760 2822.030 16.900 ;
        RECT 2466.590 16.700 2466.910 16.760 ;
        RECT 2821.710 16.700 2822.030 16.760 ;
      LAYER via ;
        RECT 2123.920 593.000 2124.180 593.260 ;
        RECT 2466.620 593.000 2466.880 593.260 ;
        RECT 2466.620 16.700 2466.880 16.960 ;
        RECT 2821.740 16.700 2822.000 16.960 ;
      LAYER met2 ;
        RECT 2122.310 600.170 2122.590 604.000 ;
        RECT 2122.310 600.030 2124.120 600.170 ;
        RECT 2122.310 600.000 2122.590 600.030 ;
        RECT 2123.980 593.290 2124.120 600.030 ;
        RECT 2123.920 592.970 2124.180 593.290 ;
        RECT 2466.620 592.970 2466.880 593.290 ;
        RECT 2466.680 16.990 2466.820 592.970 ;
        RECT 2466.620 16.670 2466.880 16.990 ;
        RECT 2821.740 16.670 2822.000 16.990 ;
        RECT 2821.800 2.400 2821.940 16.670 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2131.710 587.420 2132.030 587.480 ;
        RECT 2149.190 587.420 2149.510 587.480 ;
        RECT 2131.710 587.280 2149.510 587.420 ;
        RECT 2131.710 587.220 2132.030 587.280 ;
        RECT 2149.190 587.220 2149.510 587.280 ;
        RECT 2149.190 17.920 2149.510 17.980 ;
        RECT 2839.190 17.920 2839.510 17.980 ;
        RECT 2149.190 17.780 2839.510 17.920 ;
        RECT 2149.190 17.720 2149.510 17.780 ;
        RECT 2839.190 17.720 2839.510 17.780 ;
      LAYER via ;
        RECT 2131.740 587.220 2132.000 587.480 ;
        RECT 2149.220 587.220 2149.480 587.480 ;
        RECT 2149.220 17.720 2149.480 17.980 ;
        RECT 2839.220 17.720 2839.480 17.980 ;
      LAYER met2 ;
        RECT 2131.510 600.000 2131.790 604.000 ;
        RECT 2131.570 598.810 2131.710 600.000 ;
        RECT 2131.570 598.670 2131.940 598.810 ;
        RECT 2131.800 587.510 2131.940 598.670 ;
        RECT 2131.740 587.190 2132.000 587.510 ;
        RECT 2149.220 587.190 2149.480 587.510 ;
        RECT 2149.280 18.010 2149.420 587.190 ;
        RECT 2149.220 17.690 2149.480 18.010 ;
        RECT 2839.220 17.690 2839.480 18.010 ;
        RECT 2839.280 2.400 2839.420 17.690 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2142.290 588.100 2142.610 588.160 ;
        RECT 2480.390 588.100 2480.710 588.160 ;
        RECT 2142.290 587.960 2480.710 588.100 ;
        RECT 2142.290 587.900 2142.610 587.960 ;
        RECT 2480.390 587.900 2480.710 587.960 ;
        RECT 2480.390 20.640 2480.710 20.700 ;
        RECT 2517.650 20.640 2517.970 20.700 ;
        RECT 2480.390 20.500 2517.970 20.640 ;
        RECT 2480.390 20.440 2480.710 20.500 ;
        RECT 2517.650 20.440 2517.970 20.500 ;
        RECT 2519.030 20.640 2519.350 20.700 ;
        RECT 2857.130 20.640 2857.450 20.700 ;
        RECT 2519.030 20.500 2857.450 20.640 ;
        RECT 2519.030 20.440 2519.350 20.500 ;
        RECT 2857.130 20.440 2857.450 20.500 ;
      LAYER via ;
        RECT 2142.320 587.900 2142.580 588.160 ;
        RECT 2480.420 587.900 2480.680 588.160 ;
        RECT 2480.420 20.440 2480.680 20.700 ;
        RECT 2517.680 20.440 2517.940 20.700 ;
        RECT 2519.060 20.440 2519.320 20.700 ;
        RECT 2857.160 20.440 2857.420 20.700 ;
      LAYER met2 ;
        RECT 2140.710 600.170 2140.990 604.000 ;
        RECT 2140.710 600.030 2142.520 600.170 ;
        RECT 2140.710 600.000 2140.990 600.030 ;
        RECT 2142.380 588.190 2142.520 600.030 ;
        RECT 2142.320 587.870 2142.580 588.190 ;
        RECT 2480.420 587.870 2480.680 588.190 ;
        RECT 2480.480 20.730 2480.620 587.870 ;
        RECT 2517.740 20.730 2519.260 20.810 ;
        RECT 2480.420 20.410 2480.680 20.730 ;
        RECT 2517.680 20.670 2519.320 20.730 ;
        RECT 2517.680 20.410 2517.940 20.670 ;
        RECT 2519.060 20.410 2519.320 20.670 ;
        RECT 2857.160 20.410 2857.420 20.730 ;
        RECT 2857.220 2.400 2857.360 20.410 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2151.490 587.760 2151.810 587.820 ;
        RECT 2156.090 587.760 2156.410 587.820 ;
        RECT 2151.490 587.620 2156.410 587.760 ;
        RECT 2151.490 587.560 2151.810 587.620 ;
        RECT 2156.090 587.560 2156.410 587.620 ;
        RECT 2156.090 17.240 2156.410 17.300 ;
        RECT 2875.070 17.240 2875.390 17.300 ;
        RECT 2156.090 17.100 2875.390 17.240 ;
        RECT 2156.090 17.040 2156.410 17.100 ;
        RECT 2875.070 17.040 2875.390 17.100 ;
      LAYER via ;
        RECT 2151.520 587.560 2151.780 587.820 ;
        RECT 2156.120 587.560 2156.380 587.820 ;
        RECT 2156.120 17.040 2156.380 17.300 ;
        RECT 2875.100 17.040 2875.360 17.300 ;
      LAYER met2 ;
        RECT 2149.910 600.170 2150.190 604.000 ;
        RECT 2149.910 600.030 2151.720 600.170 ;
        RECT 2149.910 600.000 2150.190 600.030 ;
        RECT 2151.580 587.850 2151.720 600.030 ;
        RECT 2151.520 587.530 2151.780 587.850 ;
        RECT 2156.120 587.530 2156.380 587.850 ;
        RECT 2156.180 17.330 2156.320 587.530 ;
        RECT 2156.120 17.010 2156.380 17.330 ;
        RECT 2875.100 17.010 2875.360 17.330 ;
        RECT 2875.160 2.400 2875.300 17.010 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2158.850 592.180 2159.170 592.240 ;
        RECT 2501.090 592.180 2501.410 592.240 ;
        RECT 2158.850 592.040 2501.410 592.180 ;
        RECT 2158.850 591.980 2159.170 592.040 ;
        RECT 2501.090 591.980 2501.410 592.040 ;
        RECT 2501.090 20.300 2501.410 20.360 ;
        RECT 2893.010 20.300 2893.330 20.360 ;
        RECT 2501.090 20.160 2893.330 20.300 ;
        RECT 2501.090 20.100 2501.410 20.160 ;
        RECT 2893.010 20.100 2893.330 20.160 ;
      LAYER via ;
        RECT 2158.880 591.980 2159.140 592.240 ;
        RECT 2501.120 591.980 2501.380 592.240 ;
        RECT 2501.120 20.100 2501.380 20.360 ;
        RECT 2893.040 20.100 2893.300 20.360 ;
      LAYER met2 ;
        RECT 2159.110 600.000 2159.390 604.000 ;
        RECT 2159.170 598.810 2159.310 600.000 ;
        RECT 2158.940 598.670 2159.310 598.810 ;
        RECT 2158.940 592.270 2159.080 598.670 ;
        RECT 2158.880 591.950 2159.140 592.270 ;
        RECT 2501.120 591.950 2501.380 592.270 ;
        RECT 2501.180 20.390 2501.320 591.950 ;
        RECT 2501.120 20.070 2501.380 20.390 ;
        RECT 2893.040 20.070 2893.300 20.390 ;
        RECT 2893.100 2.400 2893.240 20.070 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2169.890 586.740 2170.210 586.800 ;
        RECT 2197.490 586.740 2197.810 586.800 ;
        RECT 2169.890 586.600 2197.810 586.740 ;
        RECT 2169.890 586.540 2170.210 586.600 ;
        RECT 2197.490 586.540 2197.810 586.600 ;
        RECT 2197.490 17.580 2197.810 17.640 ;
        RECT 2910.950 17.580 2911.270 17.640 ;
        RECT 2197.490 17.440 2911.270 17.580 ;
        RECT 2197.490 17.380 2197.810 17.440 ;
        RECT 2910.950 17.380 2911.270 17.440 ;
      LAYER via ;
        RECT 2169.920 586.540 2170.180 586.800 ;
        RECT 2197.520 586.540 2197.780 586.800 ;
        RECT 2197.520 17.380 2197.780 17.640 ;
        RECT 2910.980 17.380 2911.240 17.640 ;
      LAYER met2 ;
        RECT 2168.310 600.170 2168.590 604.000 ;
        RECT 2168.310 600.030 2170.120 600.170 ;
        RECT 2168.310 600.000 2168.590 600.030 ;
        RECT 2169.980 586.830 2170.120 600.030 ;
        RECT 2169.920 586.510 2170.180 586.830 ;
        RECT 2197.520 586.510 2197.780 586.830 ;
        RECT 2197.580 17.670 2197.720 586.510 ;
        RECT 2197.520 17.350 2197.780 17.670 ;
        RECT 2910.980 17.350 2911.240 17.670 ;
        RECT 2911.040 2.400 2911.180 17.350 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 858.890 39.000 859.210 39.060 ;
        RECT 1111.430 39.000 1111.750 39.060 ;
        RECT 858.890 38.860 1111.750 39.000 ;
        RECT 858.890 38.800 859.210 38.860 ;
        RECT 1111.430 38.800 1111.750 38.860 ;
      LAYER via ;
        RECT 858.920 38.800 859.180 39.060 ;
        RECT 1111.460 38.800 1111.720 39.060 ;
      LAYER met2 ;
        RECT 1112.150 600.170 1112.430 604.000 ;
        RECT 1111.520 600.030 1112.430 600.170 ;
        RECT 1111.520 39.090 1111.660 600.030 ;
        RECT 1112.150 600.000 1112.430 600.030 ;
        RECT 858.920 38.770 859.180 39.090 ;
        RECT 1111.460 38.770 1111.720 39.090 ;
        RECT 858.980 2.400 859.120 38.770 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 590.480 883.130 590.540 ;
        RECT 1119.710 590.480 1120.030 590.540 ;
        RECT 882.810 590.340 1120.030 590.480 ;
        RECT 882.810 590.280 883.130 590.340 ;
        RECT 1119.710 590.280 1120.030 590.340 ;
        RECT 876.830 20.640 877.150 20.700 ;
        RECT 882.810 20.640 883.130 20.700 ;
        RECT 876.830 20.500 883.130 20.640 ;
        RECT 876.830 20.440 877.150 20.500 ;
        RECT 882.810 20.440 883.130 20.500 ;
      LAYER via ;
        RECT 882.840 590.280 883.100 590.540 ;
        RECT 1119.740 590.280 1120.000 590.540 ;
        RECT 876.860 20.440 877.120 20.700 ;
        RECT 882.840 20.440 883.100 20.700 ;
      LAYER met2 ;
        RECT 1121.350 600.170 1121.630 604.000 ;
        RECT 1119.800 600.030 1121.630 600.170 ;
        RECT 1119.800 590.570 1119.940 600.030 ;
        RECT 1121.350 600.000 1121.630 600.030 ;
        RECT 882.840 590.250 883.100 590.570 ;
        RECT 1119.740 590.250 1120.000 590.570 ;
        RECT 882.900 20.730 883.040 590.250 ;
        RECT 876.860 20.410 877.120 20.730 ;
        RECT 882.840 20.410 883.100 20.730 ;
        RECT 876.920 2.400 877.060 20.410 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.610 590.820 896.930 590.880 ;
        RECT 1128.910 590.820 1129.230 590.880 ;
        RECT 896.610 590.680 1129.230 590.820 ;
        RECT 896.610 590.620 896.930 590.680 ;
        RECT 1128.910 590.620 1129.230 590.680 ;
        RECT 894.770 2.960 895.090 3.020 ;
        RECT 896.610 2.960 896.930 3.020 ;
        RECT 894.770 2.820 896.930 2.960 ;
        RECT 894.770 2.760 895.090 2.820 ;
        RECT 896.610 2.760 896.930 2.820 ;
      LAYER via ;
        RECT 896.640 590.620 896.900 590.880 ;
        RECT 1128.940 590.620 1129.200 590.880 ;
        RECT 894.800 2.760 895.060 3.020 ;
        RECT 896.640 2.760 896.900 3.020 ;
      LAYER met2 ;
        RECT 1130.550 600.170 1130.830 604.000 ;
        RECT 1129.000 600.030 1130.830 600.170 ;
        RECT 1129.000 590.910 1129.140 600.030 ;
        RECT 1130.550 600.000 1130.830 600.030 ;
        RECT 896.640 590.590 896.900 590.910 ;
        RECT 1128.940 590.590 1129.200 590.910 ;
        RECT 896.700 3.050 896.840 590.590 ;
        RECT 894.800 2.730 895.060 3.050 ;
        RECT 896.640 2.730 896.900 3.050 ;
        RECT 894.860 2.400 895.000 2.730 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 591.500 917.630 591.560 ;
        RECT 1138.570 591.500 1138.890 591.560 ;
        RECT 917.310 591.360 1138.890 591.500 ;
        RECT 917.310 591.300 917.630 591.360 ;
        RECT 1138.570 591.300 1138.890 591.360 ;
        RECT 912.710 20.640 913.030 20.700 ;
        RECT 917.310 20.640 917.630 20.700 ;
        RECT 912.710 20.500 917.630 20.640 ;
        RECT 912.710 20.440 913.030 20.500 ;
        RECT 917.310 20.440 917.630 20.500 ;
      LAYER via ;
        RECT 917.340 591.300 917.600 591.560 ;
        RECT 1138.600 591.300 1138.860 591.560 ;
        RECT 912.740 20.440 913.000 20.700 ;
        RECT 917.340 20.440 917.600 20.700 ;
      LAYER met2 ;
        RECT 1139.750 600.170 1140.030 604.000 ;
        RECT 1138.660 600.030 1140.030 600.170 ;
        RECT 1138.660 591.590 1138.800 600.030 ;
        RECT 1139.750 600.000 1140.030 600.030 ;
        RECT 917.340 591.270 917.600 591.590 ;
        RECT 1138.600 591.270 1138.860 591.590 ;
        RECT 917.400 20.730 917.540 591.270 ;
        RECT 912.740 20.410 913.000 20.730 ;
        RECT 917.340 20.410 917.600 20.730 ;
        RECT 912.800 2.400 912.940 20.410 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.110 592.180 931.430 592.240 ;
        RECT 1147.310 592.180 1147.630 592.240 ;
        RECT 931.110 592.040 1147.630 592.180 ;
        RECT 931.110 591.980 931.430 592.040 ;
        RECT 1147.310 591.980 1147.630 592.040 ;
        RECT 930.190 483.040 930.510 483.100 ;
        RECT 931.110 483.040 931.430 483.100 ;
        RECT 930.190 482.900 931.430 483.040 ;
        RECT 930.190 482.840 930.510 482.900 ;
        RECT 931.110 482.840 931.430 482.900 ;
        RECT 929.730 475.900 930.050 475.960 ;
        RECT 930.190 475.900 930.510 475.960 ;
        RECT 929.730 475.760 930.510 475.900 ;
        RECT 929.730 475.700 930.050 475.760 ;
        RECT 930.190 475.700 930.510 475.760 ;
        RECT 929.730 427.960 930.050 428.020 ;
        RECT 931.110 427.960 931.430 428.020 ;
        RECT 929.730 427.820 931.430 427.960 ;
        RECT 929.730 427.760 930.050 427.820 ;
        RECT 931.110 427.760 931.430 427.820 ;
        RECT 931.110 379.820 931.430 380.080 ;
        RECT 931.200 379.400 931.340 379.820 ;
        RECT 931.110 379.140 931.430 379.400 ;
        RECT 931.110 372.880 931.430 372.940 ;
        RECT 932.950 372.880 933.270 372.940 ;
        RECT 931.110 372.740 933.270 372.880 ;
        RECT 931.110 372.680 931.430 372.740 ;
        RECT 932.950 372.680 933.270 372.740 ;
        RECT 931.110 331.740 931.430 331.800 ;
        RECT 932.950 331.740 933.270 331.800 ;
        RECT 931.110 331.600 933.270 331.740 ;
        RECT 931.110 331.540 931.430 331.600 ;
        RECT 932.950 331.540 933.270 331.600 ;
        RECT 930.650 331.060 930.970 331.120 ;
        RECT 931.110 331.060 931.430 331.120 ;
        RECT 930.650 330.920 931.430 331.060 ;
        RECT 930.650 330.860 930.970 330.920 ;
        RECT 931.110 330.860 931.430 330.920 ;
        RECT 930.650 283.120 930.970 283.180 ;
        RECT 931.110 283.120 931.430 283.180 ;
        RECT 930.650 282.980 931.430 283.120 ;
        RECT 930.650 282.920 930.970 282.980 ;
        RECT 931.110 282.920 931.430 282.980 ;
        RECT 929.270 48.520 929.590 48.580 ;
        RECT 930.190 48.520 930.510 48.580 ;
        RECT 929.270 48.380 930.510 48.520 ;
        RECT 929.270 48.320 929.590 48.380 ;
        RECT 930.190 48.320 930.510 48.380 ;
      LAYER via ;
        RECT 931.140 591.980 931.400 592.240 ;
        RECT 1147.340 591.980 1147.600 592.240 ;
        RECT 930.220 482.840 930.480 483.100 ;
        RECT 931.140 482.840 931.400 483.100 ;
        RECT 929.760 475.700 930.020 475.960 ;
        RECT 930.220 475.700 930.480 475.960 ;
        RECT 929.760 427.760 930.020 428.020 ;
        RECT 931.140 427.760 931.400 428.020 ;
        RECT 931.140 379.820 931.400 380.080 ;
        RECT 931.140 379.140 931.400 379.400 ;
        RECT 931.140 372.680 931.400 372.940 ;
        RECT 932.980 372.680 933.240 372.940 ;
        RECT 931.140 331.540 931.400 331.800 ;
        RECT 932.980 331.540 933.240 331.800 ;
        RECT 930.680 330.860 930.940 331.120 ;
        RECT 931.140 330.860 931.400 331.120 ;
        RECT 930.680 282.920 930.940 283.180 ;
        RECT 931.140 282.920 931.400 283.180 ;
        RECT 929.300 48.320 929.560 48.580 ;
        RECT 930.220 48.320 930.480 48.580 ;
      LAYER met2 ;
        RECT 1148.950 600.170 1149.230 604.000 ;
        RECT 1147.400 600.030 1149.230 600.170 ;
        RECT 1147.400 592.270 1147.540 600.030 ;
        RECT 1148.950 600.000 1149.230 600.030 ;
        RECT 931.140 591.950 931.400 592.270 ;
        RECT 1147.340 591.950 1147.600 592.270 ;
        RECT 931.200 483.130 931.340 591.950 ;
        RECT 930.220 482.810 930.480 483.130 ;
        RECT 931.140 482.810 931.400 483.130 ;
        RECT 930.280 475.990 930.420 482.810 ;
        RECT 929.760 475.670 930.020 475.990 ;
        RECT 930.220 475.670 930.480 475.990 ;
        RECT 929.820 428.050 929.960 475.670 ;
        RECT 929.760 427.730 930.020 428.050 ;
        RECT 931.140 427.730 931.400 428.050 ;
        RECT 931.200 380.110 931.340 427.730 ;
        RECT 931.140 379.790 931.400 380.110 ;
        RECT 931.140 379.110 931.400 379.430 ;
        RECT 931.200 372.970 931.340 379.110 ;
        RECT 931.140 372.650 931.400 372.970 ;
        RECT 932.980 372.650 933.240 372.970 ;
        RECT 933.040 331.830 933.180 372.650 ;
        RECT 931.140 331.510 931.400 331.830 ;
        RECT 932.980 331.510 933.240 331.830 ;
        RECT 931.200 331.150 931.340 331.510 ;
        RECT 930.680 330.830 930.940 331.150 ;
        RECT 931.140 330.830 931.400 331.150 ;
        RECT 930.740 283.210 930.880 330.830 ;
        RECT 930.680 282.890 930.940 283.210 ;
        RECT 931.140 282.890 931.400 283.210 ;
        RECT 931.200 137.770 931.340 282.890 ;
        RECT 929.360 137.630 931.340 137.770 ;
        RECT 929.360 48.610 929.500 137.630 ;
        RECT 929.300 48.290 929.560 48.610 ;
        RECT 930.220 48.290 930.480 48.610 ;
        RECT 930.280 2.400 930.420 48.290 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1127.990 586.740 1128.310 586.800 ;
        RECT 1156.510 586.740 1156.830 586.800 ;
        RECT 1127.990 586.600 1156.830 586.740 ;
        RECT 1127.990 586.540 1128.310 586.600 ;
        RECT 1156.510 586.540 1156.830 586.600 ;
        RECT 948.130 20.300 948.450 20.360 ;
        RECT 1127.990 20.300 1128.310 20.360 ;
        RECT 948.130 20.160 1128.310 20.300 ;
        RECT 948.130 20.100 948.450 20.160 ;
        RECT 1127.990 20.100 1128.310 20.160 ;
      LAYER via ;
        RECT 1128.020 586.540 1128.280 586.800 ;
        RECT 1156.540 586.540 1156.800 586.800 ;
        RECT 948.160 20.100 948.420 20.360 ;
        RECT 1128.020 20.100 1128.280 20.360 ;
      LAYER met2 ;
        RECT 1158.150 600.170 1158.430 604.000 ;
        RECT 1156.600 600.030 1158.430 600.170 ;
        RECT 1156.600 586.830 1156.740 600.030 ;
        RECT 1158.150 600.000 1158.430 600.030 ;
        RECT 1128.020 586.510 1128.280 586.830 ;
        RECT 1156.540 586.510 1156.800 586.830 ;
        RECT 1128.080 20.390 1128.220 586.510 ;
        RECT 948.160 20.070 948.420 20.390 ;
        RECT 1128.020 20.070 1128.280 20.390 ;
        RECT 948.220 2.400 948.360 20.070 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.510 591.840 972.830 591.900 ;
        RECT 1166.170 591.840 1166.490 591.900 ;
        RECT 972.510 591.700 1166.490 591.840 ;
        RECT 972.510 591.640 972.830 591.700 ;
        RECT 1166.170 591.640 1166.490 591.700 ;
        RECT 966.070 16.560 966.390 16.620 ;
        RECT 972.510 16.560 972.830 16.620 ;
        RECT 966.070 16.420 972.830 16.560 ;
        RECT 966.070 16.360 966.390 16.420 ;
        RECT 972.510 16.360 972.830 16.420 ;
      LAYER via ;
        RECT 972.540 591.640 972.800 591.900 ;
        RECT 1166.200 591.640 1166.460 591.900 ;
        RECT 966.100 16.360 966.360 16.620 ;
        RECT 972.540 16.360 972.800 16.620 ;
      LAYER met2 ;
        RECT 1167.350 600.170 1167.630 604.000 ;
        RECT 1166.260 600.030 1167.630 600.170 ;
        RECT 1166.260 591.930 1166.400 600.030 ;
        RECT 1167.350 600.000 1167.630 600.030 ;
        RECT 972.540 591.610 972.800 591.930 ;
        RECT 1166.200 591.610 1166.460 591.930 ;
        RECT 972.600 16.650 972.740 591.610 ;
        RECT 966.100 16.330 966.360 16.650 ;
        RECT 972.540 16.330 972.800 16.650 ;
        RECT 966.160 2.400 966.300 16.330 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 986.310 589.460 986.630 589.520 ;
        RECT 1174.910 589.460 1175.230 589.520 ;
        RECT 986.310 589.320 1175.230 589.460 ;
        RECT 986.310 589.260 986.630 589.320 ;
        RECT 1174.910 589.260 1175.230 589.320 ;
        RECT 984.010 20.640 984.330 20.700 ;
        RECT 986.310 20.640 986.630 20.700 ;
        RECT 984.010 20.500 986.630 20.640 ;
        RECT 984.010 20.440 984.330 20.500 ;
        RECT 986.310 20.440 986.630 20.500 ;
      LAYER via ;
        RECT 986.340 589.260 986.600 589.520 ;
        RECT 1174.940 589.260 1175.200 589.520 ;
        RECT 984.040 20.440 984.300 20.700 ;
        RECT 986.340 20.440 986.600 20.700 ;
      LAYER met2 ;
        RECT 1176.550 600.170 1176.830 604.000 ;
        RECT 1175.000 600.030 1176.830 600.170 ;
        RECT 1175.000 589.550 1175.140 600.030 ;
        RECT 1176.550 600.000 1176.830 600.030 ;
        RECT 986.340 589.230 986.600 589.550 ;
        RECT 1174.940 589.230 1175.200 589.550 ;
        RECT 986.400 20.730 986.540 589.230 ;
        RECT 984.040 20.410 984.300 20.730 ;
        RECT 986.340 20.410 986.600 20.730 ;
        RECT 984.100 2.400 984.240 20.410 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.470 569.400 1007.790 569.460 ;
        RECT 1009.310 569.400 1009.630 569.460 ;
        RECT 1007.470 569.260 1009.630 569.400 ;
        RECT 1007.470 569.200 1007.790 569.260 ;
        RECT 1009.310 569.200 1009.630 569.260 ;
        RECT 662.930 43.420 663.250 43.480 ;
        RECT 1007.470 43.420 1007.790 43.480 ;
        RECT 662.930 43.280 1007.790 43.420 ;
        RECT 662.930 43.220 663.250 43.280 ;
        RECT 1007.470 43.220 1007.790 43.280 ;
      LAYER via ;
        RECT 1007.500 569.200 1007.760 569.460 ;
        RECT 1009.340 569.200 1009.600 569.460 ;
        RECT 662.960 43.220 663.220 43.480 ;
        RECT 1007.500 43.220 1007.760 43.480 ;
      LAYER met2 ;
        RECT 1010.950 600.170 1011.230 604.000 ;
        RECT 1009.400 600.030 1011.230 600.170 ;
        RECT 1009.400 569.490 1009.540 600.030 ;
        RECT 1010.950 600.000 1011.230 600.030 ;
        RECT 1007.500 569.170 1007.760 569.490 ;
        RECT 1009.340 569.170 1009.600 569.490 ;
        RECT 1007.560 43.510 1007.700 569.170 ;
        RECT 662.960 43.190 663.220 43.510 ;
        RECT 1007.500 43.190 1007.760 43.510 ;
        RECT 663.020 2.400 663.160 43.190 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1121.090 588.100 1121.410 588.160 ;
        RECT 1184.110 588.100 1184.430 588.160 ;
        RECT 1121.090 587.960 1184.430 588.100 ;
        RECT 1121.090 587.900 1121.410 587.960 ;
        RECT 1184.110 587.900 1184.430 587.960 ;
        RECT 1001.950 16.220 1002.270 16.280 ;
        RECT 1121.090 16.220 1121.410 16.280 ;
        RECT 1001.950 16.080 1121.410 16.220 ;
        RECT 1001.950 16.020 1002.270 16.080 ;
        RECT 1121.090 16.020 1121.410 16.080 ;
      LAYER via ;
        RECT 1121.120 587.900 1121.380 588.160 ;
        RECT 1184.140 587.900 1184.400 588.160 ;
        RECT 1001.980 16.020 1002.240 16.280 ;
        RECT 1121.120 16.020 1121.380 16.280 ;
      LAYER met2 ;
        RECT 1185.750 600.170 1186.030 604.000 ;
        RECT 1184.200 600.030 1186.030 600.170 ;
        RECT 1184.200 588.190 1184.340 600.030 ;
        RECT 1185.750 600.000 1186.030 600.030 ;
        RECT 1121.120 587.870 1121.380 588.190 ;
        RECT 1184.140 587.870 1184.400 588.190 ;
        RECT 1121.180 16.310 1121.320 587.870 ;
        RECT 1001.980 15.990 1002.240 16.310 ;
        RECT 1121.120 15.990 1121.380 16.310 ;
        RECT 1002.040 2.400 1002.180 15.990 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1148.690 587.420 1149.010 587.480 ;
        RECT 1194.230 587.420 1194.550 587.480 ;
        RECT 1148.690 587.280 1194.550 587.420 ;
        RECT 1148.690 587.220 1149.010 587.280 ;
        RECT 1194.230 587.220 1194.550 587.280 ;
        RECT 1019.430 20.640 1019.750 20.700 ;
        RECT 1148.690 20.640 1149.010 20.700 ;
        RECT 1019.430 20.500 1149.010 20.640 ;
        RECT 1019.430 20.440 1019.750 20.500 ;
        RECT 1148.690 20.440 1149.010 20.500 ;
      LAYER via ;
        RECT 1148.720 587.220 1148.980 587.480 ;
        RECT 1194.260 587.220 1194.520 587.480 ;
        RECT 1019.460 20.440 1019.720 20.700 ;
        RECT 1148.720 20.440 1148.980 20.700 ;
      LAYER met2 ;
        RECT 1194.950 600.170 1195.230 604.000 ;
        RECT 1194.320 600.030 1195.230 600.170 ;
        RECT 1194.320 587.510 1194.460 600.030 ;
        RECT 1194.950 600.000 1195.230 600.030 ;
        RECT 1148.720 587.190 1148.980 587.510 ;
        RECT 1194.260 587.190 1194.520 587.510 ;
        RECT 1148.780 20.730 1148.920 587.190 ;
        RECT 1019.460 20.410 1019.720 20.730 ;
        RECT 1148.720 20.410 1148.980 20.730 ;
        RECT 1019.520 2.400 1019.660 20.410 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 588.100 1186.730 588.160 ;
        RECT 1202.050 588.100 1202.370 588.160 ;
        RECT 1186.410 587.960 1202.370 588.100 ;
        RECT 1186.410 587.900 1186.730 587.960 ;
        RECT 1202.050 587.900 1202.370 587.960 ;
        RECT 1162.950 586.740 1163.270 586.800 ;
        RECT 1186.410 586.740 1186.730 586.800 ;
        RECT 1162.950 586.600 1186.730 586.740 ;
        RECT 1162.950 586.540 1163.270 586.600 ;
        RECT 1186.410 586.540 1186.730 586.600 ;
        RECT 1037.370 16.560 1037.690 16.620 ;
        RECT 1126.150 16.560 1126.470 16.620 ;
        RECT 1037.370 16.420 1126.470 16.560 ;
        RECT 1037.370 16.360 1037.690 16.420 ;
        RECT 1126.150 16.360 1126.470 16.420 ;
        RECT 1126.150 14.860 1126.470 14.920 ;
        RECT 1162.950 14.860 1163.270 14.920 ;
        RECT 1126.150 14.720 1163.270 14.860 ;
        RECT 1126.150 14.660 1126.470 14.720 ;
        RECT 1162.950 14.660 1163.270 14.720 ;
      LAYER via ;
        RECT 1186.440 587.900 1186.700 588.160 ;
        RECT 1202.080 587.900 1202.340 588.160 ;
        RECT 1162.980 586.540 1163.240 586.800 ;
        RECT 1186.440 586.540 1186.700 586.800 ;
        RECT 1037.400 16.360 1037.660 16.620 ;
        RECT 1126.180 16.360 1126.440 16.620 ;
        RECT 1126.180 14.660 1126.440 14.920 ;
        RECT 1162.980 14.660 1163.240 14.920 ;
      LAYER met2 ;
        RECT 1203.690 600.170 1203.970 604.000 ;
        RECT 1202.140 600.030 1203.970 600.170 ;
        RECT 1202.140 588.190 1202.280 600.030 ;
        RECT 1203.690 600.000 1203.970 600.030 ;
        RECT 1186.440 587.870 1186.700 588.190 ;
        RECT 1202.080 587.870 1202.340 588.190 ;
        RECT 1186.500 586.830 1186.640 587.870 ;
        RECT 1162.980 586.510 1163.240 586.830 ;
        RECT 1186.440 586.510 1186.700 586.830 ;
        RECT 1037.400 16.330 1037.660 16.650 ;
        RECT 1126.180 16.330 1126.440 16.650 ;
        RECT 1037.460 2.400 1037.600 16.330 ;
        RECT 1126.240 14.950 1126.380 16.330 ;
        RECT 1163.040 14.950 1163.180 586.510 ;
        RECT 1126.180 14.630 1126.440 14.950 ;
        RECT 1162.980 14.630 1163.240 14.950 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.990 586.740 1197.310 586.800 ;
        RECT 1211.250 586.740 1211.570 586.800 ;
        RECT 1196.990 586.600 1211.570 586.740 ;
        RECT 1196.990 586.540 1197.310 586.600 ;
        RECT 1211.250 586.540 1211.570 586.600 ;
        RECT 1055.310 19.280 1055.630 19.340 ;
        RECT 1196.990 19.280 1197.310 19.340 ;
        RECT 1055.310 19.140 1197.310 19.280 ;
        RECT 1055.310 19.080 1055.630 19.140 ;
        RECT 1196.990 19.080 1197.310 19.140 ;
      LAYER via ;
        RECT 1197.020 586.540 1197.280 586.800 ;
        RECT 1211.280 586.540 1211.540 586.800 ;
        RECT 1055.340 19.080 1055.600 19.340 ;
        RECT 1197.020 19.080 1197.280 19.340 ;
      LAYER met2 ;
        RECT 1212.890 600.170 1213.170 604.000 ;
        RECT 1211.340 600.030 1213.170 600.170 ;
        RECT 1211.340 586.830 1211.480 600.030 ;
        RECT 1212.890 600.000 1213.170 600.030 ;
        RECT 1197.020 586.510 1197.280 586.830 ;
        RECT 1211.280 586.510 1211.540 586.830 ;
        RECT 1197.080 19.370 1197.220 586.510 ;
        RECT 1055.340 19.050 1055.600 19.370 ;
        RECT 1197.020 19.050 1197.280 19.370 ;
        RECT 1055.400 2.400 1055.540 19.050 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1169.390 588.440 1169.710 588.500 ;
        RECT 1221.370 588.440 1221.690 588.500 ;
        RECT 1169.390 588.300 1221.690 588.440 ;
        RECT 1169.390 588.240 1169.710 588.300 ;
        RECT 1221.370 588.240 1221.690 588.300 ;
        RECT 1073.250 15.540 1073.570 15.600 ;
        RECT 1169.390 15.540 1169.710 15.600 ;
        RECT 1073.250 15.400 1169.710 15.540 ;
        RECT 1073.250 15.340 1073.570 15.400 ;
        RECT 1169.390 15.340 1169.710 15.400 ;
      LAYER via ;
        RECT 1169.420 588.240 1169.680 588.500 ;
        RECT 1221.400 588.240 1221.660 588.500 ;
        RECT 1073.280 15.340 1073.540 15.600 ;
        RECT 1169.420 15.340 1169.680 15.600 ;
      LAYER met2 ;
        RECT 1222.090 600.170 1222.370 604.000 ;
        RECT 1221.460 600.030 1222.370 600.170 ;
        RECT 1221.460 588.530 1221.600 600.030 ;
        RECT 1222.090 600.000 1222.370 600.030 ;
        RECT 1169.420 588.210 1169.680 588.530 ;
        RECT 1221.400 588.210 1221.660 588.530 ;
        RECT 1169.480 15.630 1169.620 588.210 ;
        RECT 1073.280 15.310 1073.540 15.630 ;
        RECT 1169.420 15.310 1169.680 15.630 ;
        RECT 1073.340 2.400 1073.480 15.310 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1090.730 17.240 1091.050 17.300 ;
        RECT 1229.190 17.240 1229.510 17.300 ;
        RECT 1090.730 17.100 1229.510 17.240 ;
        RECT 1090.730 17.040 1091.050 17.100 ;
        RECT 1229.190 17.040 1229.510 17.100 ;
      LAYER via ;
        RECT 1090.760 17.040 1091.020 17.300 ;
        RECT 1229.220 17.040 1229.480 17.300 ;
      LAYER met2 ;
        RECT 1231.290 600.170 1231.570 604.000 ;
        RECT 1229.280 600.030 1231.570 600.170 ;
        RECT 1229.280 17.330 1229.420 600.030 ;
        RECT 1231.290 600.000 1231.570 600.030 ;
        RECT 1090.760 17.010 1091.020 17.330 ;
        RECT 1229.220 17.010 1229.480 17.330 ;
        RECT 1090.820 2.400 1090.960 17.010 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1176.290 587.760 1176.610 587.820 ;
        RECT 1238.850 587.760 1239.170 587.820 ;
        RECT 1176.290 587.620 1239.170 587.760 ;
        RECT 1176.290 587.560 1176.610 587.620 ;
        RECT 1238.850 587.560 1239.170 587.620 ;
        RECT 1108.670 14.860 1108.990 14.920 ;
        RECT 1108.670 14.720 1125.920 14.860 ;
        RECT 1108.670 14.660 1108.990 14.720 ;
        RECT 1125.780 14.180 1125.920 14.720 ;
        RECT 1176.290 14.180 1176.610 14.240 ;
        RECT 1125.780 14.040 1176.610 14.180 ;
        RECT 1176.290 13.980 1176.610 14.040 ;
      LAYER via ;
        RECT 1176.320 587.560 1176.580 587.820 ;
        RECT 1238.880 587.560 1239.140 587.820 ;
        RECT 1108.700 14.660 1108.960 14.920 ;
        RECT 1176.320 13.980 1176.580 14.240 ;
      LAYER met2 ;
        RECT 1240.490 600.170 1240.770 604.000 ;
        RECT 1238.940 600.030 1240.770 600.170 ;
        RECT 1238.940 587.850 1239.080 600.030 ;
        RECT 1240.490 600.000 1240.770 600.030 ;
        RECT 1176.320 587.530 1176.580 587.850 ;
        RECT 1238.880 587.530 1239.140 587.850 ;
        RECT 1108.700 14.630 1108.960 14.950 ;
        RECT 1108.760 2.400 1108.900 14.630 ;
        RECT 1176.380 14.270 1176.520 587.530 ;
        RECT 1176.320 13.950 1176.580 14.270 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.990 593.200 1197.310 593.260 ;
        RECT 1248.970 593.200 1249.290 593.260 ;
        RECT 1196.990 593.060 1249.290 593.200 ;
        RECT 1196.990 593.000 1197.310 593.060 ;
        RECT 1248.970 593.000 1249.290 593.060 ;
        RECT 1131.210 589.800 1131.530 589.860 ;
        RECT 1196.990 589.800 1197.310 589.860 ;
        RECT 1131.210 589.660 1197.310 589.800 ;
        RECT 1131.210 589.600 1131.530 589.660 ;
        RECT 1196.990 589.600 1197.310 589.660 ;
        RECT 1126.610 16.560 1126.930 16.620 ;
        RECT 1131.210 16.560 1131.530 16.620 ;
        RECT 1126.610 16.420 1131.530 16.560 ;
        RECT 1126.610 16.360 1126.930 16.420 ;
        RECT 1131.210 16.360 1131.530 16.420 ;
      LAYER via ;
        RECT 1197.020 593.000 1197.280 593.260 ;
        RECT 1249.000 593.000 1249.260 593.260 ;
        RECT 1131.240 589.600 1131.500 589.860 ;
        RECT 1197.020 589.600 1197.280 589.860 ;
        RECT 1126.640 16.360 1126.900 16.620 ;
        RECT 1131.240 16.360 1131.500 16.620 ;
      LAYER met2 ;
        RECT 1249.690 600.170 1249.970 604.000 ;
        RECT 1249.060 600.030 1249.970 600.170 ;
        RECT 1249.060 593.290 1249.200 600.030 ;
        RECT 1249.690 600.000 1249.970 600.030 ;
        RECT 1197.020 592.970 1197.280 593.290 ;
        RECT 1249.000 592.970 1249.260 593.290 ;
        RECT 1197.080 589.890 1197.220 592.970 ;
        RECT 1131.240 589.570 1131.500 589.890 ;
        RECT 1197.020 589.570 1197.280 589.890 ;
        RECT 1131.300 16.650 1131.440 589.570 ;
        RECT 1126.640 16.330 1126.900 16.650 ;
        RECT 1131.240 16.330 1131.500 16.650 ;
        RECT 1126.700 2.400 1126.840 16.330 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1252.190 586.740 1252.510 586.800 ;
        RECT 1257.250 586.740 1257.570 586.800 ;
        RECT 1252.190 586.600 1257.570 586.740 ;
        RECT 1252.190 586.540 1252.510 586.600 ;
        RECT 1257.250 586.540 1257.570 586.600 ;
        RECT 1144.550 18.940 1144.870 19.000 ;
        RECT 1144.550 18.800 1146.620 18.940 ;
        RECT 1144.550 18.740 1144.870 18.800 ;
        RECT 1146.480 18.260 1146.620 18.800 ;
        RECT 1252.190 18.260 1252.510 18.320 ;
        RECT 1146.480 18.120 1252.510 18.260 ;
        RECT 1252.190 18.060 1252.510 18.120 ;
      LAYER via ;
        RECT 1252.220 586.540 1252.480 586.800 ;
        RECT 1257.280 586.540 1257.540 586.800 ;
        RECT 1144.580 18.740 1144.840 19.000 ;
        RECT 1252.220 18.060 1252.480 18.320 ;
      LAYER met2 ;
        RECT 1258.890 600.170 1259.170 604.000 ;
        RECT 1257.340 600.030 1259.170 600.170 ;
        RECT 1257.340 586.830 1257.480 600.030 ;
        RECT 1258.890 600.000 1259.170 600.030 ;
        RECT 1252.220 586.510 1252.480 586.830 ;
        RECT 1257.280 586.510 1257.540 586.830 ;
        RECT 1144.580 18.710 1144.840 19.030 ;
        RECT 1144.640 2.400 1144.780 18.710 ;
        RECT 1252.280 18.350 1252.420 586.510 ;
        RECT 1252.220 18.030 1252.480 18.350 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 591.160 1166.030 591.220 ;
        RECT 1266.450 591.160 1266.770 591.220 ;
        RECT 1165.710 591.020 1266.770 591.160 ;
        RECT 1165.710 590.960 1166.030 591.020 ;
        RECT 1266.450 590.960 1266.770 591.020 ;
        RECT 1162.490 20.640 1162.810 20.700 ;
        RECT 1165.710 20.640 1166.030 20.700 ;
        RECT 1162.490 20.500 1166.030 20.640 ;
        RECT 1162.490 20.440 1162.810 20.500 ;
        RECT 1165.710 20.440 1166.030 20.500 ;
      LAYER via ;
        RECT 1165.740 590.960 1166.000 591.220 ;
        RECT 1266.480 590.960 1266.740 591.220 ;
        RECT 1162.520 20.440 1162.780 20.700 ;
        RECT 1165.740 20.440 1166.000 20.700 ;
      LAYER met2 ;
        RECT 1268.090 600.170 1268.370 604.000 ;
        RECT 1266.540 600.030 1268.370 600.170 ;
        RECT 1266.540 591.250 1266.680 600.030 ;
        RECT 1268.090 600.000 1268.370 600.030 ;
        RECT 1165.740 590.930 1166.000 591.250 ;
        RECT 1266.480 590.930 1266.740 591.250 ;
        RECT 1165.800 20.730 1165.940 590.930 ;
        RECT 1162.520 20.410 1162.780 20.730 ;
        RECT 1165.740 20.410 1166.000 20.730 ;
        RECT 1162.580 2.400 1162.720 20.410 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1015.290 483.040 1015.610 483.100 ;
        RECT 1016.210 483.040 1016.530 483.100 ;
        RECT 1015.290 482.900 1016.530 483.040 ;
        RECT 1015.290 482.840 1015.610 482.900 ;
        RECT 1016.210 482.840 1016.530 482.900 ;
        RECT 1016.210 434.760 1016.530 434.820 ;
        RECT 1017.130 434.760 1017.450 434.820 ;
        RECT 1016.210 434.620 1017.450 434.760 ;
        RECT 1016.210 434.560 1016.530 434.620 ;
        RECT 1017.130 434.560 1017.450 434.620 ;
        RECT 1015.290 386.480 1015.610 386.540 ;
        RECT 1017.130 386.480 1017.450 386.540 ;
        RECT 1015.290 386.340 1017.450 386.480 ;
        RECT 1015.290 386.280 1015.610 386.340 ;
        RECT 1017.130 386.280 1017.450 386.340 ;
        RECT 1015.290 351.600 1015.610 351.860 ;
        RECT 1015.380 351.460 1015.520 351.600 ;
        RECT 1015.750 351.460 1016.070 351.520 ;
        RECT 1015.380 351.320 1016.070 351.460 ;
        RECT 1015.750 351.260 1016.070 351.320 ;
        RECT 1015.290 337.860 1015.610 337.920 ;
        RECT 1015.750 337.860 1016.070 337.920 ;
        RECT 1015.290 337.720 1016.070 337.860 ;
        RECT 1015.290 337.660 1015.610 337.720 ;
        RECT 1015.750 337.660 1016.070 337.720 ;
        RECT 1015.290 289.920 1015.610 289.980 ;
        RECT 1016.210 289.920 1016.530 289.980 ;
        RECT 1015.290 289.780 1016.530 289.920 ;
        RECT 1015.290 289.720 1015.610 289.780 ;
        RECT 1016.210 289.720 1016.530 289.780 ;
        RECT 680.410 43.080 680.730 43.140 ;
        RECT 1015.750 43.080 1016.070 43.140 ;
        RECT 680.410 42.940 1016.070 43.080 ;
        RECT 680.410 42.880 680.730 42.940 ;
        RECT 1015.750 42.880 1016.070 42.940 ;
      LAYER via ;
        RECT 1015.320 482.840 1015.580 483.100 ;
        RECT 1016.240 482.840 1016.500 483.100 ;
        RECT 1016.240 434.560 1016.500 434.820 ;
        RECT 1017.160 434.560 1017.420 434.820 ;
        RECT 1015.320 386.280 1015.580 386.540 ;
        RECT 1017.160 386.280 1017.420 386.540 ;
        RECT 1015.320 351.600 1015.580 351.860 ;
        RECT 1015.780 351.260 1016.040 351.520 ;
        RECT 1015.320 337.660 1015.580 337.920 ;
        RECT 1015.780 337.660 1016.040 337.920 ;
        RECT 1015.320 289.720 1015.580 289.980 ;
        RECT 1016.240 289.720 1016.500 289.980 ;
        RECT 680.440 42.880 680.700 43.140 ;
        RECT 1015.780 42.880 1016.040 43.140 ;
      LAYER met2 ;
        RECT 1020.150 600.170 1020.430 604.000 ;
        RECT 1018.600 600.030 1020.430 600.170 ;
        RECT 1018.600 579.885 1018.740 600.030 ;
        RECT 1020.150 600.000 1020.430 600.030 ;
        RECT 1015.310 579.515 1015.590 579.885 ;
        RECT 1018.530 579.515 1018.810 579.885 ;
        RECT 1015.380 483.130 1015.520 579.515 ;
        RECT 1015.320 482.810 1015.580 483.130 ;
        RECT 1016.240 482.810 1016.500 483.130 ;
        RECT 1016.300 434.850 1016.440 482.810 ;
        RECT 1016.240 434.530 1016.500 434.850 ;
        RECT 1017.160 434.530 1017.420 434.850 ;
        RECT 1017.220 386.570 1017.360 434.530 ;
        RECT 1015.320 386.250 1015.580 386.570 ;
        RECT 1017.160 386.250 1017.420 386.570 ;
        RECT 1015.380 351.890 1015.520 386.250 ;
        RECT 1015.320 351.570 1015.580 351.890 ;
        RECT 1015.780 351.230 1016.040 351.550 ;
        RECT 1015.840 337.950 1015.980 351.230 ;
        RECT 1015.320 337.630 1015.580 337.950 ;
        RECT 1015.780 337.630 1016.040 337.950 ;
        RECT 1015.380 290.010 1015.520 337.630 ;
        RECT 1015.320 289.690 1015.580 290.010 ;
        RECT 1016.240 289.690 1016.500 290.010 ;
        RECT 1016.300 207.130 1016.440 289.690 ;
        RECT 1015.840 206.990 1016.440 207.130 ;
        RECT 1015.840 206.450 1015.980 206.990 ;
        RECT 1015.840 206.310 1016.440 206.450 ;
        RECT 1016.300 110.400 1016.440 206.310 ;
        RECT 1015.840 110.260 1016.440 110.400 ;
        RECT 1015.840 43.170 1015.980 110.260 ;
        RECT 680.440 42.850 680.700 43.170 ;
        RECT 1015.780 42.850 1016.040 43.170 ;
        RECT 680.500 2.400 680.640 42.850 ;
        RECT 680.290 -4.800 680.850 2.400 ;
      LAYER via2 ;
        RECT 1015.310 579.560 1015.590 579.840 ;
        RECT 1018.530 579.560 1018.810 579.840 ;
      LAYER met3 ;
        RECT 1015.285 579.850 1015.615 579.865 ;
        RECT 1018.505 579.850 1018.835 579.865 ;
        RECT 1015.285 579.550 1018.835 579.850 ;
        RECT 1015.285 579.535 1015.615 579.550 ;
        RECT 1018.505 579.535 1018.835 579.550 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 592.520 1186.730 592.580 ;
        RECT 1276.570 592.520 1276.890 592.580 ;
        RECT 1186.410 592.380 1276.890 592.520 ;
        RECT 1186.410 592.320 1186.730 592.380 ;
        RECT 1276.570 592.320 1276.890 592.380 ;
        RECT 1179.970 20.640 1180.290 20.700 ;
        RECT 1186.410 20.640 1186.730 20.700 ;
        RECT 1179.970 20.500 1186.730 20.640 ;
        RECT 1179.970 20.440 1180.290 20.500 ;
        RECT 1186.410 20.440 1186.730 20.500 ;
      LAYER via ;
        RECT 1186.440 592.320 1186.700 592.580 ;
        RECT 1276.600 592.320 1276.860 592.580 ;
        RECT 1180.000 20.440 1180.260 20.700 ;
        RECT 1186.440 20.440 1186.700 20.700 ;
      LAYER met2 ;
        RECT 1277.290 600.170 1277.570 604.000 ;
        RECT 1276.660 600.030 1277.570 600.170 ;
        RECT 1276.660 592.610 1276.800 600.030 ;
        RECT 1277.290 600.000 1277.570 600.030 ;
        RECT 1186.440 592.290 1186.700 592.610 ;
        RECT 1276.600 592.290 1276.860 592.610 ;
        RECT 1186.500 588.610 1186.640 592.290 ;
        RECT 1186.500 588.470 1187.100 588.610 ;
        RECT 1186.960 585.890 1187.100 588.470 ;
        RECT 1186.500 585.750 1187.100 585.890 ;
        RECT 1186.500 20.730 1186.640 585.750 ;
        RECT 1180.000 20.410 1180.260 20.730 ;
        RECT 1186.440 20.410 1186.700 20.730 ;
        RECT 1180.060 2.400 1180.200 20.410 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 592.860 1200.530 592.920 ;
        RECT 1284.850 592.860 1285.170 592.920 ;
        RECT 1200.210 592.720 1285.170 592.860 ;
        RECT 1200.210 592.660 1200.530 592.720 ;
        RECT 1284.850 592.660 1285.170 592.720 ;
        RECT 1197.910 20.640 1198.230 20.700 ;
        RECT 1200.210 20.640 1200.530 20.700 ;
        RECT 1197.910 20.500 1200.530 20.640 ;
        RECT 1197.910 20.440 1198.230 20.500 ;
        RECT 1200.210 20.440 1200.530 20.500 ;
      LAYER via ;
        RECT 1200.240 592.660 1200.500 592.920 ;
        RECT 1284.880 592.660 1285.140 592.920 ;
        RECT 1197.940 20.440 1198.200 20.700 ;
        RECT 1200.240 20.440 1200.500 20.700 ;
      LAYER met2 ;
        RECT 1286.490 600.170 1286.770 604.000 ;
        RECT 1284.940 600.030 1286.770 600.170 ;
        RECT 1284.940 592.950 1285.080 600.030 ;
        RECT 1286.490 600.000 1286.770 600.030 ;
        RECT 1200.240 592.630 1200.500 592.950 ;
        RECT 1284.880 592.630 1285.140 592.950 ;
        RECT 1200.300 20.730 1200.440 592.630 ;
        RECT 1197.940 20.410 1198.200 20.730 ;
        RECT 1200.240 20.410 1200.500 20.730 ;
        RECT 1198.000 2.400 1198.140 20.410 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 588.100 1221.230 588.160 ;
        RECT 1294.050 588.100 1294.370 588.160 ;
        RECT 1220.910 587.960 1294.370 588.100 ;
        RECT 1220.910 587.900 1221.230 587.960 ;
        RECT 1294.050 587.900 1294.370 587.960 ;
        RECT 1215.850 20.640 1216.170 20.700 ;
        RECT 1220.910 20.640 1221.230 20.700 ;
        RECT 1215.850 20.500 1221.230 20.640 ;
        RECT 1215.850 20.440 1216.170 20.500 ;
        RECT 1220.910 20.440 1221.230 20.500 ;
      LAYER via ;
        RECT 1220.940 587.900 1221.200 588.160 ;
        RECT 1294.080 587.900 1294.340 588.160 ;
        RECT 1215.880 20.440 1216.140 20.700 ;
        RECT 1220.940 20.440 1221.200 20.700 ;
      LAYER met2 ;
        RECT 1295.690 600.170 1295.970 604.000 ;
        RECT 1294.140 600.030 1295.970 600.170 ;
        RECT 1294.140 588.190 1294.280 600.030 ;
        RECT 1295.690 600.000 1295.970 600.030 ;
        RECT 1220.940 587.870 1221.200 588.190 ;
        RECT 1294.080 587.870 1294.340 588.190 ;
        RECT 1221.000 20.730 1221.140 587.870 ;
        RECT 1215.880 20.410 1216.140 20.730 ;
        RECT 1220.940 20.410 1221.200 20.730 ;
        RECT 1215.940 2.400 1216.080 20.410 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.710 588.780 1235.030 588.840 ;
        RECT 1304.170 588.780 1304.490 588.840 ;
        RECT 1234.710 588.640 1304.490 588.780 ;
        RECT 1234.710 588.580 1235.030 588.640 ;
        RECT 1304.170 588.580 1304.490 588.640 ;
        RECT 1233.790 47.980 1234.110 48.240 ;
        RECT 1233.880 47.560 1234.020 47.980 ;
        RECT 1233.790 47.300 1234.110 47.560 ;
      LAYER via ;
        RECT 1234.740 588.580 1235.000 588.840 ;
        RECT 1304.200 588.580 1304.460 588.840 ;
        RECT 1233.820 47.980 1234.080 48.240 ;
        RECT 1233.820 47.300 1234.080 47.560 ;
      LAYER met2 ;
        RECT 1304.890 600.170 1305.170 604.000 ;
        RECT 1304.260 600.030 1305.170 600.170 ;
        RECT 1304.260 588.870 1304.400 600.030 ;
        RECT 1304.890 600.000 1305.170 600.030 ;
        RECT 1234.740 588.550 1235.000 588.870 ;
        RECT 1304.200 588.550 1304.460 588.870 ;
        RECT 1234.800 532.285 1234.940 588.550 ;
        RECT 1234.730 531.915 1235.010 532.285 ;
        RECT 1234.730 531.235 1235.010 531.605 ;
        RECT 1234.800 49.485 1234.940 531.235 ;
        RECT 1234.730 49.115 1235.010 49.485 ;
        RECT 1233.810 48.435 1234.090 48.805 ;
        RECT 1233.880 48.270 1234.020 48.435 ;
        RECT 1233.820 47.950 1234.080 48.270 ;
        RECT 1233.820 47.270 1234.080 47.590 ;
        RECT 1233.880 2.400 1234.020 47.270 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
      LAYER via2 ;
        RECT 1234.730 531.960 1235.010 532.240 ;
        RECT 1234.730 531.280 1235.010 531.560 ;
        RECT 1234.730 49.160 1235.010 49.440 ;
        RECT 1233.810 48.480 1234.090 48.760 ;
      LAYER met3 ;
        RECT 1234.705 532.250 1235.035 532.265 ;
        RECT 1234.705 531.935 1235.250 532.250 ;
        RECT 1234.950 531.585 1235.250 531.935 ;
        RECT 1234.705 531.270 1235.250 531.585 ;
        RECT 1234.705 531.255 1235.035 531.270 ;
        RECT 1234.705 49.450 1235.035 49.465 ;
        RECT 1233.110 49.150 1235.035 49.450 ;
        RECT 1233.110 48.770 1233.410 49.150 ;
        RECT 1234.705 49.135 1235.035 49.150 ;
        RECT 1233.785 48.770 1234.115 48.785 ;
        RECT 1233.110 48.470 1234.115 48.770 ;
        RECT 1233.785 48.455 1234.115 48.470 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 589.800 1255.730 589.860 ;
        RECT 1312.450 589.800 1312.770 589.860 ;
        RECT 1255.410 589.660 1312.770 589.800 ;
        RECT 1255.410 589.600 1255.730 589.660 ;
        RECT 1312.450 589.600 1312.770 589.660 ;
        RECT 1251.730 16.900 1252.050 16.960 ;
        RECT 1255.410 16.900 1255.730 16.960 ;
        RECT 1251.730 16.760 1255.730 16.900 ;
        RECT 1251.730 16.700 1252.050 16.760 ;
        RECT 1255.410 16.700 1255.730 16.760 ;
      LAYER via ;
        RECT 1255.440 589.600 1255.700 589.860 ;
        RECT 1312.480 589.600 1312.740 589.860 ;
        RECT 1251.760 16.700 1252.020 16.960 ;
        RECT 1255.440 16.700 1255.700 16.960 ;
      LAYER met2 ;
        RECT 1314.090 600.170 1314.370 604.000 ;
        RECT 1312.540 600.030 1314.370 600.170 ;
        RECT 1312.540 589.890 1312.680 600.030 ;
        RECT 1314.090 600.000 1314.370 600.030 ;
        RECT 1255.440 589.570 1255.700 589.890 ;
        RECT 1312.480 589.570 1312.740 589.890 ;
        RECT 1255.500 16.990 1255.640 589.570 ;
        RECT 1251.760 16.670 1252.020 16.990 ;
        RECT 1255.440 16.670 1255.700 16.990 ;
        RECT 1251.820 2.400 1251.960 16.670 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1268.750 590.140 1269.070 590.200 ;
        RECT 1321.650 590.140 1321.970 590.200 ;
        RECT 1268.750 590.000 1321.970 590.140 ;
        RECT 1268.750 589.940 1269.070 590.000 ;
        RECT 1321.650 589.940 1321.970 590.000 ;
        RECT 1268.750 579.600 1269.070 579.660 ;
        RECT 1269.670 579.600 1269.990 579.660 ;
        RECT 1268.750 579.460 1269.990 579.600 ;
        RECT 1268.750 579.400 1269.070 579.460 ;
        RECT 1269.670 579.400 1269.990 579.460 ;
        RECT 1268.750 531.660 1269.070 531.720 ;
        RECT 1269.670 531.660 1269.990 531.720 ;
        RECT 1268.750 531.520 1269.990 531.660 ;
        RECT 1268.750 531.460 1269.070 531.520 ;
        RECT 1269.670 531.460 1269.990 531.520 ;
        RECT 1267.830 524.180 1268.150 524.240 ;
        RECT 1268.750 524.180 1269.070 524.240 ;
        RECT 1267.830 524.040 1269.070 524.180 ;
        RECT 1267.830 523.980 1268.150 524.040 ;
        RECT 1268.750 523.980 1269.070 524.040 ;
        RECT 1267.830 476.240 1268.150 476.300 ;
        RECT 1268.750 476.240 1269.070 476.300 ;
        RECT 1267.830 476.100 1269.070 476.240 ;
        RECT 1267.830 476.040 1268.150 476.100 ;
        RECT 1268.750 476.040 1269.070 476.100 ;
        RECT 1267.830 427.620 1268.150 427.680 ;
        RECT 1268.750 427.620 1269.070 427.680 ;
        RECT 1267.830 427.480 1269.070 427.620 ;
        RECT 1267.830 427.420 1268.150 427.480 ;
        RECT 1268.750 427.420 1269.070 427.480 ;
        RECT 1267.830 379.680 1268.150 379.740 ;
        RECT 1268.750 379.680 1269.070 379.740 ;
        RECT 1267.830 379.540 1269.070 379.680 ;
        RECT 1267.830 379.480 1268.150 379.540 ;
        RECT 1268.750 379.480 1269.070 379.540 ;
        RECT 1268.290 283.120 1268.610 283.180 ;
        RECT 1268.750 283.120 1269.070 283.180 ;
        RECT 1268.290 282.980 1269.070 283.120 ;
        RECT 1268.290 282.920 1268.610 282.980 ;
        RECT 1268.750 282.920 1269.070 282.980 ;
        RECT 1268.290 241.980 1268.610 242.040 ;
        RECT 1268.750 241.980 1269.070 242.040 ;
        RECT 1268.290 241.840 1269.070 241.980 ;
        RECT 1268.290 241.780 1268.610 241.840 ;
        RECT 1268.750 241.780 1269.070 241.840 ;
        RECT 1267.370 234.500 1267.690 234.560 ;
        RECT 1268.750 234.500 1269.070 234.560 ;
        RECT 1267.370 234.360 1269.070 234.500 ;
        RECT 1267.370 234.300 1267.690 234.360 ;
        RECT 1268.750 234.300 1269.070 234.360 ;
        RECT 1267.370 186.560 1267.690 186.620 ;
        RECT 1267.830 186.560 1268.150 186.620 ;
        RECT 1267.370 186.420 1268.150 186.560 ;
        RECT 1267.370 186.360 1267.690 186.420 ;
        RECT 1267.830 186.360 1268.150 186.420 ;
        RECT 1267.830 145.420 1268.150 145.480 ;
        RECT 1268.750 145.420 1269.070 145.480 ;
        RECT 1267.830 145.280 1269.070 145.420 ;
        RECT 1267.830 145.220 1268.150 145.280 ;
        RECT 1268.750 145.220 1269.070 145.280 ;
        RECT 1267.830 137.940 1268.150 138.000 ;
        RECT 1268.750 137.940 1269.070 138.000 ;
        RECT 1267.830 137.800 1269.070 137.940 ;
        RECT 1267.830 137.740 1268.150 137.800 ;
        RECT 1268.750 137.740 1269.070 137.800 ;
        RECT 1267.370 90.000 1267.690 90.060 ;
        RECT 1267.830 90.000 1268.150 90.060 ;
        RECT 1267.370 89.860 1268.150 90.000 ;
        RECT 1267.370 89.800 1267.690 89.860 ;
        RECT 1267.830 89.800 1268.150 89.860 ;
        RECT 1267.370 48.520 1267.690 48.580 ;
        RECT 1268.290 48.520 1268.610 48.580 ;
        RECT 1267.370 48.380 1268.610 48.520 ;
        RECT 1267.370 48.320 1267.690 48.380 ;
        RECT 1268.290 48.320 1268.610 48.380 ;
        RECT 1268.290 20.300 1268.610 20.360 ;
        RECT 1268.290 20.160 1269.440 20.300 ;
        RECT 1268.290 20.100 1268.610 20.160 ;
        RECT 1269.300 20.020 1269.440 20.160 ;
        RECT 1269.210 19.760 1269.530 20.020 ;
      LAYER via ;
        RECT 1268.780 589.940 1269.040 590.200 ;
        RECT 1321.680 589.940 1321.940 590.200 ;
        RECT 1268.780 579.400 1269.040 579.660 ;
        RECT 1269.700 579.400 1269.960 579.660 ;
        RECT 1268.780 531.460 1269.040 531.720 ;
        RECT 1269.700 531.460 1269.960 531.720 ;
        RECT 1267.860 523.980 1268.120 524.240 ;
        RECT 1268.780 523.980 1269.040 524.240 ;
        RECT 1267.860 476.040 1268.120 476.300 ;
        RECT 1268.780 476.040 1269.040 476.300 ;
        RECT 1267.860 427.420 1268.120 427.680 ;
        RECT 1268.780 427.420 1269.040 427.680 ;
        RECT 1267.860 379.480 1268.120 379.740 ;
        RECT 1268.780 379.480 1269.040 379.740 ;
        RECT 1268.320 282.920 1268.580 283.180 ;
        RECT 1268.780 282.920 1269.040 283.180 ;
        RECT 1268.320 241.780 1268.580 242.040 ;
        RECT 1268.780 241.780 1269.040 242.040 ;
        RECT 1267.400 234.300 1267.660 234.560 ;
        RECT 1268.780 234.300 1269.040 234.560 ;
        RECT 1267.400 186.360 1267.660 186.620 ;
        RECT 1267.860 186.360 1268.120 186.620 ;
        RECT 1267.860 145.220 1268.120 145.480 ;
        RECT 1268.780 145.220 1269.040 145.480 ;
        RECT 1267.860 137.740 1268.120 138.000 ;
        RECT 1268.780 137.740 1269.040 138.000 ;
        RECT 1267.400 89.800 1267.660 90.060 ;
        RECT 1267.860 89.800 1268.120 90.060 ;
        RECT 1267.400 48.320 1267.660 48.580 ;
        RECT 1268.320 48.320 1268.580 48.580 ;
        RECT 1268.320 20.100 1268.580 20.360 ;
        RECT 1269.240 19.760 1269.500 20.020 ;
      LAYER met2 ;
        RECT 1323.290 600.170 1323.570 604.000 ;
        RECT 1321.740 600.030 1323.570 600.170 ;
        RECT 1321.740 590.230 1321.880 600.030 ;
        RECT 1323.290 600.000 1323.570 600.030 ;
        RECT 1268.780 589.910 1269.040 590.230 ;
        RECT 1321.680 589.910 1321.940 590.230 ;
        RECT 1268.840 579.690 1268.980 589.910 ;
        RECT 1268.780 579.370 1269.040 579.690 ;
        RECT 1269.700 579.370 1269.960 579.690 ;
        RECT 1269.760 531.750 1269.900 579.370 ;
        RECT 1268.780 531.430 1269.040 531.750 ;
        RECT 1269.700 531.430 1269.960 531.750 ;
        RECT 1268.840 524.270 1268.980 531.430 ;
        RECT 1267.860 523.950 1268.120 524.270 ;
        RECT 1268.780 523.950 1269.040 524.270 ;
        RECT 1267.920 476.330 1268.060 523.950 ;
        RECT 1267.860 476.010 1268.120 476.330 ;
        RECT 1268.780 476.010 1269.040 476.330 ;
        RECT 1268.840 427.710 1268.980 476.010 ;
        RECT 1267.860 427.390 1268.120 427.710 ;
        RECT 1268.780 427.390 1269.040 427.710 ;
        RECT 1267.920 379.770 1268.060 427.390 ;
        RECT 1267.860 379.450 1268.120 379.770 ;
        RECT 1268.780 379.450 1269.040 379.770 ;
        RECT 1268.840 283.210 1268.980 379.450 ;
        RECT 1268.320 282.890 1268.580 283.210 ;
        RECT 1268.780 282.890 1269.040 283.210 ;
        RECT 1268.380 242.070 1268.520 282.890 ;
        RECT 1268.320 241.750 1268.580 242.070 ;
        RECT 1268.780 241.750 1269.040 242.070 ;
        RECT 1268.840 234.590 1268.980 241.750 ;
        RECT 1267.400 234.270 1267.660 234.590 ;
        RECT 1268.780 234.270 1269.040 234.590 ;
        RECT 1267.460 186.650 1267.600 234.270 ;
        RECT 1267.400 186.330 1267.660 186.650 ;
        RECT 1267.860 186.330 1268.120 186.650 ;
        RECT 1267.920 145.510 1268.060 186.330 ;
        RECT 1267.860 145.190 1268.120 145.510 ;
        RECT 1268.780 145.190 1269.040 145.510 ;
        RECT 1268.840 138.030 1268.980 145.190 ;
        RECT 1267.860 137.710 1268.120 138.030 ;
        RECT 1268.780 137.710 1269.040 138.030 ;
        RECT 1267.920 90.090 1268.060 137.710 ;
        RECT 1267.400 89.770 1267.660 90.090 ;
        RECT 1267.860 89.770 1268.120 90.090 ;
        RECT 1267.460 48.610 1267.600 89.770 ;
        RECT 1267.400 48.290 1267.660 48.610 ;
        RECT 1268.320 48.290 1268.580 48.610 ;
        RECT 1268.380 20.390 1268.520 48.290 ;
        RECT 1268.320 20.070 1268.580 20.390 ;
        RECT 1269.240 19.730 1269.500 20.050 ;
        RECT 1269.300 2.400 1269.440 19.730 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 590.820 1290.230 590.880 ;
        RECT 1331.770 590.820 1332.090 590.880 ;
        RECT 1289.910 590.680 1332.090 590.820 ;
        RECT 1289.910 590.620 1290.230 590.680 ;
        RECT 1331.770 590.620 1332.090 590.680 ;
        RECT 1287.150 17.580 1287.470 17.640 ;
        RECT 1289.910 17.580 1290.230 17.640 ;
        RECT 1287.150 17.440 1290.230 17.580 ;
        RECT 1287.150 17.380 1287.470 17.440 ;
        RECT 1289.910 17.380 1290.230 17.440 ;
      LAYER via ;
        RECT 1289.940 590.620 1290.200 590.880 ;
        RECT 1331.800 590.620 1332.060 590.880 ;
        RECT 1287.180 17.380 1287.440 17.640 ;
        RECT 1289.940 17.380 1290.200 17.640 ;
      LAYER met2 ;
        RECT 1332.490 600.170 1332.770 604.000 ;
        RECT 1331.860 600.030 1332.770 600.170 ;
        RECT 1331.860 590.910 1332.000 600.030 ;
        RECT 1332.490 600.000 1332.770 600.030 ;
        RECT 1289.940 590.590 1290.200 590.910 ;
        RECT 1331.800 590.590 1332.060 590.910 ;
        RECT 1290.000 17.670 1290.140 590.590 ;
        RECT 1287.180 17.350 1287.440 17.670 ;
        RECT 1289.940 17.350 1290.200 17.670 ;
        RECT 1287.240 2.400 1287.380 17.350 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 588.780 1310.930 588.840 ;
        RECT 1340.050 588.780 1340.370 588.840 ;
        RECT 1310.610 588.640 1340.370 588.780 ;
        RECT 1310.610 588.580 1310.930 588.640 ;
        RECT 1340.050 588.580 1340.370 588.640 ;
        RECT 1305.090 16.220 1305.410 16.280 ;
        RECT 1310.610 16.220 1310.930 16.280 ;
        RECT 1305.090 16.080 1310.930 16.220 ;
        RECT 1305.090 16.020 1305.410 16.080 ;
        RECT 1310.610 16.020 1310.930 16.080 ;
      LAYER via ;
        RECT 1310.640 588.580 1310.900 588.840 ;
        RECT 1340.080 588.580 1340.340 588.840 ;
        RECT 1305.120 16.020 1305.380 16.280 ;
        RECT 1310.640 16.020 1310.900 16.280 ;
      LAYER met2 ;
        RECT 1341.690 600.170 1341.970 604.000 ;
        RECT 1340.140 600.030 1341.970 600.170 ;
        RECT 1340.140 588.870 1340.280 600.030 ;
        RECT 1341.690 600.000 1341.970 600.030 ;
        RECT 1310.640 588.550 1310.900 588.870 ;
        RECT 1340.080 588.550 1340.340 588.870 ;
        RECT 1310.700 16.310 1310.840 588.550 ;
        RECT 1305.120 15.990 1305.380 16.310 ;
        RECT 1310.640 15.990 1310.900 16.310 ;
        RECT 1305.180 2.400 1305.320 15.990 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.410 589.800 1324.730 589.860 ;
        RECT 1349.250 589.800 1349.570 589.860 ;
        RECT 1324.410 589.660 1349.570 589.800 ;
        RECT 1324.410 589.600 1324.730 589.660 ;
        RECT 1349.250 589.600 1349.570 589.660 ;
      LAYER via ;
        RECT 1324.440 589.600 1324.700 589.860 ;
        RECT 1349.280 589.600 1349.540 589.860 ;
      LAYER met2 ;
        RECT 1350.890 600.170 1351.170 604.000 ;
        RECT 1349.340 600.030 1351.170 600.170 ;
        RECT 1349.340 589.890 1349.480 600.030 ;
        RECT 1350.890 600.000 1351.170 600.030 ;
        RECT 1324.440 589.570 1324.700 589.890 ;
        RECT 1349.280 589.570 1349.540 589.890 ;
        RECT 1324.500 17.410 1324.640 589.570 ;
        RECT 1323.120 17.270 1324.640 17.410 ;
        RECT 1323.120 2.400 1323.260 17.270 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1345.110 587.080 1345.430 587.140 ;
        RECT 1359.370 587.080 1359.690 587.140 ;
        RECT 1345.110 586.940 1359.690 587.080 ;
        RECT 1345.110 586.880 1345.430 586.940 ;
        RECT 1359.370 586.880 1359.690 586.940 ;
        RECT 1340.510 17.580 1340.830 17.640 ;
        RECT 1345.110 17.580 1345.430 17.640 ;
        RECT 1340.510 17.440 1345.430 17.580 ;
        RECT 1340.510 17.380 1340.830 17.440 ;
        RECT 1345.110 17.380 1345.430 17.440 ;
      LAYER via ;
        RECT 1345.140 586.880 1345.400 587.140 ;
        RECT 1359.400 586.880 1359.660 587.140 ;
        RECT 1340.540 17.380 1340.800 17.640 ;
        RECT 1345.140 17.380 1345.400 17.640 ;
      LAYER met2 ;
        RECT 1360.090 600.170 1360.370 604.000 ;
        RECT 1359.460 600.030 1360.370 600.170 ;
        RECT 1359.460 587.170 1359.600 600.030 ;
        RECT 1360.090 600.000 1360.370 600.030 ;
        RECT 1345.140 586.850 1345.400 587.170 ;
        RECT 1359.400 586.850 1359.660 587.170 ;
        RECT 1345.200 17.670 1345.340 586.850 ;
        RECT 1340.540 17.350 1340.800 17.670 ;
        RECT 1345.140 17.350 1345.400 17.670 ;
        RECT 1340.600 2.400 1340.740 17.350 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 698.350 45.120 698.670 45.180 ;
        RECT 1028.630 45.120 1028.950 45.180 ;
        RECT 698.350 44.980 1028.950 45.120 ;
        RECT 698.350 44.920 698.670 44.980 ;
        RECT 1028.630 44.920 1028.950 44.980 ;
      LAYER via ;
        RECT 698.380 44.920 698.640 45.180 ;
        RECT 1028.660 44.920 1028.920 45.180 ;
      LAYER met2 ;
        RECT 1029.350 600.170 1029.630 604.000 ;
        RECT 1028.720 600.030 1029.630 600.170 ;
        RECT 1028.720 45.210 1028.860 600.030 ;
        RECT 1029.350 600.000 1029.630 600.030 ;
        RECT 698.380 44.890 698.640 45.210 ;
        RECT 1028.660 44.890 1028.920 45.210 ;
        RECT 698.440 2.400 698.580 44.890 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1362.590 587.080 1362.910 587.140 ;
        RECT 1367.650 587.080 1367.970 587.140 ;
        RECT 1362.590 586.940 1367.970 587.080 ;
        RECT 1362.590 586.880 1362.910 586.940 ;
        RECT 1367.650 586.880 1367.970 586.940 ;
        RECT 1358.450 17.580 1358.770 17.640 ;
        RECT 1362.590 17.580 1362.910 17.640 ;
        RECT 1358.450 17.440 1362.910 17.580 ;
        RECT 1358.450 17.380 1358.770 17.440 ;
        RECT 1362.590 17.380 1362.910 17.440 ;
      LAYER via ;
        RECT 1362.620 586.880 1362.880 587.140 ;
        RECT 1367.680 586.880 1367.940 587.140 ;
        RECT 1358.480 17.380 1358.740 17.640 ;
        RECT 1362.620 17.380 1362.880 17.640 ;
      LAYER met2 ;
        RECT 1369.290 600.170 1369.570 604.000 ;
        RECT 1367.740 600.030 1369.570 600.170 ;
        RECT 1367.740 587.170 1367.880 600.030 ;
        RECT 1369.290 600.000 1369.570 600.030 ;
        RECT 1362.620 586.850 1362.880 587.170 ;
        RECT 1367.680 586.850 1367.940 587.170 ;
        RECT 1362.680 17.670 1362.820 586.850 ;
        RECT 1358.480 17.350 1358.740 17.670 ;
        RECT 1362.620 17.350 1362.880 17.670 ;
        RECT 1358.540 2.400 1358.680 17.350 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1372.250 483.040 1372.570 483.100 ;
        RECT 1373.630 483.040 1373.950 483.100 ;
        RECT 1372.250 482.900 1373.950 483.040 ;
        RECT 1372.250 482.840 1372.570 482.900 ;
        RECT 1373.630 482.840 1373.950 482.900 ;
        RECT 1373.170 434.760 1373.490 434.820 ;
        RECT 1374.090 434.760 1374.410 434.820 ;
        RECT 1373.170 434.620 1374.410 434.760 ;
        RECT 1373.170 434.560 1373.490 434.620 ;
        RECT 1374.090 434.560 1374.410 434.620 ;
        RECT 1373.630 362.340 1373.950 362.400 ;
        RECT 1375.470 362.340 1375.790 362.400 ;
        RECT 1373.630 362.200 1375.790 362.340 ;
        RECT 1373.630 362.140 1373.950 362.200 ;
        RECT 1375.470 362.140 1375.790 362.200 ;
        RECT 1374.550 338.200 1374.870 338.260 ;
        RECT 1375.470 338.200 1375.790 338.260 ;
        RECT 1374.550 338.060 1375.790 338.200 ;
        RECT 1374.550 338.000 1374.870 338.060 ;
        RECT 1375.470 338.000 1375.790 338.060 ;
        RECT 1373.630 265.780 1373.950 265.840 ;
        RECT 1375.470 265.780 1375.790 265.840 ;
        RECT 1373.630 265.640 1375.790 265.780 ;
        RECT 1373.630 265.580 1373.950 265.640 ;
        RECT 1375.470 265.580 1375.790 265.640 ;
        RECT 1374.550 241.640 1374.870 241.700 ;
        RECT 1375.470 241.640 1375.790 241.700 ;
        RECT 1374.550 241.500 1375.790 241.640 ;
        RECT 1374.550 241.440 1374.870 241.500 ;
        RECT 1375.470 241.440 1375.790 241.500 ;
        RECT 1373.630 193.020 1373.950 193.080 ;
        RECT 1375.470 193.020 1375.790 193.080 ;
        RECT 1373.630 192.880 1375.790 193.020 ;
        RECT 1373.630 192.820 1373.950 192.880 ;
        RECT 1375.470 192.820 1375.790 192.880 ;
        RECT 1374.550 145.080 1374.870 145.140 ;
        RECT 1375.470 145.080 1375.790 145.140 ;
        RECT 1374.550 144.940 1375.790 145.080 ;
        RECT 1374.550 144.880 1374.870 144.940 ;
        RECT 1375.470 144.880 1375.790 144.940 ;
        RECT 1375.010 48.520 1375.330 48.580 ;
        RECT 1376.390 48.520 1376.710 48.580 ;
        RECT 1375.010 48.380 1376.710 48.520 ;
        RECT 1375.010 48.320 1375.330 48.380 ;
        RECT 1376.390 48.320 1376.710 48.380 ;
        RECT 1376.390 2.960 1376.710 3.020 ;
        RECT 1376.850 2.960 1377.170 3.020 ;
        RECT 1376.390 2.820 1377.170 2.960 ;
        RECT 1376.390 2.760 1376.710 2.820 ;
        RECT 1376.850 2.760 1377.170 2.820 ;
      LAYER via ;
        RECT 1372.280 482.840 1372.540 483.100 ;
        RECT 1373.660 482.840 1373.920 483.100 ;
        RECT 1373.200 434.560 1373.460 434.820 ;
        RECT 1374.120 434.560 1374.380 434.820 ;
        RECT 1373.660 362.140 1373.920 362.400 ;
        RECT 1375.500 362.140 1375.760 362.400 ;
        RECT 1374.580 338.000 1374.840 338.260 ;
        RECT 1375.500 338.000 1375.760 338.260 ;
        RECT 1373.660 265.580 1373.920 265.840 ;
        RECT 1375.500 265.580 1375.760 265.840 ;
        RECT 1374.580 241.440 1374.840 241.700 ;
        RECT 1375.500 241.440 1375.760 241.700 ;
        RECT 1373.660 192.820 1373.920 193.080 ;
        RECT 1375.500 192.820 1375.760 193.080 ;
        RECT 1374.580 144.880 1374.840 145.140 ;
        RECT 1375.500 144.880 1375.760 145.140 ;
        RECT 1375.040 48.320 1375.300 48.580 ;
        RECT 1376.420 48.320 1376.680 48.580 ;
        RECT 1376.420 2.760 1376.680 3.020 ;
        RECT 1376.880 2.760 1377.140 3.020 ;
      LAYER met2 ;
        RECT 1378.490 600.850 1378.770 604.000 ;
        RECT 1376.020 600.710 1378.770 600.850 ;
        RECT 1376.020 545.770 1376.160 600.710 ;
        RECT 1378.490 600.000 1378.770 600.710 ;
        RECT 1374.640 545.630 1376.160 545.770 ;
        RECT 1374.640 545.090 1374.780 545.630 ;
        RECT 1374.180 544.950 1374.780 545.090 ;
        RECT 1374.180 497.490 1374.320 544.950 ;
        RECT 1374.180 497.350 1374.780 497.490 ;
        RECT 1374.640 484.005 1374.780 497.350 ;
        RECT 1374.570 483.635 1374.850 484.005 ;
        RECT 1372.280 482.810 1372.540 483.130 ;
        RECT 1373.650 482.955 1373.930 483.325 ;
        RECT 1373.660 482.810 1373.920 482.955 ;
        RECT 1372.340 435.045 1372.480 482.810 ;
        RECT 1372.270 434.675 1372.550 435.045 ;
        RECT 1373.190 434.675 1373.470 435.045 ;
        RECT 1373.200 434.530 1373.460 434.675 ;
        RECT 1374.120 434.530 1374.380 434.850 ;
        RECT 1374.180 399.570 1374.320 434.530 ;
        RECT 1373.720 399.430 1374.320 399.570 ;
        RECT 1373.720 362.430 1373.860 399.430 ;
        RECT 1373.660 362.110 1373.920 362.430 ;
        RECT 1375.500 362.110 1375.760 362.430 ;
        RECT 1375.560 338.290 1375.700 362.110 ;
        RECT 1374.580 337.970 1374.840 338.290 ;
        RECT 1375.500 337.970 1375.760 338.290 ;
        RECT 1374.640 303.690 1374.780 337.970 ;
        RECT 1373.720 303.550 1374.780 303.690 ;
        RECT 1373.720 265.870 1373.860 303.550 ;
        RECT 1373.660 265.550 1373.920 265.870 ;
        RECT 1375.500 265.550 1375.760 265.870 ;
        RECT 1375.560 241.730 1375.700 265.550 ;
        RECT 1374.580 241.410 1374.840 241.730 ;
        RECT 1375.500 241.410 1375.760 241.730 ;
        RECT 1374.640 207.130 1374.780 241.410 ;
        RECT 1373.720 206.990 1374.780 207.130 ;
        RECT 1373.720 193.110 1373.860 206.990 ;
        RECT 1373.660 192.790 1373.920 193.110 ;
        RECT 1375.500 192.790 1375.760 193.110 ;
        RECT 1375.560 145.170 1375.700 192.790 ;
        RECT 1374.580 144.850 1374.840 145.170 ;
        RECT 1375.500 144.850 1375.760 145.170 ;
        RECT 1374.640 110.570 1374.780 144.850 ;
        RECT 1373.720 110.430 1374.780 110.570 ;
        RECT 1373.720 73.170 1373.860 110.430 ;
        RECT 1373.720 73.030 1375.240 73.170 ;
        RECT 1375.100 48.610 1375.240 73.030 ;
        RECT 1375.040 48.290 1375.300 48.610 ;
        RECT 1376.420 48.290 1376.680 48.610 ;
        RECT 1376.480 48.010 1376.620 48.290 ;
        RECT 1376.480 47.870 1377.080 48.010 ;
        RECT 1376.940 3.050 1377.080 47.870 ;
        RECT 1376.420 2.730 1376.680 3.050 ;
        RECT 1376.880 2.730 1377.140 3.050 ;
        RECT 1376.480 2.400 1376.620 2.730 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
      LAYER via2 ;
        RECT 1374.570 483.680 1374.850 483.960 ;
        RECT 1373.650 483.000 1373.930 483.280 ;
        RECT 1372.270 434.720 1372.550 435.000 ;
        RECT 1373.190 434.720 1373.470 435.000 ;
      LAYER met3 ;
        RECT 1374.545 483.970 1374.875 483.985 ;
        RECT 1373.870 483.670 1374.875 483.970 ;
        RECT 1373.870 483.305 1374.170 483.670 ;
        RECT 1374.545 483.655 1374.875 483.670 ;
        RECT 1373.625 482.990 1374.170 483.305 ;
        RECT 1373.625 482.975 1373.955 482.990 ;
        RECT 1372.245 435.010 1372.575 435.025 ;
        RECT 1373.165 435.010 1373.495 435.025 ;
        RECT 1372.245 434.710 1373.495 435.010 ;
        RECT 1372.245 434.695 1372.575 434.710 ;
        RECT 1373.165 434.695 1373.495 434.710 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1389.270 588.780 1389.590 588.840 ;
        RECT 1393.410 588.780 1393.730 588.840 ;
        RECT 1389.270 588.640 1393.730 588.780 ;
        RECT 1389.270 588.580 1389.590 588.640 ;
        RECT 1393.410 588.580 1393.730 588.640 ;
      LAYER via ;
        RECT 1389.300 588.580 1389.560 588.840 ;
        RECT 1393.440 588.580 1393.700 588.840 ;
      LAYER met2 ;
        RECT 1387.690 600.170 1387.970 604.000 ;
        RECT 1387.690 600.030 1389.500 600.170 ;
        RECT 1387.690 600.000 1387.970 600.030 ;
        RECT 1389.360 588.870 1389.500 600.030 ;
        RECT 1389.300 588.550 1389.560 588.870 ;
        RECT 1393.440 588.550 1393.700 588.870 ;
        RECT 1393.500 20.810 1393.640 588.550 ;
        RECT 1393.500 20.670 1394.560 20.810 ;
        RECT 1394.420 2.400 1394.560 20.670 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1398.470 586.740 1398.790 586.800 ;
        RECT 1400.310 586.740 1400.630 586.800 ;
        RECT 1398.470 586.600 1400.630 586.740 ;
        RECT 1398.470 586.540 1398.790 586.600 ;
        RECT 1400.310 586.540 1400.630 586.600 ;
        RECT 1399.850 20.300 1400.170 20.360 ;
        RECT 1412.270 20.300 1412.590 20.360 ;
        RECT 1399.850 20.160 1412.590 20.300 ;
        RECT 1399.850 20.100 1400.170 20.160 ;
        RECT 1412.270 20.100 1412.590 20.160 ;
      LAYER via ;
        RECT 1398.500 586.540 1398.760 586.800 ;
        RECT 1400.340 586.540 1400.600 586.800 ;
        RECT 1399.880 20.100 1400.140 20.360 ;
        RECT 1412.300 20.100 1412.560 20.360 ;
      LAYER met2 ;
        RECT 1396.890 600.170 1397.170 604.000 ;
        RECT 1396.890 600.030 1398.700 600.170 ;
        RECT 1396.890 600.000 1397.170 600.030 ;
        RECT 1398.560 586.830 1398.700 600.030 ;
        RECT 1398.500 586.510 1398.760 586.830 ;
        RECT 1400.340 586.510 1400.600 586.830 ;
        RECT 1400.400 56.170 1400.540 586.510 ;
        RECT 1399.940 56.030 1400.540 56.170 ;
        RECT 1399.940 20.390 1400.080 56.030 ;
        RECT 1399.880 20.070 1400.140 20.390 ;
        RECT 1412.300 20.070 1412.560 20.390 ;
        RECT 1412.360 2.400 1412.500 20.070 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1406.750 15.880 1407.070 15.940 ;
        RECT 1429.750 15.880 1430.070 15.940 ;
        RECT 1406.750 15.740 1430.070 15.880 ;
        RECT 1406.750 15.680 1407.070 15.740 ;
        RECT 1429.750 15.680 1430.070 15.740 ;
      LAYER via ;
        RECT 1406.780 15.680 1407.040 15.940 ;
        RECT 1429.780 15.680 1430.040 15.940 ;
      LAYER met2 ;
        RECT 1406.090 600.170 1406.370 604.000 ;
        RECT 1406.090 600.030 1406.980 600.170 ;
        RECT 1406.090 600.000 1406.370 600.030 ;
        RECT 1406.840 15.970 1406.980 600.030 ;
        RECT 1406.780 15.650 1407.040 15.970 ;
        RECT 1429.780 15.650 1430.040 15.970 ;
        RECT 1429.840 2.400 1429.980 15.650 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1416.870 586.740 1417.190 586.800 ;
        RECT 1420.090 586.740 1420.410 586.800 ;
        RECT 1416.870 586.600 1420.410 586.740 ;
        RECT 1416.870 586.540 1417.190 586.600 ;
        RECT 1420.090 586.540 1420.410 586.600 ;
        RECT 1420.550 20.640 1420.870 20.700 ;
        RECT 1447.690 20.640 1448.010 20.700 ;
        RECT 1420.550 20.500 1448.010 20.640 ;
        RECT 1420.550 20.440 1420.870 20.500 ;
        RECT 1447.690 20.440 1448.010 20.500 ;
      LAYER via ;
        RECT 1416.900 586.540 1417.160 586.800 ;
        RECT 1420.120 586.540 1420.380 586.800 ;
        RECT 1420.580 20.440 1420.840 20.700 ;
        RECT 1447.720 20.440 1447.980 20.700 ;
      LAYER met2 ;
        RECT 1415.290 600.170 1415.570 604.000 ;
        RECT 1415.290 600.030 1417.100 600.170 ;
        RECT 1415.290 600.000 1415.570 600.030 ;
        RECT 1416.960 586.830 1417.100 600.030 ;
        RECT 1416.900 586.510 1417.160 586.830 ;
        RECT 1420.120 586.510 1420.380 586.830 ;
        RECT 1420.180 582.490 1420.320 586.510 ;
        RECT 1420.180 582.350 1420.780 582.490 ;
        RECT 1420.640 20.730 1420.780 582.350 ;
        RECT 1420.580 20.410 1420.840 20.730 ;
        RECT 1447.720 20.410 1447.980 20.730 ;
        RECT 1447.780 2.400 1447.920 20.410 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1426.070 586.740 1426.390 586.800 ;
        RECT 1427.910 586.740 1428.230 586.800 ;
        RECT 1426.070 586.600 1428.230 586.740 ;
        RECT 1426.070 586.540 1426.390 586.600 ;
        RECT 1427.910 586.540 1428.230 586.600 ;
        RECT 1427.910 19.280 1428.230 19.340 ;
        RECT 1465.630 19.280 1465.950 19.340 ;
        RECT 1427.910 19.140 1465.950 19.280 ;
        RECT 1427.910 19.080 1428.230 19.140 ;
        RECT 1465.630 19.080 1465.950 19.140 ;
      LAYER via ;
        RECT 1426.100 586.540 1426.360 586.800 ;
        RECT 1427.940 586.540 1428.200 586.800 ;
        RECT 1427.940 19.080 1428.200 19.340 ;
        RECT 1465.660 19.080 1465.920 19.340 ;
      LAYER met2 ;
        RECT 1424.490 600.170 1424.770 604.000 ;
        RECT 1424.490 600.030 1426.300 600.170 ;
        RECT 1424.490 600.000 1424.770 600.030 ;
        RECT 1426.160 586.830 1426.300 600.030 ;
        RECT 1426.100 586.510 1426.360 586.830 ;
        RECT 1427.940 586.510 1428.200 586.830 ;
        RECT 1428.000 19.370 1428.140 586.510 ;
        RECT 1427.940 19.050 1428.200 19.370 ;
        RECT 1465.660 19.050 1465.920 19.370 ;
        RECT 1465.720 2.400 1465.860 19.050 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.350 17.920 1434.670 17.980 ;
        RECT 1483.570 17.920 1483.890 17.980 ;
        RECT 1434.350 17.780 1483.890 17.920 ;
        RECT 1434.350 17.720 1434.670 17.780 ;
        RECT 1483.570 17.720 1483.890 17.780 ;
      LAYER via ;
        RECT 1434.380 17.720 1434.640 17.980 ;
        RECT 1483.600 17.720 1483.860 17.980 ;
      LAYER met2 ;
        RECT 1433.690 600.170 1433.970 604.000 ;
        RECT 1433.690 600.030 1434.580 600.170 ;
        RECT 1433.690 600.000 1433.970 600.030 ;
        RECT 1434.440 18.010 1434.580 600.030 ;
        RECT 1434.380 17.690 1434.640 18.010 ;
        RECT 1483.600 17.690 1483.860 18.010 ;
        RECT 1483.660 2.400 1483.800 17.690 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1444.470 586.740 1444.790 586.800 ;
        RECT 1447.690 586.740 1448.010 586.800 ;
        RECT 1444.470 586.600 1448.010 586.740 ;
        RECT 1444.470 586.540 1444.790 586.600 ;
        RECT 1447.690 586.540 1448.010 586.600 ;
        RECT 1448.150 16.900 1448.470 16.960 ;
        RECT 1501.510 16.900 1501.830 16.960 ;
        RECT 1448.150 16.760 1501.830 16.900 ;
        RECT 1448.150 16.700 1448.470 16.760 ;
        RECT 1501.510 16.700 1501.830 16.760 ;
      LAYER via ;
        RECT 1444.500 586.540 1444.760 586.800 ;
        RECT 1447.720 586.540 1447.980 586.800 ;
        RECT 1448.180 16.700 1448.440 16.960 ;
        RECT 1501.540 16.700 1501.800 16.960 ;
      LAYER met2 ;
        RECT 1442.890 600.170 1443.170 604.000 ;
        RECT 1442.890 600.030 1444.700 600.170 ;
        RECT 1442.890 600.000 1443.170 600.030 ;
        RECT 1444.560 586.830 1444.700 600.030 ;
        RECT 1444.500 586.510 1444.760 586.830 ;
        RECT 1447.720 586.510 1447.980 586.830 ;
        RECT 1447.780 582.490 1447.920 586.510 ;
        RECT 1447.780 582.350 1448.380 582.490 ;
        RECT 1448.240 16.990 1448.380 582.350 ;
        RECT 1448.180 16.670 1448.440 16.990 ;
        RECT 1501.540 16.670 1501.800 16.990 ;
        RECT 1501.600 2.400 1501.740 16.670 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.510 20.300 1455.830 20.360 ;
        RECT 1518.990 20.300 1519.310 20.360 ;
        RECT 1455.510 20.160 1519.310 20.300 ;
        RECT 1455.510 20.100 1455.830 20.160 ;
        RECT 1518.990 20.100 1519.310 20.160 ;
      LAYER via ;
        RECT 1455.540 20.100 1455.800 20.360 ;
        RECT 1519.020 20.100 1519.280 20.360 ;
      LAYER met2 ;
        RECT 1452.090 600.170 1452.370 604.000 ;
        RECT 1452.090 600.030 1454.360 600.170 ;
        RECT 1452.090 600.000 1452.370 600.030 ;
        RECT 1454.220 583.170 1454.360 600.030 ;
        RECT 1454.220 583.030 1455.740 583.170 ;
        RECT 1455.600 20.390 1455.740 583.030 ;
        RECT 1455.540 20.070 1455.800 20.390 ;
        RECT 1519.020 20.070 1519.280 20.390 ;
        RECT 1519.080 2.400 1519.220 20.070 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 716.290 47.840 716.610 47.900 ;
        RECT 1035.530 47.840 1035.850 47.900 ;
        RECT 716.290 47.700 1035.850 47.840 ;
        RECT 716.290 47.640 716.610 47.700 ;
        RECT 1035.530 47.640 1035.850 47.700 ;
      LAYER via ;
        RECT 716.320 47.640 716.580 47.900 ;
        RECT 1035.560 47.640 1035.820 47.900 ;
      LAYER met2 ;
        RECT 1038.550 600.170 1038.830 604.000 ;
        RECT 1036.540 600.030 1038.830 600.170 ;
        RECT 1036.540 583.170 1036.680 600.030 ;
        RECT 1038.550 600.000 1038.830 600.030 ;
        RECT 1035.620 583.030 1036.680 583.170 ;
        RECT 1035.620 47.930 1035.760 583.030 ;
        RECT 716.320 47.610 716.580 47.930 ;
        RECT 1035.560 47.610 1035.820 47.930 ;
        RECT 716.380 2.400 716.520 47.610 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1462.410 17.240 1462.730 17.300 ;
        RECT 1536.930 17.240 1537.250 17.300 ;
        RECT 1462.410 17.100 1537.250 17.240 ;
        RECT 1462.410 17.040 1462.730 17.100 ;
        RECT 1536.930 17.040 1537.250 17.100 ;
      LAYER via ;
        RECT 1462.440 17.040 1462.700 17.300 ;
        RECT 1536.960 17.040 1537.220 17.300 ;
      LAYER met2 ;
        RECT 1461.290 600.170 1461.570 604.000 ;
        RECT 1461.290 600.030 1462.640 600.170 ;
        RECT 1461.290 600.000 1461.570 600.030 ;
        RECT 1462.500 17.330 1462.640 600.030 ;
        RECT 1462.440 17.010 1462.700 17.330 ;
        RECT 1536.960 17.010 1537.220 17.330 ;
        RECT 1537.020 2.400 1537.160 17.010 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1471.610 586.740 1471.930 586.800 ;
        RECT 1476.210 586.740 1476.530 586.800 ;
        RECT 1471.610 586.600 1476.530 586.740 ;
        RECT 1471.610 586.540 1471.930 586.600 ;
        RECT 1476.210 586.540 1476.530 586.600 ;
        RECT 1476.210 19.280 1476.530 19.340 ;
        RECT 1554.870 19.280 1555.190 19.340 ;
        RECT 1476.210 19.140 1555.190 19.280 ;
        RECT 1476.210 19.080 1476.530 19.140 ;
        RECT 1554.870 19.080 1555.190 19.140 ;
      LAYER via ;
        RECT 1471.640 586.540 1471.900 586.800 ;
        RECT 1476.240 586.540 1476.500 586.800 ;
        RECT 1476.240 19.080 1476.500 19.340 ;
        RECT 1554.900 19.080 1555.160 19.340 ;
      LAYER met2 ;
        RECT 1470.030 600.170 1470.310 604.000 ;
        RECT 1470.030 600.030 1471.840 600.170 ;
        RECT 1470.030 600.000 1470.310 600.030 ;
        RECT 1471.700 586.830 1471.840 600.030 ;
        RECT 1471.640 586.510 1471.900 586.830 ;
        RECT 1476.240 586.510 1476.500 586.830 ;
        RECT 1476.300 19.370 1476.440 586.510 ;
        RECT 1476.240 19.050 1476.500 19.370 ;
        RECT 1554.900 19.050 1555.160 19.370 ;
        RECT 1554.960 2.400 1555.100 19.050 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1480.810 589.120 1481.130 589.180 ;
        RECT 1480.810 588.980 1511.400 589.120 ;
        RECT 1480.810 588.920 1481.130 588.980 ;
        RECT 1511.260 588.440 1511.400 588.980 ;
        RECT 1511.260 588.300 1517.380 588.440 ;
        RECT 1517.240 587.420 1517.380 588.300 ;
        RECT 1517.240 587.280 1539.000 587.420 ;
        RECT 1538.860 586.740 1539.000 587.280 ;
        RECT 1562.690 586.740 1563.010 586.800 ;
        RECT 1538.860 586.600 1563.010 586.740 ;
        RECT 1562.690 586.540 1563.010 586.600 ;
        RECT 1562.690 20.640 1563.010 20.700 ;
        RECT 1572.810 20.640 1573.130 20.700 ;
        RECT 1562.690 20.500 1573.130 20.640 ;
        RECT 1562.690 20.440 1563.010 20.500 ;
        RECT 1572.810 20.440 1573.130 20.500 ;
      LAYER via ;
        RECT 1480.840 588.920 1481.100 589.180 ;
        RECT 1562.720 586.540 1562.980 586.800 ;
        RECT 1562.720 20.440 1562.980 20.700 ;
        RECT 1572.840 20.440 1573.100 20.700 ;
      LAYER met2 ;
        RECT 1479.230 600.170 1479.510 604.000 ;
        RECT 1479.230 600.030 1481.040 600.170 ;
        RECT 1479.230 600.000 1479.510 600.030 ;
        RECT 1480.900 589.210 1481.040 600.030 ;
        RECT 1480.840 588.890 1481.100 589.210 ;
        RECT 1562.720 586.510 1562.980 586.830 ;
        RECT 1562.780 20.730 1562.920 586.510 ;
        RECT 1562.720 20.410 1562.980 20.730 ;
        RECT 1572.840 20.410 1573.100 20.730 ;
        RECT 1572.900 2.400 1573.040 20.410 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 17.920 1490.330 17.980 ;
        RECT 1590.290 17.920 1590.610 17.980 ;
        RECT 1490.010 17.780 1590.610 17.920 ;
        RECT 1490.010 17.720 1490.330 17.780 ;
        RECT 1590.290 17.720 1590.610 17.780 ;
      LAYER via ;
        RECT 1490.040 17.720 1490.300 17.980 ;
        RECT 1590.320 17.720 1590.580 17.980 ;
      LAYER met2 ;
        RECT 1488.430 600.170 1488.710 604.000 ;
        RECT 1488.430 600.030 1490.240 600.170 ;
        RECT 1488.430 600.000 1488.710 600.030 ;
        RECT 1490.100 18.010 1490.240 600.030 ;
        RECT 1490.040 17.690 1490.300 18.010 ;
        RECT 1590.320 17.690 1590.580 18.010 ;
        RECT 1590.380 2.400 1590.520 17.690 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1499.210 586.740 1499.530 586.800 ;
        RECT 1503.810 586.740 1504.130 586.800 ;
        RECT 1499.210 586.600 1504.130 586.740 ;
        RECT 1499.210 586.540 1499.530 586.600 ;
        RECT 1503.810 586.540 1504.130 586.600 ;
        RECT 1547.970 18.940 1548.290 19.000 ;
        RECT 1608.230 18.940 1608.550 19.000 ;
        RECT 1547.970 18.800 1608.550 18.940 ;
        RECT 1547.970 18.740 1548.290 18.800 ;
        RECT 1608.230 18.740 1608.550 18.800 ;
        RECT 1503.810 16.900 1504.130 16.960 ;
        RECT 1547.970 16.900 1548.290 16.960 ;
        RECT 1503.810 16.760 1548.290 16.900 ;
        RECT 1503.810 16.700 1504.130 16.760 ;
        RECT 1547.970 16.700 1548.290 16.760 ;
      LAYER via ;
        RECT 1499.240 586.540 1499.500 586.800 ;
        RECT 1503.840 586.540 1504.100 586.800 ;
        RECT 1548.000 18.740 1548.260 19.000 ;
        RECT 1608.260 18.740 1608.520 19.000 ;
        RECT 1503.840 16.700 1504.100 16.960 ;
        RECT 1548.000 16.700 1548.260 16.960 ;
      LAYER met2 ;
        RECT 1497.630 600.170 1497.910 604.000 ;
        RECT 1497.630 600.030 1499.440 600.170 ;
        RECT 1497.630 600.000 1497.910 600.030 ;
        RECT 1499.300 586.830 1499.440 600.030 ;
        RECT 1499.240 586.510 1499.500 586.830 ;
        RECT 1503.840 586.510 1504.100 586.830 ;
        RECT 1503.900 16.990 1504.040 586.510 ;
        RECT 1548.000 18.710 1548.260 19.030 ;
        RECT 1608.260 18.710 1608.520 19.030 ;
        RECT 1548.060 16.990 1548.200 18.710 ;
        RECT 1503.840 16.670 1504.100 16.990 ;
        RECT 1548.000 16.670 1548.260 16.990 ;
        RECT 1608.320 2.400 1608.460 18.710 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1508.410 586.740 1508.730 586.800 ;
        RECT 1514.390 586.740 1514.710 586.800 ;
        RECT 1508.410 586.600 1514.710 586.740 ;
        RECT 1508.410 586.540 1508.730 586.600 ;
        RECT 1514.390 586.540 1514.710 586.600 ;
        RECT 1514.390 18.940 1514.710 19.000 ;
        RECT 1514.390 18.800 1540.840 18.940 ;
        RECT 1514.390 18.740 1514.710 18.800 ;
        RECT 1540.700 18.600 1540.840 18.800 ;
        RECT 1626.170 18.600 1626.490 18.660 ;
        RECT 1540.700 18.460 1626.490 18.600 ;
        RECT 1626.170 18.400 1626.490 18.460 ;
      LAYER via ;
        RECT 1508.440 586.540 1508.700 586.800 ;
        RECT 1514.420 586.540 1514.680 586.800 ;
        RECT 1514.420 18.740 1514.680 19.000 ;
        RECT 1626.200 18.400 1626.460 18.660 ;
      LAYER met2 ;
        RECT 1506.830 600.170 1507.110 604.000 ;
        RECT 1506.830 600.030 1508.640 600.170 ;
        RECT 1506.830 600.000 1507.110 600.030 ;
        RECT 1508.500 586.830 1508.640 600.030 ;
        RECT 1508.440 586.510 1508.700 586.830 ;
        RECT 1514.420 586.510 1514.680 586.830 ;
        RECT 1514.480 19.030 1514.620 586.510 ;
        RECT 1514.420 18.710 1514.680 19.030 ;
        RECT 1626.200 18.370 1626.460 18.690 ;
        RECT 1626.260 2.400 1626.400 18.370 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.150 587.080 1517.470 587.140 ;
        RECT 1528.190 587.080 1528.510 587.140 ;
        RECT 1517.150 586.940 1528.510 587.080 ;
        RECT 1517.150 586.880 1517.470 586.940 ;
        RECT 1528.190 586.880 1528.510 586.940 ;
        RECT 1528.190 18.260 1528.510 18.320 ;
        RECT 1644.110 18.260 1644.430 18.320 ;
        RECT 1528.190 18.120 1644.430 18.260 ;
        RECT 1528.190 18.060 1528.510 18.120 ;
        RECT 1644.110 18.060 1644.430 18.120 ;
      LAYER via ;
        RECT 1517.180 586.880 1517.440 587.140 ;
        RECT 1528.220 586.880 1528.480 587.140 ;
        RECT 1528.220 18.060 1528.480 18.320 ;
        RECT 1644.140 18.060 1644.400 18.320 ;
      LAYER met2 ;
        RECT 1516.030 600.170 1516.310 604.000 ;
        RECT 1516.030 600.030 1517.380 600.170 ;
        RECT 1516.030 600.000 1516.310 600.030 ;
        RECT 1517.240 587.170 1517.380 600.030 ;
        RECT 1517.180 586.850 1517.440 587.170 ;
        RECT 1528.220 586.850 1528.480 587.170 ;
        RECT 1528.280 18.350 1528.420 586.850 ;
        RECT 1528.220 18.030 1528.480 18.350 ;
        RECT 1644.140 18.030 1644.400 18.350 ;
        RECT 1644.200 2.400 1644.340 18.030 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1526.810 588.440 1527.130 588.500 ;
        RECT 1563.150 588.440 1563.470 588.500 ;
        RECT 1526.810 588.300 1563.470 588.440 ;
        RECT 1526.810 588.240 1527.130 588.300 ;
        RECT 1563.150 588.240 1563.470 588.300 ;
        RECT 1563.150 19.620 1563.470 19.680 ;
        RECT 1662.050 19.620 1662.370 19.680 ;
        RECT 1563.150 19.480 1662.370 19.620 ;
        RECT 1563.150 19.420 1563.470 19.480 ;
        RECT 1662.050 19.420 1662.370 19.480 ;
      LAYER via ;
        RECT 1526.840 588.240 1527.100 588.500 ;
        RECT 1563.180 588.240 1563.440 588.500 ;
        RECT 1563.180 19.420 1563.440 19.680 ;
        RECT 1662.080 19.420 1662.340 19.680 ;
      LAYER met2 ;
        RECT 1525.230 600.170 1525.510 604.000 ;
        RECT 1525.230 600.030 1527.040 600.170 ;
        RECT 1525.230 600.000 1525.510 600.030 ;
        RECT 1526.900 588.530 1527.040 600.030 ;
        RECT 1526.840 588.210 1527.100 588.530 ;
        RECT 1563.180 588.210 1563.440 588.530 ;
        RECT 1563.240 19.710 1563.380 588.210 ;
        RECT 1563.180 19.390 1563.440 19.710 ;
        RECT 1662.080 19.390 1662.340 19.710 ;
        RECT 1662.140 2.400 1662.280 19.390 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1536.010 587.760 1536.330 587.820 ;
        RECT 1536.010 587.620 1539.460 587.760 ;
        RECT 1536.010 587.560 1536.330 587.620 ;
        RECT 1539.320 587.420 1539.460 587.620 ;
        RECT 1570.510 587.420 1570.830 587.480 ;
        RECT 1539.320 587.280 1570.830 587.420 ;
        RECT 1570.510 587.220 1570.830 587.280 ;
        RECT 1570.050 579.600 1570.370 579.660 ;
        RECT 1570.510 579.600 1570.830 579.660 ;
        RECT 1570.050 579.460 1570.830 579.600 ;
        RECT 1570.050 579.400 1570.370 579.460 ;
        RECT 1570.510 579.400 1570.830 579.460 ;
        RECT 1570.510 545.260 1570.830 545.320 ;
        RECT 1570.140 545.120 1570.830 545.260 ;
        RECT 1570.140 544.980 1570.280 545.120 ;
        RECT 1570.510 545.060 1570.830 545.120 ;
        RECT 1570.050 544.720 1570.370 544.980 ;
        RECT 1569.590 496.980 1569.910 497.040 ;
        RECT 1570.510 496.980 1570.830 497.040 ;
        RECT 1569.590 496.840 1570.830 496.980 ;
        RECT 1569.590 496.780 1569.910 496.840 ;
        RECT 1570.510 496.780 1570.830 496.840 ;
        RECT 1569.590 427.620 1569.910 427.680 ;
        RECT 1570.050 427.620 1570.370 427.680 ;
        RECT 1569.590 427.480 1570.370 427.620 ;
        RECT 1569.590 427.420 1569.910 427.480 ;
        RECT 1570.050 427.420 1570.370 427.480 ;
        RECT 1570.050 420.820 1570.370 420.880 ;
        RECT 1570.970 420.820 1571.290 420.880 ;
        RECT 1570.050 420.680 1571.290 420.820 ;
        RECT 1570.050 420.620 1570.370 420.680 ;
        RECT 1570.970 420.620 1571.290 420.680 ;
        RECT 1570.050 289.720 1570.370 289.980 ;
        RECT 1570.140 289.300 1570.280 289.720 ;
        RECT 1570.050 289.040 1570.370 289.300 ;
        RECT 1570.050 255.380 1570.370 255.640 ;
        RECT 1570.140 254.960 1570.280 255.380 ;
        RECT 1570.050 254.700 1570.370 254.960 ;
        RECT 1568.670 217.500 1568.990 217.560 ;
        RECT 1570.050 217.500 1570.370 217.560 ;
        RECT 1568.670 217.360 1570.370 217.500 ;
        RECT 1568.670 217.300 1568.990 217.360 ;
        RECT 1570.050 217.300 1570.370 217.360 ;
        RECT 1568.670 193.360 1568.990 193.420 ;
        RECT 1569.590 193.360 1569.910 193.420 ;
        RECT 1568.670 193.220 1569.910 193.360 ;
        RECT 1568.670 193.160 1568.990 193.220 ;
        RECT 1569.590 193.160 1569.910 193.220 ;
        RECT 1568.210 144.400 1568.530 144.460 ;
        RECT 1569.590 144.400 1569.910 144.460 ;
        RECT 1568.210 144.260 1569.910 144.400 ;
        RECT 1568.210 144.200 1568.530 144.260 ;
        RECT 1569.590 144.200 1569.910 144.260 ;
        RECT 1568.210 96.800 1568.530 96.860 ;
        RECT 1569.590 96.800 1569.910 96.860 ;
        RECT 1568.210 96.660 1569.910 96.800 ;
        RECT 1568.210 96.600 1568.530 96.660 ;
        RECT 1569.590 96.600 1569.910 96.660 ;
        RECT 1569.590 19.280 1569.910 19.340 ;
        RECT 1679.530 19.280 1679.850 19.340 ;
        RECT 1569.590 19.140 1679.850 19.280 ;
        RECT 1569.590 19.080 1569.910 19.140 ;
        RECT 1679.530 19.080 1679.850 19.140 ;
      LAYER via ;
        RECT 1536.040 587.560 1536.300 587.820 ;
        RECT 1570.540 587.220 1570.800 587.480 ;
        RECT 1570.080 579.400 1570.340 579.660 ;
        RECT 1570.540 579.400 1570.800 579.660 ;
        RECT 1570.540 545.060 1570.800 545.320 ;
        RECT 1570.080 544.720 1570.340 544.980 ;
        RECT 1569.620 496.780 1569.880 497.040 ;
        RECT 1570.540 496.780 1570.800 497.040 ;
        RECT 1569.620 427.420 1569.880 427.680 ;
        RECT 1570.080 427.420 1570.340 427.680 ;
        RECT 1570.080 420.620 1570.340 420.880 ;
        RECT 1571.000 420.620 1571.260 420.880 ;
        RECT 1570.080 289.720 1570.340 289.980 ;
        RECT 1570.080 289.040 1570.340 289.300 ;
        RECT 1570.080 255.380 1570.340 255.640 ;
        RECT 1570.080 254.700 1570.340 254.960 ;
        RECT 1568.700 217.300 1568.960 217.560 ;
        RECT 1570.080 217.300 1570.340 217.560 ;
        RECT 1568.700 193.160 1568.960 193.420 ;
        RECT 1569.620 193.160 1569.880 193.420 ;
        RECT 1568.240 144.200 1568.500 144.460 ;
        RECT 1569.620 144.200 1569.880 144.460 ;
        RECT 1568.240 96.600 1568.500 96.860 ;
        RECT 1569.620 96.600 1569.880 96.860 ;
        RECT 1569.620 19.080 1569.880 19.340 ;
        RECT 1679.560 19.080 1679.820 19.340 ;
      LAYER met2 ;
        RECT 1534.430 600.170 1534.710 604.000 ;
        RECT 1534.430 600.030 1536.240 600.170 ;
        RECT 1534.430 600.000 1534.710 600.030 ;
        RECT 1536.100 587.850 1536.240 600.030 ;
        RECT 1536.040 587.530 1536.300 587.850 ;
        RECT 1570.540 587.190 1570.800 587.510 ;
        RECT 1570.600 579.770 1570.740 587.190 ;
        RECT 1570.140 579.690 1570.740 579.770 ;
        RECT 1570.080 579.630 1570.800 579.690 ;
        RECT 1570.080 579.370 1570.340 579.630 ;
        RECT 1570.540 579.370 1570.800 579.630 ;
        RECT 1570.140 579.215 1570.280 579.370 ;
        RECT 1570.600 545.350 1570.740 579.370 ;
        RECT 1570.540 545.030 1570.800 545.350 ;
        RECT 1570.080 544.690 1570.340 545.010 ;
        RECT 1570.140 531.490 1570.280 544.690 ;
        RECT 1570.140 531.350 1570.740 531.490 ;
        RECT 1570.600 497.070 1570.740 531.350 ;
        RECT 1569.620 496.750 1569.880 497.070 ;
        RECT 1570.540 496.750 1570.800 497.070 ;
        RECT 1569.680 427.710 1569.820 496.750 ;
        RECT 1569.620 427.390 1569.880 427.710 ;
        RECT 1570.080 427.390 1570.340 427.710 ;
        RECT 1570.140 420.910 1570.280 427.390 ;
        RECT 1570.080 420.590 1570.340 420.910 ;
        RECT 1571.000 420.590 1571.260 420.910 ;
        RECT 1571.060 337.010 1571.200 420.590 ;
        RECT 1570.140 336.870 1571.200 337.010 ;
        RECT 1570.140 290.010 1570.280 336.870 ;
        RECT 1570.080 289.690 1570.340 290.010 ;
        RECT 1570.080 289.010 1570.340 289.330 ;
        RECT 1570.140 255.670 1570.280 289.010 ;
        RECT 1570.080 255.350 1570.340 255.670 ;
        RECT 1570.080 254.670 1570.340 254.990 ;
        RECT 1570.140 217.590 1570.280 254.670 ;
        RECT 1568.700 217.270 1568.960 217.590 ;
        RECT 1570.080 217.270 1570.340 217.590 ;
        RECT 1568.760 193.450 1568.900 217.270 ;
        RECT 1568.700 193.130 1568.960 193.450 ;
        RECT 1569.620 193.130 1569.880 193.450 ;
        RECT 1569.680 144.490 1569.820 193.130 ;
        RECT 1568.240 144.170 1568.500 144.490 ;
        RECT 1569.620 144.170 1569.880 144.490 ;
        RECT 1568.300 96.890 1568.440 144.170 ;
        RECT 1568.240 96.570 1568.500 96.890 ;
        RECT 1569.620 96.570 1569.880 96.890 ;
        RECT 1569.680 19.370 1569.820 96.570 ;
        RECT 1569.620 19.050 1569.880 19.370 ;
        RECT 1679.560 19.050 1679.820 19.370 ;
        RECT 1679.620 2.400 1679.760 19.050 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.470 17.240 1697.790 17.300 ;
        RECT 1583.480 17.100 1697.790 17.240 ;
        RECT 1545.210 16.220 1545.530 16.280 ;
        RECT 1583.480 16.220 1583.620 17.100 ;
        RECT 1697.470 17.040 1697.790 17.100 ;
        RECT 1545.210 16.080 1583.620 16.220 ;
        RECT 1545.210 16.020 1545.530 16.080 ;
      LAYER via ;
        RECT 1545.240 16.020 1545.500 16.280 ;
        RECT 1697.500 17.040 1697.760 17.300 ;
      LAYER met2 ;
        RECT 1543.630 600.170 1543.910 604.000 ;
        RECT 1543.630 600.030 1545.440 600.170 ;
        RECT 1543.630 600.000 1543.910 600.030 ;
        RECT 1545.300 16.310 1545.440 600.030 ;
        RECT 1697.500 17.010 1697.760 17.330 ;
        RECT 1545.240 15.990 1545.500 16.310 ;
        RECT 1697.560 2.400 1697.700 17.010 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1042.430 583.340 1042.750 583.400 ;
        RECT 1046.110 583.340 1046.430 583.400 ;
        RECT 1042.430 583.200 1046.430 583.340 ;
        RECT 1042.430 583.140 1042.750 583.200 ;
        RECT 1046.110 583.140 1046.430 583.200 ;
        RECT 810.590 22.680 810.910 22.740 ;
        RECT 1042.430 22.680 1042.750 22.740 ;
        RECT 810.590 22.540 1042.750 22.680 ;
        RECT 810.590 22.480 810.910 22.540 ;
        RECT 1042.430 22.480 1042.750 22.540 ;
        RECT 734.230 17.580 734.550 17.640 ;
        RECT 810.590 17.580 810.910 17.640 ;
        RECT 734.230 17.440 810.910 17.580 ;
        RECT 734.230 17.380 734.550 17.440 ;
        RECT 810.590 17.380 810.910 17.440 ;
      LAYER via ;
        RECT 1042.460 583.140 1042.720 583.400 ;
        RECT 1046.140 583.140 1046.400 583.400 ;
        RECT 810.620 22.480 810.880 22.740 ;
        RECT 1042.460 22.480 1042.720 22.740 ;
        RECT 734.260 17.380 734.520 17.640 ;
        RECT 810.620 17.380 810.880 17.640 ;
      LAYER met2 ;
        RECT 1047.750 600.170 1048.030 604.000 ;
        RECT 1046.200 600.030 1048.030 600.170 ;
        RECT 1046.200 583.430 1046.340 600.030 ;
        RECT 1047.750 600.000 1048.030 600.030 ;
        RECT 1042.460 583.110 1042.720 583.430 ;
        RECT 1046.140 583.110 1046.400 583.430 ;
        RECT 1042.520 22.770 1042.660 583.110 ;
        RECT 810.620 22.450 810.880 22.770 ;
        RECT 1042.460 22.450 1042.720 22.770 ;
        RECT 810.680 17.670 810.820 22.450 ;
        RECT 734.260 17.350 734.520 17.670 ;
        RECT 810.620 17.350 810.880 17.670 ;
        RECT 734.320 2.400 734.460 17.350 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1554.410 587.080 1554.730 587.140 ;
        RECT 1576.490 587.080 1576.810 587.140 ;
        RECT 1554.410 586.940 1576.810 587.080 ;
        RECT 1554.410 586.880 1554.730 586.940 ;
        RECT 1576.490 586.880 1576.810 586.940 ;
        RECT 1576.490 17.580 1576.810 17.640 ;
        RECT 1715.410 17.580 1715.730 17.640 ;
        RECT 1576.490 17.440 1715.730 17.580 ;
        RECT 1576.490 17.380 1576.810 17.440 ;
        RECT 1715.410 17.380 1715.730 17.440 ;
      LAYER via ;
        RECT 1554.440 586.880 1554.700 587.140 ;
        RECT 1576.520 586.880 1576.780 587.140 ;
        RECT 1576.520 17.380 1576.780 17.640 ;
        RECT 1715.440 17.380 1715.700 17.640 ;
      LAYER met2 ;
        RECT 1552.830 600.170 1553.110 604.000 ;
        RECT 1552.830 600.030 1554.640 600.170 ;
        RECT 1552.830 600.000 1553.110 600.030 ;
        RECT 1554.500 587.170 1554.640 600.030 ;
        RECT 1554.440 586.850 1554.700 587.170 ;
        RECT 1576.520 586.850 1576.780 587.170 ;
        RECT 1576.580 17.670 1576.720 586.850 ;
        RECT 1576.520 17.350 1576.780 17.670 ;
        RECT 1715.440 17.350 1715.700 17.670 ;
        RECT 1715.500 2.400 1715.640 17.350 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1563.610 588.440 1563.930 588.500 ;
        RECT 1596.730 588.440 1597.050 588.500 ;
        RECT 1563.610 588.300 1597.050 588.440 ;
        RECT 1563.610 588.240 1563.930 588.300 ;
        RECT 1596.730 588.240 1597.050 588.300 ;
        RECT 1597.190 16.220 1597.510 16.280 ;
        RECT 1733.350 16.220 1733.670 16.280 ;
        RECT 1597.190 16.080 1733.670 16.220 ;
        RECT 1597.190 16.020 1597.510 16.080 ;
        RECT 1733.350 16.020 1733.670 16.080 ;
      LAYER via ;
        RECT 1563.640 588.240 1563.900 588.500 ;
        RECT 1596.760 588.240 1597.020 588.500 ;
        RECT 1597.220 16.020 1597.480 16.280 ;
        RECT 1733.380 16.020 1733.640 16.280 ;
      LAYER met2 ;
        RECT 1562.030 600.170 1562.310 604.000 ;
        RECT 1562.030 600.030 1563.840 600.170 ;
        RECT 1562.030 600.000 1562.310 600.030 ;
        RECT 1563.700 588.530 1563.840 600.030 ;
        RECT 1563.640 588.210 1563.900 588.530 ;
        RECT 1596.760 588.210 1597.020 588.530 ;
        RECT 1596.820 585.890 1596.960 588.210 ;
        RECT 1596.820 585.750 1597.420 585.890 ;
        RECT 1597.280 16.310 1597.420 585.750 ;
        RECT 1597.220 15.990 1597.480 16.310 ;
        RECT 1733.380 15.990 1733.640 16.310 ;
        RECT 1733.440 2.400 1733.580 15.990 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.810 589.460 1573.130 589.520 ;
        RECT 1610.990 589.460 1611.310 589.520 ;
        RECT 1572.810 589.320 1611.310 589.460 ;
        RECT 1572.810 589.260 1573.130 589.320 ;
        RECT 1610.990 589.260 1611.310 589.320 ;
        RECT 1610.990 15.880 1611.310 15.940 ;
        RECT 1751.290 15.880 1751.610 15.940 ;
        RECT 1610.990 15.740 1751.610 15.880 ;
        RECT 1610.990 15.680 1611.310 15.740 ;
        RECT 1751.290 15.680 1751.610 15.740 ;
      LAYER via ;
        RECT 1572.840 589.260 1573.100 589.520 ;
        RECT 1611.020 589.260 1611.280 589.520 ;
        RECT 1611.020 15.680 1611.280 15.940 ;
        RECT 1751.320 15.680 1751.580 15.940 ;
      LAYER met2 ;
        RECT 1571.230 600.170 1571.510 604.000 ;
        RECT 1571.230 600.030 1573.040 600.170 ;
        RECT 1571.230 600.000 1571.510 600.030 ;
        RECT 1572.900 589.550 1573.040 600.030 ;
        RECT 1572.840 589.230 1573.100 589.550 ;
        RECT 1611.020 589.230 1611.280 589.550 ;
        RECT 1611.080 15.970 1611.220 589.230 ;
        RECT 1611.020 15.650 1611.280 15.970 ;
        RECT 1751.320 15.650 1751.580 15.970 ;
        RECT 1751.380 2.400 1751.520 15.650 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1659.290 589.460 1659.610 589.520 ;
        RECT 1611.540 589.320 1659.610 589.460 ;
        RECT 1582.010 589.120 1582.330 589.180 ;
        RECT 1611.540 589.120 1611.680 589.320 ;
        RECT 1659.290 589.260 1659.610 589.320 ;
        RECT 1582.010 588.980 1611.680 589.120 ;
        RECT 1582.010 588.920 1582.330 588.980 ;
        RECT 1659.290 15.540 1659.610 15.600 ;
        RECT 1768.770 15.540 1769.090 15.600 ;
        RECT 1659.290 15.400 1769.090 15.540 ;
        RECT 1659.290 15.340 1659.610 15.400 ;
        RECT 1768.770 15.340 1769.090 15.400 ;
      LAYER via ;
        RECT 1582.040 588.920 1582.300 589.180 ;
        RECT 1659.320 589.260 1659.580 589.520 ;
        RECT 1659.320 15.340 1659.580 15.600 ;
        RECT 1768.800 15.340 1769.060 15.600 ;
      LAYER met2 ;
        RECT 1580.430 600.170 1580.710 604.000 ;
        RECT 1580.430 600.030 1582.240 600.170 ;
        RECT 1580.430 600.000 1580.710 600.030 ;
        RECT 1582.100 589.210 1582.240 600.030 ;
        RECT 1659.320 589.230 1659.580 589.550 ;
        RECT 1582.040 588.890 1582.300 589.210 ;
        RECT 1659.380 15.630 1659.520 589.230 ;
        RECT 1659.320 15.310 1659.580 15.630 ;
        RECT 1768.800 15.310 1769.060 15.630 ;
        RECT 1768.860 2.400 1769.000 15.310 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1591.210 586.740 1591.530 586.800 ;
        RECT 1593.510 586.740 1593.830 586.800 ;
        RECT 1591.210 586.600 1593.830 586.740 ;
        RECT 1591.210 586.540 1591.530 586.600 ;
        RECT 1593.510 586.540 1593.830 586.600 ;
        RECT 1593.510 17.920 1593.830 17.980 ;
        RECT 1786.710 17.920 1787.030 17.980 ;
        RECT 1593.510 17.780 1787.030 17.920 ;
        RECT 1593.510 17.720 1593.830 17.780 ;
        RECT 1786.710 17.720 1787.030 17.780 ;
      LAYER via ;
        RECT 1591.240 586.540 1591.500 586.800 ;
        RECT 1593.540 586.540 1593.800 586.800 ;
        RECT 1593.540 17.720 1593.800 17.980 ;
        RECT 1786.740 17.720 1787.000 17.980 ;
      LAYER met2 ;
        RECT 1589.630 600.170 1589.910 604.000 ;
        RECT 1589.630 600.030 1591.440 600.170 ;
        RECT 1589.630 600.000 1589.910 600.030 ;
        RECT 1591.300 586.830 1591.440 600.030 ;
        RECT 1591.240 586.510 1591.500 586.830 ;
        RECT 1593.540 586.510 1593.800 586.830 ;
        RECT 1593.600 18.010 1593.740 586.510 ;
        RECT 1593.540 17.690 1593.800 18.010 ;
        RECT 1786.740 17.690 1787.000 18.010 ;
        RECT 1786.800 2.400 1786.940 17.690 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.410 588.440 1600.730 588.500 ;
        RECT 1600.410 588.300 1622.720 588.440 ;
        RECT 1600.410 588.240 1600.730 588.300 ;
        RECT 1622.580 588.100 1622.720 588.300 ;
        RECT 1659.750 588.100 1660.070 588.160 ;
        RECT 1622.580 587.960 1660.070 588.100 ;
        RECT 1659.750 587.900 1660.070 587.960 ;
        RECT 1659.750 16.560 1660.070 16.620 ;
        RECT 1804.650 16.560 1804.970 16.620 ;
        RECT 1659.750 16.420 1804.970 16.560 ;
        RECT 1659.750 16.360 1660.070 16.420 ;
        RECT 1804.650 16.360 1804.970 16.420 ;
      LAYER via ;
        RECT 1600.440 588.240 1600.700 588.500 ;
        RECT 1659.780 587.900 1660.040 588.160 ;
        RECT 1659.780 16.360 1660.040 16.620 ;
        RECT 1804.680 16.360 1804.940 16.620 ;
      LAYER met2 ;
        RECT 1598.830 600.170 1599.110 604.000 ;
        RECT 1598.830 600.030 1600.640 600.170 ;
        RECT 1598.830 600.000 1599.110 600.030 ;
        RECT 1600.500 588.530 1600.640 600.030 ;
        RECT 1600.440 588.210 1600.700 588.530 ;
        RECT 1659.780 587.870 1660.040 588.190 ;
        RECT 1659.840 16.650 1659.980 587.870 ;
        RECT 1659.780 16.330 1660.040 16.650 ;
        RECT 1804.680 16.330 1804.940 16.650 ;
        RECT 1804.740 2.400 1804.880 16.330 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1609.610 588.780 1609.930 588.840 ;
        RECT 1789.930 588.780 1790.250 588.840 ;
        RECT 1609.610 588.640 1790.250 588.780 ;
        RECT 1609.610 588.580 1609.930 588.640 ;
        RECT 1789.930 588.580 1790.250 588.640 ;
        RECT 1790.390 17.920 1790.710 17.980 ;
        RECT 1822.590 17.920 1822.910 17.980 ;
        RECT 1790.390 17.780 1822.910 17.920 ;
        RECT 1790.390 17.720 1790.710 17.780 ;
        RECT 1822.590 17.720 1822.910 17.780 ;
      LAYER via ;
        RECT 1609.640 588.580 1609.900 588.840 ;
        RECT 1789.960 588.580 1790.220 588.840 ;
        RECT 1790.420 17.720 1790.680 17.980 ;
        RECT 1822.620 17.720 1822.880 17.980 ;
      LAYER met2 ;
        RECT 1608.030 600.170 1608.310 604.000 ;
        RECT 1608.030 600.030 1609.840 600.170 ;
        RECT 1608.030 600.000 1608.310 600.030 ;
        RECT 1609.700 588.870 1609.840 600.030 ;
        RECT 1609.640 588.550 1609.900 588.870 ;
        RECT 1789.960 588.550 1790.220 588.870 ;
        RECT 1790.020 585.890 1790.160 588.550 ;
        RECT 1790.020 585.750 1790.620 585.890 ;
        RECT 1790.480 18.010 1790.620 585.750 ;
        RECT 1790.420 17.690 1790.680 18.010 ;
        RECT 1822.620 17.690 1822.880 18.010 ;
        RECT 1822.680 2.400 1822.820 17.690 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1618.810 586.740 1619.130 586.800 ;
        RECT 1621.110 586.740 1621.430 586.800 ;
        RECT 1618.810 586.600 1621.430 586.740 ;
        RECT 1618.810 586.540 1619.130 586.600 ;
        RECT 1621.110 586.540 1621.430 586.600 ;
        RECT 1621.110 20.640 1621.430 20.700 ;
        RECT 1840.070 20.640 1840.390 20.700 ;
        RECT 1621.110 20.500 1840.390 20.640 ;
        RECT 1621.110 20.440 1621.430 20.500 ;
        RECT 1840.070 20.440 1840.390 20.500 ;
      LAYER via ;
        RECT 1618.840 586.540 1619.100 586.800 ;
        RECT 1621.140 586.540 1621.400 586.800 ;
        RECT 1621.140 20.440 1621.400 20.700 ;
        RECT 1840.100 20.440 1840.360 20.700 ;
      LAYER met2 ;
        RECT 1617.230 600.170 1617.510 604.000 ;
        RECT 1617.230 600.030 1619.040 600.170 ;
        RECT 1617.230 600.000 1617.510 600.030 ;
        RECT 1618.900 586.830 1619.040 600.030 ;
        RECT 1618.840 586.510 1619.100 586.830 ;
        RECT 1621.140 586.510 1621.400 586.830 ;
        RECT 1621.200 20.730 1621.340 586.510 ;
        RECT 1621.140 20.410 1621.400 20.730 ;
        RECT 1840.100 20.410 1840.360 20.730 ;
        RECT 1840.160 2.400 1840.300 20.410 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1628.010 20.300 1628.330 20.360 ;
        RECT 1858.010 20.300 1858.330 20.360 ;
        RECT 1628.010 20.160 1858.330 20.300 ;
        RECT 1628.010 20.100 1628.330 20.160 ;
        RECT 1858.010 20.100 1858.330 20.160 ;
      LAYER via ;
        RECT 1628.040 20.100 1628.300 20.360 ;
        RECT 1858.040 20.100 1858.300 20.360 ;
      LAYER met2 ;
        RECT 1626.430 600.170 1626.710 604.000 ;
        RECT 1626.430 600.030 1628.240 600.170 ;
        RECT 1626.430 600.000 1626.710 600.030 ;
        RECT 1628.100 20.390 1628.240 600.030 ;
        RECT 1628.040 20.070 1628.300 20.390 ;
        RECT 1858.040 20.070 1858.300 20.390 ;
        RECT 1858.100 2.400 1858.240 20.070 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1637.210 587.420 1637.530 587.480 ;
        RECT 1673.090 587.420 1673.410 587.480 ;
        RECT 1637.210 587.280 1673.410 587.420 ;
        RECT 1637.210 587.220 1637.530 587.280 ;
        RECT 1673.090 587.220 1673.410 587.280 ;
        RECT 1673.090 16.900 1673.410 16.960 ;
        RECT 1875.950 16.900 1876.270 16.960 ;
        RECT 1673.090 16.760 1876.270 16.900 ;
        RECT 1673.090 16.700 1673.410 16.760 ;
        RECT 1875.950 16.700 1876.270 16.760 ;
      LAYER via ;
        RECT 1637.240 587.220 1637.500 587.480 ;
        RECT 1673.120 587.220 1673.380 587.480 ;
        RECT 1673.120 16.700 1673.380 16.960 ;
        RECT 1875.980 16.700 1876.240 16.960 ;
      LAYER met2 ;
        RECT 1635.630 600.170 1635.910 604.000 ;
        RECT 1635.630 600.030 1637.440 600.170 ;
        RECT 1635.630 600.000 1635.910 600.030 ;
        RECT 1637.300 587.510 1637.440 600.030 ;
        RECT 1637.240 587.190 1637.500 587.510 ;
        RECT 1673.120 587.190 1673.380 587.510 ;
        RECT 1673.180 16.990 1673.320 587.190 ;
        RECT 1673.120 16.670 1673.380 16.990 ;
        RECT 1875.980 16.670 1876.240 16.990 ;
        RECT 1876.040 2.400 1876.180 16.670 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 752.170 30.840 752.490 30.900 ;
        RECT 1056.230 30.840 1056.550 30.900 ;
        RECT 752.170 30.700 1056.550 30.840 ;
        RECT 752.170 30.640 752.490 30.700 ;
        RECT 1056.230 30.640 1056.550 30.700 ;
      LAYER via ;
        RECT 752.200 30.640 752.460 30.900 ;
        RECT 1056.260 30.640 1056.520 30.900 ;
      LAYER met2 ;
        RECT 1056.950 600.170 1057.230 604.000 ;
        RECT 1056.320 600.030 1057.230 600.170 ;
        RECT 1056.320 30.930 1056.460 600.030 ;
        RECT 1056.950 600.000 1057.230 600.030 ;
        RECT 752.200 30.610 752.460 30.930 ;
        RECT 1056.260 30.610 1056.520 30.930 ;
        RECT 752.260 2.400 752.400 30.610 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1646.410 586.740 1646.730 586.800 ;
        RECT 1648.710 586.740 1649.030 586.800 ;
        RECT 1646.410 586.600 1649.030 586.740 ;
        RECT 1646.410 586.540 1646.730 586.600 ;
        RECT 1648.710 586.540 1649.030 586.600 ;
        RECT 1648.710 19.960 1649.030 20.020 ;
        RECT 1893.890 19.960 1894.210 20.020 ;
        RECT 1648.710 19.820 1894.210 19.960 ;
        RECT 1648.710 19.760 1649.030 19.820 ;
        RECT 1893.890 19.760 1894.210 19.820 ;
      LAYER via ;
        RECT 1646.440 586.540 1646.700 586.800 ;
        RECT 1648.740 586.540 1649.000 586.800 ;
        RECT 1648.740 19.760 1649.000 20.020 ;
        RECT 1893.920 19.760 1894.180 20.020 ;
      LAYER met2 ;
        RECT 1644.830 600.170 1645.110 604.000 ;
        RECT 1644.830 600.030 1646.640 600.170 ;
        RECT 1644.830 600.000 1645.110 600.030 ;
        RECT 1646.500 586.830 1646.640 600.030 ;
        RECT 1646.440 586.510 1646.700 586.830 ;
        RECT 1648.740 586.510 1649.000 586.830 ;
        RECT 1648.800 20.050 1648.940 586.510 ;
        RECT 1648.740 19.730 1649.000 20.050 ;
        RECT 1893.920 19.730 1894.180 20.050 ;
        RECT 1893.980 2.400 1894.120 19.730 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1655.610 589.120 1655.930 589.180 ;
        RECT 1686.890 589.120 1687.210 589.180 ;
        RECT 1655.610 588.980 1687.210 589.120 ;
        RECT 1655.610 588.920 1655.930 588.980 ;
        RECT 1686.890 588.920 1687.210 588.980 ;
        RECT 1686.890 15.200 1687.210 15.260 ;
        RECT 1911.830 15.200 1912.150 15.260 ;
        RECT 1686.890 15.060 1912.150 15.200 ;
        RECT 1686.890 15.000 1687.210 15.060 ;
        RECT 1911.830 15.000 1912.150 15.060 ;
      LAYER via ;
        RECT 1655.640 588.920 1655.900 589.180 ;
        RECT 1686.920 588.920 1687.180 589.180 ;
        RECT 1686.920 15.000 1687.180 15.260 ;
        RECT 1911.860 15.000 1912.120 15.260 ;
      LAYER met2 ;
        RECT 1654.030 600.170 1654.310 604.000 ;
        RECT 1654.030 600.030 1655.840 600.170 ;
        RECT 1654.030 600.000 1654.310 600.030 ;
        RECT 1655.700 589.210 1655.840 600.030 ;
        RECT 1655.640 588.890 1655.900 589.210 ;
        RECT 1686.920 588.890 1687.180 589.210 ;
        RECT 1686.980 15.290 1687.120 588.890 ;
        RECT 1686.920 14.970 1687.180 15.290 ;
        RECT 1911.860 14.970 1912.120 15.290 ;
        RECT 1911.920 2.400 1912.060 14.970 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1664.810 587.080 1665.130 587.140 ;
        RECT 1669.410 587.080 1669.730 587.140 ;
        RECT 1664.810 586.940 1669.730 587.080 ;
        RECT 1664.810 586.880 1665.130 586.940 ;
        RECT 1669.410 586.880 1669.730 586.940 ;
        RECT 1669.410 18.940 1669.730 19.000 ;
        RECT 1929.310 18.940 1929.630 19.000 ;
        RECT 1669.410 18.800 1929.630 18.940 ;
        RECT 1669.410 18.740 1669.730 18.800 ;
        RECT 1929.310 18.740 1929.630 18.800 ;
      LAYER via ;
        RECT 1664.840 586.880 1665.100 587.140 ;
        RECT 1669.440 586.880 1669.700 587.140 ;
        RECT 1669.440 18.740 1669.700 19.000 ;
        RECT 1929.340 18.740 1929.600 19.000 ;
      LAYER met2 ;
        RECT 1663.230 600.170 1663.510 604.000 ;
        RECT 1663.230 600.030 1665.040 600.170 ;
        RECT 1663.230 600.000 1663.510 600.030 ;
        RECT 1664.900 587.170 1665.040 600.030 ;
        RECT 1664.840 586.850 1665.100 587.170 ;
        RECT 1669.440 586.850 1669.700 587.170 ;
        RECT 1669.500 19.030 1669.640 586.850 ;
        RECT 1669.440 18.710 1669.700 19.030 ;
        RECT 1929.340 18.710 1929.600 19.030 ;
        RECT 1929.400 2.400 1929.540 18.710 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1674.010 587.080 1674.330 587.140 ;
        RECT 1693.790 587.080 1694.110 587.140 ;
        RECT 1674.010 586.940 1694.110 587.080 ;
        RECT 1674.010 586.880 1674.330 586.940 ;
        RECT 1693.790 586.880 1694.110 586.940 ;
        RECT 1693.790 19.620 1694.110 19.680 ;
        RECT 1947.250 19.620 1947.570 19.680 ;
        RECT 1693.790 19.480 1947.570 19.620 ;
        RECT 1693.790 19.420 1694.110 19.480 ;
        RECT 1947.250 19.420 1947.570 19.480 ;
      LAYER via ;
        RECT 1674.040 586.880 1674.300 587.140 ;
        RECT 1693.820 586.880 1694.080 587.140 ;
        RECT 1693.820 19.420 1694.080 19.680 ;
        RECT 1947.280 19.420 1947.540 19.680 ;
      LAYER met2 ;
        RECT 1672.430 600.170 1672.710 604.000 ;
        RECT 1672.430 600.030 1674.240 600.170 ;
        RECT 1672.430 600.000 1672.710 600.030 ;
        RECT 1674.100 587.170 1674.240 600.030 ;
        RECT 1674.040 586.850 1674.300 587.170 ;
        RECT 1693.820 586.850 1694.080 587.170 ;
        RECT 1693.880 19.710 1694.020 586.850 ;
        RECT 1693.820 19.390 1694.080 19.710 ;
        RECT 1947.280 19.390 1947.540 19.710 ;
        RECT 1947.340 2.400 1947.480 19.390 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.210 587.420 1683.530 587.480 ;
        RECT 1705.750 587.420 1706.070 587.480 ;
        RECT 1683.210 587.280 1706.070 587.420 ;
        RECT 1683.210 587.220 1683.530 587.280 ;
        RECT 1705.750 587.220 1706.070 587.280 ;
        RECT 1706.210 579.600 1706.530 579.660 ;
        RECT 1707.130 579.600 1707.450 579.660 ;
        RECT 1706.210 579.460 1707.450 579.600 ;
        RECT 1706.210 579.400 1706.530 579.460 ;
        RECT 1707.130 579.400 1707.450 579.460 ;
        RECT 1707.130 531.320 1707.450 531.380 ;
        RECT 1707.590 531.320 1707.910 531.380 ;
        RECT 1707.130 531.180 1707.910 531.320 ;
        RECT 1707.130 531.120 1707.450 531.180 ;
        RECT 1707.590 531.120 1707.910 531.180 ;
        RECT 1707.590 483.180 1707.910 483.440 ;
        RECT 1707.130 483.040 1707.450 483.100 ;
        RECT 1707.680 483.040 1707.820 483.180 ;
        RECT 1707.130 482.900 1707.820 483.040 ;
        RECT 1707.130 482.840 1707.450 482.900 ;
        RECT 1707.130 476.240 1707.450 476.300 ;
        RECT 1707.590 476.240 1707.910 476.300 ;
        RECT 1707.130 476.100 1707.910 476.240 ;
        RECT 1707.130 476.040 1707.450 476.100 ;
        RECT 1707.590 476.040 1707.910 476.100 ;
        RECT 1706.670 448.700 1706.990 448.760 ;
        RECT 1707.590 448.700 1707.910 448.760 ;
        RECT 1706.670 448.560 1707.910 448.700 ;
        RECT 1706.670 448.500 1706.990 448.560 ;
        RECT 1707.590 448.500 1707.910 448.560 ;
        RECT 1708.510 379.680 1708.830 379.740 ;
        RECT 1709.430 379.680 1709.750 379.740 ;
        RECT 1708.510 379.540 1709.750 379.680 ;
        RECT 1708.510 379.480 1708.830 379.540 ;
        RECT 1709.430 379.480 1709.750 379.540 ;
        RECT 1707.590 338.200 1707.910 338.260 ;
        RECT 1709.430 338.200 1709.750 338.260 ;
        RECT 1707.590 338.060 1709.750 338.200 ;
        RECT 1707.590 338.000 1707.910 338.060 ;
        RECT 1709.430 338.000 1709.750 338.060 ;
        RECT 1706.210 234.840 1706.530 234.900 ;
        RECT 1706.670 234.840 1706.990 234.900 ;
        RECT 1706.210 234.700 1706.990 234.840 ;
        RECT 1706.210 234.640 1706.530 234.700 ;
        RECT 1706.670 234.640 1706.990 234.700 ;
        RECT 1706.210 234.160 1706.530 234.220 ;
        RECT 1707.130 234.160 1707.450 234.220 ;
        RECT 1706.210 234.020 1707.450 234.160 ;
        RECT 1706.210 233.960 1706.530 234.020 ;
        RECT 1707.130 233.960 1707.450 234.020 ;
        RECT 1707.590 110.400 1707.910 110.460 ;
        RECT 1708.510 110.400 1708.830 110.460 ;
        RECT 1707.590 110.260 1708.830 110.400 ;
        RECT 1707.590 110.200 1707.910 110.260 ;
        RECT 1708.510 110.200 1708.830 110.260 ;
        RECT 1708.510 19.280 1708.830 19.340 ;
        RECT 1965.190 19.280 1965.510 19.340 ;
        RECT 1708.510 19.140 1965.510 19.280 ;
        RECT 1708.510 19.080 1708.830 19.140 ;
        RECT 1965.190 19.080 1965.510 19.140 ;
      LAYER via ;
        RECT 1683.240 587.220 1683.500 587.480 ;
        RECT 1705.780 587.220 1706.040 587.480 ;
        RECT 1706.240 579.400 1706.500 579.660 ;
        RECT 1707.160 579.400 1707.420 579.660 ;
        RECT 1707.160 531.120 1707.420 531.380 ;
        RECT 1707.620 531.120 1707.880 531.380 ;
        RECT 1707.620 483.180 1707.880 483.440 ;
        RECT 1707.160 482.840 1707.420 483.100 ;
        RECT 1707.160 476.040 1707.420 476.300 ;
        RECT 1707.620 476.040 1707.880 476.300 ;
        RECT 1706.700 448.500 1706.960 448.760 ;
        RECT 1707.620 448.500 1707.880 448.760 ;
        RECT 1708.540 379.480 1708.800 379.740 ;
        RECT 1709.460 379.480 1709.720 379.740 ;
        RECT 1707.620 338.000 1707.880 338.260 ;
        RECT 1709.460 338.000 1709.720 338.260 ;
        RECT 1706.240 234.640 1706.500 234.900 ;
        RECT 1706.700 234.640 1706.960 234.900 ;
        RECT 1706.240 233.960 1706.500 234.220 ;
        RECT 1707.160 233.960 1707.420 234.220 ;
        RECT 1707.620 110.200 1707.880 110.460 ;
        RECT 1708.540 110.200 1708.800 110.460 ;
        RECT 1708.540 19.080 1708.800 19.340 ;
        RECT 1965.220 19.080 1965.480 19.340 ;
      LAYER met2 ;
        RECT 1681.630 600.170 1681.910 604.000 ;
        RECT 1681.630 600.030 1683.440 600.170 ;
        RECT 1681.630 600.000 1681.910 600.030 ;
        RECT 1683.300 587.510 1683.440 600.030 ;
        RECT 1683.240 587.190 1683.500 587.510 ;
        RECT 1705.780 587.190 1706.040 587.510 ;
        RECT 1705.840 580.450 1705.980 587.190 ;
        RECT 1705.840 580.310 1706.210 580.450 ;
        RECT 1706.070 579.770 1706.210 580.310 ;
        RECT 1706.070 579.690 1706.440 579.770 ;
        RECT 1706.070 579.630 1706.500 579.690 ;
        RECT 1706.240 579.370 1706.500 579.630 ;
        RECT 1707.160 579.370 1707.420 579.690 ;
        RECT 1706.300 579.215 1706.440 579.370 ;
        RECT 1707.220 531.410 1707.360 579.370 ;
        RECT 1707.160 531.090 1707.420 531.410 ;
        RECT 1707.620 531.090 1707.880 531.410 ;
        RECT 1707.680 483.470 1707.820 531.090 ;
        RECT 1707.620 483.150 1707.880 483.470 ;
        RECT 1707.160 482.810 1707.420 483.130 ;
        RECT 1707.220 476.330 1707.360 482.810 ;
        RECT 1707.160 476.010 1707.420 476.330 ;
        RECT 1707.620 476.010 1707.880 476.330 ;
        RECT 1707.680 448.790 1707.820 476.010 ;
        RECT 1706.700 448.530 1706.960 448.790 ;
        RECT 1707.620 448.530 1707.880 448.790 ;
        RECT 1706.700 448.470 1707.880 448.530 ;
        RECT 1706.760 448.390 1707.820 448.470 ;
        RECT 1707.680 403.650 1707.820 448.390 ;
        RECT 1707.680 403.510 1708.740 403.650 ;
        RECT 1708.600 379.770 1708.740 403.510 ;
        RECT 1708.540 379.450 1708.800 379.770 ;
        RECT 1709.460 379.450 1709.720 379.770 ;
        RECT 1709.520 338.290 1709.660 379.450 ;
        RECT 1707.620 337.970 1707.880 338.290 ;
        RECT 1709.460 337.970 1709.720 338.290 ;
        RECT 1707.680 303.690 1707.820 337.970 ;
        RECT 1706.760 303.550 1707.820 303.690 ;
        RECT 1706.760 234.930 1706.900 303.550 ;
        RECT 1706.240 234.610 1706.500 234.930 ;
        RECT 1706.700 234.610 1706.960 234.930 ;
        RECT 1706.300 234.250 1706.440 234.610 ;
        RECT 1706.240 233.930 1706.500 234.250 ;
        RECT 1707.160 233.930 1707.420 234.250 ;
        RECT 1707.220 110.570 1707.360 233.930 ;
        RECT 1707.220 110.490 1707.820 110.570 ;
        RECT 1707.220 110.430 1707.880 110.490 ;
        RECT 1707.620 110.170 1707.880 110.430 ;
        RECT 1708.540 110.170 1708.800 110.490 ;
        RECT 1708.600 60.250 1708.740 110.170 ;
        RECT 1708.600 60.110 1709.200 60.250 ;
        RECT 1709.060 58.890 1709.200 60.110 ;
        RECT 1708.600 58.750 1709.200 58.890 ;
        RECT 1708.600 19.370 1708.740 58.750 ;
        RECT 1708.540 19.050 1708.800 19.370 ;
        RECT 1965.220 19.050 1965.480 19.370 ;
        RECT 1965.280 2.400 1965.420 19.050 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1692.410 591.840 1692.730 591.900 ;
        RECT 1981.290 591.840 1981.610 591.900 ;
        RECT 1692.410 591.700 1981.610 591.840 ;
        RECT 1692.410 591.640 1692.730 591.700 ;
        RECT 1981.290 591.640 1981.610 591.700 ;
      LAYER via ;
        RECT 1692.440 591.640 1692.700 591.900 ;
        RECT 1981.320 591.640 1981.580 591.900 ;
      LAYER met2 ;
        RECT 1690.830 600.170 1691.110 604.000 ;
        RECT 1690.830 600.030 1692.640 600.170 ;
        RECT 1690.830 600.000 1691.110 600.030 ;
        RECT 1692.500 591.930 1692.640 600.030 ;
        RECT 1692.440 591.610 1692.700 591.930 ;
        RECT 1981.320 591.610 1981.580 591.930 ;
        RECT 1981.380 3.130 1981.520 591.610 ;
        RECT 1981.380 2.990 1983.360 3.130 ;
        RECT 1983.220 2.400 1983.360 2.990 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1701.610 587.080 1701.930 587.140 ;
        RECT 1714.490 587.080 1714.810 587.140 ;
        RECT 1701.610 586.940 1714.810 587.080 ;
        RECT 1701.610 586.880 1701.930 586.940 ;
        RECT 1714.490 586.880 1714.810 586.940 ;
        RECT 1714.490 18.600 1714.810 18.660 ;
        RECT 2001.070 18.600 2001.390 18.660 ;
        RECT 1714.490 18.460 2001.390 18.600 ;
        RECT 1714.490 18.400 1714.810 18.460 ;
        RECT 2001.070 18.400 2001.390 18.460 ;
      LAYER via ;
        RECT 1701.640 586.880 1701.900 587.140 ;
        RECT 1714.520 586.880 1714.780 587.140 ;
        RECT 1714.520 18.400 1714.780 18.660 ;
        RECT 2001.100 18.400 2001.360 18.660 ;
      LAYER met2 ;
        RECT 1700.030 600.170 1700.310 604.000 ;
        RECT 1700.030 600.030 1701.840 600.170 ;
        RECT 1700.030 600.000 1700.310 600.030 ;
        RECT 1701.700 587.170 1701.840 600.030 ;
        RECT 1701.640 586.850 1701.900 587.170 ;
        RECT 1714.520 586.850 1714.780 587.170 ;
        RECT 1714.580 18.690 1714.720 586.850 ;
        RECT 1714.520 18.370 1714.780 18.690 ;
        RECT 2001.100 18.370 2001.360 18.690 ;
        RECT 2001.160 2.400 2001.300 18.370 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 592.520 1711.130 592.580 ;
        RECT 2004.750 592.520 2005.070 592.580 ;
        RECT 1710.810 592.380 2005.070 592.520 ;
        RECT 1710.810 592.320 1711.130 592.380 ;
        RECT 2004.750 592.320 2005.070 592.380 ;
        RECT 2002.910 531.320 2003.230 531.380 ;
        RECT 2004.290 531.320 2004.610 531.380 ;
        RECT 2002.910 531.180 2004.610 531.320 ;
        RECT 2002.910 531.120 2003.230 531.180 ;
        RECT 2004.290 531.120 2004.610 531.180 ;
        RECT 2002.910 483.380 2003.230 483.440 ;
        RECT 2003.830 483.380 2004.150 483.440 ;
        RECT 2002.910 483.240 2004.150 483.380 ;
        RECT 2002.910 483.180 2003.230 483.240 ;
        RECT 2003.830 483.180 2004.150 483.240 ;
        RECT 2003.830 458.900 2004.150 458.960 ;
        RECT 2005.210 458.900 2005.530 458.960 ;
        RECT 2003.830 458.760 2005.530 458.900 ;
        RECT 2003.830 458.700 2004.150 458.760 ;
        RECT 2005.210 458.700 2005.530 458.760 ;
        RECT 2003.830 427.620 2004.150 427.680 ;
        RECT 2004.750 427.620 2005.070 427.680 ;
        RECT 2003.830 427.480 2005.070 427.620 ;
        RECT 2003.830 427.420 2004.150 427.480 ;
        RECT 2004.750 427.420 2005.070 427.480 ;
        RECT 2004.750 352.140 2005.070 352.200 ;
        RECT 2004.750 352.000 2005.440 352.140 ;
        RECT 2004.750 351.940 2005.070 352.000 ;
        RECT 2005.300 351.860 2005.440 352.000 ;
        RECT 2005.210 351.600 2005.530 351.860 ;
        RECT 2004.750 338.200 2005.070 338.260 ;
        RECT 2005.210 338.200 2005.530 338.260 ;
        RECT 2004.750 338.060 2005.530 338.200 ;
        RECT 2004.750 338.000 2005.070 338.060 ;
        RECT 2005.210 338.000 2005.530 338.060 ;
        RECT 2003.830 283.120 2004.150 283.180 ;
        RECT 2004.750 283.120 2005.070 283.180 ;
        RECT 2003.830 282.980 2005.070 283.120 ;
        RECT 2003.830 282.920 2004.150 282.980 ;
        RECT 2004.750 282.920 2005.070 282.980 ;
        RECT 2002.910 193.020 2003.230 193.080 ;
        RECT 2003.830 193.020 2004.150 193.080 ;
        RECT 2002.910 192.880 2004.150 193.020 ;
        RECT 2002.910 192.820 2003.230 192.880 ;
        RECT 2003.830 192.820 2004.150 192.880 ;
        RECT 2002.910 145.080 2003.230 145.140 ;
        RECT 2004.290 145.080 2004.610 145.140 ;
        RECT 2002.910 144.940 2004.610 145.080 ;
        RECT 2002.910 144.880 2003.230 144.940 ;
        RECT 2004.290 144.880 2004.610 144.940 ;
        RECT 2003.830 96.460 2004.150 96.520 ;
        RECT 2005.210 96.460 2005.530 96.520 ;
        RECT 2003.830 96.320 2005.530 96.460 ;
        RECT 2003.830 96.260 2004.150 96.320 ;
        RECT 2005.210 96.260 2005.530 96.320 ;
        RECT 2003.830 48.520 2004.150 48.580 ;
        RECT 2004.750 48.520 2005.070 48.580 ;
        RECT 2003.830 48.380 2005.070 48.520 ;
        RECT 2003.830 48.320 2004.150 48.380 ;
        RECT 2004.750 48.320 2005.070 48.380 ;
        RECT 2004.750 3.980 2005.070 4.040 ;
        RECT 2018.550 3.980 2018.870 4.040 ;
        RECT 2004.750 3.840 2018.870 3.980 ;
        RECT 2004.750 3.780 2005.070 3.840 ;
        RECT 2018.550 3.780 2018.870 3.840 ;
      LAYER via ;
        RECT 1710.840 592.320 1711.100 592.580 ;
        RECT 2004.780 592.320 2005.040 592.580 ;
        RECT 2002.940 531.120 2003.200 531.380 ;
        RECT 2004.320 531.120 2004.580 531.380 ;
        RECT 2002.940 483.180 2003.200 483.440 ;
        RECT 2003.860 483.180 2004.120 483.440 ;
        RECT 2003.860 458.700 2004.120 458.960 ;
        RECT 2005.240 458.700 2005.500 458.960 ;
        RECT 2003.860 427.420 2004.120 427.680 ;
        RECT 2004.780 427.420 2005.040 427.680 ;
        RECT 2004.780 351.940 2005.040 352.200 ;
        RECT 2005.240 351.600 2005.500 351.860 ;
        RECT 2004.780 338.000 2005.040 338.260 ;
        RECT 2005.240 338.000 2005.500 338.260 ;
        RECT 2003.860 282.920 2004.120 283.180 ;
        RECT 2004.780 282.920 2005.040 283.180 ;
        RECT 2002.940 192.820 2003.200 193.080 ;
        RECT 2003.860 192.820 2004.120 193.080 ;
        RECT 2002.940 144.880 2003.200 145.140 ;
        RECT 2004.320 144.880 2004.580 145.140 ;
        RECT 2003.860 96.260 2004.120 96.520 ;
        RECT 2005.240 96.260 2005.500 96.520 ;
        RECT 2003.860 48.320 2004.120 48.580 ;
        RECT 2004.780 48.320 2005.040 48.580 ;
        RECT 2004.780 3.780 2005.040 4.040 ;
        RECT 2018.580 3.780 2018.840 4.040 ;
      LAYER met2 ;
        RECT 1709.230 600.170 1709.510 604.000 ;
        RECT 1709.230 600.030 1711.040 600.170 ;
        RECT 1709.230 600.000 1709.510 600.030 ;
        RECT 1710.900 592.610 1711.040 600.030 ;
        RECT 1710.840 592.290 1711.100 592.610 ;
        RECT 2004.780 592.290 2005.040 592.610 ;
        RECT 2004.840 545.090 2004.980 592.290 ;
        RECT 2004.380 544.950 2004.980 545.090 ;
        RECT 2004.380 531.410 2004.520 544.950 ;
        RECT 2002.940 531.090 2003.200 531.410 ;
        RECT 2004.320 531.090 2004.580 531.410 ;
        RECT 2003.000 483.470 2003.140 531.090 ;
        RECT 2002.940 483.150 2003.200 483.470 ;
        RECT 2003.860 483.150 2004.120 483.470 ;
        RECT 2003.920 458.990 2004.060 483.150 ;
        RECT 2003.860 458.670 2004.120 458.990 ;
        RECT 2005.240 458.670 2005.500 458.990 ;
        RECT 2005.300 434.930 2005.440 458.670 ;
        RECT 2004.840 434.790 2005.440 434.930 ;
        RECT 2004.840 427.710 2004.980 434.790 ;
        RECT 2003.860 427.390 2004.120 427.710 ;
        RECT 2004.780 427.390 2005.040 427.710 ;
        RECT 2003.920 385.290 2004.060 427.390 ;
        RECT 2003.920 385.150 2004.980 385.290 ;
        RECT 2004.840 352.230 2004.980 385.150 ;
        RECT 2004.780 351.910 2005.040 352.230 ;
        RECT 2005.240 351.570 2005.500 351.890 ;
        RECT 2005.300 338.290 2005.440 351.570 ;
        RECT 2004.780 337.970 2005.040 338.290 ;
        RECT 2005.240 337.970 2005.500 338.290 ;
        RECT 2004.840 283.210 2004.980 337.970 ;
        RECT 2003.860 282.890 2004.120 283.210 ;
        RECT 2004.780 282.890 2005.040 283.210 ;
        RECT 2003.920 193.110 2004.060 282.890 ;
        RECT 2002.940 192.790 2003.200 193.110 ;
        RECT 2003.860 192.790 2004.120 193.110 ;
        RECT 2003.000 145.170 2003.140 192.790 ;
        RECT 2002.940 144.850 2003.200 145.170 ;
        RECT 2004.320 144.850 2004.580 145.170 ;
        RECT 2004.380 110.570 2004.520 144.850 ;
        RECT 2004.380 110.430 2005.440 110.570 ;
        RECT 2005.300 96.550 2005.440 110.430 ;
        RECT 2003.860 96.230 2004.120 96.550 ;
        RECT 2005.240 96.230 2005.500 96.550 ;
        RECT 2003.920 48.610 2004.060 96.230 ;
        RECT 2003.860 48.290 2004.120 48.610 ;
        RECT 2004.780 48.290 2005.040 48.610 ;
        RECT 2004.840 4.070 2004.980 48.290 ;
        RECT 2004.780 3.750 2005.040 4.070 ;
        RECT 2018.580 3.750 2018.840 4.070 ;
        RECT 2018.640 2.400 2018.780 3.750 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1720.010 587.080 1720.330 587.140 ;
        RECT 1728.290 587.080 1728.610 587.140 ;
        RECT 1720.010 586.940 1728.610 587.080 ;
        RECT 1720.010 586.880 1720.330 586.940 ;
        RECT 1728.290 586.880 1728.610 586.940 ;
        RECT 1728.290 18.260 1728.610 18.320 ;
        RECT 2036.490 18.260 2036.810 18.320 ;
        RECT 1728.290 18.120 2036.810 18.260 ;
        RECT 1728.290 18.060 1728.610 18.120 ;
        RECT 2036.490 18.060 2036.810 18.120 ;
      LAYER via ;
        RECT 1720.040 586.880 1720.300 587.140 ;
        RECT 1728.320 586.880 1728.580 587.140 ;
        RECT 1728.320 18.060 1728.580 18.320 ;
        RECT 2036.520 18.060 2036.780 18.320 ;
      LAYER met2 ;
        RECT 1718.430 600.170 1718.710 604.000 ;
        RECT 1718.430 600.030 1720.240 600.170 ;
        RECT 1718.430 600.000 1718.710 600.030 ;
        RECT 1720.100 587.170 1720.240 600.030 ;
        RECT 1720.040 586.850 1720.300 587.170 ;
        RECT 1728.320 586.850 1728.580 587.170 ;
        RECT 1728.380 18.350 1728.520 586.850 ;
        RECT 1728.320 18.030 1728.580 18.350 ;
        RECT 2036.520 18.030 2036.780 18.350 ;
        RECT 2036.580 2.400 2036.720 18.030 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1729.210 589.460 1729.530 589.520 ;
        RECT 2038.790 589.460 2039.110 589.520 ;
        RECT 1729.210 589.320 2039.110 589.460 ;
        RECT 1729.210 589.260 1729.530 589.320 ;
        RECT 2038.790 589.260 2039.110 589.320 ;
        RECT 2038.790 18.260 2039.110 18.320 ;
        RECT 2054.430 18.260 2054.750 18.320 ;
        RECT 2038.790 18.120 2054.750 18.260 ;
        RECT 2038.790 18.060 2039.110 18.120 ;
        RECT 2054.430 18.060 2054.750 18.120 ;
      LAYER via ;
        RECT 1729.240 589.260 1729.500 589.520 ;
        RECT 2038.820 589.260 2039.080 589.520 ;
        RECT 2038.820 18.060 2039.080 18.320 ;
        RECT 2054.460 18.060 2054.720 18.320 ;
      LAYER met2 ;
        RECT 1727.630 600.170 1727.910 604.000 ;
        RECT 1727.630 600.030 1729.440 600.170 ;
        RECT 1727.630 600.000 1727.910 600.030 ;
        RECT 1729.300 589.550 1729.440 600.030 ;
        RECT 1729.240 589.230 1729.500 589.550 ;
        RECT 2038.820 589.230 2039.080 589.550 ;
        RECT 2038.880 18.350 2039.020 589.230 ;
        RECT 2038.820 18.030 2039.080 18.350 ;
        RECT 2054.460 18.030 2054.720 18.350 ;
        RECT 2054.520 2.400 2054.660 18.030 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1062.670 583.000 1062.990 583.060 ;
        RECT 1064.510 583.000 1064.830 583.060 ;
        RECT 1062.670 582.860 1064.830 583.000 ;
        RECT 1062.670 582.800 1062.990 582.860 ;
        RECT 1064.510 582.800 1064.830 582.860 ;
        RECT 769.650 31.180 769.970 31.240 ;
        RECT 1062.670 31.180 1062.990 31.240 ;
        RECT 769.650 31.040 1062.990 31.180 ;
        RECT 769.650 30.980 769.970 31.040 ;
        RECT 1062.670 30.980 1062.990 31.040 ;
      LAYER via ;
        RECT 1062.700 582.800 1062.960 583.060 ;
        RECT 1064.540 582.800 1064.800 583.060 ;
        RECT 769.680 30.980 769.940 31.240 ;
        RECT 1062.700 30.980 1062.960 31.240 ;
      LAYER met2 ;
        RECT 1066.150 600.170 1066.430 604.000 ;
        RECT 1064.600 600.030 1066.430 600.170 ;
        RECT 1064.600 583.090 1064.740 600.030 ;
        RECT 1066.150 600.000 1066.430 600.030 ;
        RECT 1062.700 582.770 1062.960 583.090 ;
        RECT 1064.540 582.770 1064.800 583.090 ;
        RECT 1062.760 31.270 1062.900 582.770 ;
        RECT 769.680 30.950 769.940 31.270 ;
        RECT 1062.700 30.950 1062.960 31.270 ;
        RECT 769.740 2.400 769.880 30.950 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1737.950 587.080 1738.270 587.140 ;
        RECT 1748.990 587.080 1749.310 587.140 ;
        RECT 1737.950 586.940 1749.310 587.080 ;
        RECT 1737.950 586.880 1738.270 586.940 ;
        RECT 1748.990 586.880 1749.310 586.940 ;
        RECT 1748.990 17.580 1749.310 17.640 ;
        RECT 2072.370 17.580 2072.690 17.640 ;
        RECT 1748.990 17.440 2072.690 17.580 ;
        RECT 1748.990 17.380 1749.310 17.440 ;
        RECT 2072.370 17.380 2072.690 17.440 ;
      LAYER via ;
        RECT 1737.980 586.880 1738.240 587.140 ;
        RECT 1749.020 586.880 1749.280 587.140 ;
        RECT 1749.020 17.380 1749.280 17.640 ;
        RECT 2072.400 17.380 2072.660 17.640 ;
      LAYER met2 ;
        RECT 1736.370 600.170 1736.650 604.000 ;
        RECT 1736.370 600.030 1738.180 600.170 ;
        RECT 1736.370 600.000 1736.650 600.030 ;
        RECT 1738.040 587.170 1738.180 600.030 ;
        RECT 1737.980 586.850 1738.240 587.170 ;
        RECT 1749.020 586.850 1749.280 587.170 ;
        RECT 1749.080 17.670 1749.220 586.850 ;
        RECT 1749.020 17.350 1749.280 17.670 ;
        RECT 2072.400 17.350 2072.660 17.670 ;
        RECT 2072.460 2.400 2072.600 17.350 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1747.150 593.200 1747.470 593.260 ;
        RECT 2084.790 593.200 2085.110 593.260 ;
        RECT 1747.150 593.060 2085.110 593.200 ;
        RECT 1747.150 593.000 1747.470 593.060 ;
        RECT 2084.790 593.000 2085.110 593.060 ;
        RECT 2084.790 2.960 2085.110 3.020 ;
        RECT 2089.850 2.960 2090.170 3.020 ;
        RECT 2084.790 2.820 2090.170 2.960 ;
        RECT 2084.790 2.760 2085.110 2.820 ;
        RECT 2089.850 2.760 2090.170 2.820 ;
      LAYER via ;
        RECT 1747.180 593.000 1747.440 593.260 ;
        RECT 2084.820 593.000 2085.080 593.260 ;
        RECT 2084.820 2.760 2085.080 3.020 ;
        RECT 2089.880 2.760 2090.140 3.020 ;
      LAYER met2 ;
        RECT 1745.570 600.170 1745.850 604.000 ;
        RECT 1745.570 600.030 1747.380 600.170 ;
        RECT 1745.570 600.000 1745.850 600.030 ;
        RECT 1747.240 593.290 1747.380 600.030 ;
        RECT 1747.180 592.970 1747.440 593.290 ;
        RECT 2084.820 592.970 2085.080 593.290 ;
        RECT 2084.880 3.050 2085.020 592.970 ;
        RECT 2084.820 2.730 2085.080 3.050 ;
        RECT 2089.880 2.730 2090.140 3.050 ;
        RECT 2089.940 2.400 2090.080 2.730 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1756.350 586.740 1756.670 586.800 ;
        RECT 1762.330 586.740 1762.650 586.800 ;
        RECT 1756.350 586.600 1762.650 586.740 ;
        RECT 1756.350 586.540 1756.670 586.600 ;
        RECT 1762.330 586.540 1762.650 586.600 ;
        RECT 1762.330 17.240 1762.650 17.300 ;
        RECT 2107.790 17.240 2108.110 17.300 ;
        RECT 1762.330 17.100 2108.110 17.240 ;
        RECT 1762.330 17.040 1762.650 17.100 ;
        RECT 2107.790 17.040 2108.110 17.100 ;
      LAYER via ;
        RECT 1756.380 586.540 1756.640 586.800 ;
        RECT 1762.360 586.540 1762.620 586.800 ;
        RECT 1762.360 17.040 1762.620 17.300 ;
        RECT 2107.820 17.040 2108.080 17.300 ;
      LAYER met2 ;
        RECT 1754.770 600.170 1755.050 604.000 ;
        RECT 1754.770 600.030 1756.580 600.170 ;
        RECT 1754.770 600.000 1755.050 600.030 ;
        RECT 1756.440 586.830 1756.580 600.030 ;
        RECT 1756.380 586.510 1756.640 586.830 ;
        RECT 1762.360 586.510 1762.620 586.830 ;
        RECT 1762.420 585.890 1762.560 586.510 ;
        RECT 1762.420 585.750 1763.020 585.890 ;
        RECT 1762.880 29.650 1763.020 585.750 ;
        RECT 1762.420 29.510 1763.020 29.650 ;
        RECT 1762.420 17.330 1762.560 29.510 ;
        RECT 1762.360 17.010 1762.620 17.330 ;
        RECT 2107.820 17.010 2108.080 17.330 ;
        RECT 2107.880 2.400 2108.020 17.010 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1765.550 588.100 1765.870 588.160 ;
        RECT 2126.650 588.100 2126.970 588.160 ;
        RECT 1765.550 587.960 2126.970 588.100 ;
        RECT 1765.550 587.900 1765.870 587.960 ;
        RECT 2126.650 587.900 2126.970 587.960 ;
        RECT 2125.730 2.960 2126.050 3.020 ;
        RECT 2126.650 2.960 2126.970 3.020 ;
        RECT 2125.730 2.820 2126.970 2.960 ;
        RECT 2125.730 2.760 2126.050 2.820 ;
        RECT 2126.650 2.760 2126.970 2.820 ;
      LAYER via ;
        RECT 1765.580 587.900 1765.840 588.160 ;
        RECT 2126.680 587.900 2126.940 588.160 ;
        RECT 2125.760 2.760 2126.020 3.020 ;
        RECT 2126.680 2.760 2126.940 3.020 ;
      LAYER met2 ;
        RECT 1763.970 600.170 1764.250 604.000 ;
        RECT 1763.970 600.030 1765.780 600.170 ;
        RECT 1763.970 600.000 1764.250 600.030 ;
        RECT 1765.640 588.190 1765.780 600.030 ;
        RECT 1765.580 587.870 1765.840 588.190 ;
        RECT 2126.680 587.870 2126.940 588.190 ;
        RECT 2126.740 3.050 2126.880 587.870 ;
        RECT 2125.760 2.730 2126.020 3.050 ;
        RECT 2126.680 2.730 2126.940 3.050 ;
        RECT 2125.820 2.400 2125.960 2.730 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1774.750 590.480 1775.070 590.540 ;
        RECT 1824.890 590.480 1825.210 590.540 ;
        RECT 1774.750 590.340 1825.210 590.480 ;
        RECT 1774.750 590.280 1775.070 590.340 ;
        RECT 1824.890 590.280 1825.210 590.340 ;
        RECT 1824.890 17.920 1825.210 17.980 ;
        RECT 2143.670 17.920 2143.990 17.980 ;
        RECT 1824.890 17.780 2143.990 17.920 ;
        RECT 1824.890 17.720 1825.210 17.780 ;
        RECT 2143.670 17.720 2143.990 17.780 ;
      LAYER via ;
        RECT 1774.780 590.280 1775.040 590.540 ;
        RECT 1824.920 590.280 1825.180 590.540 ;
        RECT 1824.920 17.720 1825.180 17.980 ;
        RECT 2143.700 17.720 2143.960 17.980 ;
      LAYER met2 ;
        RECT 1773.170 600.170 1773.450 604.000 ;
        RECT 1773.170 600.030 1774.980 600.170 ;
        RECT 1773.170 600.000 1773.450 600.030 ;
        RECT 1774.840 590.570 1774.980 600.030 ;
        RECT 1774.780 590.250 1775.040 590.570 ;
        RECT 1824.920 590.250 1825.180 590.570 ;
        RECT 1824.980 18.010 1825.120 590.250 ;
        RECT 1824.920 17.690 1825.180 18.010 ;
        RECT 2143.700 17.690 2143.960 18.010 ;
        RECT 2143.760 2.400 2143.900 17.690 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1783.950 591.160 1784.270 591.220 ;
        RECT 1783.950 591.020 1825.580 591.160 ;
        RECT 1783.950 590.960 1784.270 591.020 ;
        RECT 1825.440 590.480 1825.580 591.020 ;
        RECT 1825.440 590.340 1861.460 590.480 ;
        RECT 1861.320 590.140 1861.460 590.340 ;
        RECT 1873.190 590.140 1873.510 590.200 ;
        RECT 1861.320 590.000 1873.510 590.140 ;
        RECT 1873.190 589.940 1873.510 590.000 ;
        RECT 1873.190 15.540 1873.510 15.600 ;
        RECT 2161.610 15.540 2161.930 15.600 ;
        RECT 1873.190 15.400 2161.930 15.540 ;
        RECT 1873.190 15.340 1873.510 15.400 ;
        RECT 2161.610 15.340 2161.930 15.400 ;
      LAYER via ;
        RECT 1783.980 590.960 1784.240 591.220 ;
        RECT 1873.220 589.940 1873.480 590.200 ;
        RECT 1873.220 15.340 1873.480 15.600 ;
        RECT 2161.640 15.340 2161.900 15.600 ;
      LAYER met2 ;
        RECT 1782.370 600.170 1782.650 604.000 ;
        RECT 1782.370 600.030 1784.180 600.170 ;
        RECT 1782.370 600.000 1782.650 600.030 ;
        RECT 1784.040 591.250 1784.180 600.030 ;
        RECT 1783.980 590.930 1784.240 591.250 ;
        RECT 1873.220 589.910 1873.480 590.230 ;
        RECT 1873.280 15.630 1873.420 589.910 ;
        RECT 1873.220 15.310 1873.480 15.630 ;
        RECT 2161.640 15.310 2161.900 15.630 ;
        RECT 2161.700 2.400 2161.840 15.310 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 36.280 1793.930 36.340 ;
        RECT 2179.090 36.280 2179.410 36.340 ;
        RECT 1793.610 36.140 2179.410 36.280 ;
        RECT 1793.610 36.080 1793.930 36.140 ;
        RECT 2179.090 36.080 2179.410 36.140 ;
      LAYER via ;
        RECT 1793.640 36.080 1793.900 36.340 ;
        RECT 2179.120 36.080 2179.380 36.340 ;
      LAYER met2 ;
        RECT 1791.570 600.170 1791.850 604.000 ;
        RECT 1791.570 600.030 1793.840 600.170 ;
        RECT 1791.570 600.000 1791.850 600.030 ;
        RECT 1793.700 36.370 1793.840 600.030 ;
        RECT 1793.640 36.050 1793.900 36.370 ;
        RECT 2179.120 36.050 2179.380 36.370 ;
        RECT 2179.180 2.400 2179.320 36.050 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.440 588.980 1849.960 589.120 ;
        RECT 1802.350 588.440 1802.670 588.500 ;
        RECT 1848.440 588.440 1848.580 588.980 ;
        RECT 1802.350 588.300 1848.580 588.440 ;
        RECT 1849.820 588.440 1849.960 588.980 ;
        RECT 1973.470 588.580 1973.790 588.840 ;
        RECT 1974.390 588.780 1974.710 588.840 ;
        RECT 1974.390 588.640 2022.000 588.780 ;
        RECT 1974.390 588.580 1974.710 588.640 ;
        RECT 1901.250 588.440 1901.570 588.500 ;
        RECT 1849.820 588.300 1901.570 588.440 ;
        RECT 1802.350 588.240 1802.670 588.300 ;
        RECT 1901.250 588.240 1901.570 588.300 ;
        RECT 1966.110 588.440 1966.430 588.500 ;
        RECT 1973.560 588.440 1973.700 588.580 ;
        RECT 2021.860 588.500 2022.000 588.640 ;
        RECT 1966.110 588.300 1973.700 588.440 ;
        RECT 1966.110 588.240 1966.430 588.300 ;
        RECT 2021.770 588.240 2022.090 588.500 ;
        RECT 1901.250 587.420 1901.570 587.480 ;
        RECT 1918.270 587.420 1918.590 587.480 ;
        RECT 1901.250 587.280 1918.590 587.420 ;
        RECT 1901.250 587.220 1901.570 587.280 ;
        RECT 1918.270 587.220 1918.590 587.280 ;
        RECT 2021.770 586.060 2022.090 586.120 ;
        RECT 2052.590 586.060 2052.910 586.120 ;
        RECT 2021.770 585.920 2052.910 586.060 ;
        RECT 2021.770 585.860 2022.090 585.920 ;
        RECT 2052.590 585.860 2052.910 585.920 ;
        RECT 2052.590 15.200 2052.910 15.260 ;
        RECT 2197.030 15.200 2197.350 15.260 ;
        RECT 2052.590 15.060 2197.350 15.200 ;
        RECT 2052.590 15.000 2052.910 15.060 ;
        RECT 2197.030 15.000 2197.350 15.060 ;
      LAYER via ;
        RECT 1802.380 588.240 1802.640 588.500 ;
        RECT 1973.500 588.580 1973.760 588.840 ;
        RECT 1974.420 588.580 1974.680 588.840 ;
        RECT 1901.280 588.240 1901.540 588.500 ;
        RECT 1966.140 588.240 1966.400 588.500 ;
        RECT 2021.800 588.240 2022.060 588.500 ;
        RECT 1901.280 587.220 1901.540 587.480 ;
        RECT 1918.300 587.220 1918.560 587.480 ;
        RECT 2021.800 585.860 2022.060 586.120 ;
        RECT 2052.620 585.860 2052.880 586.120 ;
        RECT 2052.620 15.000 2052.880 15.260 ;
        RECT 2197.060 15.000 2197.320 15.260 ;
      LAYER met2 ;
        RECT 1800.770 600.170 1801.050 604.000 ;
        RECT 1800.770 600.030 1802.580 600.170 ;
        RECT 1800.770 600.000 1801.050 600.030 ;
        RECT 1802.440 588.530 1802.580 600.030 ;
        RECT 1973.500 588.610 1973.760 588.870 ;
        RECT 1974.420 588.610 1974.680 588.870 ;
        RECT 1973.500 588.550 1974.680 588.610 ;
        RECT 1802.380 588.210 1802.640 588.530 ;
        RECT 1901.280 588.210 1901.540 588.530 ;
        RECT 1966.140 588.210 1966.400 588.530 ;
        RECT 1973.560 588.470 1974.620 588.550 ;
        RECT 2021.800 588.210 2022.060 588.530 ;
        RECT 1901.340 587.510 1901.480 588.210 ;
        RECT 1966.200 588.045 1966.340 588.210 ;
        RECT 1966.130 587.675 1966.410 588.045 ;
        RECT 1901.280 587.190 1901.540 587.510 ;
        RECT 1918.300 587.365 1918.560 587.510 ;
        RECT 1918.290 586.995 1918.570 587.365 ;
        RECT 2021.860 586.150 2022.000 588.210 ;
        RECT 2021.800 585.830 2022.060 586.150 ;
        RECT 2052.620 585.830 2052.880 586.150 ;
        RECT 2052.680 15.290 2052.820 585.830 ;
        RECT 2052.620 14.970 2052.880 15.290 ;
        RECT 2197.060 14.970 2197.320 15.290 ;
        RECT 2197.120 2.400 2197.260 14.970 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
      LAYER via2 ;
        RECT 1966.130 587.720 1966.410 588.000 ;
        RECT 1918.290 587.040 1918.570 587.320 ;
      LAYER met3 ;
        RECT 1966.105 588.010 1966.435 588.025 ;
        RECT 1918.510 587.710 1966.435 588.010 ;
        RECT 1918.510 587.345 1918.810 587.710 ;
        RECT 1966.105 587.695 1966.435 587.710 ;
        RECT 1918.265 587.030 1918.810 587.345 ;
        RECT 1918.265 587.015 1918.595 587.030 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1811.550 591.500 1811.870 591.560 ;
        RECT 2214.970 591.500 2215.290 591.560 ;
        RECT 1811.550 591.360 2215.290 591.500 ;
        RECT 1811.550 591.300 1811.870 591.360 ;
        RECT 2214.970 591.300 2215.290 591.360 ;
      LAYER via ;
        RECT 1811.580 591.300 1811.840 591.560 ;
        RECT 2215.000 591.300 2215.260 591.560 ;
      LAYER met2 ;
        RECT 1809.970 600.170 1810.250 604.000 ;
        RECT 1809.970 600.030 1811.780 600.170 ;
        RECT 1809.970 600.000 1810.250 600.030 ;
        RECT 1811.640 591.590 1811.780 600.030 ;
        RECT 1811.580 591.270 1811.840 591.590 ;
        RECT 2215.000 591.270 2215.260 591.590 ;
        RECT 2215.060 2.400 2215.200 591.270 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1820.290 592.860 1820.610 592.920 ;
        RECT 1900.790 592.860 1901.110 592.920 ;
        RECT 1820.290 592.720 1901.110 592.860 ;
        RECT 1820.290 592.660 1820.610 592.720 ;
        RECT 1900.790 592.660 1901.110 592.720 ;
        RECT 1900.790 15.880 1901.110 15.940 ;
        RECT 2232.910 15.880 2233.230 15.940 ;
        RECT 1900.790 15.740 2233.230 15.880 ;
        RECT 1900.790 15.680 1901.110 15.740 ;
        RECT 2232.910 15.680 2233.230 15.740 ;
      LAYER via ;
        RECT 1820.320 592.660 1820.580 592.920 ;
        RECT 1900.820 592.660 1901.080 592.920 ;
        RECT 1900.820 15.680 1901.080 15.940 ;
        RECT 2232.940 15.680 2233.200 15.940 ;
      LAYER met2 ;
        RECT 1819.170 600.170 1819.450 604.000 ;
        RECT 1819.170 600.030 1820.520 600.170 ;
        RECT 1819.170 600.000 1819.450 600.030 ;
        RECT 1820.380 592.950 1820.520 600.030 ;
        RECT 1820.320 592.630 1820.580 592.950 ;
        RECT 1900.820 592.630 1901.080 592.950 ;
        RECT 1900.880 15.970 1901.020 592.630 ;
        RECT 1900.820 15.650 1901.080 15.970 ;
        RECT 2232.940 15.650 2233.200 15.970 ;
        RECT 2233.000 2.400 2233.140 15.650 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1070.030 583.000 1070.350 583.060 ;
        RECT 1073.710 583.000 1074.030 583.060 ;
        RECT 1070.030 582.860 1074.030 583.000 ;
        RECT 1070.030 582.800 1070.350 582.860 ;
        RECT 1073.710 582.800 1074.030 582.860 ;
        RECT 787.590 31.860 787.910 31.920 ;
        RECT 1070.030 31.860 1070.350 31.920 ;
        RECT 787.590 31.720 1070.350 31.860 ;
        RECT 787.590 31.660 787.910 31.720 ;
        RECT 1070.030 31.660 1070.350 31.720 ;
      LAYER via ;
        RECT 1070.060 582.800 1070.320 583.060 ;
        RECT 1073.740 582.800 1074.000 583.060 ;
        RECT 787.620 31.660 787.880 31.920 ;
        RECT 1070.060 31.660 1070.320 31.920 ;
      LAYER met2 ;
        RECT 1075.350 600.170 1075.630 604.000 ;
        RECT 1073.800 600.030 1075.630 600.170 ;
        RECT 1073.800 583.090 1073.940 600.030 ;
        RECT 1075.350 600.000 1075.630 600.030 ;
        RECT 1070.060 582.770 1070.320 583.090 ;
        RECT 1073.740 582.770 1074.000 583.090 ;
        RECT 1070.120 31.950 1070.260 582.770 ;
        RECT 787.620 31.630 787.880 31.950 ;
        RECT 1070.060 31.630 1070.320 31.950 ;
        RECT 787.680 2.400 787.820 31.630 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1829.950 591.160 1830.270 591.220 ;
        RECT 2249.470 591.160 2249.790 591.220 ;
        RECT 1829.950 591.020 2249.790 591.160 ;
        RECT 1829.950 590.960 1830.270 591.020 ;
        RECT 2249.470 590.960 2249.790 591.020 ;
      LAYER via ;
        RECT 1829.980 590.960 1830.240 591.220 ;
        RECT 2249.500 590.960 2249.760 591.220 ;
      LAYER met2 ;
        RECT 1828.370 600.170 1828.650 604.000 ;
        RECT 1828.370 600.030 1830.180 600.170 ;
        RECT 1828.370 600.000 1828.650 600.030 ;
        RECT 1830.040 591.250 1830.180 600.030 ;
        RECT 1829.980 590.930 1830.240 591.250 ;
        RECT 2249.500 590.930 2249.760 591.250 ;
        RECT 2249.560 3.130 2249.700 590.930 ;
        RECT 2249.560 2.990 2251.080 3.130 ;
        RECT 2250.940 2.400 2251.080 2.990 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1839.150 587.080 1839.470 587.140 ;
        RECT 1845.590 587.080 1845.910 587.140 ;
        RECT 1839.150 586.940 1845.910 587.080 ;
        RECT 1839.150 586.880 1839.470 586.940 ;
        RECT 1845.590 586.880 1845.910 586.940 ;
        RECT 1845.590 16.560 1845.910 16.620 ;
        RECT 2268.330 16.560 2268.650 16.620 ;
        RECT 1845.590 16.420 2268.650 16.560 ;
        RECT 1845.590 16.360 1845.910 16.420 ;
        RECT 2268.330 16.360 2268.650 16.420 ;
      LAYER via ;
        RECT 1839.180 586.880 1839.440 587.140 ;
        RECT 1845.620 586.880 1845.880 587.140 ;
        RECT 1845.620 16.360 1845.880 16.620 ;
        RECT 2268.360 16.360 2268.620 16.620 ;
      LAYER met2 ;
        RECT 1837.570 600.170 1837.850 604.000 ;
        RECT 1837.570 600.030 1839.380 600.170 ;
        RECT 1837.570 600.000 1837.850 600.030 ;
        RECT 1839.240 587.170 1839.380 600.030 ;
        RECT 1839.180 586.850 1839.440 587.170 ;
        RECT 1845.620 586.850 1845.880 587.170 ;
        RECT 1845.680 16.650 1845.820 586.850 ;
        RECT 1845.620 16.330 1845.880 16.650 ;
        RECT 2268.360 16.330 2268.620 16.650 ;
        RECT 2268.420 2.400 2268.560 16.330 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.350 592.180 1848.670 592.240 ;
        RECT 1873.190 592.180 1873.510 592.240 ;
        RECT 1848.350 592.040 1873.510 592.180 ;
        RECT 1848.350 591.980 1848.670 592.040 ;
        RECT 1873.190 591.980 1873.510 592.040 ;
        RECT 1873.190 590.820 1873.510 590.880 ;
        RECT 2283.970 590.820 2284.290 590.880 ;
        RECT 1873.190 590.680 2284.290 590.820 ;
        RECT 1873.190 590.620 1873.510 590.680 ;
        RECT 2283.970 590.620 2284.290 590.680 ;
        RECT 2283.970 2.960 2284.290 3.020 ;
        RECT 2286.270 2.960 2286.590 3.020 ;
        RECT 2283.970 2.820 2286.590 2.960 ;
        RECT 2283.970 2.760 2284.290 2.820 ;
        RECT 2286.270 2.760 2286.590 2.820 ;
      LAYER via ;
        RECT 1848.380 591.980 1848.640 592.240 ;
        RECT 1873.220 591.980 1873.480 592.240 ;
        RECT 1873.220 590.620 1873.480 590.880 ;
        RECT 2284.000 590.620 2284.260 590.880 ;
        RECT 2284.000 2.760 2284.260 3.020 ;
        RECT 2286.300 2.760 2286.560 3.020 ;
      LAYER met2 ;
        RECT 1846.770 600.170 1847.050 604.000 ;
        RECT 1846.770 600.030 1848.580 600.170 ;
        RECT 1846.770 600.000 1847.050 600.030 ;
        RECT 1848.440 592.270 1848.580 600.030 ;
        RECT 1848.380 591.950 1848.640 592.270 ;
        RECT 1873.220 591.950 1873.480 592.270 ;
        RECT 1873.280 590.910 1873.420 591.950 ;
        RECT 1873.220 590.590 1873.480 590.910 ;
        RECT 2284.000 590.590 2284.260 590.910 ;
        RECT 2284.060 3.050 2284.200 590.590 ;
        RECT 2284.000 2.730 2284.260 3.050 ;
        RECT 2286.300 2.730 2286.560 3.050 ;
        RECT 2286.360 2.400 2286.500 2.730 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1857.550 587.080 1857.870 587.140 ;
        RECT 1886.990 587.080 1887.310 587.140 ;
        RECT 1857.550 586.940 1887.310 587.080 ;
        RECT 1857.550 586.880 1857.870 586.940 ;
        RECT 1886.990 586.880 1887.310 586.940 ;
        RECT 1886.990 16.220 1887.310 16.280 ;
        RECT 2304.210 16.220 2304.530 16.280 ;
        RECT 1886.990 16.080 2304.530 16.220 ;
        RECT 1886.990 16.020 1887.310 16.080 ;
        RECT 2304.210 16.020 2304.530 16.080 ;
      LAYER via ;
        RECT 1857.580 586.880 1857.840 587.140 ;
        RECT 1887.020 586.880 1887.280 587.140 ;
        RECT 1887.020 16.020 1887.280 16.280 ;
        RECT 2304.240 16.020 2304.500 16.280 ;
      LAYER met2 ;
        RECT 1855.970 600.170 1856.250 604.000 ;
        RECT 1855.970 600.030 1857.780 600.170 ;
        RECT 1855.970 600.000 1856.250 600.030 ;
        RECT 1857.640 587.170 1857.780 600.030 ;
        RECT 1857.580 586.850 1857.840 587.170 ;
        RECT 1887.020 586.850 1887.280 587.170 ;
        RECT 1887.080 16.310 1887.220 586.850 ;
        RECT 1887.020 15.990 1887.280 16.310 ;
        RECT 2304.240 15.990 2304.500 16.310 ;
        RECT 2304.300 2.400 2304.440 15.990 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1866.750 590.480 1867.070 590.540 ;
        RECT 2318.470 590.480 2318.790 590.540 ;
        RECT 1866.750 590.340 2318.790 590.480 ;
        RECT 1866.750 590.280 1867.070 590.340 ;
        RECT 2318.470 590.280 2318.790 590.340 ;
      LAYER via ;
        RECT 1866.780 590.280 1867.040 590.540 ;
        RECT 2318.500 590.280 2318.760 590.540 ;
      LAYER met2 ;
        RECT 1865.170 600.170 1865.450 604.000 ;
        RECT 1865.170 600.030 1866.980 600.170 ;
        RECT 1865.170 600.000 1865.450 600.030 ;
        RECT 1866.840 590.570 1866.980 600.030 ;
        RECT 1866.780 590.250 1867.040 590.570 ;
        RECT 2318.500 590.250 2318.760 590.570 ;
        RECT 2318.560 17.410 2318.700 590.250 ;
        RECT 2318.560 17.270 2322.380 17.410 ;
        RECT 2322.240 2.400 2322.380 17.270 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.410 16.900 1876.730 16.960 ;
        RECT 2339.630 16.900 2339.950 16.960 ;
        RECT 1876.410 16.760 2339.950 16.900 ;
        RECT 1876.410 16.700 1876.730 16.760 ;
        RECT 2339.630 16.700 2339.950 16.760 ;
      LAYER via ;
        RECT 1876.440 16.700 1876.700 16.960 ;
        RECT 2339.660 16.700 2339.920 16.960 ;
      LAYER met2 ;
        RECT 1874.370 600.170 1874.650 604.000 ;
        RECT 1874.370 600.030 1876.640 600.170 ;
        RECT 1874.370 600.000 1874.650 600.030 ;
        RECT 1876.500 16.990 1876.640 600.030 ;
        RECT 1876.440 16.670 1876.700 16.990 ;
        RECT 2339.660 16.670 2339.920 16.990 ;
        RECT 2339.720 2.400 2339.860 16.670 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1885.150 590.140 1885.470 590.200 ;
        RECT 2352.970 590.140 2353.290 590.200 ;
        RECT 1885.150 590.000 2353.290 590.140 ;
        RECT 1885.150 589.940 1885.470 590.000 ;
        RECT 2352.970 589.940 2353.290 590.000 ;
      LAYER via ;
        RECT 1885.180 589.940 1885.440 590.200 ;
        RECT 2353.000 589.940 2353.260 590.200 ;
      LAYER met2 ;
        RECT 1883.570 600.170 1883.850 604.000 ;
        RECT 1883.570 600.030 1885.380 600.170 ;
        RECT 1883.570 600.000 1883.850 600.030 ;
        RECT 1885.240 590.230 1885.380 600.030 ;
        RECT 1885.180 589.910 1885.440 590.230 ;
        RECT 2353.000 589.910 2353.260 590.230 ;
        RECT 2353.060 16.730 2353.200 589.910 ;
        RECT 2353.060 16.590 2357.800 16.730 ;
        RECT 2357.660 2.400 2357.800 16.590 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1894.350 586.740 1894.670 586.800 ;
        RECT 1897.110 586.740 1897.430 586.800 ;
        RECT 1894.350 586.600 1897.430 586.740 ;
        RECT 1894.350 586.540 1894.670 586.600 ;
        RECT 1897.110 586.540 1897.430 586.600 ;
        RECT 1897.110 20.640 1897.430 20.700 ;
        RECT 2375.510 20.640 2375.830 20.700 ;
        RECT 1897.110 20.500 2375.830 20.640 ;
        RECT 1897.110 20.440 1897.430 20.500 ;
        RECT 2375.510 20.440 2375.830 20.500 ;
      LAYER via ;
        RECT 1894.380 586.540 1894.640 586.800 ;
        RECT 1897.140 586.540 1897.400 586.800 ;
        RECT 1897.140 20.440 1897.400 20.700 ;
        RECT 2375.540 20.440 2375.800 20.700 ;
      LAYER met2 ;
        RECT 1892.770 600.170 1893.050 604.000 ;
        RECT 1892.770 600.030 1894.580 600.170 ;
        RECT 1892.770 600.000 1893.050 600.030 ;
        RECT 1894.440 586.830 1894.580 600.030 ;
        RECT 1894.380 586.510 1894.640 586.830 ;
        RECT 1897.140 586.510 1897.400 586.830 ;
        RECT 1897.200 20.730 1897.340 586.510 ;
        RECT 1897.140 20.410 1897.400 20.730 ;
        RECT 2375.540 20.410 2375.800 20.730 ;
        RECT 2375.600 2.400 2375.740 20.410 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1903.550 589.800 1903.870 589.860 ;
        RECT 2387.470 589.800 2387.790 589.860 ;
        RECT 1903.550 589.660 2387.790 589.800 ;
        RECT 1903.550 589.600 1903.870 589.660 ;
        RECT 2387.470 589.600 2387.790 589.660 ;
        RECT 2387.470 20.640 2387.790 20.700 ;
        RECT 2393.450 20.640 2393.770 20.700 ;
        RECT 2387.470 20.500 2393.770 20.640 ;
        RECT 2387.470 20.440 2387.790 20.500 ;
        RECT 2393.450 20.440 2393.770 20.500 ;
      LAYER via ;
        RECT 1903.580 589.600 1903.840 589.860 ;
        RECT 2387.500 589.600 2387.760 589.860 ;
        RECT 2387.500 20.440 2387.760 20.700 ;
        RECT 2393.480 20.440 2393.740 20.700 ;
      LAYER met2 ;
        RECT 1901.970 600.170 1902.250 604.000 ;
        RECT 1901.970 600.030 1903.780 600.170 ;
        RECT 1901.970 600.000 1902.250 600.030 ;
        RECT 1903.640 589.890 1903.780 600.030 ;
        RECT 1903.580 589.570 1903.840 589.890 ;
        RECT 2387.500 589.570 2387.760 589.890 ;
        RECT 2387.560 20.730 2387.700 589.570 ;
        RECT 2387.500 20.410 2387.760 20.730 ;
        RECT 2393.480 20.410 2393.740 20.730 ;
        RECT 2393.540 2.400 2393.680 20.410 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1912.750 586.740 1913.070 586.800 ;
        RECT 1917.810 586.740 1918.130 586.800 ;
        RECT 1912.750 586.600 1918.130 586.740 ;
        RECT 1912.750 586.540 1913.070 586.600 ;
        RECT 1917.810 586.540 1918.130 586.600 ;
        RECT 1917.350 20.300 1917.670 20.360 ;
        RECT 2411.390 20.300 2411.710 20.360 ;
        RECT 1917.350 20.160 2411.710 20.300 ;
        RECT 1917.350 20.100 1917.670 20.160 ;
        RECT 2411.390 20.100 2411.710 20.160 ;
      LAYER via ;
        RECT 1912.780 586.540 1913.040 586.800 ;
        RECT 1917.840 586.540 1918.100 586.800 ;
        RECT 1917.380 20.100 1917.640 20.360 ;
        RECT 2411.420 20.100 2411.680 20.360 ;
      LAYER met2 ;
        RECT 1911.170 600.170 1911.450 604.000 ;
        RECT 1911.170 600.030 1912.980 600.170 ;
        RECT 1911.170 600.000 1911.450 600.030 ;
        RECT 1912.840 586.830 1912.980 600.030 ;
        RECT 1912.780 586.510 1913.040 586.830 ;
        RECT 1917.840 586.510 1918.100 586.830 ;
        RECT 1917.900 29.650 1918.040 586.510 ;
        RECT 1917.440 29.510 1918.040 29.650 ;
        RECT 1917.440 20.390 1917.580 29.510 ;
        RECT 1917.380 20.070 1917.640 20.390 ;
        RECT 2411.420 20.070 2411.680 20.390 ;
        RECT 2411.480 2.400 2411.620 20.070 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 805.530 31.520 805.850 31.580 ;
        RECT 1083.830 31.520 1084.150 31.580 ;
        RECT 805.530 31.380 1084.150 31.520 ;
        RECT 805.530 31.320 805.850 31.380 ;
        RECT 1083.830 31.320 1084.150 31.380 ;
      LAYER via ;
        RECT 805.560 31.320 805.820 31.580 ;
        RECT 1083.860 31.320 1084.120 31.580 ;
      LAYER met2 ;
        RECT 1084.550 600.170 1084.830 604.000 ;
        RECT 1083.920 600.030 1084.830 600.170 ;
        RECT 1083.920 31.610 1084.060 600.030 ;
        RECT 1084.550 600.000 1084.830 600.030 ;
        RECT 805.560 31.290 805.820 31.610 ;
        RECT 1083.860 31.290 1084.120 31.610 ;
        RECT 805.620 2.400 805.760 31.290 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 37.980 3.150 38.040 ;
        RECT 669.830 37.980 670.150 38.040 ;
        RECT 2.830 37.840 670.150 37.980 ;
        RECT 2.830 37.780 3.150 37.840 ;
        RECT 669.830 37.780 670.150 37.840 ;
      LAYER via ;
        RECT 2.860 37.780 3.120 38.040 ;
        RECT 669.860 37.780 670.120 38.040 ;
      LAYER met2 ;
        RECT 671.470 600.170 671.750 604.000 ;
        RECT 669.920 600.030 671.750 600.170 ;
        RECT 669.920 38.070 670.060 600.030 ;
        RECT 671.470 600.000 671.750 600.030 ;
        RECT 2.860 37.750 3.120 38.070 ;
        RECT 669.860 37.750 670.120 38.070 ;
        RECT 2.920 2.400 3.060 37.750 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 669.370 569.400 669.690 569.460 ;
        RECT 672.590 569.400 672.910 569.460 ;
        RECT 669.370 569.260 672.910 569.400 ;
        RECT 669.370 569.200 669.690 569.260 ;
        RECT 672.590 569.200 672.910 569.260 ;
        RECT 8.350 38.660 8.670 38.720 ;
        RECT 669.370 38.660 669.690 38.720 ;
        RECT 8.350 38.520 669.690 38.660 ;
        RECT 8.350 38.460 8.670 38.520 ;
        RECT 669.370 38.460 669.690 38.520 ;
      LAYER via ;
        RECT 669.400 569.200 669.660 569.460 ;
        RECT 672.620 569.200 672.880 569.460 ;
        RECT 8.380 38.460 8.640 38.720 ;
        RECT 669.400 38.460 669.660 38.720 ;
      LAYER met2 ;
        RECT 674.230 600.170 674.510 604.000 ;
        RECT 672.680 600.030 674.510 600.170 ;
        RECT 672.680 569.490 672.820 600.030 ;
        RECT 674.230 600.000 674.510 600.030 ;
        RECT 669.400 569.170 669.660 569.490 ;
        RECT 672.620 569.170 672.880 569.490 ;
        RECT 669.460 38.750 669.600 569.170 ;
        RECT 8.380 38.430 8.640 38.750 ;
        RECT 669.400 38.430 669.660 38.750 ;
        RECT 8.440 2.400 8.580 38.430 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 38.320 14.650 38.380 ;
        RECT 676.730 38.320 677.050 38.380 ;
        RECT 14.330 38.180 677.050 38.320 ;
        RECT 14.330 38.120 14.650 38.180 ;
        RECT 676.730 38.120 677.050 38.180 ;
      LAYER via ;
        RECT 14.360 38.120 14.620 38.380 ;
        RECT 676.760 38.120 677.020 38.380 ;
      LAYER met2 ;
        RECT 677.450 600.170 677.730 604.000 ;
        RECT 676.820 600.030 677.730 600.170 ;
        RECT 676.820 38.410 676.960 600.030 ;
        RECT 677.450 600.000 677.730 600.030 ;
        RECT 14.360 38.090 14.620 38.410 ;
        RECT 676.760 38.090 677.020 38.410 ;
        RECT 14.420 2.400 14.560 38.090 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 683.170 569.060 683.490 569.120 ;
        RECT 687.770 569.060 688.090 569.120 ;
        RECT 683.170 568.920 688.090 569.060 ;
        RECT 683.170 568.860 683.490 568.920 ;
        RECT 687.770 568.860 688.090 568.920 ;
        RECT 38.250 39.000 38.570 39.060 ;
        RECT 683.170 39.000 683.490 39.060 ;
        RECT 38.250 38.860 683.490 39.000 ;
        RECT 38.250 38.800 38.570 38.860 ;
        RECT 683.170 38.800 683.490 38.860 ;
      LAYER via ;
        RECT 683.200 568.860 683.460 569.120 ;
        RECT 687.800 568.860 688.060 569.120 ;
        RECT 38.280 38.800 38.540 39.060 ;
        RECT 683.200 38.800 683.460 39.060 ;
      LAYER met2 ;
        RECT 689.410 600.170 689.690 604.000 ;
        RECT 687.860 600.030 689.690 600.170 ;
        RECT 687.860 569.150 688.000 600.030 ;
        RECT 689.410 600.000 689.690 600.030 ;
        RECT 683.200 568.830 683.460 569.150 ;
        RECT 687.800 568.830 688.060 569.150 ;
        RECT 683.260 39.090 683.400 568.830 ;
        RECT 38.280 38.770 38.540 39.090 ;
        RECT 683.200 38.770 683.460 39.090 ;
        RECT 38.340 2.400 38.480 38.770 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 240.650 39.340 240.970 39.400 ;
        RECT 794.030 39.340 794.350 39.400 ;
        RECT 240.650 39.200 794.350 39.340 ;
        RECT 240.650 39.140 240.970 39.200 ;
        RECT 794.030 39.140 794.350 39.200 ;
      LAYER via ;
        RECT 240.680 39.140 240.940 39.400 ;
        RECT 794.060 39.140 794.320 39.400 ;
      LAYER met2 ;
        RECT 793.830 600.000 794.110 604.000 ;
        RECT 793.890 598.810 794.030 600.000 ;
        RECT 793.890 598.670 794.260 598.810 ;
        RECT 794.120 39.430 794.260 598.670 ;
        RECT 240.680 39.110 240.940 39.430 ;
        RECT 794.060 39.110 794.320 39.430 ;
        RECT 240.740 2.400 240.880 39.110 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 46.480 258.450 46.540 ;
        RECT 800.930 46.480 801.250 46.540 ;
        RECT 258.130 46.340 801.250 46.480 ;
        RECT 258.130 46.280 258.450 46.340 ;
        RECT 800.930 46.280 801.250 46.340 ;
      LAYER via ;
        RECT 258.160 46.280 258.420 46.540 ;
        RECT 800.960 46.280 801.220 46.540 ;
      LAYER met2 ;
        RECT 803.030 600.170 803.310 604.000 ;
        RECT 801.020 600.030 803.310 600.170 ;
        RECT 801.020 46.570 801.160 600.030 ;
        RECT 803.030 600.000 803.310 600.030 ;
        RECT 258.160 46.250 258.420 46.570 ;
        RECT 800.960 46.250 801.220 46.570 ;
        RECT 258.220 2.400 258.360 46.250 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 808.290 572.460 808.610 572.520 ;
        RECT 809.210 572.460 809.530 572.520 ;
        RECT 808.290 572.320 809.530 572.460 ;
        RECT 808.290 572.260 808.610 572.320 ;
        RECT 809.210 572.260 809.530 572.320 ;
        RECT 808.290 524.520 808.610 524.580 ;
        RECT 809.210 524.520 809.530 524.580 ;
        RECT 808.290 524.380 809.530 524.520 ;
        RECT 808.290 524.320 808.610 524.380 ;
        RECT 809.210 524.320 809.530 524.380 ;
        RECT 807.830 338.200 808.150 338.260 ;
        RECT 808.290 338.200 808.610 338.260 ;
        RECT 807.830 338.060 808.610 338.200 ;
        RECT 807.830 338.000 808.150 338.060 ;
        RECT 808.290 338.000 808.610 338.060 ;
        RECT 807.830 241.640 808.150 241.700 ;
        RECT 808.750 241.640 809.070 241.700 ;
        RECT 807.830 241.500 809.070 241.640 ;
        RECT 807.830 241.440 808.150 241.500 ;
        RECT 808.750 241.440 809.070 241.500 ;
        RECT 807.830 193.360 808.150 193.420 ;
        RECT 808.290 193.360 808.610 193.420 ;
        RECT 807.830 193.220 808.610 193.360 ;
        RECT 807.830 193.160 808.150 193.220 ;
        RECT 808.290 193.160 808.610 193.220 ;
        RECT 808.290 145.420 808.610 145.480 ;
        RECT 807.920 145.280 808.610 145.420 ;
        RECT 807.920 145.140 808.060 145.280 ;
        RECT 808.290 145.220 808.610 145.280 ;
        RECT 807.830 144.880 808.150 145.140 ;
        RECT 807.830 96.800 808.150 96.860 ;
        RECT 808.290 96.800 808.610 96.860 ;
        RECT 807.830 96.660 808.610 96.800 ;
        RECT 807.830 96.600 808.150 96.660 ;
        RECT 808.290 96.600 808.610 96.660 ;
        RECT 774.250 89.660 774.570 89.720 ;
        RECT 808.290 89.660 808.610 89.720 ;
        RECT 774.250 89.520 808.610 89.660 ;
        RECT 774.250 89.460 774.570 89.520 ;
        RECT 808.290 89.460 808.610 89.520 ;
        RECT 276.070 46.820 276.390 46.880 ;
        RECT 774.250 46.820 774.570 46.880 ;
        RECT 276.070 46.680 774.570 46.820 ;
        RECT 276.070 46.620 276.390 46.680 ;
        RECT 774.250 46.620 774.570 46.680 ;
      LAYER via ;
        RECT 808.320 572.260 808.580 572.520 ;
        RECT 809.240 572.260 809.500 572.520 ;
        RECT 808.320 524.320 808.580 524.580 ;
        RECT 809.240 524.320 809.500 524.580 ;
        RECT 807.860 338.000 808.120 338.260 ;
        RECT 808.320 338.000 808.580 338.260 ;
        RECT 807.860 241.440 808.120 241.700 ;
        RECT 808.780 241.440 809.040 241.700 ;
        RECT 807.860 193.160 808.120 193.420 ;
        RECT 808.320 193.160 808.580 193.420 ;
        RECT 808.320 145.220 808.580 145.480 ;
        RECT 807.860 144.880 808.120 145.140 ;
        RECT 807.860 96.600 808.120 96.860 ;
        RECT 808.320 96.600 808.580 96.860 ;
        RECT 774.280 89.460 774.540 89.720 ;
        RECT 808.320 89.460 808.580 89.720 ;
        RECT 276.100 46.620 276.360 46.880 ;
        RECT 774.280 46.620 774.540 46.880 ;
      LAYER met2 ;
        RECT 812.230 600.850 812.510 604.000 ;
        RECT 809.760 600.710 812.510 600.850 ;
        RECT 809.760 596.770 809.900 600.710 ;
        RECT 812.230 600.000 812.510 600.710 ;
        RECT 808.380 596.630 809.900 596.770 ;
        RECT 808.380 572.550 808.520 596.630 ;
        RECT 808.320 572.230 808.580 572.550 ;
        RECT 809.240 572.230 809.500 572.550 ;
        RECT 809.300 524.610 809.440 572.230 ;
        RECT 808.320 524.290 808.580 524.610 ;
        RECT 809.240 524.290 809.500 524.610 ;
        RECT 808.380 400.930 808.520 524.290 ;
        RECT 808.380 400.790 808.980 400.930 ;
        RECT 808.840 399.570 808.980 400.790 ;
        RECT 808.380 399.430 808.980 399.570 ;
        RECT 808.380 338.290 808.520 399.430 ;
        RECT 807.860 337.970 808.120 338.290 ;
        RECT 808.320 337.970 808.580 338.290 ;
        RECT 807.920 307.090 808.060 337.970 ;
        RECT 807.920 306.950 808.980 307.090 ;
        RECT 808.840 303.010 808.980 306.950 ;
        RECT 808.380 302.870 808.980 303.010 ;
        RECT 808.380 266.290 808.520 302.870 ;
        RECT 808.380 266.150 808.980 266.290 ;
        RECT 808.840 241.730 808.980 266.150 ;
        RECT 807.860 241.410 808.120 241.730 ;
        RECT 808.780 241.410 809.040 241.730 ;
        RECT 807.920 193.450 808.060 241.410 ;
        RECT 807.860 193.130 808.120 193.450 ;
        RECT 808.320 193.130 808.580 193.450 ;
        RECT 808.380 145.510 808.520 193.130 ;
        RECT 808.320 145.190 808.580 145.510 ;
        RECT 807.860 144.850 808.120 145.170 ;
        RECT 807.920 96.890 808.060 144.850 ;
        RECT 807.860 96.570 808.120 96.890 ;
        RECT 808.320 96.570 808.580 96.890 ;
        RECT 808.380 89.750 808.520 96.570 ;
        RECT 774.280 89.430 774.540 89.750 ;
        RECT 808.320 89.430 808.580 89.750 ;
        RECT 774.340 46.910 774.480 89.430 ;
        RECT 276.100 46.590 276.360 46.910 ;
        RECT 774.280 46.590 774.540 46.910 ;
        RECT 276.160 2.400 276.300 46.590 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 47.160 294.330 47.220 ;
        RECT 821.630 47.160 821.950 47.220 ;
        RECT 294.010 47.020 821.950 47.160 ;
        RECT 294.010 46.960 294.330 47.020 ;
        RECT 821.630 46.960 821.950 47.020 ;
      LAYER via ;
        RECT 294.040 46.960 294.300 47.220 ;
        RECT 821.660 46.960 821.920 47.220 ;
      LAYER met2 ;
        RECT 821.430 600.000 821.710 604.000 ;
        RECT 821.490 598.810 821.630 600.000 ;
        RECT 821.490 598.670 821.860 598.810 ;
        RECT 821.720 47.250 821.860 598.670 ;
        RECT 294.040 46.930 294.300 47.250 ;
        RECT 821.660 46.930 821.920 47.250 ;
        RECT 294.100 2.400 294.240 46.930 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 47.500 312.270 47.560 ;
        RECT 828.530 47.500 828.850 47.560 ;
        RECT 311.950 47.360 828.850 47.500 ;
        RECT 311.950 47.300 312.270 47.360 ;
        RECT 828.530 47.300 828.850 47.360 ;
      LAYER via ;
        RECT 311.980 47.300 312.240 47.560 ;
        RECT 828.560 47.300 828.820 47.560 ;
      LAYER met2 ;
        RECT 830.630 600.170 830.910 604.000 ;
        RECT 828.620 600.030 830.910 600.170 ;
        RECT 828.620 47.590 828.760 600.030 ;
        RECT 830.630 600.000 830.910 600.030 ;
        RECT 311.980 47.270 312.240 47.590 ;
        RECT 828.560 47.270 828.820 47.590 ;
        RECT 312.040 2.400 312.180 47.270 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.970 569.400 835.290 569.460 ;
        RECT 838.190 569.400 838.510 569.460 ;
        RECT 834.970 569.260 838.510 569.400 ;
        RECT 834.970 569.200 835.290 569.260 ;
        RECT 838.190 569.200 838.510 569.260 ;
        RECT 329.890 26.080 330.210 26.140 ;
        RECT 834.970 26.080 835.290 26.140 ;
        RECT 329.890 25.940 835.290 26.080 ;
        RECT 329.890 25.880 330.210 25.940 ;
        RECT 834.970 25.880 835.290 25.940 ;
      LAYER via ;
        RECT 835.000 569.200 835.260 569.460 ;
        RECT 838.220 569.200 838.480 569.460 ;
        RECT 329.920 25.880 330.180 26.140 ;
        RECT 835.000 25.880 835.260 26.140 ;
      LAYER met2 ;
        RECT 839.830 600.170 840.110 604.000 ;
        RECT 838.280 600.030 840.110 600.170 ;
        RECT 838.280 569.490 838.420 600.030 ;
        RECT 839.830 600.000 840.110 600.030 ;
        RECT 835.000 569.170 835.260 569.490 ;
        RECT 838.220 569.170 838.480 569.490 ;
        RECT 835.060 26.170 835.200 569.170 ;
        RECT 329.920 25.850 330.180 26.170 ;
        RECT 835.000 25.850 835.260 26.170 ;
        RECT 329.980 2.400 330.120 25.850 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 26.420 347.690 26.480 ;
        RECT 849.690 26.420 850.010 26.480 ;
        RECT 347.370 26.280 850.010 26.420 ;
        RECT 347.370 26.220 347.690 26.280 ;
        RECT 849.690 26.220 850.010 26.280 ;
      LAYER via ;
        RECT 347.400 26.220 347.660 26.480 ;
        RECT 849.720 26.220 849.980 26.480 ;
      LAYER met2 ;
        RECT 848.570 600.170 848.850 604.000 ;
        RECT 848.570 600.030 849.920 600.170 ;
        RECT 848.570 600.000 848.850 600.030 ;
        RECT 849.780 26.510 849.920 600.030 ;
        RECT 347.400 26.190 347.660 26.510 ;
        RECT 849.720 26.190 849.980 26.510 ;
        RECT 347.460 2.400 347.600 26.190 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 26.760 365.630 26.820 ;
        RECT 856.130 26.760 856.450 26.820 ;
        RECT 365.310 26.620 856.450 26.760 ;
        RECT 365.310 26.560 365.630 26.620 ;
        RECT 856.130 26.560 856.450 26.620 ;
      LAYER via ;
        RECT 365.340 26.560 365.600 26.820 ;
        RECT 856.160 26.560 856.420 26.820 ;
      LAYER met2 ;
        RECT 857.770 600.170 858.050 604.000 ;
        RECT 856.220 600.030 858.050 600.170 ;
        RECT 856.220 26.850 856.360 600.030 ;
        RECT 857.770 600.000 858.050 600.030 ;
        RECT 365.340 26.530 365.600 26.850 ;
        RECT 856.160 26.530 856.420 26.850 ;
        RECT 365.400 2.400 365.540 26.530 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.570 545.600 862.890 545.660 ;
        RECT 865.330 545.600 865.650 545.660 ;
        RECT 862.570 545.460 865.650 545.600 ;
        RECT 862.570 545.400 862.890 545.460 ;
        RECT 865.330 545.400 865.650 545.460 ;
        RECT 383.250 27.100 383.570 27.160 ;
        RECT 862.570 27.100 862.890 27.160 ;
        RECT 383.250 26.960 862.890 27.100 ;
        RECT 383.250 26.900 383.570 26.960 ;
        RECT 862.570 26.900 862.890 26.960 ;
      LAYER via ;
        RECT 862.600 545.400 862.860 545.660 ;
        RECT 865.360 545.400 865.620 545.660 ;
        RECT 383.280 26.900 383.540 27.160 ;
        RECT 862.600 26.900 862.860 27.160 ;
      LAYER met2 ;
        RECT 866.970 600.170 867.250 604.000 ;
        RECT 865.420 600.030 867.250 600.170 ;
        RECT 865.420 545.690 865.560 600.030 ;
        RECT 866.970 600.000 867.250 600.030 ;
        RECT 862.600 545.370 862.860 545.690 ;
        RECT 865.360 545.370 865.620 545.690 ;
        RECT 862.660 27.190 862.800 545.370 ;
        RECT 383.280 26.870 383.540 27.190 ;
        RECT 862.600 26.870 862.860 27.190 ;
        RECT 383.340 2.400 383.480 26.870 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 27.440 401.510 27.500 ;
        RECT 877.290 27.440 877.610 27.500 ;
        RECT 401.190 27.300 877.610 27.440 ;
        RECT 401.190 27.240 401.510 27.300 ;
        RECT 877.290 27.240 877.610 27.300 ;
      LAYER via ;
        RECT 401.220 27.240 401.480 27.500 ;
        RECT 877.320 27.240 877.580 27.500 ;
      LAYER met2 ;
        RECT 876.170 600.170 876.450 604.000 ;
        RECT 876.170 600.030 877.520 600.170 ;
        RECT 876.170 600.000 876.450 600.030 ;
        RECT 877.380 27.530 877.520 600.030 ;
        RECT 401.220 27.210 401.480 27.530 ;
        RECT 877.320 27.210 877.580 27.530 ;
        RECT 401.280 2.400 401.420 27.210 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 697.430 569.400 697.750 569.460 ;
        RECT 700.190 569.400 700.510 569.460 ;
        RECT 697.430 569.260 700.510 569.400 ;
        RECT 697.430 569.200 697.750 569.260 ;
        RECT 700.190 569.200 700.510 569.260 ;
        RECT 62.170 24.040 62.490 24.100 ;
        RECT 697.430 24.040 697.750 24.100 ;
        RECT 62.170 23.900 697.750 24.040 ;
        RECT 62.170 23.840 62.490 23.900 ;
        RECT 697.430 23.840 697.750 23.900 ;
      LAYER via ;
        RECT 697.460 569.200 697.720 569.460 ;
        RECT 700.220 569.200 700.480 569.460 ;
        RECT 62.200 23.840 62.460 24.100 ;
        RECT 697.460 23.840 697.720 24.100 ;
      LAYER met2 ;
        RECT 701.830 600.170 702.110 604.000 ;
        RECT 700.280 600.030 702.110 600.170 ;
        RECT 700.280 569.490 700.420 600.030 ;
        RECT 701.830 600.000 702.110 600.030 ;
        RECT 697.460 569.170 697.720 569.490 ;
        RECT 700.220 569.170 700.480 569.490 ;
        RECT 697.520 24.130 697.660 569.170 ;
        RECT 62.200 23.810 62.460 24.130 ;
        RECT 697.460 23.810 697.720 24.130 ;
        RECT 62.260 2.400 62.400 23.810 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 23.700 419.450 23.760 ;
        RECT 883.730 23.700 884.050 23.760 ;
        RECT 419.130 23.560 884.050 23.700 ;
        RECT 419.130 23.500 419.450 23.560 ;
        RECT 883.730 23.500 884.050 23.560 ;
      LAYER via ;
        RECT 419.160 23.500 419.420 23.760 ;
        RECT 883.760 23.500 884.020 23.760 ;
      LAYER met2 ;
        RECT 885.370 600.170 885.650 604.000 ;
        RECT 883.820 600.030 885.650 600.170 ;
        RECT 883.820 23.790 883.960 600.030 ;
        RECT 885.370 600.000 885.650 600.030 ;
        RECT 419.160 23.470 419.420 23.790 ;
        RECT 883.760 23.470 884.020 23.790 ;
        RECT 419.220 2.400 419.360 23.470 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 890.170 569.400 890.490 569.460 ;
        RECT 892.930 569.400 893.250 569.460 ;
        RECT 890.170 569.260 893.250 569.400 ;
        RECT 890.170 569.200 890.490 569.260 ;
        RECT 892.930 569.200 893.250 569.260 ;
        RECT 436.610 23.020 436.930 23.080 ;
        RECT 890.170 23.020 890.490 23.080 ;
        RECT 436.610 22.880 890.490 23.020 ;
        RECT 436.610 22.820 436.930 22.880 ;
        RECT 890.170 22.820 890.490 22.880 ;
      LAYER via ;
        RECT 890.200 569.200 890.460 569.460 ;
        RECT 892.960 569.200 893.220 569.460 ;
        RECT 436.640 22.820 436.900 23.080 ;
        RECT 890.200 22.820 890.460 23.080 ;
      LAYER met2 ;
        RECT 894.570 600.170 894.850 604.000 ;
        RECT 893.020 600.030 894.850 600.170 ;
        RECT 893.020 569.490 893.160 600.030 ;
        RECT 894.570 600.000 894.850 600.030 ;
        RECT 890.200 569.170 890.460 569.490 ;
        RECT 892.960 569.170 893.220 569.490 ;
        RECT 890.260 23.110 890.400 569.170 ;
        RECT 436.640 22.790 436.900 23.110 ;
        RECT 890.200 22.790 890.460 23.110 ;
        RECT 436.700 2.400 436.840 22.790 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 23.360 454.870 23.420 ;
        RECT 904.430 23.360 904.750 23.420 ;
        RECT 454.550 23.220 904.750 23.360 ;
        RECT 454.550 23.160 454.870 23.220 ;
        RECT 904.430 23.160 904.750 23.220 ;
      LAYER via ;
        RECT 454.580 23.160 454.840 23.420 ;
        RECT 904.460 23.160 904.720 23.420 ;
      LAYER met2 ;
        RECT 903.770 600.170 904.050 604.000 ;
        RECT 903.770 600.030 904.660 600.170 ;
        RECT 903.770 600.000 904.050 600.030 ;
        RECT 904.520 23.450 904.660 600.030 ;
        RECT 454.580 23.130 454.840 23.450 ;
        RECT 904.460 23.130 904.720 23.450 ;
        RECT 454.640 2.400 454.780 23.130 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 48.180 472.810 48.240 ;
        RECT 911.330 48.180 911.650 48.240 ;
        RECT 472.490 48.040 911.650 48.180 ;
        RECT 472.490 47.980 472.810 48.040 ;
        RECT 911.330 47.980 911.650 48.040 ;
      LAYER via ;
        RECT 472.520 47.980 472.780 48.240 ;
        RECT 911.360 47.980 911.620 48.240 ;
      LAYER met2 ;
        RECT 912.970 600.170 913.250 604.000 ;
        RECT 911.420 600.030 913.250 600.170 ;
        RECT 911.420 48.270 911.560 600.030 ;
        RECT 912.970 600.000 913.250 600.030 ;
        RECT 472.520 47.950 472.780 48.270 ;
        RECT 911.360 47.950 911.620 48.270 ;
        RECT 472.580 2.400 472.720 47.950 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 918.230 386.480 918.550 386.540 ;
        RECT 918.690 386.480 919.010 386.540 ;
        RECT 918.230 386.340 919.010 386.480 ;
        RECT 918.230 386.280 918.550 386.340 ;
        RECT 918.690 386.280 919.010 386.340 ;
        RECT 918.690 283.120 919.010 283.180 ;
        RECT 919.150 283.120 919.470 283.180 ;
        RECT 918.690 282.980 919.470 283.120 ;
        RECT 918.690 282.920 919.010 282.980 ;
        RECT 919.150 282.920 919.470 282.980 ;
        RECT 916.850 138.280 917.170 138.340 ;
        RECT 919.150 138.280 919.470 138.340 ;
        RECT 916.850 138.140 919.470 138.280 ;
        RECT 916.850 138.080 917.170 138.140 ;
        RECT 919.150 138.080 919.470 138.140 ;
        RECT 918.690 96.460 919.010 96.520 ;
        RECT 919.610 96.460 919.930 96.520 ;
        RECT 918.690 96.320 919.930 96.460 ;
        RECT 918.690 96.260 919.010 96.320 ;
        RECT 919.610 96.260 919.930 96.320 ;
        RECT 918.230 48.180 918.550 48.240 ;
        RECT 919.150 48.180 919.470 48.240 ;
        RECT 918.230 48.040 919.470 48.180 ;
        RECT 918.230 47.980 918.550 48.040 ;
        RECT 919.150 47.980 919.470 48.040 ;
        RECT 490.430 44.440 490.750 44.500 ;
        RECT 919.150 44.440 919.470 44.500 ;
        RECT 490.430 44.300 919.470 44.440 ;
        RECT 490.430 44.240 490.750 44.300 ;
        RECT 919.150 44.240 919.470 44.300 ;
      LAYER via ;
        RECT 918.260 386.280 918.520 386.540 ;
        RECT 918.720 386.280 918.980 386.540 ;
        RECT 918.720 282.920 918.980 283.180 ;
        RECT 919.180 282.920 919.440 283.180 ;
        RECT 916.880 138.080 917.140 138.340 ;
        RECT 919.180 138.080 919.440 138.340 ;
        RECT 918.720 96.260 918.980 96.520 ;
        RECT 919.640 96.260 919.900 96.520 ;
        RECT 918.260 47.980 918.520 48.240 ;
        RECT 919.180 47.980 919.440 48.240 ;
        RECT 490.460 44.240 490.720 44.500 ;
        RECT 919.180 44.240 919.440 44.500 ;
      LAYER met2 ;
        RECT 922.170 600.170 922.450 604.000 ;
        RECT 920.160 600.030 922.450 600.170 ;
        RECT 920.160 596.770 920.300 600.030 ;
        RECT 922.170 600.000 922.450 600.030 ;
        RECT 918.780 596.630 920.300 596.770 ;
        RECT 918.780 545.770 918.920 596.630 ;
        RECT 918.780 545.630 919.380 545.770 ;
        RECT 919.240 545.090 919.380 545.630 ;
        RECT 918.780 544.950 919.380 545.090 ;
        RECT 918.780 458.730 918.920 544.950 ;
        RECT 918.320 458.590 918.920 458.730 ;
        RECT 918.320 386.570 918.460 458.590 ;
        RECT 918.260 386.250 918.520 386.570 ;
        RECT 918.720 386.250 918.980 386.570 ;
        RECT 918.780 283.210 918.920 386.250 ;
        RECT 918.720 282.890 918.980 283.210 ;
        RECT 919.180 282.890 919.440 283.210 ;
        RECT 919.240 241.810 919.380 282.890 ;
        RECT 919.240 241.670 919.840 241.810 ;
        RECT 919.700 241.130 919.840 241.670 ;
        RECT 918.780 240.990 919.840 241.130 ;
        RECT 916.870 185.795 917.150 186.165 ;
        RECT 918.250 186.050 918.530 186.165 ;
        RECT 918.780 186.050 918.920 240.990 ;
        RECT 918.250 185.910 918.920 186.050 ;
        RECT 918.250 185.795 918.530 185.910 ;
        RECT 916.940 138.370 917.080 185.795 ;
        RECT 916.880 138.050 917.140 138.370 ;
        RECT 919.180 138.050 919.440 138.370 ;
        RECT 919.240 96.970 919.380 138.050 ;
        RECT 918.780 96.830 919.380 96.970 ;
        RECT 918.780 96.550 918.920 96.830 ;
        RECT 918.720 96.230 918.980 96.550 ;
        RECT 919.640 96.230 919.900 96.550 ;
        RECT 919.700 49.485 919.840 96.230 ;
        RECT 919.630 49.115 919.910 49.485 ;
        RECT 918.250 48.435 918.530 48.805 ;
        RECT 918.320 48.270 918.460 48.435 ;
        RECT 918.260 47.950 918.520 48.270 ;
        RECT 919.180 47.950 919.440 48.270 ;
        RECT 919.240 44.530 919.380 47.950 ;
        RECT 490.460 44.210 490.720 44.530 ;
        RECT 919.180 44.210 919.440 44.530 ;
        RECT 490.520 2.400 490.660 44.210 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 916.870 185.840 917.150 186.120 ;
        RECT 918.250 185.840 918.530 186.120 ;
        RECT 919.630 49.160 919.910 49.440 ;
        RECT 918.250 48.480 918.530 48.760 ;
      LAYER met3 ;
        RECT 916.845 186.130 917.175 186.145 ;
        RECT 918.225 186.130 918.555 186.145 ;
        RECT 916.845 185.830 918.555 186.130 ;
        RECT 916.845 185.815 917.175 185.830 ;
        RECT 918.225 185.815 918.555 185.830 ;
        RECT 919.605 49.450 919.935 49.465 ;
        RECT 917.550 49.150 919.935 49.450 ;
        RECT 917.550 48.770 917.850 49.150 ;
        RECT 919.605 49.135 919.935 49.150 ;
        RECT 918.225 48.770 918.555 48.785 ;
        RECT 917.550 48.470 918.555 48.770 ;
        RECT 918.225 48.455 918.555 48.470 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 932.030 379.820 932.350 380.080 ;
        RECT 932.120 379.400 932.260 379.820 ;
        RECT 932.030 379.140 932.350 379.400 ;
        RECT 507.910 34.240 508.230 34.300 ;
        RECT 932.030 34.240 932.350 34.300 ;
        RECT 507.910 34.100 932.350 34.240 ;
        RECT 507.910 34.040 508.230 34.100 ;
        RECT 932.030 34.040 932.350 34.100 ;
      LAYER via ;
        RECT 932.060 379.820 932.320 380.080 ;
        RECT 932.060 379.140 932.320 379.400 ;
        RECT 507.940 34.040 508.200 34.300 ;
        RECT 932.060 34.040 932.320 34.300 ;
      LAYER met2 ;
        RECT 931.370 600.170 931.650 604.000 ;
        RECT 931.370 600.030 932.260 600.170 ;
        RECT 931.370 600.000 931.650 600.030 ;
        RECT 932.120 380.110 932.260 600.030 ;
        RECT 932.060 379.790 932.320 380.110 ;
        RECT 932.060 379.110 932.320 379.430 ;
        RECT 932.120 34.330 932.260 379.110 ;
        RECT 507.940 34.010 508.200 34.330 ;
        RECT 932.060 34.010 932.320 34.330 ;
        RECT 508.000 2.400 508.140 34.010 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 30.160 526.170 30.220 ;
        RECT 938.470 30.160 938.790 30.220 ;
        RECT 525.850 30.020 938.790 30.160 ;
        RECT 525.850 29.960 526.170 30.020 ;
        RECT 938.470 29.960 938.790 30.020 ;
      LAYER via ;
        RECT 525.880 29.960 526.140 30.220 ;
        RECT 938.500 29.960 938.760 30.220 ;
      LAYER met2 ;
        RECT 940.570 600.170 940.850 604.000 ;
        RECT 938.560 600.030 940.850 600.170 ;
        RECT 938.560 30.250 938.700 600.030 ;
        RECT 940.570 600.000 940.850 600.030 ;
        RECT 525.880 29.930 526.140 30.250 ;
        RECT 938.500 29.930 938.760 30.250 ;
        RECT 525.940 2.400 526.080 29.930 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 945.370 572.460 945.690 572.520 ;
        RECT 946.290 572.460 946.610 572.520 ;
        RECT 945.370 572.320 946.610 572.460 ;
        RECT 945.370 572.260 945.690 572.320 ;
        RECT 946.290 572.260 946.610 572.320 ;
        RECT 945.370 524.860 945.690 524.920 ;
        RECT 945.830 524.860 946.150 524.920 ;
        RECT 945.370 524.720 946.150 524.860 ;
        RECT 945.370 524.660 945.690 524.720 ;
        RECT 945.830 524.660 946.150 524.720 ;
        RECT 945.830 517.380 946.150 517.440 ;
        RECT 947.670 517.380 947.990 517.440 ;
        RECT 945.830 517.240 947.990 517.380 ;
        RECT 945.830 517.180 946.150 517.240 ;
        RECT 947.670 517.180 947.990 517.240 ;
        RECT 946.750 475.560 947.070 475.620 ;
        RECT 947.670 475.560 947.990 475.620 ;
        RECT 946.750 475.420 947.990 475.560 ;
        RECT 946.750 475.360 947.070 475.420 ;
        RECT 947.670 475.360 947.990 475.420 ;
        RECT 946.290 427.960 946.610 428.020 ;
        RECT 946.750 427.960 947.070 428.020 ;
        RECT 946.290 427.820 947.070 427.960 ;
        RECT 946.290 427.760 946.610 427.820 ;
        RECT 946.750 427.760 947.070 427.820 ;
        RECT 945.370 386.480 945.690 386.540 ;
        RECT 946.290 386.480 946.610 386.540 ;
        RECT 945.370 386.340 946.610 386.480 ;
        RECT 945.370 386.280 945.690 386.340 ;
        RECT 946.290 386.280 946.610 386.340 ;
        RECT 945.370 379.340 945.690 379.400 ;
        RECT 945.830 379.340 946.150 379.400 ;
        RECT 945.370 379.200 946.150 379.340 ;
        RECT 945.370 379.140 945.690 379.200 ;
        RECT 945.830 379.140 946.150 379.200 ;
        RECT 945.830 351.940 946.150 352.200 ;
        RECT 945.920 351.520 946.060 351.940 ;
        RECT 945.830 351.260 946.150 351.520 ;
        RECT 945.830 303.520 946.150 303.580 ;
        RECT 946.750 303.520 947.070 303.580 ;
        RECT 945.830 303.380 947.070 303.520 ;
        RECT 945.830 303.320 946.150 303.380 ;
        RECT 946.750 303.320 947.070 303.380 ;
        RECT 946.750 255.380 947.070 255.640 ;
        RECT 946.840 254.960 946.980 255.380 ;
        RECT 946.750 254.700 947.070 254.960 ;
        RECT 945.370 193.360 945.690 193.420 ;
        RECT 946.750 193.360 947.070 193.420 ;
        RECT 945.370 193.220 947.070 193.360 ;
        RECT 945.370 193.160 945.690 193.220 ;
        RECT 946.750 193.160 947.070 193.220 ;
        RECT 543.790 29.480 544.110 29.540 ;
        RECT 946.750 29.480 947.070 29.540 ;
        RECT 543.790 29.340 947.070 29.480 ;
        RECT 543.790 29.280 544.110 29.340 ;
        RECT 946.750 29.280 947.070 29.340 ;
      LAYER via ;
        RECT 945.400 572.260 945.660 572.520 ;
        RECT 946.320 572.260 946.580 572.520 ;
        RECT 945.400 524.660 945.660 524.920 ;
        RECT 945.860 524.660 946.120 524.920 ;
        RECT 945.860 517.180 946.120 517.440 ;
        RECT 947.700 517.180 947.960 517.440 ;
        RECT 946.780 475.360 947.040 475.620 ;
        RECT 947.700 475.360 947.960 475.620 ;
        RECT 946.320 427.760 946.580 428.020 ;
        RECT 946.780 427.760 947.040 428.020 ;
        RECT 945.400 386.280 945.660 386.540 ;
        RECT 946.320 386.280 946.580 386.540 ;
        RECT 945.400 379.140 945.660 379.400 ;
        RECT 945.860 379.140 946.120 379.400 ;
        RECT 945.860 351.940 946.120 352.200 ;
        RECT 945.860 351.260 946.120 351.520 ;
        RECT 945.860 303.320 946.120 303.580 ;
        RECT 946.780 303.320 947.040 303.580 ;
        RECT 946.780 255.380 947.040 255.640 ;
        RECT 946.780 254.700 947.040 254.960 ;
        RECT 945.400 193.160 945.660 193.420 ;
        RECT 946.780 193.160 947.040 193.420 ;
        RECT 543.820 29.280 544.080 29.540 ;
        RECT 946.780 29.280 947.040 29.540 ;
      LAYER met2 ;
        RECT 949.770 600.170 950.050 604.000 ;
        RECT 948.220 600.030 950.050 600.170 ;
        RECT 948.220 596.770 948.360 600.030 ;
        RECT 949.770 600.000 950.050 600.030 ;
        RECT 946.380 596.630 948.360 596.770 ;
        RECT 946.380 572.550 946.520 596.630 ;
        RECT 945.400 572.230 945.660 572.550 ;
        RECT 946.320 572.230 946.580 572.550 ;
        RECT 945.460 524.950 945.600 572.230 ;
        RECT 945.400 524.630 945.660 524.950 ;
        RECT 945.860 524.630 946.120 524.950 ;
        RECT 945.920 517.470 946.060 524.630 ;
        RECT 945.860 517.150 946.120 517.470 ;
        RECT 947.700 517.150 947.960 517.470 ;
        RECT 947.760 475.650 947.900 517.150 ;
        RECT 946.780 475.330 947.040 475.650 ;
        RECT 947.700 475.330 947.960 475.650 ;
        RECT 946.840 428.050 946.980 475.330 ;
        RECT 946.320 427.730 946.580 428.050 ;
        RECT 946.780 427.730 947.040 428.050 ;
        RECT 946.380 386.570 946.520 427.730 ;
        RECT 945.400 386.250 945.660 386.570 ;
        RECT 946.320 386.250 946.580 386.570 ;
        RECT 945.460 379.430 945.600 386.250 ;
        RECT 945.400 379.110 945.660 379.430 ;
        RECT 945.860 379.110 946.120 379.430 ;
        RECT 945.920 352.230 946.060 379.110 ;
        RECT 945.860 351.910 946.120 352.230 ;
        RECT 945.860 351.230 946.120 351.550 ;
        RECT 945.920 303.610 946.060 351.230 ;
        RECT 945.860 303.290 946.120 303.610 ;
        RECT 946.780 303.290 947.040 303.610 ;
        RECT 946.840 255.670 946.980 303.290 ;
        RECT 946.780 255.350 947.040 255.670 ;
        RECT 946.780 254.670 947.040 254.990 ;
        RECT 946.840 193.450 946.980 254.670 ;
        RECT 945.400 193.130 945.660 193.450 ;
        RECT 946.780 193.130 947.040 193.450 ;
        RECT 945.460 145.365 945.600 193.130 ;
        RECT 945.390 144.995 945.670 145.365 ;
        RECT 946.770 144.315 947.050 144.685 ;
        RECT 946.840 29.570 946.980 144.315 ;
        RECT 543.820 29.250 544.080 29.570 ;
        RECT 946.780 29.250 947.040 29.570 ;
        RECT 543.880 2.400 544.020 29.250 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 945.390 145.040 945.670 145.320 ;
        RECT 946.770 144.360 947.050 144.640 ;
      LAYER met3 ;
        RECT 945.365 145.330 945.695 145.345 ;
        RECT 945.365 145.030 946.370 145.330 ;
        RECT 945.365 145.015 945.695 145.030 ;
        RECT 946.070 144.650 946.370 145.030 ;
        RECT 946.745 144.650 947.075 144.665 ;
        RECT 946.070 144.350 947.075 144.650 ;
        RECT 946.745 144.335 947.075 144.350 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 29.140 562.050 29.200 ;
        RECT 959.630 29.140 959.950 29.200 ;
        RECT 561.730 29.000 959.950 29.140 ;
        RECT 561.730 28.940 562.050 29.000 ;
        RECT 959.630 28.940 959.950 29.000 ;
      LAYER via ;
        RECT 561.760 28.940 562.020 29.200 ;
        RECT 959.660 28.940 959.920 29.200 ;
      LAYER met2 ;
        RECT 958.970 600.170 959.250 604.000 ;
        RECT 958.970 600.030 959.860 600.170 ;
        RECT 958.970 600.000 959.250 600.030 ;
        RECT 959.720 29.230 959.860 600.030 ;
        RECT 561.760 28.910 562.020 29.230 ;
        RECT 959.660 28.910 959.920 29.230 ;
        RECT 561.820 2.400 561.960 28.910 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 580.130 28.800 580.450 28.860 ;
        RECT 966.070 28.800 966.390 28.860 ;
        RECT 580.130 28.660 966.390 28.800 ;
        RECT 580.130 28.600 580.450 28.660 ;
        RECT 966.070 28.600 966.390 28.660 ;
      LAYER via ;
        RECT 580.160 28.600 580.420 28.860 ;
        RECT 966.100 28.600 966.360 28.860 ;
      LAYER met2 ;
        RECT 968.170 600.170 968.450 604.000 ;
        RECT 966.160 600.030 968.450 600.170 ;
        RECT 966.160 28.890 966.300 600.030 ;
        RECT 968.170 600.000 968.450 600.030 ;
        RECT 580.160 28.570 580.420 28.890 ;
        RECT 966.100 28.570 966.360 28.890 ;
        RECT 580.220 14.690 580.360 28.570 ;
        RECT 579.760 14.550 580.360 14.690 ;
        RECT 579.760 2.400 579.900 14.550 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1901.710 2533.240 1902.030 2533.300 ;
        RECT 1903.090 2533.240 1903.410 2533.300 ;
        RECT 1901.710 2533.100 1903.410 2533.240 ;
        RECT 1901.710 2533.040 1902.030 2533.100 ;
        RECT 1903.090 2533.040 1903.410 2533.100 ;
        RECT 654.190 2501.960 654.510 2502.020 ;
        RECT 1903.090 2501.960 1903.410 2502.020 ;
        RECT 654.190 2501.820 1903.410 2501.960 ;
        RECT 654.190 2501.760 654.510 2501.820 ;
        RECT 1903.090 2501.760 1903.410 2501.820 ;
        RECT 654.190 595.580 654.510 595.640 ;
        RECT 711.230 595.580 711.550 595.640 ;
        RECT 712.610 595.580 712.930 595.640 ;
        RECT 654.190 595.440 712.930 595.580 ;
        RECT 654.190 595.380 654.510 595.440 ;
        RECT 711.230 595.380 711.550 595.440 ;
        RECT 712.610 595.380 712.930 595.440 ;
        RECT 86.090 24.380 86.410 24.440 ;
        RECT 711.230 24.380 711.550 24.440 ;
        RECT 86.090 24.240 711.550 24.380 ;
        RECT 86.090 24.180 86.410 24.240 ;
        RECT 711.230 24.180 711.550 24.240 ;
      LAYER via ;
        RECT 1901.740 2533.040 1902.000 2533.300 ;
        RECT 1903.120 2533.040 1903.380 2533.300 ;
        RECT 654.220 2501.760 654.480 2502.020 ;
        RECT 1903.120 2501.760 1903.380 2502.020 ;
        RECT 654.220 595.380 654.480 595.640 ;
        RECT 711.260 595.380 711.520 595.640 ;
        RECT 712.640 595.380 712.900 595.640 ;
        RECT 86.120 24.180 86.380 24.440 ;
        RECT 711.260 24.180 711.520 24.440 ;
      LAYER met2 ;
        RECT 1901.730 2705.195 1902.010 2705.565 ;
        RECT 1901.800 2533.330 1901.940 2705.195 ;
        RECT 1901.740 2533.010 1902.000 2533.330 ;
        RECT 1903.120 2533.010 1903.380 2533.330 ;
        RECT 1903.180 2502.050 1903.320 2533.010 ;
        RECT 654.220 2501.730 654.480 2502.050 ;
        RECT 1903.120 2501.730 1903.380 2502.050 ;
        RECT 654.280 595.670 654.420 2501.730 ;
        RECT 714.250 600.170 714.530 604.000 ;
        RECT 712.700 600.030 714.530 600.170 ;
        RECT 712.700 595.670 712.840 600.030 ;
        RECT 714.250 600.000 714.530 600.030 ;
        RECT 654.220 595.350 654.480 595.670 ;
        RECT 711.260 595.350 711.520 595.670 ;
        RECT 712.640 595.350 712.900 595.670 ;
        RECT 711.320 24.470 711.460 595.350 ;
        RECT 86.120 24.150 86.380 24.470 ;
        RECT 711.260 24.150 711.520 24.470 ;
        RECT 86.180 2.400 86.320 24.150 ;
        RECT 85.970 -4.800 86.530 2.400 ;
      LAYER via2 ;
        RECT 1901.730 2705.240 1902.010 2705.520 ;
      LAYER met3 ;
        RECT 1885.335 2707.080 1889.335 2707.360 ;
        RECT 1885.335 2706.760 1889.370 2707.080 ;
        RECT 1889.070 2705.530 1889.370 2706.760 ;
        RECT 1901.705 2705.530 1902.035 2705.545 ;
        RECT 1889.070 2705.230 1902.035 2705.530 ;
        RECT 1901.705 2705.215 1902.035 2705.230 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.970 569.400 973.290 569.460 ;
        RECT 975.730 569.400 976.050 569.460 ;
        RECT 972.970 569.260 976.050 569.400 ;
        RECT 972.970 569.200 973.290 569.260 ;
        RECT 975.730 569.200 976.050 569.260 ;
        RECT 597.150 28.460 597.470 28.520 ;
        RECT 973.430 28.460 973.750 28.520 ;
        RECT 597.150 28.320 973.750 28.460 ;
        RECT 597.150 28.260 597.470 28.320 ;
        RECT 973.430 28.260 973.750 28.320 ;
      LAYER via ;
        RECT 973.000 569.200 973.260 569.460 ;
        RECT 975.760 569.200 976.020 569.460 ;
        RECT 597.180 28.260 597.440 28.520 ;
        RECT 973.460 28.260 973.720 28.520 ;
      LAYER met2 ;
        RECT 977.370 600.170 977.650 604.000 ;
        RECT 975.820 600.030 977.650 600.170 ;
        RECT 975.820 569.490 975.960 600.030 ;
        RECT 977.370 600.000 977.650 600.030 ;
        RECT 973.000 569.170 973.260 569.490 ;
        RECT 975.760 569.170 976.020 569.490 ;
        RECT 973.060 33.730 973.200 569.170 ;
        RECT 973.060 33.590 973.660 33.730 ;
        RECT 973.520 28.550 973.660 33.590 ;
        RECT 597.180 28.230 597.440 28.550 ;
        RECT 973.460 28.230 973.720 28.550 ;
        RECT 597.240 2.400 597.380 28.230 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 28.120 615.410 28.180 ;
        RECT 987.690 28.120 988.010 28.180 ;
        RECT 615.090 27.980 988.010 28.120 ;
        RECT 615.090 27.920 615.410 27.980 ;
        RECT 987.690 27.920 988.010 27.980 ;
      LAYER via ;
        RECT 615.120 27.920 615.380 28.180 ;
        RECT 987.720 27.920 987.980 28.180 ;
      LAYER met2 ;
        RECT 986.570 600.170 986.850 604.000 ;
        RECT 986.570 600.030 987.920 600.170 ;
        RECT 986.570 600.000 986.850 600.030 ;
        RECT 987.780 28.210 987.920 600.030 ;
        RECT 615.120 27.890 615.380 28.210 ;
        RECT 987.720 27.890 987.980 28.210 ;
        RECT 615.180 2.400 615.320 27.890 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 647.290 2815.440 647.610 2815.500 ;
        RECT 1483.570 2815.440 1483.890 2815.500 ;
        RECT 647.290 2815.300 1483.890 2815.440 ;
        RECT 647.290 2815.240 647.610 2815.300 ;
        RECT 1483.570 2815.240 1483.890 2815.300 ;
        RECT 647.290 594.560 647.610 594.620 ;
        RECT 725.030 594.560 725.350 594.620 ;
        RECT 647.290 594.420 725.350 594.560 ;
        RECT 647.290 594.360 647.610 594.420 ;
        RECT 725.030 594.360 725.350 594.420 ;
        RECT 724.570 579.600 724.890 579.660 ;
        RECT 726.410 579.600 726.730 579.660 ;
        RECT 724.570 579.460 726.730 579.600 ;
        RECT 724.570 579.400 724.890 579.460 ;
        RECT 726.410 579.400 726.730 579.460 ;
        RECT 724.110 427.620 724.430 427.680 ;
        RECT 725.490 427.620 725.810 427.680 ;
        RECT 724.110 427.480 725.810 427.620 ;
        RECT 724.110 427.420 724.430 427.480 ;
        RECT 725.490 427.420 725.810 427.480 ;
        RECT 724.110 379.680 724.430 379.740 ;
        RECT 725.030 379.680 725.350 379.740 ;
        RECT 724.110 379.540 725.350 379.680 ;
        RECT 724.110 379.480 724.430 379.540 ;
        RECT 725.030 379.480 725.350 379.540 ;
        RECT 724.110 331.400 724.430 331.460 ;
        RECT 725.490 331.400 725.810 331.460 ;
        RECT 724.110 331.260 725.810 331.400 ;
        RECT 724.110 331.200 724.430 331.260 ;
        RECT 725.490 331.200 725.810 331.260 ;
        RECT 725.490 283.120 725.810 283.180 ;
        RECT 725.950 283.120 726.270 283.180 ;
        RECT 725.490 282.980 726.270 283.120 ;
        RECT 725.490 282.920 725.810 282.980 ;
        RECT 725.950 282.920 726.270 282.980 ;
        RECT 725.950 255.580 726.270 255.640 ;
        RECT 725.580 255.440 726.270 255.580 ;
        RECT 725.580 255.300 725.720 255.440 ;
        RECT 725.950 255.380 726.270 255.440 ;
        RECT 725.490 255.040 725.810 255.300 ;
        RECT 725.030 96.460 725.350 96.520 ;
        RECT 725.950 96.460 726.270 96.520 ;
        RECT 725.030 96.320 726.270 96.460 ;
        RECT 725.030 96.260 725.350 96.320 ;
        RECT 725.950 96.260 726.270 96.320 ;
        RECT 109.550 24.720 109.870 24.780 ;
        RECT 725.030 24.720 725.350 24.780 ;
        RECT 109.550 24.580 725.350 24.720 ;
        RECT 109.550 24.520 109.870 24.580 ;
        RECT 725.030 24.520 725.350 24.580 ;
      LAYER via ;
        RECT 647.320 2815.240 647.580 2815.500 ;
        RECT 1483.600 2815.240 1483.860 2815.500 ;
        RECT 647.320 594.360 647.580 594.620 ;
        RECT 725.060 594.360 725.320 594.620 ;
        RECT 724.600 579.400 724.860 579.660 ;
        RECT 726.440 579.400 726.700 579.660 ;
        RECT 724.140 427.420 724.400 427.680 ;
        RECT 725.520 427.420 725.780 427.680 ;
        RECT 724.140 379.480 724.400 379.740 ;
        RECT 725.060 379.480 725.320 379.740 ;
        RECT 724.140 331.200 724.400 331.460 ;
        RECT 725.520 331.200 725.780 331.460 ;
        RECT 725.520 282.920 725.780 283.180 ;
        RECT 725.980 282.920 726.240 283.180 ;
        RECT 725.980 255.380 726.240 255.640 ;
        RECT 725.520 255.040 725.780 255.300 ;
        RECT 725.060 96.260 725.320 96.520 ;
        RECT 725.980 96.260 726.240 96.520 ;
        RECT 109.580 24.520 109.840 24.780 ;
        RECT 725.060 24.520 725.320 24.780 ;
      LAYER met2 ;
        RECT 1483.590 2816.035 1483.870 2816.405 ;
        RECT 1483.660 2815.530 1483.800 2816.035 ;
        RECT 647.320 2815.210 647.580 2815.530 ;
        RECT 1483.600 2815.210 1483.860 2815.530 ;
        RECT 647.380 594.650 647.520 2815.210 ;
        RECT 726.210 600.170 726.490 604.000 ;
        RECT 725.120 600.030 726.490 600.170 ;
        RECT 725.120 594.650 725.260 600.030 ;
        RECT 726.210 600.000 726.490 600.030 ;
        RECT 647.320 594.330 647.580 594.650 ;
        RECT 725.060 594.330 725.320 594.650 ;
        RECT 725.120 579.770 725.260 594.330 ;
        RECT 724.660 579.690 725.260 579.770 ;
        RECT 724.600 579.630 725.260 579.690 ;
        RECT 724.600 579.370 724.860 579.630 ;
        RECT 726.440 579.370 726.700 579.690 ;
        RECT 724.660 579.215 724.800 579.370 ;
        RECT 726.500 531.605 726.640 579.370 ;
        RECT 725.510 531.235 725.790 531.605 ;
        RECT 726.430 531.235 726.710 531.605 ;
        RECT 725.580 427.710 725.720 531.235 ;
        RECT 724.140 427.390 724.400 427.710 ;
        RECT 725.520 427.390 725.780 427.710 ;
        RECT 724.200 379.770 724.340 427.390 ;
        RECT 724.140 379.450 724.400 379.770 ;
        RECT 725.060 379.450 725.320 379.770 ;
        RECT 725.120 379.285 725.260 379.450 ;
        RECT 724.130 378.915 724.410 379.285 ;
        RECT 725.050 378.915 725.330 379.285 ;
        RECT 724.200 331.490 724.340 378.915 ;
        RECT 724.140 331.170 724.400 331.490 ;
        RECT 725.520 331.170 725.780 331.490 ;
        RECT 725.580 331.005 725.720 331.170 ;
        RECT 725.510 330.635 725.790 331.005 ;
        RECT 725.970 329.955 726.250 330.325 ;
        RECT 726.040 283.210 726.180 329.955 ;
        RECT 725.520 282.890 725.780 283.210 ;
        RECT 725.980 282.890 726.240 283.210 ;
        RECT 725.580 269.010 725.720 282.890 ;
        RECT 725.580 268.870 726.180 269.010 ;
        RECT 726.040 255.670 726.180 268.870 ;
        RECT 725.980 255.350 726.240 255.670 ;
        RECT 725.520 255.010 725.780 255.330 ;
        RECT 725.580 207.810 725.720 255.010 ;
        RECT 724.660 207.670 725.720 207.810 ;
        RECT 724.660 179.930 724.800 207.670 ;
        RECT 724.660 179.790 725.720 179.930 ;
        RECT 725.580 179.250 725.720 179.790 ;
        RECT 724.200 179.110 725.720 179.250 ;
        RECT 724.200 155.450 724.340 179.110 ;
        RECT 724.200 155.310 724.800 155.450 ;
        RECT 724.660 96.970 724.800 155.310 ;
        RECT 724.660 96.830 725.260 96.970 ;
        RECT 725.120 96.550 725.260 96.830 ;
        RECT 725.060 96.230 725.320 96.550 ;
        RECT 725.980 96.230 726.240 96.550 ;
        RECT 726.040 60.930 726.180 96.230 ;
        RECT 725.120 60.790 726.180 60.930 ;
        RECT 725.120 24.810 725.260 60.790 ;
        RECT 109.580 24.490 109.840 24.810 ;
        RECT 725.060 24.490 725.320 24.810 ;
        RECT 109.640 2.400 109.780 24.490 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 1483.590 2816.080 1483.870 2816.360 ;
        RECT 725.510 531.280 725.790 531.560 ;
        RECT 726.430 531.280 726.710 531.560 ;
        RECT 724.130 378.960 724.410 379.240 ;
        RECT 725.050 378.960 725.330 379.240 ;
        RECT 725.510 330.680 725.790 330.960 ;
        RECT 725.970 330.000 726.250 330.280 ;
      LAYER met3 ;
        RECT 1500.000 2818.600 1504.000 2818.880 ;
        RECT 1499.910 2818.280 1504.000 2818.600 ;
        RECT 1483.565 2816.370 1483.895 2816.385 ;
        RECT 1499.910 2816.370 1500.210 2818.280 ;
        RECT 1483.565 2816.070 1500.210 2816.370 ;
        RECT 1483.565 2816.055 1483.895 2816.070 ;
        RECT 725.485 531.570 725.815 531.585 ;
        RECT 726.405 531.570 726.735 531.585 ;
        RECT 725.485 531.270 726.735 531.570 ;
        RECT 725.485 531.255 725.815 531.270 ;
        RECT 726.405 531.255 726.735 531.270 ;
        RECT 724.105 379.250 724.435 379.265 ;
        RECT 725.025 379.250 725.355 379.265 ;
        RECT 724.105 378.950 725.355 379.250 ;
        RECT 724.105 378.935 724.435 378.950 ;
        RECT 725.025 378.935 725.355 378.950 ;
        RECT 725.485 330.970 725.815 330.985 ;
        RECT 725.485 330.670 726.490 330.970 ;
        RECT 725.485 330.655 725.815 330.670 ;
        RECT 726.190 330.305 726.490 330.670 ;
        RECT 725.945 329.990 726.490 330.305 ;
        RECT 725.945 329.975 726.275 329.990 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 655.110 2916.420 655.430 2916.480 ;
        RECT 1747.610 2916.420 1747.930 2916.480 ;
        RECT 655.110 2916.280 1747.930 2916.420 ;
        RECT 655.110 2916.220 655.430 2916.280 ;
        RECT 1747.610 2916.220 1747.930 2916.280 ;
        RECT 655.110 722.200 655.430 722.460 ;
        RECT 655.200 720.760 655.340 722.200 ;
        RECT 655.110 720.500 655.430 720.760 ;
        RECT 655.110 594.220 655.430 594.280 ;
        RECT 738.830 594.220 739.150 594.280 ;
        RECT 655.110 594.080 739.150 594.220 ;
        RECT 655.110 594.020 655.430 594.080 ;
        RECT 738.830 594.020 739.150 594.080 ;
        RECT 133.470 25.060 133.790 25.120 ;
        RECT 738.830 25.060 739.150 25.120 ;
        RECT 133.470 24.920 739.150 25.060 ;
        RECT 133.470 24.860 133.790 24.920 ;
        RECT 738.830 24.860 739.150 24.920 ;
      LAYER via ;
        RECT 655.140 2916.220 655.400 2916.480 ;
        RECT 1747.640 2916.220 1747.900 2916.480 ;
        RECT 655.140 722.200 655.400 722.460 ;
        RECT 655.140 720.500 655.400 720.760 ;
        RECT 655.140 594.020 655.400 594.280 ;
        RECT 738.860 594.020 739.120 594.280 ;
        RECT 133.500 24.860 133.760 25.120 ;
        RECT 738.860 24.860 739.120 25.120 ;
      LAYER met2 ;
        RECT 655.140 2916.190 655.400 2916.510 ;
        RECT 1747.640 2916.190 1747.900 2916.510 ;
        RECT 655.200 722.490 655.340 2916.190 ;
        RECT 1747.700 2900.055 1747.840 2916.190 ;
        RECT 1747.570 2896.055 1747.850 2900.055 ;
        RECT 655.140 722.170 655.400 722.490 ;
        RECT 655.140 720.470 655.400 720.790 ;
        RECT 655.200 594.310 655.340 720.470 ;
        RECT 738.630 600.000 738.910 604.000 ;
        RECT 738.690 598.810 738.830 600.000 ;
        RECT 738.690 598.670 739.060 598.810 ;
        RECT 738.920 594.310 739.060 598.670 ;
        RECT 655.140 593.990 655.400 594.310 ;
        RECT 738.860 593.990 739.120 594.310 ;
        RECT 738.920 25.150 739.060 593.990 ;
        RECT 133.500 24.830 133.760 25.150 ;
        RECT 738.860 24.830 739.120 25.150 ;
        RECT 133.560 2.400 133.700 24.830 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 646.830 2502.300 647.150 2502.360 ;
        RECT 1886.990 2502.300 1887.310 2502.360 ;
        RECT 646.830 2502.160 1887.310 2502.300 ;
        RECT 646.830 2502.100 647.150 2502.160 ;
        RECT 1886.990 2502.100 1887.310 2502.160 ;
        RECT 646.830 593.880 647.150 593.940 ;
        RECT 745.270 593.880 745.590 593.940 ;
        RECT 646.830 593.740 745.590 593.880 ;
        RECT 646.830 593.680 647.150 593.740 ;
        RECT 745.270 593.680 745.590 593.740 ;
        RECT 151.410 25.400 151.730 25.460 ;
        RECT 745.270 25.400 745.590 25.460 ;
        RECT 151.410 25.260 745.590 25.400 ;
        RECT 151.410 25.200 151.730 25.260 ;
        RECT 745.270 25.200 745.590 25.260 ;
      LAYER via ;
        RECT 646.860 2502.100 647.120 2502.360 ;
        RECT 1887.020 2502.100 1887.280 2502.360 ;
        RECT 646.860 593.680 647.120 593.940 ;
        RECT 745.300 593.680 745.560 593.940 ;
        RECT 151.440 25.200 151.700 25.460 ;
        RECT 745.300 25.200 745.560 25.460 ;
      LAYER met2 ;
        RECT 1887.010 2860.235 1887.290 2860.605 ;
        RECT 1887.080 2502.390 1887.220 2860.235 ;
        RECT 646.860 2502.070 647.120 2502.390 ;
        RECT 1887.020 2502.070 1887.280 2502.390 ;
        RECT 646.920 593.970 647.060 2502.070 ;
        RECT 747.830 600.170 748.110 604.000 ;
        RECT 745.360 600.030 748.110 600.170 ;
        RECT 745.360 593.970 745.500 600.030 ;
        RECT 747.830 600.000 748.110 600.030 ;
        RECT 646.860 593.650 647.120 593.970 ;
        RECT 745.300 593.650 745.560 593.970 ;
        RECT 745.360 25.490 745.500 593.650 ;
        RECT 151.440 25.170 151.700 25.490 ;
        RECT 745.300 25.170 745.560 25.490 ;
        RECT 151.500 2.400 151.640 25.170 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 1887.010 2860.280 1887.290 2860.560 ;
      LAYER met3 ;
        RECT 1885.335 2863.160 1889.335 2863.760 ;
        RECT 1887.230 2860.585 1887.530 2863.160 ;
        RECT 1886.985 2860.270 1887.530 2860.585 ;
        RECT 1886.985 2860.255 1887.315 2860.270 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 753.550 476.240 753.870 476.300 ;
        RECT 754.930 476.240 755.250 476.300 ;
        RECT 753.550 476.100 755.250 476.240 ;
        RECT 753.550 476.040 753.870 476.100 ;
        RECT 754.930 476.040 755.250 476.100 ;
        RECT 752.630 458.900 752.950 458.960 ;
        RECT 753.550 458.900 753.870 458.960 ;
        RECT 752.630 458.760 753.870 458.900 ;
        RECT 752.630 458.700 752.950 458.760 ;
        RECT 753.550 458.700 753.870 458.760 ;
        RECT 752.630 144.740 752.950 144.800 ;
        RECT 753.090 144.740 753.410 144.800 ;
        RECT 752.630 144.600 753.410 144.740 ;
        RECT 752.630 144.540 752.950 144.600 ;
        RECT 753.090 144.540 753.410 144.600 ;
        RECT 169.350 45.800 169.670 45.860 ;
        RECT 753.090 45.800 753.410 45.860 ;
        RECT 169.350 45.660 753.410 45.800 ;
        RECT 169.350 45.600 169.670 45.660 ;
        RECT 753.090 45.600 753.410 45.660 ;
      LAYER via ;
        RECT 753.580 476.040 753.840 476.300 ;
        RECT 754.960 476.040 755.220 476.300 ;
        RECT 752.660 458.700 752.920 458.960 ;
        RECT 753.580 458.700 753.840 458.960 ;
        RECT 752.660 144.540 752.920 144.800 ;
        RECT 753.120 144.540 753.380 144.800 ;
        RECT 169.380 45.600 169.640 45.860 ;
        RECT 753.120 45.600 753.380 45.860 ;
      LAYER met2 ;
        RECT 757.030 601.530 757.310 604.000 ;
        RECT 755.480 601.390 757.310 601.530 ;
        RECT 755.480 579.770 755.620 601.390 ;
        RECT 757.030 600.000 757.310 601.390 ;
        RECT 755.020 579.630 755.620 579.770 ;
        RECT 755.020 476.330 755.160 579.630 ;
        RECT 753.580 476.010 753.840 476.330 ;
        RECT 754.960 476.010 755.220 476.330 ;
        RECT 753.640 458.990 753.780 476.010 ;
        RECT 752.660 458.670 752.920 458.990 ;
        RECT 753.580 458.670 753.840 458.990 ;
        RECT 752.720 144.830 752.860 458.670 ;
        RECT 752.660 144.510 752.920 144.830 ;
        RECT 753.120 144.510 753.380 144.830 ;
        RECT 753.180 45.890 753.320 144.510 ;
        RECT 169.380 45.570 169.640 45.890 ;
        RECT 753.120 45.570 753.380 45.890 ;
        RECT 169.440 2.400 169.580 45.570 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 25.740 187.150 25.800 ;
        RECT 766.890 25.740 767.210 25.800 ;
        RECT 186.830 25.600 767.210 25.740 ;
        RECT 186.830 25.540 187.150 25.600 ;
        RECT 766.890 25.540 767.210 25.600 ;
      LAYER via ;
        RECT 186.860 25.540 187.120 25.800 ;
        RECT 766.920 25.540 767.180 25.800 ;
      LAYER met2 ;
        RECT 766.230 600.170 766.510 604.000 ;
        RECT 766.230 600.030 767.120 600.170 ;
        RECT 766.230 600.000 766.510 600.030 ;
        RECT 766.980 25.830 767.120 600.030 ;
        RECT 186.860 25.510 187.120 25.830 ;
        RECT 766.920 25.510 767.180 25.830 ;
        RECT 186.920 2.400 187.060 25.510 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 46.140 205.090 46.200 ;
        RECT 772.870 46.140 773.190 46.200 ;
        RECT 204.770 46.000 773.190 46.140 ;
        RECT 204.770 45.940 205.090 46.000 ;
        RECT 772.870 45.940 773.190 46.000 ;
      LAYER via ;
        RECT 204.800 45.940 205.060 46.200 ;
        RECT 772.900 45.940 773.160 46.200 ;
      LAYER met2 ;
        RECT 775.430 600.170 775.710 604.000 ;
        RECT 772.960 600.030 775.710 600.170 ;
        RECT 772.960 46.230 773.100 600.030 ;
        RECT 775.430 600.000 775.710 600.030 ;
        RECT 204.800 45.910 205.060 46.230 ;
        RECT 772.900 45.910 773.160 46.230 ;
        RECT 204.860 2.400 205.000 45.910 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 780.690 531.320 781.010 531.380 ;
        RECT 782.530 531.320 782.850 531.380 ;
        RECT 780.690 531.180 782.850 531.320 ;
        RECT 780.690 531.120 781.010 531.180 ;
        RECT 782.530 531.120 782.850 531.180 ;
        RECT 780.230 144.740 780.550 144.800 ;
        RECT 780.690 144.740 781.010 144.800 ;
        RECT 780.230 144.600 781.010 144.740 ;
        RECT 780.230 144.540 780.550 144.600 ;
        RECT 780.690 144.540 781.010 144.600 ;
        RECT 222.710 32.200 223.030 32.260 ;
        RECT 780.690 32.200 781.010 32.260 ;
        RECT 222.710 32.060 781.010 32.200 ;
        RECT 222.710 32.000 223.030 32.060 ;
        RECT 780.690 32.000 781.010 32.060 ;
      LAYER via ;
        RECT 780.720 531.120 780.980 531.380 ;
        RECT 782.560 531.120 782.820 531.380 ;
        RECT 780.260 144.540 780.520 144.800 ;
        RECT 780.720 144.540 780.980 144.800 ;
        RECT 222.740 32.000 223.000 32.260 ;
        RECT 780.720 32.000 780.980 32.260 ;
      LAYER met2 ;
        RECT 784.630 601.530 784.910 604.000 ;
        RECT 783.080 601.390 784.910 601.530 ;
        RECT 783.080 586.570 783.220 601.390 ;
        RECT 784.630 600.000 784.910 601.390 ;
        RECT 782.620 586.430 783.220 586.570 ;
        RECT 782.620 531.410 782.760 586.430 ;
        RECT 780.720 531.090 780.980 531.410 ;
        RECT 782.560 531.090 782.820 531.410 ;
        RECT 780.780 403.650 780.920 531.090 ;
        RECT 780.320 403.510 780.920 403.650 ;
        RECT 780.320 144.830 780.460 403.510 ;
        RECT 780.260 144.510 780.520 144.830 ;
        RECT 780.720 144.510 780.980 144.830 ;
        RECT 780.780 32.290 780.920 144.510 ;
        RECT 222.740 31.970 223.000 32.290 ;
        RECT 780.720 31.970 780.980 32.290 ;
        RECT 222.800 2.400 222.940 31.970 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 676.270 569.400 676.590 569.460 ;
        RECT 678.570 569.400 678.890 569.460 ;
        RECT 676.270 569.260 678.890 569.400 ;
        RECT 676.270 569.200 676.590 569.260 ;
        RECT 678.570 569.200 678.890 569.260 ;
        RECT 20.310 30.840 20.630 30.900 ;
        RECT 676.270 30.840 676.590 30.900 ;
        RECT 20.310 30.700 676.590 30.840 ;
        RECT 20.310 30.640 20.630 30.700 ;
        RECT 676.270 30.640 676.590 30.700 ;
      LAYER via ;
        RECT 676.300 569.200 676.560 569.460 ;
        RECT 678.600 569.200 678.860 569.460 ;
        RECT 20.340 30.640 20.600 30.900 ;
        RECT 676.300 30.640 676.560 30.900 ;
      LAYER met2 ;
        RECT 680.210 600.170 680.490 604.000 ;
        RECT 678.660 600.030 680.490 600.170 ;
        RECT 678.660 569.490 678.800 600.030 ;
        RECT 680.210 600.000 680.490 600.030 ;
        RECT 676.300 569.170 676.560 569.490 ;
        RECT 678.600 569.170 678.860 569.490 ;
        RECT 676.360 30.930 676.500 569.170 ;
        RECT 20.340 30.610 20.600 30.930 ;
        RECT 676.300 30.610 676.560 30.930 ;
        RECT 20.400 2.400 20.540 30.610 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.570 2504.340 517.890 2504.400 ;
        RECT 524.010 2504.340 524.330 2504.400 ;
        RECT 1888.370 2504.340 1888.690 2504.400 ;
        RECT 517.570 2504.200 1888.690 2504.340 ;
        RECT 517.570 2504.140 517.890 2504.200 ;
        RECT 524.010 2504.140 524.330 2504.200 ;
        RECT 1888.370 2504.140 1888.690 2504.200 ;
        RECT 350.590 2038.880 350.910 2038.940 ;
        RECT 524.010 2038.880 524.330 2038.940 ;
        RECT 2083.870 2038.880 2084.190 2038.940 ;
        RECT 350.590 2038.740 2084.190 2038.880 ;
        RECT 350.590 2038.680 350.910 2038.740 ;
        RECT 524.010 2038.680 524.330 2038.740 ;
        RECT 2083.870 2038.680 2084.190 2038.740 ;
        RECT 349.210 593.200 349.530 593.260 ;
        RECT 351.510 593.200 351.830 593.260 ;
        RECT 690.990 593.200 691.310 593.260 ;
        RECT 349.210 593.060 691.310 593.200 ;
        RECT 349.210 593.000 349.530 593.060 ;
        RECT 351.510 593.000 351.830 593.060 ;
        RECT 690.990 593.000 691.310 593.060 ;
        RECT 47.910 589.800 48.230 589.860 ;
        RECT 349.210 589.800 349.530 589.860 ;
        RECT 47.910 589.660 349.530 589.800 ;
        RECT 47.910 589.600 48.230 589.660 ;
        RECT 349.210 589.600 349.530 589.660 ;
        RECT 44.230 17.580 44.550 17.640 ;
        RECT 47.910 17.580 48.230 17.640 ;
        RECT 44.230 17.440 48.230 17.580 ;
        RECT 44.230 17.380 44.550 17.440 ;
        RECT 47.910 17.380 48.230 17.440 ;
      LAYER via ;
        RECT 517.600 2504.140 517.860 2504.400 ;
        RECT 524.040 2504.140 524.300 2504.400 ;
        RECT 1888.400 2504.140 1888.660 2504.400 ;
        RECT 350.620 2038.680 350.880 2038.940 ;
        RECT 524.040 2038.680 524.300 2038.940 ;
        RECT 2083.900 2038.680 2084.160 2038.940 ;
        RECT 349.240 593.000 349.500 593.260 ;
        RECT 351.540 593.000 351.800 593.260 ;
        RECT 691.020 593.000 691.280 593.260 ;
        RECT 47.940 589.600 48.200 589.860 ;
        RECT 349.240 589.600 349.500 589.860 ;
        RECT 44.260 17.380 44.520 17.640 ;
        RECT 47.940 17.380 48.200 17.640 ;
      LAYER met2 ;
        RECT 519.330 2600.730 519.610 2604.000 ;
        RECT 517.660 2600.590 519.610 2600.730 ;
        RECT 517.660 2504.430 517.800 2600.590 ;
        RECT 519.330 2600.000 519.610 2600.590 ;
        RECT 1888.390 2595.715 1888.670 2596.085 ;
        RECT 1888.460 2504.430 1888.600 2595.715 ;
        RECT 517.600 2504.110 517.860 2504.430 ;
        RECT 524.040 2504.110 524.300 2504.430 ;
        RECT 1888.400 2504.110 1888.660 2504.430 ;
        RECT 524.100 2038.970 524.240 2504.110 ;
        RECT 350.620 2038.650 350.880 2038.970 ;
        RECT 524.040 2038.650 524.300 2038.970 ;
        RECT 2083.900 2038.650 2084.160 2038.970 ;
        RECT 350.680 1851.485 350.820 2038.650 ;
        RECT 2083.960 1873.245 2084.100 2038.650 ;
        RECT 2083.890 1872.875 2084.170 1873.245 ;
        RECT 350.610 1851.115 350.890 1851.485 ;
        RECT 351.530 1851.115 351.810 1851.485 ;
        RECT 351.600 593.290 351.740 1851.115 ;
        RECT 692.630 600.170 692.910 604.000 ;
        RECT 691.080 600.030 692.910 600.170 ;
        RECT 691.080 593.290 691.220 600.030 ;
        RECT 692.630 600.000 692.910 600.030 ;
        RECT 349.240 592.970 349.500 593.290 ;
        RECT 351.540 592.970 351.800 593.290 ;
        RECT 691.020 592.970 691.280 593.290 ;
        RECT 349.300 589.890 349.440 592.970 ;
        RECT 47.940 589.570 48.200 589.890 ;
        RECT 349.240 589.570 349.500 589.890 ;
        RECT 48.000 17.670 48.140 589.570 ;
        RECT 44.260 17.350 44.520 17.670 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 44.320 2.400 44.460 17.350 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 1888.390 2595.760 1888.670 2596.040 ;
        RECT 2083.890 1872.920 2084.170 1873.200 ;
        RECT 350.610 1851.160 350.890 1851.440 ;
        RECT 351.530 1851.160 351.810 1851.440 ;
      LAYER met3 ;
        RECT 1885.335 2596.600 1889.335 2597.200 ;
        RECT 1888.150 2596.065 1888.450 2596.600 ;
        RECT 1888.150 2595.750 1888.695 2596.065 ;
        RECT 1888.365 2595.735 1888.695 2595.750 ;
        RECT 2083.865 1873.210 2084.195 1873.225 ;
        RECT 2075.830 1872.910 2084.195 1873.210 ;
        RECT 2075.830 1870.320 2076.130 1872.910 ;
        RECT 2083.865 1872.895 2084.195 1872.910 ;
        RECT 2072.375 1869.720 2076.375 1870.320 ;
        RECT 350.585 1851.450 350.915 1851.465 ;
        RECT 351.505 1851.450 351.835 1851.465 ;
        RECT 360.000 1851.450 364.000 1851.600 ;
        RECT 350.585 1851.150 364.000 1851.450 ;
        RECT 350.585 1851.135 350.915 1851.150 ;
        RECT 351.505 1851.135 351.835 1851.150 ;
        RECT 360.000 1851.000 364.000 1851.150 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1501.050 2897.380 1501.370 2897.440 ;
        RECT 1554.870 2897.380 1555.190 2897.440 ;
        RECT 1501.050 2897.240 1555.190 2897.380 ;
        RECT 1501.050 2897.180 1501.370 2897.240 ;
        RECT 1554.870 2897.180 1555.190 2897.240 ;
        RECT 1501.050 2895.340 1501.370 2895.400 ;
        RECT 1485.500 2895.200 1501.370 2895.340 ;
        RECT 651.890 2895.000 652.210 2895.060 ;
        RECT 762.750 2895.000 763.070 2895.060 ;
        RECT 859.350 2895.000 859.670 2895.060 ;
        RECT 955.950 2895.000 956.270 2895.060 ;
        RECT 1052.550 2895.000 1052.870 2895.060 ;
        RECT 1149.150 2895.000 1149.470 2895.060 ;
        RECT 1245.750 2895.000 1246.070 2895.060 ;
        RECT 1342.350 2895.000 1342.670 2895.060 ;
        RECT 651.890 2894.860 763.070 2895.000 ;
        RECT 651.890 2894.800 652.210 2894.860 ;
        RECT 762.750 2894.800 763.070 2894.860 ;
        RECT 810.680 2894.860 859.670 2895.000 ;
        RECT 762.750 2893.980 763.070 2894.040 ;
        RECT 762.750 2893.840 786.440 2893.980 ;
        RECT 762.750 2893.780 763.070 2893.840 ;
        RECT 786.300 2893.640 786.440 2893.840 ;
        RECT 810.680 2893.640 810.820 2894.860 ;
        RECT 859.350 2894.800 859.670 2894.860 ;
        RECT 907.280 2894.860 956.270 2895.000 ;
        RECT 859.350 2893.980 859.670 2894.040 ;
        RECT 859.350 2893.840 883.040 2893.980 ;
        RECT 859.350 2893.780 859.670 2893.840 ;
        RECT 786.300 2893.500 810.820 2893.640 ;
        RECT 882.900 2893.640 883.040 2893.840 ;
        RECT 907.280 2893.640 907.420 2894.860 ;
        RECT 955.950 2894.800 956.270 2894.860 ;
        RECT 1003.880 2894.860 1052.870 2895.000 ;
        RECT 955.950 2893.980 956.270 2894.040 ;
        RECT 955.950 2893.840 979.640 2893.980 ;
        RECT 955.950 2893.780 956.270 2893.840 ;
        RECT 882.900 2893.500 907.420 2893.640 ;
        RECT 979.500 2893.640 979.640 2893.840 ;
        RECT 1003.880 2893.640 1004.020 2894.860 ;
        RECT 1052.550 2894.800 1052.870 2894.860 ;
        RECT 1100.480 2894.860 1149.470 2895.000 ;
        RECT 1052.550 2893.980 1052.870 2894.040 ;
        RECT 1052.550 2893.840 1076.240 2893.980 ;
        RECT 1052.550 2893.780 1052.870 2893.840 ;
        RECT 979.500 2893.500 1004.020 2893.640 ;
        RECT 1076.100 2893.640 1076.240 2893.840 ;
        RECT 1100.480 2893.640 1100.620 2894.860 ;
        RECT 1149.150 2894.800 1149.470 2894.860 ;
        RECT 1197.080 2894.860 1246.070 2895.000 ;
        RECT 1149.150 2893.980 1149.470 2894.040 ;
        RECT 1149.150 2893.840 1172.840 2893.980 ;
        RECT 1149.150 2893.780 1149.470 2893.840 ;
        RECT 1076.100 2893.500 1100.620 2893.640 ;
        RECT 1172.700 2893.640 1172.840 2893.840 ;
        RECT 1197.080 2893.640 1197.220 2894.860 ;
        RECT 1245.750 2894.800 1246.070 2894.860 ;
        RECT 1293.680 2894.860 1342.670 2895.000 ;
        RECT 1245.750 2893.980 1246.070 2894.040 ;
        RECT 1245.750 2893.840 1269.440 2893.980 ;
        RECT 1245.750 2893.780 1246.070 2893.840 ;
        RECT 1172.700 2893.500 1197.220 2893.640 ;
        RECT 1269.300 2893.640 1269.440 2893.840 ;
        RECT 1293.680 2893.640 1293.820 2894.860 ;
        RECT 1342.350 2894.800 1342.670 2894.860 ;
        RECT 1414.570 2895.000 1414.890 2895.060 ;
        RECT 1485.500 2895.000 1485.640 2895.200 ;
        RECT 1501.050 2895.140 1501.370 2895.200 ;
        RECT 1414.570 2894.860 1485.640 2895.000 ;
        RECT 1414.570 2894.800 1414.890 2894.860 ;
        RECT 1342.350 2893.980 1342.670 2894.040 ;
        RECT 1414.570 2893.980 1414.890 2894.040 ;
        RECT 1342.350 2893.840 1366.040 2893.980 ;
        RECT 1342.350 2893.780 1342.670 2893.840 ;
        RECT 1269.300 2893.500 1293.820 2893.640 ;
        RECT 1365.900 2893.640 1366.040 2893.840 ;
        RECT 1366.360 2893.840 1414.890 2893.980 ;
        RECT 1366.360 2893.640 1366.500 2893.840 ;
        RECT 1414.570 2893.780 1414.890 2893.840 ;
        RECT 1365.900 2893.500 1366.500 2893.640 ;
        RECT 446.730 2594.440 447.050 2594.500 ;
        RECT 612.790 2594.440 613.110 2594.500 ;
        RECT 446.730 2594.300 613.110 2594.440 ;
        RECT 446.730 2594.240 447.050 2594.300 ;
        RECT 612.790 2594.240 613.110 2594.300 ;
        RECT 614.170 2594.440 614.490 2594.500 ;
        RECT 648.670 2594.440 648.990 2594.500 ;
        RECT 614.170 2594.300 648.990 2594.440 ;
        RECT 614.170 2594.240 614.490 2594.300 ;
        RECT 648.670 2594.240 648.990 2594.300 ;
        RECT 648.670 2592.740 648.990 2592.800 ;
        RECT 651.890 2592.740 652.210 2592.800 ;
        RECT 648.670 2592.600 652.210 2592.740 ;
        RECT 648.670 2592.540 648.990 2592.600 ;
        RECT 651.890 2592.540 652.210 2592.600 ;
        RECT 648.670 1752.940 648.990 1753.000 ;
        RECT 652.350 1752.940 652.670 1753.000 ;
        RECT 648.670 1752.800 652.670 1752.940 ;
        RECT 648.670 1752.740 648.990 1752.800 ;
        RECT 652.350 1752.740 652.670 1752.800 ;
        RECT 652.350 1703.300 652.670 1703.360 ;
        RECT 1907.690 1703.300 1908.010 1703.360 ;
        RECT 652.350 1703.160 1908.010 1703.300 ;
        RECT 652.350 1703.100 652.670 1703.160 ;
        RECT 1907.690 1703.100 1908.010 1703.160 ;
        RECT 686.940 588.300 688.000 588.440 ;
        RECT 652.350 588.100 652.670 588.160 ;
        RECT 686.940 588.100 687.080 588.300 ;
        RECT 652.350 587.960 687.080 588.100 ;
        RECT 687.860 588.100 688.000 588.300 ;
        RECT 794.950 588.100 795.270 588.160 ;
        RECT 687.860 587.960 795.270 588.100 ;
        RECT 652.350 587.900 652.670 587.960 ;
        RECT 794.950 587.900 795.270 587.960 ;
        RECT 246.630 22.680 246.950 22.740 ;
        RECT 652.350 22.680 652.670 22.740 ;
        RECT 246.630 22.540 652.670 22.680 ;
        RECT 246.630 22.480 246.950 22.540 ;
        RECT 652.350 22.480 652.670 22.540 ;
      LAYER via ;
        RECT 1501.080 2897.180 1501.340 2897.440 ;
        RECT 1554.900 2897.180 1555.160 2897.440 ;
        RECT 651.920 2894.800 652.180 2895.060 ;
        RECT 762.780 2894.800 763.040 2895.060 ;
        RECT 762.780 2893.780 763.040 2894.040 ;
        RECT 859.380 2894.800 859.640 2895.060 ;
        RECT 859.380 2893.780 859.640 2894.040 ;
        RECT 955.980 2894.800 956.240 2895.060 ;
        RECT 955.980 2893.780 956.240 2894.040 ;
        RECT 1052.580 2894.800 1052.840 2895.060 ;
        RECT 1052.580 2893.780 1052.840 2894.040 ;
        RECT 1149.180 2894.800 1149.440 2895.060 ;
        RECT 1149.180 2893.780 1149.440 2894.040 ;
        RECT 1245.780 2894.800 1246.040 2895.060 ;
        RECT 1245.780 2893.780 1246.040 2894.040 ;
        RECT 1342.380 2894.800 1342.640 2895.060 ;
        RECT 1414.600 2894.800 1414.860 2895.060 ;
        RECT 1501.080 2895.140 1501.340 2895.400 ;
        RECT 1342.380 2893.780 1342.640 2894.040 ;
        RECT 1414.600 2893.780 1414.860 2894.040 ;
        RECT 446.760 2594.240 447.020 2594.500 ;
        RECT 612.820 2594.240 613.080 2594.500 ;
        RECT 614.200 2594.240 614.460 2594.500 ;
        RECT 648.700 2594.240 648.960 2594.500 ;
        RECT 648.700 2592.540 648.960 2592.800 ;
        RECT 651.920 2592.540 652.180 2592.800 ;
        RECT 648.700 1752.740 648.960 1753.000 ;
        RECT 652.380 1752.740 652.640 1753.000 ;
        RECT 652.380 1703.100 652.640 1703.360 ;
        RECT 1907.720 1703.100 1907.980 1703.360 ;
        RECT 652.380 587.900 652.640 588.160 ;
        RECT 794.980 587.900 795.240 588.160 ;
        RECT 246.660 22.480 246.920 22.740 ;
        RECT 652.380 22.480 652.640 22.740 ;
      LAYER met2 ;
        RECT 1501.080 2897.150 1501.340 2897.470 ;
        RECT 1554.900 2897.210 1555.160 2897.470 ;
        RECT 1556.210 2897.210 1556.490 2900.055 ;
        RECT 1554.900 2897.150 1556.490 2897.210 ;
        RECT 1501.140 2895.430 1501.280 2897.150 ;
        RECT 1554.960 2897.070 1556.490 2897.150 ;
        RECT 1556.210 2896.055 1556.490 2897.070 ;
        RECT 1501.080 2895.110 1501.340 2895.430 ;
        RECT 651.920 2894.770 652.180 2895.090 ;
        RECT 762.780 2894.770 763.040 2895.090 ;
        RECT 859.380 2894.770 859.640 2895.090 ;
        RECT 955.980 2894.770 956.240 2895.090 ;
        RECT 1052.580 2894.770 1052.840 2895.090 ;
        RECT 1149.180 2894.770 1149.440 2895.090 ;
        RECT 1245.780 2894.770 1246.040 2895.090 ;
        RECT 1342.380 2894.770 1342.640 2895.090 ;
        RECT 1414.600 2894.770 1414.860 2895.090 ;
        RECT 446.650 2600.660 446.930 2604.000 ;
        RECT 446.650 2600.000 446.960 2600.660 ;
        RECT 446.820 2594.530 446.960 2600.000 ;
        RECT 446.760 2594.210 447.020 2594.530 ;
        RECT 612.820 2594.210 613.080 2594.530 ;
        RECT 614.200 2594.210 614.460 2594.530 ;
        RECT 648.700 2594.210 648.960 2594.530 ;
        RECT 612.880 2593.930 613.020 2594.210 ;
        RECT 614.260 2593.930 614.400 2594.210 ;
        RECT 612.880 2593.790 614.400 2593.930 ;
        RECT 648.760 2592.830 648.900 2594.210 ;
        RECT 651.980 2592.830 652.120 2894.770 ;
        RECT 762.840 2894.070 762.980 2894.770 ;
        RECT 859.440 2894.070 859.580 2894.770 ;
        RECT 956.040 2894.070 956.180 2894.770 ;
        RECT 1052.640 2894.070 1052.780 2894.770 ;
        RECT 1149.240 2894.070 1149.380 2894.770 ;
        RECT 1245.840 2894.070 1245.980 2894.770 ;
        RECT 1342.440 2894.070 1342.580 2894.770 ;
        RECT 1414.660 2894.070 1414.800 2894.770 ;
        RECT 762.780 2893.750 763.040 2894.070 ;
        RECT 859.380 2893.750 859.640 2894.070 ;
        RECT 955.980 2893.750 956.240 2894.070 ;
        RECT 1052.580 2893.750 1052.840 2894.070 ;
        RECT 1149.180 2893.750 1149.440 2894.070 ;
        RECT 1245.780 2893.750 1246.040 2894.070 ;
        RECT 1342.380 2893.750 1342.640 2894.070 ;
        RECT 1414.600 2893.750 1414.860 2894.070 ;
        RECT 648.700 2592.510 648.960 2592.830 ;
        RECT 651.920 2592.510 652.180 2592.830 ;
        RECT 648.760 1754.925 648.900 2592.510 ;
        RECT 1907.710 1836.835 1907.990 1837.205 ;
        RECT 648.690 1754.555 648.970 1754.925 ;
        RECT 648.760 1753.030 648.900 1754.555 ;
        RECT 648.700 1752.710 648.960 1753.030 ;
        RECT 652.380 1752.710 652.640 1753.030 ;
        RECT 652.440 1703.390 652.580 1752.710 ;
        RECT 1907.780 1703.390 1907.920 1836.835 ;
        RECT 652.380 1703.070 652.640 1703.390 ;
        RECT 1907.720 1703.070 1907.980 1703.390 ;
        RECT 652.440 588.190 652.580 1703.070 ;
        RECT 796.590 600.170 796.870 604.000 ;
        RECT 795.040 600.030 796.870 600.170 ;
        RECT 795.040 588.190 795.180 600.030 ;
        RECT 796.590 600.000 796.870 600.030 ;
        RECT 652.380 587.870 652.640 588.190 ;
        RECT 794.980 587.870 795.240 588.190 ;
        RECT 652.440 22.770 652.580 587.870 ;
        RECT 246.660 22.450 246.920 22.770 ;
        RECT 652.380 22.450 652.640 22.770 ;
        RECT 246.720 2.400 246.860 22.450 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 1907.710 1836.880 1907.990 1837.160 ;
        RECT 648.690 1754.600 648.970 1754.880 ;
      LAYER met3 ;
        RECT 1920.000 1838.440 1924.000 1839.040 ;
        RECT 1907.685 1837.170 1908.015 1837.185 ;
        RECT 1920.350 1837.170 1920.650 1838.440 ;
        RECT 1907.685 1836.870 1920.650 1837.170 ;
        RECT 1907.685 1836.855 1908.015 1836.870 ;
        RECT 627.030 1754.890 631.030 1755.040 ;
        RECT 648.665 1754.890 648.995 1754.905 ;
        RECT 627.030 1754.590 648.995 1754.890 ;
        RECT 627.030 1754.440 631.030 1754.590 ;
        RECT 648.665 1754.575 648.995 1754.590 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1525.430 2898.060 1525.750 2898.120 ;
        RECT 1576.030 2898.060 1576.350 2898.120 ;
        RECT 1525.430 2897.920 1576.350 2898.060 ;
        RECT 1525.430 2897.860 1525.750 2897.920 ;
        RECT 1576.030 2897.860 1576.350 2897.920 ;
        RECT 1525.430 2896.700 1525.750 2896.760 ;
        RECT 1525.060 2896.560 1525.750 2896.700 ;
        RECT 1497.830 2896.020 1498.150 2896.080 ;
        RECT 1525.060 2896.020 1525.200 2896.560 ;
        RECT 1525.430 2896.500 1525.750 2896.560 ;
        RECT 1497.830 2895.880 1525.200 2896.020 ;
        RECT 1497.830 2895.820 1498.150 2895.880 ;
        RECT 1485.870 2895.000 1486.190 2895.060 ;
        RECT 1497.830 2895.000 1498.150 2895.060 ;
        RECT 1485.870 2894.860 1498.150 2895.000 ;
        RECT 1485.870 2894.800 1486.190 2894.860 ;
        RECT 1497.830 2894.800 1498.150 2894.860 ;
        RECT 737.910 2894.660 738.230 2894.720 ;
        RECT 761.370 2894.660 761.690 2894.720 ;
        RECT 857.970 2894.660 858.290 2894.720 ;
        RECT 954.570 2894.660 954.890 2894.720 ;
        RECT 1051.170 2894.660 1051.490 2894.720 ;
        RECT 1147.770 2894.660 1148.090 2894.720 ;
        RECT 1244.370 2894.660 1244.690 2894.720 ;
        RECT 1340.510 2894.660 1340.830 2894.720 ;
        RECT 737.910 2894.520 761.690 2894.660 ;
        RECT 737.910 2894.460 738.230 2894.520 ;
        RECT 761.370 2894.460 761.690 2894.520 ;
        RECT 811.140 2894.520 858.290 2894.660 ;
        RECT 613.710 2893.640 614.030 2893.700 ;
        RECT 737.910 2893.640 738.230 2893.700 ;
        RECT 613.710 2893.500 642.000 2893.640 ;
        RECT 613.710 2893.440 614.030 2893.500 ;
        RECT 641.860 2893.300 642.000 2893.500 ;
        RECT 690.160 2893.500 738.230 2893.640 ;
        RECT 690.160 2893.300 690.300 2893.500 ;
        RECT 737.910 2893.440 738.230 2893.500 ;
        RECT 641.860 2893.160 690.300 2893.300 ;
        RECT 761.370 2893.300 761.690 2893.360 ;
        RECT 811.140 2893.300 811.280 2894.520 ;
        RECT 857.970 2894.460 858.290 2894.520 ;
        RECT 907.740 2894.520 954.890 2894.660 ;
        RECT 761.370 2893.160 811.280 2893.300 ;
        RECT 857.970 2893.300 858.290 2893.360 ;
        RECT 907.740 2893.300 907.880 2894.520 ;
        RECT 954.570 2894.460 954.890 2894.520 ;
        RECT 1004.340 2894.520 1051.490 2894.660 ;
        RECT 857.970 2893.160 907.880 2893.300 ;
        RECT 954.570 2893.300 954.890 2893.360 ;
        RECT 1004.340 2893.300 1004.480 2894.520 ;
        RECT 1051.170 2894.460 1051.490 2894.520 ;
        RECT 1100.940 2894.520 1148.090 2894.660 ;
        RECT 954.570 2893.160 1004.480 2893.300 ;
        RECT 1051.170 2893.300 1051.490 2893.360 ;
        RECT 1100.940 2893.300 1101.080 2894.520 ;
        RECT 1147.770 2894.460 1148.090 2894.520 ;
        RECT 1197.540 2894.520 1244.690 2894.660 ;
        RECT 1051.170 2893.160 1101.080 2893.300 ;
        RECT 1147.770 2893.300 1148.090 2893.360 ;
        RECT 1197.540 2893.300 1197.680 2894.520 ;
        RECT 1244.370 2894.460 1244.690 2894.520 ;
        RECT 1294.140 2894.520 1340.830 2894.660 ;
        RECT 1147.770 2893.160 1197.680 2893.300 ;
        RECT 1244.370 2893.300 1244.690 2893.360 ;
        RECT 1294.140 2893.300 1294.280 2894.520 ;
        RECT 1340.510 2894.460 1340.830 2894.520 ;
        RECT 1390.190 2894.320 1390.510 2894.380 ;
        RECT 1390.190 2894.180 1437.800 2894.320 ;
        RECT 1390.190 2894.120 1390.510 2894.180 ;
        RECT 1244.370 2893.160 1294.280 2893.300 ;
        RECT 1340.510 2893.300 1340.830 2893.360 ;
        RECT 1390.190 2893.300 1390.510 2893.360 ;
        RECT 1340.510 2893.160 1390.510 2893.300 ;
        RECT 1437.660 2893.300 1437.800 2894.180 ;
        RECT 1485.870 2893.300 1486.190 2893.360 ;
        RECT 1437.660 2893.160 1486.190 2893.300 ;
        RECT 761.370 2893.100 761.690 2893.160 ;
        RECT 857.970 2893.100 858.290 2893.160 ;
        RECT 954.570 2893.100 954.890 2893.160 ;
        RECT 1051.170 2893.100 1051.490 2893.160 ;
        RECT 1147.770 2893.100 1148.090 2893.160 ;
        RECT 1244.370 2893.100 1244.690 2893.160 ;
        RECT 1340.510 2893.100 1340.830 2893.160 ;
        RECT 1390.190 2893.100 1390.510 2893.160 ;
        RECT 1485.870 2893.100 1486.190 2893.160 ;
        RECT 638.550 2594.100 638.870 2594.160 ;
        RECT 614.260 2593.960 638.870 2594.100 ;
        RECT 496.410 2593.760 496.730 2593.820 ;
        RECT 458.780 2593.620 496.730 2593.760 ;
        RECT 432.930 2593.420 433.250 2593.480 ;
        RECT 432.930 2593.280 447.880 2593.420 ;
        RECT 432.930 2593.220 433.250 2593.280 ;
        RECT 447.740 2593.080 447.880 2593.280 ;
        RECT 458.780 2593.080 458.920 2593.620 ;
        RECT 496.410 2593.560 496.730 2593.620 ;
        RECT 496.870 2593.760 497.190 2593.820 ;
        RECT 612.330 2593.760 612.650 2593.820 ;
        RECT 614.260 2593.760 614.400 2593.960 ;
        RECT 638.550 2593.900 638.870 2593.960 ;
        RECT 496.870 2593.620 524.700 2593.760 ;
        RECT 611.895 2593.620 614.400 2593.760 ;
        RECT 496.870 2593.560 497.190 2593.620 ;
        RECT 524.560 2593.420 524.700 2593.620 ;
        RECT 612.330 2593.560 612.650 2593.620 ;
        RECT 545.170 2593.420 545.490 2593.480 ;
        RECT 524.560 2593.280 545.490 2593.420 ;
        RECT 545.170 2593.220 545.490 2593.280 ;
        RECT 545.630 2593.420 545.950 2593.480 ;
        RECT 545.630 2593.280 579.900 2593.420 ;
        RECT 545.630 2593.220 545.950 2593.280 ;
        RECT 447.740 2592.940 458.920 2593.080 ;
        RECT 579.760 2593.080 579.900 2593.280 ;
        RECT 612.420 2593.080 612.560 2593.560 ;
        RECT 579.760 2592.940 612.560 2593.080 ;
        RECT 638.550 1703.640 638.870 1703.700 ;
        RECT 1908.150 1703.640 1908.470 1703.700 ;
        RECT 638.550 1703.500 1908.470 1703.640 ;
        RECT 638.550 1703.440 638.870 1703.500 ;
        RECT 1908.150 1703.440 1908.470 1703.500 ;
        RECT 613.250 1689.360 613.570 1689.420 ;
        RECT 638.550 1689.360 638.870 1689.420 ;
        RECT 613.250 1689.220 638.870 1689.360 ;
        RECT 613.250 1689.160 613.570 1689.220 ;
        RECT 638.550 1689.160 638.870 1689.220 ;
        RECT 612.790 1607.760 613.110 1607.820 ;
        RECT 613.710 1607.760 614.030 1607.820 ;
        RECT 612.790 1607.620 614.030 1607.760 ;
        RECT 612.790 1607.560 613.110 1607.620 ;
        RECT 613.710 1607.560 614.030 1607.620 ;
        RECT 612.330 1593.820 612.650 1593.880 ;
        RECT 613.710 1593.820 614.030 1593.880 ;
        RECT 612.330 1593.680 614.030 1593.820 ;
        RECT 612.330 1593.620 612.650 1593.680 ;
        RECT 613.710 1593.620 614.030 1593.680 ;
        RECT 612.330 1545.880 612.650 1545.940 ;
        RECT 613.250 1545.880 613.570 1545.940 ;
        RECT 612.330 1545.740 613.570 1545.880 ;
        RECT 612.330 1545.680 612.650 1545.740 ;
        RECT 613.250 1545.680 613.570 1545.740 ;
        RECT 612.790 1124.620 613.110 1124.680 ;
        RECT 613.710 1124.620 614.030 1124.680 ;
        RECT 612.790 1124.480 614.030 1124.620 ;
        RECT 612.790 1124.420 613.110 1124.480 ;
        RECT 613.710 1124.420 614.030 1124.480 ;
        RECT 613.710 1077.020 614.030 1077.080 ;
        RECT 613.340 1076.880 614.030 1077.020 ;
        RECT 613.340 1076.400 613.480 1076.880 ;
        RECT 613.710 1076.820 614.030 1076.880 ;
        RECT 613.250 1076.140 613.570 1076.400 ;
        RECT 613.710 979.440 614.030 979.500 ;
        RECT 614.630 979.440 614.950 979.500 ;
        RECT 613.710 979.300 614.950 979.440 ;
        RECT 613.710 979.240 614.030 979.300 ;
        RECT 614.630 979.240 614.950 979.300 ;
        RECT 613.710 883.560 614.030 883.620 ;
        RECT 613.340 883.420 614.030 883.560 ;
        RECT 613.340 882.940 613.480 883.420 ;
        RECT 613.710 883.360 614.030 883.420 ;
        RECT 613.250 882.680 613.570 882.940 ;
        RECT 612.790 807.400 613.110 807.460 ;
        RECT 613.710 807.400 614.030 807.460 ;
        RECT 612.790 807.260 614.030 807.400 ;
        RECT 612.790 807.200 613.110 807.260 ;
        RECT 613.710 807.200 614.030 807.260 ;
        RECT 612.790 737.700 613.110 737.760 ;
        RECT 613.710 737.700 614.030 737.760 ;
        RECT 612.790 737.560 614.030 737.700 ;
        RECT 612.790 737.500 613.110 737.560 ;
        RECT 613.710 737.500 614.030 737.560 ;
        RECT 612.790 689.900 613.110 690.160 ;
        RECT 612.880 689.420 613.020 689.900 ;
        RECT 613.250 689.420 613.570 689.480 ;
        RECT 612.880 689.280 613.570 689.420 ;
        RECT 613.250 689.220 613.570 689.280 ;
        RECT 610.490 589.120 610.810 589.180 ;
        RECT 613.250 589.120 613.570 589.180 ;
        RECT 804.150 589.120 804.470 589.180 ;
        RECT 610.490 588.980 804.470 589.120 ;
        RECT 610.490 588.920 610.810 588.980 ;
        RECT 613.250 588.920 613.570 588.980 ;
        RECT 804.150 588.920 804.470 588.980 ;
        RECT 264.110 22.340 264.430 22.400 ;
        RECT 610.490 22.340 610.810 22.400 ;
        RECT 264.110 22.200 610.810 22.340 ;
        RECT 264.110 22.140 264.430 22.200 ;
        RECT 610.490 22.140 610.810 22.200 ;
      LAYER via ;
        RECT 1525.460 2897.860 1525.720 2898.120 ;
        RECT 1576.060 2897.860 1576.320 2898.120 ;
        RECT 1497.860 2895.820 1498.120 2896.080 ;
        RECT 1525.460 2896.500 1525.720 2896.760 ;
        RECT 1485.900 2894.800 1486.160 2895.060 ;
        RECT 1497.860 2894.800 1498.120 2895.060 ;
        RECT 737.940 2894.460 738.200 2894.720 ;
        RECT 761.400 2894.460 761.660 2894.720 ;
        RECT 613.740 2893.440 614.000 2893.700 ;
        RECT 737.940 2893.440 738.200 2893.700 ;
        RECT 761.400 2893.100 761.660 2893.360 ;
        RECT 858.000 2894.460 858.260 2894.720 ;
        RECT 858.000 2893.100 858.260 2893.360 ;
        RECT 954.600 2894.460 954.860 2894.720 ;
        RECT 954.600 2893.100 954.860 2893.360 ;
        RECT 1051.200 2894.460 1051.460 2894.720 ;
        RECT 1051.200 2893.100 1051.460 2893.360 ;
        RECT 1147.800 2894.460 1148.060 2894.720 ;
        RECT 1147.800 2893.100 1148.060 2893.360 ;
        RECT 1244.400 2894.460 1244.660 2894.720 ;
        RECT 1244.400 2893.100 1244.660 2893.360 ;
        RECT 1340.540 2894.460 1340.800 2894.720 ;
        RECT 1390.220 2894.120 1390.480 2894.380 ;
        RECT 1340.540 2893.100 1340.800 2893.360 ;
        RECT 1390.220 2893.100 1390.480 2893.360 ;
        RECT 1485.900 2893.100 1486.160 2893.360 ;
        RECT 432.960 2593.220 433.220 2593.480 ;
        RECT 496.440 2593.560 496.700 2593.820 ;
        RECT 496.900 2593.560 497.160 2593.820 ;
        RECT 612.360 2593.560 612.620 2593.820 ;
        RECT 638.580 2593.900 638.840 2594.160 ;
        RECT 545.200 2593.220 545.460 2593.480 ;
        RECT 545.660 2593.220 545.920 2593.480 ;
        RECT 638.580 1703.440 638.840 1703.700 ;
        RECT 1908.180 1703.440 1908.440 1703.700 ;
        RECT 613.280 1689.160 613.540 1689.420 ;
        RECT 638.580 1689.160 638.840 1689.420 ;
        RECT 612.820 1607.560 613.080 1607.820 ;
        RECT 613.740 1607.560 614.000 1607.820 ;
        RECT 612.360 1593.620 612.620 1593.880 ;
        RECT 613.740 1593.620 614.000 1593.880 ;
        RECT 612.360 1545.680 612.620 1545.940 ;
        RECT 613.280 1545.680 613.540 1545.940 ;
        RECT 612.820 1124.420 613.080 1124.680 ;
        RECT 613.740 1124.420 614.000 1124.680 ;
        RECT 613.740 1076.820 614.000 1077.080 ;
        RECT 613.280 1076.140 613.540 1076.400 ;
        RECT 613.740 979.240 614.000 979.500 ;
        RECT 614.660 979.240 614.920 979.500 ;
        RECT 613.740 883.360 614.000 883.620 ;
        RECT 613.280 882.680 613.540 882.940 ;
        RECT 612.820 807.200 613.080 807.460 ;
        RECT 613.740 807.200 614.000 807.460 ;
        RECT 612.820 737.500 613.080 737.760 ;
        RECT 613.740 737.500 614.000 737.760 ;
        RECT 612.820 689.900 613.080 690.160 ;
        RECT 613.280 689.220 613.540 689.480 ;
        RECT 610.520 588.920 610.780 589.180 ;
        RECT 613.280 588.920 613.540 589.180 ;
        RECT 804.180 588.920 804.440 589.180 ;
        RECT 264.140 22.140 264.400 22.400 ;
        RECT 610.520 22.140 610.780 22.400 ;
      LAYER met2 ;
        RECT 1525.460 2897.830 1525.720 2898.150 ;
        RECT 1576.060 2897.890 1576.320 2898.150 ;
        RECT 1577.370 2897.890 1577.650 2900.055 ;
        RECT 1576.060 2897.830 1577.650 2897.890 ;
        RECT 1525.520 2896.790 1525.660 2897.830 ;
        RECT 1576.120 2897.750 1577.650 2897.830 ;
        RECT 1525.460 2896.470 1525.720 2896.790 ;
        RECT 1497.860 2895.790 1498.120 2896.110 ;
        RECT 1577.370 2896.055 1577.650 2897.750 ;
        RECT 1497.920 2895.090 1498.060 2895.790 ;
        RECT 1485.900 2894.770 1486.160 2895.090 ;
        RECT 1497.860 2894.770 1498.120 2895.090 ;
        RECT 737.940 2894.430 738.200 2894.750 ;
        RECT 761.400 2894.430 761.660 2894.750 ;
        RECT 858.000 2894.430 858.260 2894.750 ;
        RECT 954.600 2894.430 954.860 2894.750 ;
        RECT 1051.200 2894.430 1051.460 2894.750 ;
        RECT 1147.800 2894.430 1148.060 2894.750 ;
        RECT 1244.400 2894.430 1244.660 2894.750 ;
        RECT 1340.540 2894.430 1340.800 2894.750 ;
        RECT 738.000 2893.730 738.140 2894.430 ;
        RECT 613.740 2893.410 614.000 2893.730 ;
        RECT 737.940 2893.410 738.200 2893.730 ;
        RECT 432.850 2600.660 433.130 2604.000 ;
        RECT 432.850 2600.000 433.160 2600.660 ;
        RECT 433.020 2593.510 433.160 2600.000 ;
        RECT 613.800 2598.690 613.940 2893.410 ;
        RECT 761.460 2893.390 761.600 2894.430 ;
        RECT 858.060 2893.390 858.200 2894.430 ;
        RECT 954.660 2893.390 954.800 2894.430 ;
        RECT 1051.260 2893.390 1051.400 2894.430 ;
        RECT 1147.860 2893.390 1148.000 2894.430 ;
        RECT 1244.460 2893.390 1244.600 2894.430 ;
        RECT 1340.600 2893.390 1340.740 2894.430 ;
        RECT 1390.220 2894.090 1390.480 2894.410 ;
        RECT 1390.280 2893.390 1390.420 2894.090 ;
        RECT 1485.960 2893.390 1486.100 2894.770 ;
        RECT 761.400 2893.070 761.660 2893.390 ;
        RECT 858.000 2893.070 858.260 2893.390 ;
        RECT 954.600 2893.070 954.860 2893.390 ;
        RECT 1051.200 2893.070 1051.460 2893.390 ;
        RECT 1147.800 2893.070 1148.060 2893.390 ;
        RECT 1244.400 2893.070 1244.660 2893.390 ;
        RECT 1340.540 2893.070 1340.800 2893.390 ;
        RECT 1390.220 2893.070 1390.480 2893.390 ;
        RECT 1485.900 2893.070 1486.160 2893.390 ;
        RECT 612.420 2598.550 613.940 2598.690 ;
        RECT 496.500 2593.850 497.100 2593.930 ;
        RECT 612.420 2593.850 612.560 2598.550 ;
        RECT 638.580 2593.870 638.840 2594.190 ;
        RECT 496.440 2593.790 497.160 2593.850 ;
        RECT 496.440 2593.530 496.700 2593.790 ;
        RECT 496.900 2593.530 497.160 2593.790 ;
        RECT 612.360 2593.530 612.620 2593.850 ;
        RECT 432.960 2593.190 433.220 2593.510 ;
        RECT 545.200 2593.250 545.460 2593.510 ;
        RECT 545.660 2593.250 545.920 2593.510 ;
        RECT 545.200 2593.190 545.920 2593.250 ;
        RECT 545.260 2593.110 545.860 2593.190 ;
        RECT 613.090 1700.410 613.370 1704.000 ;
        RECT 638.640 1703.730 638.780 2593.870 ;
        RECT 1908.170 1801.475 1908.450 1801.845 ;
        RECT 1908.240 1703.730 1908.380 1801.475 ;
        RECT 638.580 1703.410 638.840 1703.730 ;
        RECT 1908.180 1703.410 1908.440 1703.730 ;
        RECT 613.090 1700.000 613.480 1700.410 ;
        RECT 613.340 1689.450 613.480 1700.000 ;
        RECT 638.640 1689.450 638.780 1703.410 ;
        RECT 613.280 1689.130 613.540 1689.450 ;
        RECT 638.580 1689.130 638.840 1689.450 ;
        RECT 613.340 1607.930 613.480 1689.130 ;
        RECT 612.880 1607.850 613.480 1607.930 ;
        RECT 612.820 1607.790 613.480 1607.850 ;
        RECT 612.820 1607.530 613.080 1607.790 ;
        RECT 613.740 1607.530 614.000 1607.850 ;
        RECT 612.880 1607.375 613.020 1607.530 ;
        RECT 613.800 1593.910 613.940 1607.530 ;
        RECT 612.360 1593.590 612.620 1593.910 ;
        RECT 613.740 1593.590 614.000 1593.910 ;
        RECT 612.420 1545.970 612.560 1593.590 ;
        RECT 612.360 1545.650 612.620 1545.970 ;
        RECT 613.280 1545.650 613.540 1545.970 ;
        RECT 613.340 1511.200 613.480 1545.650 ;
        RECT 612.880 1511.060 613.480 1511.200 ;
        RECT 612.880 1510.690 613.020 1511.060 ;
        RECT 612.880 1510.550 613.480 1510.690 ;
        RECT 613.340 1462.920 613.480 1510.550 ;
        RECT 613.340 1462.780 613.940 1462.920 ;
        RECT 613.800 1462.410 613.940 1462.780 ;
        RECT 613.340 1462.270 613.940 1462.410 ;
        RECT 613.340 1414.810 613.480 1462.270 ;
        RECT 612.880 1414.670 613.480 1414.810 ;
        RECT 612.880 1414.130 613.020 1414.670 ;
        RECT 612.880 1413.990 613.480 1414.130 ;
        RECT 613.340 1366.530 613.480 1413.990 ;
        RECT 613.340 1366.390 613.940 1366.530 ;
        RECT 613.800 1365.850 613.940 1366.390 ;
        RECT 613.340 1365.710 613.940 1365.850 ;
        RECT 613.340 1318.250 613.480 1365.710 ;
        RECT 612.880 1318.110 613.480 1318.250 ;
        RECT 612.880 1317.570 613.020 1318.110 ;
        RECT 612.880 1317.430 613.480 1317.570 ;
        RECT 613.340 1269.970 613.480 1317.430 ;
        RECT 613.340 1269.830 613.940 1269.970 ;
        RECT 613.800 1269.290 613.940 1269.830 ;
        RECT 613.340 1269.150 613.940 1269.290 ;
        RECT 613.340 1221.690 613.480 1269.150 ;
        RECT 612.880 1221.550 613.480 1221.690 ;
        RECT 612.880 1221.010 613.020 1221.550 ;
        RECT 612.880 1220.870 613.480 1221.010 ;
        RECT 613.340 1173.410 613.480 1220.870 ;
        RECT 613.340 1173.270 613.940 1173.410 ;
        RECT 613.800 1172.730 613.940 1173.270 ;
        RECT 613.340 1172.590 613.940 1172.730 ;
        RECT 613.340 1125.130 613.480 1172.590 ;
        RECT 612.880 1124.990 613.480 1125.130 ;
        RECT 612.880 1124.710 613.020 1124.990 ;
        RECT 612.820 1124.390 613.080 1124.710 ;
        RECT 613.740 1124.390 614.000 1124.710 ;
        RECT 613.800 1077.110 613.940 1124.390 ;
        RECT 613.740 1076.790 614.000 1077.110 ;
        RECT 613.280 1076.110 613.540 1076.430 ;
        RECT 613.340 1062.685 613.480 1076.110 ;
        RECT 613.270 1062.315 613.550 1062.685 ;
        RECT 614.190 1062.315 614.470 1062.685 ;
        RECT 614.260 1027.210 614.400 1062.315 ;
        RECT 613.340 1027.070 614.400 1027.210 ;
        RECT 613.340 1014.405 613.480 1027.070 ;
        RECT 613.270 1014.035 613.550 1014.405 ;
        RECT 614.650 1014.035 614.930 1014.405 ;
        RECT 614.720 979.530 614.860 1014.035 ;
        RECT 613.740 979.210 614.000 979.530 ;
        RECT 614.660 979.210 614.920 979.530 ;
        RECT 613.800 932.010 613.940 979.210 ;
        RECT 612.880 931.870 613.940 932.010 ;
        RECT 612.880 931.330 613.020 931.870 ;
        RECT 612.880 931.190 613.480 931.330 ;
        RECT 613.340 917.730 613.480 931.190 ;
        RECT 613.340 917.590 613.940 917.730 ;
        RECT 613.800 883.650 613.940 917.590 ;
        RECT 613.740 883.330 614.000 883.650 ;
        RECT 613.280 882.650 613.540 882.970 ;
        RECT 613.340 835.450 613.480 882.650 ;
        RECT 612.880 835.310 613.480 835.450 ;
        RECT 612.880 807.490 613.020 835.310 ;
        RECT 612.820 807.170 613.080 807.490 ;
        RECT 613.740 807.170 614.000 807.490 ;
        RECT 613.800 737.790 613.940 807.170 ;
        RECT 612.820 737.470 613.080 737.790 ;
        RECT 613.740 737.470 614.000 737.790 ;
        RECT 612.880 690.190 613.020 737.470 ;
        RECT 612.820 689.870 613.080 690.190 ;
        RECT 613.280 689.190 613.540 689.510 ;
        RECT 613.340 589.210 613.480 689.190 ;
        RECT 805.790 600.170 806.070 604.000 ;
        RECT 804.240 600.030 806.070 600.170 ;
        RECT 804.240 589.210 804.380 600.030 ;
        RECT 805.790 600.000 806.070 600.030 ;
        RECT 610.520 588.890 610.780 589.210 ;
        RECT 613.280 588.890 613.540 589.210 ;
        RECT 804.180 588.890 804.440 589.210 ;
        RECT 610.580 22.430 610.720 588.890 ;
        RECT 264.140 22.110 264.400 22.430 ;
        RECT 610.520 22.110 610.780 22.430 ;
        RECT 264.200 2.400 264.340 22.110 ;
        RECT 263.990 -4.800 264.550 2.400 ;
      LAYER via2 ;
        RECT 1908.170 1801.520 1908.450 1801.800 ;
        RECT 613.270 1062.360 613.550 1062.640 ;
        RECT 614.190 1062.360 614.470 1062.640 ;
        RECT 613.270 1014.080 613.550 1014.360 ;
        RECT 614.650 1014.080 614.930 1014.360 ;
      LAYER met3 ;
        RECT 1920.000 1804.440 1924.000 1805.040 ;
        RECT 1908.145 1801.810 1908.475 1801.825 ;
        RECT 1920.350 1801.810 1920.650 1804.440 ;
        RECT 1908.145 1801.510 1920.650 1801.810 ;
        RECT 1908.145 1801.495 1908.475 1801.510 ;
        RECT 613.245 1062.650 613.575 1062.665 ;
        RECT 614.165 1062.650 614.495 1062.665 ;
        RECT 613.245 1062.350 614.495 1062.650 ;
        RECT 613.245 1062.335 613.575 1062.350 ;
        RECT 614.165 1062.335 614.495 1062.350 ;
        RECT 613.245 1014.370 613.575 1014.385 ;
        RECT 614.625 1014.370 614.955 1014.385 ;
        RECT 613.245 1014.070 614.955 1014.370 ;
        RECT 613.245 1014.055 613.575 1014.070 ;
        RECT 614.625 1014.055 614.955 1014.070 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 2767.160 562.050 2767.220 ;
        RECT 580.130 2767.160 580.450 2767.220 ;
        RECT 561.730 2767.020 580.450 2767.160 ;
        RECT 561.730 2766.960 562.050 2767.020 ;
        RECT 580.130 2766.960 580.450 2767.020 ;
        RECT 580.130 2490.400 580.450 2490.460 ;
        RECT 1736.570 2490.400 1736.890 2490.460 ;
        RECT 580.130 2490.260 1736.890 2490.400 ;
        RECT 580.130 2490.200 580.450 2490.260 ;
        RECT 1736.570 2490.200 1736.890 2490.260 ;
        RECT 544.710 2488.020 545.030 2488.080 ;
        RECT 580.130 2488.020 580.450 2488.080 ;
        RECT 544.710 2487.880 580.450 2488.020 ;
        RECT 544.710 2487.820 545.030 2487.880 ;
        RECT 580.130 2487.820 580.450 2487.880 ;
        RECT 483.070 1979.380 483.390 1979.440 ;
        RECT 418.760 1979.240 483.390 1979.380 ;
        RECT 357.950 1978.700 358.270 1978.760 ;
        RECT 418.760 1978.700 418.900 1979.240 ;
        RECT 483.070 1979.180 483.390 1979.240 ;
        RECT 357.950 1978.560 418.900 1978.700 ;
        RECT 496.410 1978.700 496.730 1978.760 ;
        RECT 544.710 1978.700 545.030 1978.760 ;
        RECT 629.350 1978.700 629.670 1978.760 ;
        RECT 496.410 1978.560 629.670 1978.700 ;
        RECT 357.950 1978.500 358.270 1978.560 ;
        RECT 496.410 1978.500 496.730 1978.560 ;
        RECT 544.710 1978.500 545.030 1978.560 ;
        RECT 629.350 1978.500 629.670 1978.560 ;
        RECT 282.510 591.500 282.830 591.560 ;
        RECT 629.350 591.500 629.670 591.560 ;
        RECT 634.410 591.500 634.730 591.560 ;
        RECT 282.510 591.360 634.730 591.500 ;
        RECT 282.510 591.300 282.830 591.360 ;
        RECT 629.350 591.300 629.670 591.360 ;
        RECT 634.410 591.300 634.730 591.360 ;
        RECT 634.410 588.780 634.730 588.840 ;
        RECT 814.270 588.780 814.590 588.840 ;
        RECT 634.410 588.640 814.590 588.780 ;
        RECT 634.410 588.580 634.730 588.640 ;
        RECT 814.270 588.580 814.590 588.640 ;
      LAYER via ;
        RECT 561.760 2766.960 562.020 2767.220 ;
        RECT 580.160 2766.960 580.420 2767.220 ;
        RECT 580.160 2490.200 580.420 2490.460 ;
        RECT 1736.600 2490.200 1736.860 2490.460 ;
        RECT 544.740 2487.820 545.000 2488.080 ;
        RECT 580.160 2487.820 580.420 2488.080 ;
        RECT 357.980 1978.500 358.240 1978.760 ;
        RECT 483.100 1979.180 483.360 1979.440 ;
        RECT 496.440 1978.500 496.700 1978.760 ;
        RECT 544.740 1978.500 545.000 1978.760 ;
        RECT 629.380 1978.500 629.640 1978.760 ;
        RECT 282.540 591.300 282.800 591.560 ;
        RECT 629.380 591.300 629.640 591.560 ;
        RECT 634.440 591.300 634.700 591.560 ;
        RECT 634.440 588.580 634.700 588.840 ;
        RECT 814.300 588.580 814.560 588.840 ;
      LAYER met2 ;
        RECT 561.760 2766.930 562.020 2767.250 ;
        RECT 580.160 2766.930 580.420 2767.250 ;
        RECT 561.820 2759.520 561.960 2766.930 ;
        RECT 561.650 2759.100 561.960 2759.520 ;
        RECT 561.650 2755.520 561.930 2759.100 ;
        RECT 580.220 2490.490 580.360 2766.930 ;
        RECT 1736.530 2500.000 1736.810 2504.000 ;
        RECT 1736.660 2490.490 1736.800 2500.000 ;
        RECT 580.160 2490.170 580.420 2490.490 ;
        RECT 1736.600 2490.170 1736.860 2490.490 ;
        RECT 580.220 2488.110 580.360 2490.170 ;
        RECT 544.740 2487.790 545.000 2488.110 ;
        RECT 580.160 2487.790 580.420 2488.110 ;
        RECT 483.100 1979.325 483.360 1979.470 ;
        RECT 483.090 1978.955 483.370 1979.325 ;
        RECT 496.430 1978.955 496.710 1979.325 ;
        RECT 496.500 1978.790 496.640 1978.955 ;
        RECT 544.800 1978.790 544.940 2487.790 ;
        RECT 357.980 1978.470 358.240 1978.790 ;
        RECT 496.440 1978.470 496.700 1978.790 ;
        RECT 544.740 1978.470 545.000 1978.790 ;
        RECT 629.380 1978.470 629.640 1978.790 ;
        RECT 358.040 1814.765 358.180 1978.470 ;
        RECT 357.970 1814.395 358.250 1814.765 ;
        RECT 629.440 591.590 629.580 1978.470 ;
        RECT 814.990 600.170 815.270 604.000 ;
        RECT 814.360 600.030 815.270 600.170 ;
        RECT 282.540 591.270 282.800 591.590 ;
        RECT 629.380 591.270 629.640 591.590 ;
        RECT 634.440 591.270 634.700 591.590 ;
        RECT 282.600 24.210 282.740 591.270 ;
        RECT 634.500 588.870 634.640 591.270 ;
        RECT 814.360 588.870 814.500 600.030 ;
        RECT 814.990 600.000 815.270 600.030 ;
        RECT 634.440 588.550 634.700 588.870 ;
        RECT 814.300 588.550 814.560 588.870 ;
        RECT 282.140 24.070 282.740 24.210 ;
        RECT 282.140 2.400 282.280 24.070 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 483.090 1979.000 483.370 1979.280 ;
        RECT 496.430 1979.000 496.710 1979.280 ;
        RECT 357.970 1814.440 358.250 1814.720 ;
      LAYER met3 ;
        RECT 483.065 1979.290 483.395 1979.305 ;
        RECT 496.405 1979.290 496.735 1979.305 ;
        RECT 483.065 1978.990 496.735 1979.290 ;
        RECT 483.065 1978.975 483.395 1978.990 ;
        RECT 496.405 1978.975 496.735 1978.990 ;
        RECT 357.945 1814.730 358.275 1814.745 ;
        RECT 360.000 1814.730 364.000 1814.880 ;
        RECT 357.945 1814.430 364.000 1814.730 ;
        RECT 357.945 1814.415 358.275 1814.430 ;
        RECT 360.000 1814.280 364.000 1814.430 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.970 2487.340 559.290 2487.400 ;
        RECT 629.810 2487.340 630.130 2487.400 ;
        RECT 1863.530 2487.340 1863.850 2487.400 ;
        RECT 558.970 2487.200 1863.850 2487.340 ;
        RECT 558.970 2487.140 559.290 2487.200 ;
        RECT 629.810 2487.140 630.130 2487.200 ;
        RECT 1863.530 2487.140 1863.850 2487.200 ;
        RECT 413.610 1683.580 413.930 1683.640 ;
        RECT 629.810 1683.580 630.130 1683.640 ;
        RECT 413.610 1683.440 630.130 1683.580 ;
        RECT 413.610 1683.380 413.930 1683.440 ;
        RECT 629.810 1683.380 630.130 1683.440 ;
        RECT 413.610 592.520 413.930 592.580 ;
        RECT 822.550 592.520 822.870 592.580 ;
        RECT 413.610 592.380 822.870 592.520 ;
        RECT 413.610 592.320 413.930 592.380 ;
        RECT 822.550 592.320 822.870 592.380 ;
        RECT 303.210 590.140 303.530 590.200 ;
        RECT 413.610 590.140 413.930 590.200 ;
        RECT 303.210 590.000 413.930 590.140 ;
        RECT 303.210 589.940 303.530 590.000 ;
        RECT 413.610 589.940 413.930 590.000 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 559.000 2487.140 559.260 2487.400 ;
        RECT 629.840 2487.140 630.100 2487.400 ;
        RECT 1863.560 2487.140 1863.820 2487.400 ;
        RECT 413.640 1683.380 413.900 1683.640 ;
        RECT 629.840 1683.380 630.100 1683.640 ;
        RECT 413.640 592.320 413.900 592.580 ;
        RECT 822.580 592.320 822.840 592.580 ;
        RECT 303.240 589.940 303.500 590.200 ;
        RECT 413.640 589.940 413.900 590.200 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 562.570 2600.730 562.850 2604.000 ;
        RECT 559.060 2600.590 562.850 2600.730 ;
        RECT 559.060 2487.430 559.200 2600.590 ;
        RECT 562.570 2600.000 562.850 2600.590 ;
        RECT 1863.490 2500.000 1863.770 2504.000 ;
        RECT 1863.620 2487.430 1863.760 2500.000 ;
        RECT 559.000 2487.110 559.260 2487.430 ;
        RECT 629.840 2487.110 630.100 2487.430 ;
        RECT 1863.560 2487.110 1863.820 2487.430 ;
        RECT 412.530 1700.410 412.810 1704.000 ;
        RECT 412.530 1700.270 413.840 1700.410 ;
        RECT 412.530 1700.000 412.810 1700.270 ;
        RECT 413.700 1683.670 413.840 1700.270 ;
        RECT 629.900 1683.670 630.040 2487.110 ;
        RECT 413.640 1683.350 413.900 1683.670 ;
        RECT 629.840 1683.350 630.100 1683.670 ;
        RECT 413.700 592.610 413.840 1683.350 ;
        RECT 824.190 600.170 824.470 604.000 ;
        RECT 822.640 600.030 824.470 600.170 ;
        RECT 822.640 592.610 822.780 600.030 ;
        RECT 824.190 600.000 824.470 600.030 ;
        RECT 413.640 592.290 413.900 592.610 ;
        RECT 822.580 592.290 822.840 592.610 ;
        RECT 413.700 590.230 413.840 592.290 ;
        RECT 303.240 589.910 303.500 590.230 ;
        RECT 413.640 589.910 413.900 590.230 ;
        RECT 303.300 16.990 303.440 589.910 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1653.770 2898.060 1654.090 2898.120 ;
        RECT 1674.010 2898.060 1674.330 2898.120 ;
        RECT 1653.770 2897.920 1674.330 2898.060 ;
        RECT 1653.770 2897.860 1654.090 2897.920 ;
        RECT 1674.010 2897.860 1674.330 2897.920 ;
        RECT 1653.770 2896.500 1654.090 2896.760 ;
        RECT 1674.010 2896.500 1674.330 2896.760 ;
        RECT 1821.210 2896.500 1821.530 2896.760 ;
        RECT 1653.860 2893.640 1654.000 2896.500 ;
        RECT 1611.540 2893.500 1654.000 2893.640 ;
        RECT 1567.840 2892.140 1572.120 2892.280 ;
        RECT 646.370 2891.940 646.690 2892.000 ;
        RECT 1567.840 2891.940 1567.980 2892.140 ;
        RECT 646.370 2891.800 1567.980 2891.940 ;
        RECT 646.370 2891.740 646.690 2891.800 ;
        RECT 1571.980 2891.260 1572.120 2892.140 ;
        RECT 1611.540 2891.260 1611.680 2893.500 ;
        RECT 1571.980 2891.120 1611.680 2891.260 ;
        RECT 1674.100 2890.920 1674.240 2896.500 ;
        RECT 1821.300 2891.940 1821.440 2896.500 ;
        RECT 1696.180 2891.800 1821.440 2891.940 ;
        RECT 1696.180 2891.260 1696.320 2891.800 ;
        RECT 1693.880 2891.120 1696.320 2891.260 ;
        RECT 1674.100 2890.780 1674.700 2890.920 ;
        RECT 1674.560 2890.240 1674.700 2890.780 ;
        RECT 1693.880 2890.580 1694.020 2891.120 ;
        RECT 1675.940 2890.440 1694.020 2890.580 ;
        RECT 1675.940 2890.240 1676.080 2890.440 ;
        RECT 1674.560 2890.100 1676.080 2890.240 ;
        RECT 593.010 2625.380 593.330 2625.440 ;
        RECT 641.770 2625.380 642.090 2625.440 ;
        RECT 646.370 2625.380 646.690 2625.440 ;
        RECT 593.010 2625.240 646.690 2625.380 ;
        RECT 593.010 2625.180 593.330 2625.240 ;
        RECT 641.770 2625.180 642.090 2625.240 ;
        RECT 646.370 2625.180 646.690 2625.240 ;
        RECT 645.450 1870.580 645.770 1870.640 ;
        RECT 644.160 1870.440 645.770 1870.580 ;
        RECT 644.160 1870.300 644.300 1870.440 ;
        RECT 645.450 1870.380 645.770 1870.440 ;
        RECT 644.070 1870.040 644.390 1870.300 ;
        RECT 644.070 1801.220 644.390 1801.280 ;
        RECT 645.450 1801.220 645.770 1801.280 ;
        RECT 644.070 1801.080 645.770 1801.220 ;
        RECT 644.070 1801.020 644.390 1801.080 ;
        RECT 645.450 1801.020 645.770 1801.080 ;
        RECT 643.610 1739.000 643.930 1739.060 ;
        RECT 645.450 1739.000 645.770 1739.060 ;
        RECT 643.610 1738.860 645.770 1739.000 ;
        RECT 643.610 1738.800 643.930 1738.860 ;
        RECT 645.450 1738.800 645.770 1738.860 ;
        RECT 643.610 1727.780 643.930 1727.840 ;
        RECT 645.450 1727.780 645.770 1727.840 ;
        RECT 643.610 1727.640 645.770 1727.780 ;
        RECT 643.610 1727.580 643.930 1727.640 ;
        RECT 645.450 1727.580 645.770 1727.640 ;
        RECT 643.610 1680.180 643.930 1680.240 ;
        RECT 645.450 1680.180 645.770 1680.240 ;
        RECT 643.610 1680.040 645.770 1680.180 ;
        RECT 643.610 1679.980 643.930 1680.040 ;
        RECT 645.450 1679.980 645.770 1680.040 ;
        RECT 643.610 1635.300 643.930 1635.360 ;
        RECT 645.450 1635.300 645.770 1635.360 ;
        RECT 643.610 1635.160 645.770 1635.300 ;
        RECT 643.610 1635.100 643.930 1635.160 ;
        RECT 645.450 1635.100 645.770 1635.160 ;
        RECT 643.610 1558.120 643.930 1558.180 ;
        RECT 645.450 1558.120 645.770 1558.180 ;
        RECT 643.610 1557.980 645.770 1558.120 ;
        RECT 643.610 1557.920 643.930 1557.980 ;
        RECT 645.450 1557.920 645.770 1557.980 ;
        RECT 643.610 1535.340 643.930 1535.400 ;
        RECT 645.450 1535.340 645.770 1535.400 ;
        RECT 643.610 1535.200 645.770 1535.340 ;
        RECT 643.610 1535.140 643.930 1535.200 ;
        RECT 645.450 1535.140 645.770 1535.200 ;
        RECT 643.610 1487.060 643.930 1487.120 ;
        RECT 645.450 1487.060 645.770 1487.120 ;
        RECT 643.610 1486.920 645.770 1487.060 ;
        RECT 643.610 1486.860 643.930 1486.920 ;
        RECT 645.450 1486.860 645.770 1486.920 ;
        RECT 643.610 1438.780 643.930 1438.840 ;
        RECT 645.450 1438.780 645.770 1438.840 ;
        RECT 643.610 1438.640 645.770 1438.780 ;
        RECT 643.610 1438.580 643.930 1438.640 ;
        RECT 645.450 1438.580 645.770 1438.640 ;
        RECT 643.610 1371.460 643.930 1371.520 ;
        RECT 645.450 1371.460 645.770 1371.520 ;
        RECT 643.610 1371.320 645.770 1371.460 ;
        RECT 643.610 1371.260 643.930 1371.320 ;
        RECT 645.450 1371.260 645.770 1371.320 ;
        RECT 643.610 1342.220 643.930 1342.280 ;
        RECT 645.450 1342.220 645.770 1342.280 ;
        RECT 643.610 1342.080 645.770 1342.220 ;
        RECT 643.610 1342.020 643.930 1342.080 ;
        RECT 645.450 1342.020 645.770 1342.080 ;
        RECT 643.610 1293.940 643.930 1294.000 ;
        RECT 645.450 1293.940 645.770 1294.000 ;
        RECT 643.610 1293.800 645.770 1293.940 ;
        RECT 643.610 1293.740 643.930 1293.800 ;
        RECT 645.450 1293.740 645.770 1293.800 ;
        RECT 643.610 1245.660 643.930 1245.720 ;
        RECT 645.450 1245.660 645.770 1245.720 ;
        RECT 643.610 1245.520 645.770 1245.660 ;
        RECT 643.610 1245.460 643.930 1245.520 ;
        RECT 645.450 1245.460 645.770 1245.520 ;
        RECT 643.610 1197.380 643.930 1197.440 ;
        RECT 645.450 1197.380 645.770 1197.440 ;
        RECT 643.610 1197.240 645.770 1197.380 ;
        RECT 643.610 1197.180 643.930 1197.240 ;
        RECT 645.450 1197.180 645.770 1197.240 ;
        RECT 643.610 1148.760 643.930 1148.820 ;
        RECT 645.450 1148.760 645.770 1148.820 ;
        RECT 643.610 1148.620 645.770 1148.760 ;
        RECT 643.610 1148.560 643.930 1148.620 ;
        RECT 645.450 1148.560 645.770 1148.620 ;
        RECT 643.610 1100.480 643.930 1100.540 ;
        RECT 645.450 1100.480 645.770 1100.540 ;
        RECT 643.610 1100.340 645.770 1100.480 ;
        RECT 643.610 1100.280 643.930 1100.340 ;
        RECT 645.450 1100.280 645.770 1100.340 ;
        RECT 643.610 1052.200 643.930 1052.260 ;
        RECT 645.450 1052.200 645.770 1052.260 ;
        RECT 643.610 1052.060 645.770 1052.200 ;
        RECT 643.610 1052.000 643.930 1052.060 ;
        RECT 645.450 1052.000 645.770 1052.060 ;
        RECT 643.610 978.080 643.930 978.140 ;
        RECT 645.450 978.080 645.770 978.140 ;
        RECT 643.610 977.940 645.770 978.080 ;
        RECT 643.610 977.880 643.930 977.940 ;
        RECT 645.450 977.880 645.770 977.940 ;
        RECT 643.610 955.640 643.930 955.700 ;
        RECT 645.450 955.640 645.770 955.700 ;
        RECT 643.610 955.500 645.770 955.640 ;
        RECT 643.610 955.440 643.930 955.500 ;
        RECT 645.450 955.440 645.770 955.500 ;
        RECT 643.610 886.960 643.930 887.020 ;
        RECT 645.450 886.960 645.770 887.020 ;
        RECT 643.610 886.820 645.770 886.960 ;
        RECT 643.610 886.760 643.930 886.820 ;
        RECT 645.450 886.760 645.770 886.820 ;
        RECT 643.610 878.120 643.930 878.180 ;
        RECT 645.450 878.120 645.770 878.180 ;
        RECT 643.610 877.980 645.770 878.120 ;
        RECT 643.610 877.920 643.930 877.980 ;
        RECT 645.450 877.920 645.770 877.980 ;
        RECT 643.610 810.800 643.930 810.860 ;
        RECT 645.450 810.800 645.770 810.860 ;
        RECT 643.610 810.660 645.770 810.800 ;
        RECT 643.610 810.600 643.930 810.660 ;
        RECT 645.450 810.600 645.770 810.660 ;
        RECT 643.610 749.260 643.930 749.320 ;
        RECT 645.450 749.260 645.770 749.320 ;
        RECT 643.610 749.120 645.770 749.260 ;
        RECT 643.610 749.060 643.930 749.120 ;
        RECT 645.450 749.060 645.770 749.120 ;
        RECT 644.070 717.640 644.390 717.700 ;
        RECT 645.450 717.640 645.770 717.700 ;
        RECT 644.070 717.500 645.770 717.640 ;
        RECT 644.070 717.440 644.390 717.500 ;
        RECT 645.450 717.440 645.770 717.500 ;
        RECT 644.070 676.160 644.390 676.220 ;
        RECT 645.450 676.160 645.770 676.220 ;
        RECT 644.070 676.020 645.770 676.160 ;
        RECT 644.070 675.960 644.390 676.020 ;
        RECT 645.450 675.960 645.770 676.020 ;
        RECT 644.070 652.020 644.390 652.080 ;
        RECT 645.450 652.020 645.770 652.080 ;
        RECT 644.070 651.880 645.770 652.020 ;
        RECT 644.070 651.820 644.390 651.880 ;
        RECT 645.450 651.820 645.770 651.880 ;
        RECT 644.070 627.880 644.390 627.940 ;
        RECT 645.450 627.880 645.770 627.940 ;
        RECT 644.070 627.740 645.770 627.880 ;
        RECT 644.070 627.680 644.390 627.740 ;
        RECT 645.450 627.680 645.770 627.740 ;
        RECT 688.230 588.440 688.550 588.500 ;
        RECT 831.290 588.440 831.610 588.500 ;
        RECT 688.230 588.300 831.610 588.440 ;
        RECT 688.230 588.240 688.550 588.300 ;
        RECT 831.290 588.240 831.610 588.300 ;
        RECT 644.070 587.760 644.390 587.820 ;
        RECT 688.230 587.760 688.550 587.820 ;
        RECT 644.070 587.620 688.550 587.760 ;
        RECT 644.070 587.560 644.390 587.620 ;
        RECT 688.230 587.560 688.550 587.620 ;
        RECT 643.610 579.600 643.930 579.660 ;
        RECT 644.990 579.600 645.310 579.660 ;
        RECT 643.610 579.460 645.310 579.600 ;
        RECT 643.610 579.400 643.930 579.460 ;
        RECT 644.990 579.400 645.310 579.460 ;
        RECT 644.530 386.140 644.850 386.200 ;
        RECT 644.990 386.140 645.310 386.200 ;
        RECT 644.530 386.000 645.310 386.140 ;
        RECT 644.530 385.940 644.850 386.000 ;
        RECT 644.990 385.940 645.310 386.000 ;
        RECT 644.070 337.860 644.390 337.920 ;
        RECT 645.450 337.860 645.770 337.920 ;
        RECT 644.070 337.720 645.770 337.860 ;
        RECT 644.070 337.660 644.390 337.720 ;
        RECT 645.450 337.660 645.770 337.720 ;
        RECT 644.070 303.520 644.390 303.580 ;
        RECT 645.450 303.520 645.770 303.580 ;
        RECT 644.070 303.380 645.770 303.520 ;
        RECT 644.070 303.320 644.390 303.380 ;
        RECT 645.450 303.320 645.770 303.380 ;
        RECT 645.450 241.640 645.770 241.700 ;
        RECT 645.080 241.500 645.770 241.640 ;
        RECT 645.080 241.360 645.220 241.500 ;
        RECT 645.450 241.440 645.770 241.500 ;
        RECT 644.990 241.100 645.310 241.360 ;
        RECT 645.450 234.300 645.770 234.560 ;
        RECT 645.540 233.880 645.680 234.300 ;
        RECT 645.450 233.620 645.770 233.880 ;
        RECT 644.070 169.220 644.390 169.280 ;
        RECT 645.450 169.220 645.770 169.280 ;
        RECT 644.070 169.080 645.770 169.220 ;
        RECT 644.070 169.020 644.390 169.080 ;
        RECT 645.450 169.020 645.770 169.080 ;
        RECT 643.610 96.460 643.930 96.520 ;
        RECT 645.450 96.460 645.770 96.520 ;
        RECT 643.610 96.320 645.770 96.460 ;
        RECT 643.610 96.260 643.930 96.320 ;
        RECT 645.450 96.260 645.770 96.320 ;
        RECT 643.610 48.520 643.930 48.580 ;
        RECT 644.530 48.520 644.850 48.580 ;
        RECT 643.610 48.380 644.850 48.520 ;
        RECT 643.610 48.320 643.930 48.380 ;
        RECT 644.530 48.320 644.850 48.380 ;
        RECT 317.930 36.280 318.250 36.340 ;
        RECT 644.530 36.280 644.850 36.340 ;
        RECT 317.930 36.140 644.850 36.280 ;
        RECT 317.930 36.080 318.250 36.140 ;
        RECT 644.530 36.080 644.850 36.140 ;
      LAYER via ;
        RECT 1653.800 2897.860 1654.060 2898.120 ;
        RECT 1674.040 2897.860 1674.300 2898.120 ;
        RECT 1653.800 2896.500 1654.060 2896.760 ;
        RECT 1674.040 2896.500 1674.300 2896.760 ;
        RECT 1821.240 2896.500 1821.500 2896.760 ;
        RECT 646.400 2891.740 646.660 2892.000 ;
        RECT 593.040 2625.180 593.300 2625.440 ;
        RECT 641.800 2625.180 642.060 2625.440 ;
        RECT 646.400 2625.180 646.660 2625.440 ;
        RECT 645.480 1870.380 645.740 1870.640 ;
        RECT 644.100 1870.040 644.360 1870.300 ;
        RECT 644.100 1801.020 644.360 1801.280 ;
        RECT 645.480 1801.020 645.740 1801.280 ;
        RECT 643.640 1738.800 643.900 1739.060 ;
        RECT 645.480 1738.800 645.740 1739.060 ;
        RECT 643.640 1727.580 643.900 1727.840 ;
        RECT 645.480 1727.580 645.740 1727.840 ;
        RECT 643.640 1679.980 643.900 1680.240 ;
        RECT 645.480 1679.980 645.740 1680.240 ;
        RECT 643.640 1635.100 643.900 1635.360 ;
        RECT 645.480 1635.100 645.740 1635.360 ;
        RECT 643.640 1557.920 643.900 1558.180 ;
        RECT 645.480 1557.920 645.740 1558.180 ;
        RECT 643.640 1535.140 643.900 1535.400 ;
        RECT 645.480 1535.140 645.740 1535.400 ;
        RECT 643.640 1486.860 643.900 1487.120 ;
        RECT 645.480 1486.860 645.740 1487.120 ;
        RECT 643.640 1438.580 643.900 1438.840 ;
        RECT 645.480 1438.580 645.740 1438.840 ;
        RECT 643.640 1371.260 643.900 1371.520 ;
        RECT 645.480 1371.260 645.740 1371.520 ;
        RECT 643.640 1342.020 643.900 1342.280 ;
        RECT 645.480 1342.020 645.740 1342.280 ;
        RECT 643.640 1293.740 643.900 1294.000 ;
        RECT 645.480 1293.740 645.740 1294.000 ;
        RECT 643.640 1245.460 643.900 1245.720 ;
        RECT 645.480 1245.460 645.740 1245.720 ;
        RECT 643.640 1197.180 643.900 1197.440 ;
        RECT 645.480 1197.180 645.740 1197.440 ;
        RECT 643.640 1148.560 643.900 1148.820 ;
        RECT 645.480 1148.560 645.740 1148.820 ;
        RECT 643.640 1100.280 643.900 1100.540 ;
        RECT 645.480 1100.280 645.740 1100.540 ;
        RECT 643.640 1052.000 643.900 1052.260 ;
        RECT 645.480 1052.000 645.740 1052.260 ;
        RECT 643.640 977.880 643.900 978.140 ;
        RECT 645.480 977.880 645.740 978.140 ;
        RECT 643.640 955.440 643.900 955.700 ;
        RECT 645.480 955.440 645.740 955.700 ;
        RECT 643.640 886.760 643.900 887.020 ;
        RECT 645.480 886.760 645.740 887.020 ;
        RECT 643.640 877.920 643.900 878.180 ;
        RECT 645.480 877.920 645.740 878.180 ;
        RECT 643.640 810.600 643.900 810.860 ;
        RECT 645.480 810.600 645.740 810.860 ;
        RECT 643.640 749.060 643.900 749.320 ;
        RECT 645.480 749.060 645.740 749.320 ;
        RECT 644.100 717.440 644.360 717.700 ;
        RECT 645.480 717.440 645.740 717.700 ;
        RECT 644.100 675.960 644.360 676.220 ;
        RECT 645.480 675.960 645.740 676.220 ;
        RECT 644.100 651.820 644.360 652.080 ;
        RECT 645.480 651.820 645.740 652.080 ;
        RECT 644.100 627.680 644.360 627.940 ;
        RECT 645.480 627.680 645.740 627.940 ;
        RECT 688.260 588.240 688.520 588.500 ;
        RECT 831.320 588.240 831.580 588.500 ;
        RECT 644.100 587.560 644.360 587.820 ;
        RECT 688.260 587.560 688.520 587.820 ;
        RECT 643.640 579.400 643.900 579.660 ;
        RECT 645.020 579.400 645.280 579.660 ;
        RECT 644.560 385.940 644.820 386.200 ;
        RECT 645.020 385.940 645.280 386.200 ;
        RECT 644.100 337.660 644.360 337.920 ;
        RECT 645.480 337.660 645.740 337.920 ;
        RECT 644.100 303.320 644.360 303.580 ;
        RECT 645.480 303.320 645.740 303.580 ;
        RECT 645.480 241.440 645.740 241.700 ;
        RECT 645.020 241.100 645.280 241.360 ;
        RECT 645.480 234.300 645.740 234.560 ;
        RECT 645.480 233.620 645.740 233.880 ;
        RECT 644.100 169.020 644.360 169.280 ;
        RECT 645.480 169.020 645.740 169.280 ;
        RECT 643.640 96.260 643.900 96.520 ;
        RECT 645.480 96.260 645.740 96.520 ;
        RECT 643.640 48.320 643.900 48.580 ;
        RECT 644.560 48.320 644.820 48.580 ;
        RECT 317.960 36.080 318.220 36.340 ;
        RECT 644.560 36.080 644.820 36.340 ;
      LAYER met2 ;
        RECT 1653.800 2897.830 1654.060 2898.150 ;
        RECT 1674.040 2897.830 1674.300 2898.150 ;
        RECT 1653.860 2896.790 1654.000 2897.830 ;
        RECT 1674.100 2896.790 1674.240 2897.830 ;
        RECT 1653.800 2896.470 1654.060 2896.790 ;
        RECT 1674.040 2896.470 1674.300 2896.790 ;
        RECT 1821.240 2896.530 1821.500 2896.790 ;
        RECT 1822.090 2896.530 1822.370 2900.055 ;
        RECT 1821.240 2896.470 1822.370 2896.530 ;
        RECT 1821.300 2896.390 1822.370 2896.470 ;
        RECT 1822.090 2896.055 1822.370 2896.390 ;
        RECT 646.400 2891.710 646.660 2892.030 ;
        RECT 593.030 2625.635 593.310 2626.005 ;
        RECT 593.100 2625.470 593.240 2625.635 ;
        RECT 646.460 2625.470 646.600 2891.710 ;
        RECT 593.040 2625.150 593.300 2625.470 ;
        RECT 641.800 2625.150 642.060 2625.470 ;
        RECT 646.400 2625.150 646.660 2625.470 ;
        RECT 641.860 2621.130 642.000 2625.150 ;
        RECT 641.860 2620.990 642.920 2621.130 ;
        RECT 642.780 1939.885 642.920 2620.990 ;
        RECT 642.710 1939.515 642.990 1939.885 ;
        RECT 645.470 1939.515 645.750 1939.885 ;
        RECT 645.540 1870.670 645.680 1939.515 ;
        RECT 645.480 1870.350 645.740 1870.670 ;
        RECT 644.100 1870.010 644.360 1870.330 ;
        RECT 644.160 1801.310 644.300 1870.010 ;
        RECT 644.100 1800.990 644.360 1801.310 ;
        RECT 645.480 1800.990 645.740 1801.310 ;
        RECT 645.540 1739.090 645.680 1800.990 ;
        RECT 643.640 1738.770 643.900 1739.090 ;
        RECT 645.480 1738.770 645.740 1739.090 ;
        RECT 643.700 1727.870 643.840 1738.770 ;
        RECT 643.640 1727.550 643.900 1727.870 ;
        RECT 645.480 1727.550 645.740 1727.870 ;
        RECT 645.540 1680.270 645.680 1727.550 ;
        RECT 643.640 1679.950 643.900 1680.270 ;
        RECT 645.480 1679.950 645.740 1680.270 ;
        RECT 643.700 1635.390 643.840 1679.950 ;
        RECT 643.640 1635.070 643.900 1635.390 ;
        RECT 645.480 1635.070 645.740 1635.390 ;
        RECT 645.540 1558.210 645.680 1635.070 ;
        RECT 643.640 1557.890 643.900 1558.210 ;
        RECT 645.480 1557.890 645.740 1558.210 ;
        RECT 643.700 1535.430 643.840 1557.890 ;
        RECT 643.640 1535.110 643.900 1535.430 ;
        RECT 645.480 1535.110 645.740 1535.430 ;
        RECT 645.540 1487.150 645.680 1535.110 ;
        RECT 643.640 1486.830 643.900 1487.150 ;
        RECT 645.480 1486.830 645.740 1487.150 ;
        RECT 643.700 1438.870 643.840 1486.830 ;
        RECT 643.640 1438.550 643.900 1438.870 ;
        RECT 645.480 1438.550 645.740 1438.870 ;
        RECT 645.540 1371.550 645.680 1438.550 ;
        RECT 643.640 1371.230 643.900 1371.550 ;
        RECT 645.480 1371.230 645.740 1371.550 ;
        RECT 643.700 1342.310 643.840 1371.230 ;
        RECT 643.640 1341.990 643.900 1342.310 ;
        RECT 645.480 1341.990 645.740 1342.310 ;
        RECT 645.540 1294.030 645.680 1341.990 ;
        RECT 643.640 1293.710 643.900 1294.030 ;
        RECT 645.480 1293.710 645.740 1294.030 ;
        RECT 643.700 1245.750 643.840 1293.710 ;
        RECT 643.640 1245.430 643.900 1245.750 ;
        RECT 645.480 1245.430 645.740 1245.750 ;
        RECT 645.540 1197.470 645.680 1245.430 ;
        RECT 643.640 1197.150 643.900 1197.470 ;
        RECT 645.480 1197.150 645.740 1197.470 ;
        RECT 643.700 1148.850 643.840 1197.150 ;
        RECT 643.640 1148.530 643.900 1148.850 ;
        RECT 645.480 1148.530 645.740 1148.850 ;
        RECT 645.540 1100.570 645.680 1148.530 ;
        RECT 643.640 1100.250 643.900 1100.570 ;
        RECT 645.480 1100.250 645.740 1100.570 ;
        RECT 643.700 1052.290 643.840 1100.250 ;
        RECT 643.640 1051.970 643.900 1052.290 ;
        RECT 645.480 1051.970 645.740 1052.290 ;
        RECT 645.540 978.170 645.680 1051.970 ;
        RECT 643.640 977.850 643.900 978.170 ;
        RECT 645.480 977.850 645.740 978.170 ;
        RECT 643.700 955.730 643.840 977.850 ;
        RECT 643.640 955.410 643.900 955.730 ;
        RECT 645.480 955.410 645.740 955.730 ;
        RECT 645.540 887.050 645.680 955.410 ;
        RECT 643.640 886.730 643.900 887.050 ;
        RECT 645.480 886.730 645.740 887.050 ;
        RECT 643.700 878.210 643.840 886.730 ;
        RECT 643.640 877.890 643.900 878.210 ;
        RECT 645.480 877.890 645.740 878.210 ;
        RECT 645.540 810.890 645.680 877.890 ;
        RECT 643.640 810.570 643.900 810.890 ;
        RECT 645.480 810.570 645.740 810.890 ;
        RECT 643.700 749.350 643.840 810.570 ;
        RECT 643.640 749.030 643.900 749.350 ;
        RECT 645.480 749.030 645.740 749.350 ;
        RECT 645.540 717.730 645.680 749.030 ;
        RECT 644.100 717.410 644.360 717.730 ;
        RECT 645.480 717.410 645.740 717.730 ;
        RECT 644.160 676.250 644.300 717.410 ;
        RECT 644.100 675.930 644.360 676.250 ;
        RECT 645.480 675.930 645.740 676.250 ;
        RECT 645.540 652.110 645.680 675.930 ;
        RECT 644.100 651.790 644.360 652.110 ;
        RECT 645.480 651.790 645.740 652.110 ;
        RECT 644.160 628.165 644.300 651.790 ;
        RECT 644.090 627.795 644.370 628.165 ;
        RECT 645.470 627.795 645.750 628.165 ;
        RECT 644.100 627.650 644.360 627.795 ;
        RECT 645.480 627.650 645.740 627.795 ;
        RECT 644.160 587.850 644.300 627.650 ;
        RECT 833.390 600.170 833.670 604.000 ;
        RECT 831.380 600.030 833.670 600.170 ;
        RECT 831.380 588.530 831.520 600.030 ;
        RECT 833.390 600.000 833.670 600.030 ;
        RECT 688.260 588.210 688.520 588.530 ;
        RECT 831.320 588.210 831.580 588.530 ;
        RECT 688.320 587.850 688.460 588.210 ;
        RECT 644.100 587.530 644.360 587.850 ;
        RECT 688.260 587.530 688.520 587.850 ;
        RECT 644.160 579.885 644.300 587.530 ;
        RECT 643.640 579.370 643.900 579.690 ;
        RECT 644.090 579.515 644.370 579.885 ;
        RECT 645.010 579.515 645.290 579.885 ;
        RECT 645.020 579.370 645.280 579.515 ;
        RECT 643.700 531.605 643.840 579.370 ;
        RECT 643.630 531.235 643.910 531.605 ;
        RECT 644.550 531.235 644.830 531.605 ;
        RECT 644.620 495.450 644.760 531.235 ;
        RECT 644.620 495.310 645.680 495.450 ;
        RECT 645.540 448.530 645.680 495.310 ;
        RECT 644.620 448.390 645.680 448.530 ;
        RECT 644.620 399.570 644.760 448.390 ;
        RECT 644.620 399.430 645.220 399.570 ;
        RECT 645.080 386.230 645.220 399.430 ;
        RECT 644.560 385.910 644.820 386.230 ;
        RECT 645.020 385.910 645.280 386.230 ;
        RECT 644.620 339.165 644.760 385.910 ;
        RECT 644.550 338.795 644.830 339.165 ;
        RECT 645.470 338.115 645.750 338.485 ;
        RECT 645.540 337.950 645.680 338.115 ;
        RECT 644.100 337.630 644.360 337.950 ;
        RECT 645.480 337.630 645.740 337.950 ;
        RECT 644.160 303.610 644.300 337.630 ;
        RECT 644.100 303.290 644.360 303.610 ;
        RECT 645.480 303.290 645.740 303.610 ;
        RECT 645.540 290.090 645.680 303.290 ;
        RECT 645.080 289.950 645.680 290.090 ;
        RECT 645.080 266.290 645.220 289.950 ;
        RECT 645.080 266.150 645.680 266.290 ;
        RECT 645.540 241.730 645.680 266.150 ;
        RECT 645.480 241.410 645.740 241.730 ;
        RECT 645.020 241.070 645.280 241.390 ;
        RECT 645.080 235.010 645.220 241.070 ;
        RECT 645.080 234.870 645.680 235.010 ;
        RECT 645.540 234.590 645.680 234.870 ;
        RECT 645.480 234.270 645.740 234.590 ;
        RECT 645.480 233.590 645.740 233.910 ;
        RECT 645.540 169.310 645.680 233.590 ;
        RECT 644.100 168.990 644.360 169.310 ;
        RECT 645.480 168.990 645.740 169.310 ;
        RECT 644.160 158.170 644.300 168.990 ;
        RECT 644.160 158.030 644.760 158.170 ;
        RECT 644.620 110.570 644.760 158.030 ;
        RECT 644.620 110.430 645.680 110.570 ;
        RECT 645.540 96.550 645.680 110.430 ;
        RECT 643.640 96.230 643.900 96.550 ;
        RECT 645.480 96.230 645.740 96.550 ;
        RECT 643.700 48.610 643.840 96.230 ;
        RECT 643.640 48.290 643.900 48.610 ;
        RECT 644.560 48.290 644.820 48.610 ;
        RECT 644.620 36.370 644.760 48.290 ;
        RECT 317.960 36.050 318.220 36.370 ;
        RECT 644.560 36.050 644.820 36.370 ;
        RECT 318.020 2.400 318.160 36.050 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 593.030 2625.680 593.310 2625.960 ;
        RECT 642.710 1939.560 642.990 1939.840 ;
        RECT 645.470 1939.560 645.750 1939.840 ;
        RECT 644.090 627.840 644.370 628.120 ;
        RECT 645.470 627.840 645.750 628.120 ;
        RECT 644.090 579.560 644.370 579.840 ;
        RECT 645.010 579.560 645.290 579.840 ;
        RECT 643.630 531.280 643.910 531.560 ;
        RECT 644.550 531.280 644.830 531.560 ;
        RECT 644.550 338.840 644.830 339.120 ;
        RECT 645.470 338.160 645.750 338.440 ;
      LAYER met3 ;
        RECT 574.800 2625.970 578.800 2626.480 ;
        RECT 593.005 2625.970 593.335 2625.985 ;
        RECT 574.800 2625.880 593.335 2625.970 ;
        RECT 578.070 2625.670 593.335 2625.880 ;
        RECT 593.005 2625.655 593.335 2625.670 ;
        RECT 627.030 1939.850 631.030 1940.000 ;
        RECT 642.685 1939.850 643.015 1939.865 ;
        RECT 645.445 1939.850 645.775 1939.865 ;
        RECT 627.030 1939.550 645.775 1939.850 ;
        RECT 627.030 1939.400 631.030 1939.550 ;
        RECT 642.685 1939.535 643.015 1939.550 ;
        RECT 645.445 1939.535 645.775 1939.550 ;
        RECT 644.065 628.130 644.395 628.145 ;
        RECT 645.445 628.130 645.775 628.145 ;
        RECT 644.065 627.830 645.775 628.130 ;
        RECT 644.065 627.815 644.395 627.830 ;
        RECT 645.445 627.815 645.775 627.830 ;
        RECT 644.065 579.850 644.395 579.865 ;
        RECT 644.985 579.850 645.315 579.865 ;
        RECT 644.065 579.550 645.315 579.850 ;
        RECT 644.065 579.535 644.395 579.550 ;
        RECT 644.985 579.535 645.315 579.550 ;
        RECT 643.605 531.570 643.935 531.585 ;
        RECT 644.525 531.570 644.855 531.585 ;
        RECT 643.605 531.270 644.855 531.570 ;
        RECT 643.605 531.255 643.935 531.270 ;
        RECT 644.525 531.255 644.855 531.270 ;
        RECT 644.525 339.130 644.855 339.145 ;
        RECT 644.525 338.830 646.450 339.130 ;
        RECT 644.525 338.815 644.855 338.830 ;
        RECT 645.445 338.450 645.775 338.465 ;
        RECT 646.150 338.450 646.450 338.830 ;
        RECT 645.445 338.150 646.450 338.450 ;
        RECT 645.445 338.135 645.775 338.150 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 2504.680 482.930 2504.740 ;
        RECT 1901.710 2504.680 1902.030 2504.740 ;
        RECT 482.610 2504.540 1902.030 2504.680 ;
        RECT 482.610 2504.480 482.930 2504.540 ;
        RECT 1901.710 2504.480 1902.030 2504.540 ;
        RECT 351.510 2501.280 351.830 2501.340 ;
        RECT 476.170 2501.280 476.490 2501.340 ;
        RECT 482.610 2501.280 482.930 2501.340 ;
        RECT 351.510 2501.140 482.930 2501.280 ;
        RECT 351.510 2501.080 351.830 2501.140 ;
        RECT 476.170 2501.080 476.490 2501.140 ;
        RECT 482.610 2501.080 482.930 2501.140 ;
        RECT 337.710 587.420 338.030 587.480 ;
        RECT 355.190 587.420 355.510 587.480 ;
        RECT 841.870 587.420 842.190 587.480 ;
        RECT 337.710 587.280 842.190 587.420 ;
        RECT 337.710 587.220 338.030 587.280 ;
        RECT 355.190 587.220 355.510 587.280 ;
        RECT 841.870 587.220 842.190 587.280 ;
      LAYER via ;
        RECT 482.640 2504.480 482.900 2504.740 ;
        RECT 1901.740 2504.480 1902.000 2504.740 ;
        RECT 351.540 2501.080 351.800 2501.340 ;
        RECT 476.200 2501.080 476.460 2501.340 ;
        RECT 482.640 2501.080 482.900 2501.340 ;
        RECT 337.740 587.220 338.000 587.480 ;
        RECT 355.220 587.220 355.480 587.480 ;
        RECT 841.900 587.220 842.160 587.480 ;
      LAYER met2 ;
        RECT 476.090 2600.660 476.370 2604.000 ;
        RECT 476.090 2600.000 476.400 2600.660 ;
        RECT 476.260 2501.370 476.400 2600.000 ;
        RECT 1901.730 2532.475 1902.010 2532.845 ;
        RECT 1901.800 2504.770 1901.940 2532.475 ;
        RECT 482.640 2504.450 482.900 2504.770 ;
        RECT 1901.740 2504.450 1902.000 2504.770 ;
        RECT 482.700 2501.370 482.840 2504.450 ;
        RECT 351.540 2501.050 351.800 2501.370 ;
        RECT 476.200 2501.050 476.460 2501.370 ;
        RECT 482.640 2501.050 482.900 2501.370 ;
        RECT 351.600 1889.565 351.740 2501.050 ;
        RECT 351.530 1889.195 351.810 1889.565 ;
        RECT 355.210 1889.195 355.490 1889.565 ;
        RECT 355.280 587.510 355.420 1889.195 ;
        RECT 842.590 600.170 842.870 604.000 ;
        RECT 841.960 600.030 842.870 600.170 ;
        RECT 841.960 587.510 842.100 600.030 ;
        RECT 842.590 600.000 842.870 600.030 ;
        RECT 337.740 587.190 338.000 587.510 ;
        RECT 355.220 587.190 355.480 587.510 ;
        RECT 841.900 587.190 842.160 587.510 ;
        RECT 337.800 24.210 337.940 587.190 ;
        RECT 335.960 24.070 337.940 24.210 ;
        RECT 335.960 2.400 336.100 24.070 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 1901.730 2532.520 1902.010 2532.800 ;
        RECT 351.530 1889.240 351.810 1889.520 ;
        RECT 355.210 1889.240 355.490 1889.520 ;
      LAYER met3 ;
        RECT 1885.335 2534.360 1889.335 2534.640 ;
        RECT 1885.335 2534.040 1889.370 2534.360 ;
        RECT 1889.070 2532.810 1889.370 2534.040 ;
        RECT 1901.705 2532.810 1902.035 2532.825 ;
        RECT 1889.070 2532.510 1902.035 2532.810 ;
        RECT 1901.705 2532.495 1902.035 2532.510 ;
        RECT 351.505 1889.530 351.835 1889.545 ;
        RECT 355.185 1889.530 355.515 1889.545 ;
        RECT 360.000 1889.530 364.000 1889.680 ;
        RECT 351.505 1889.230 364.000 1889.530 ;
        RECT 351.505 1889.215 351.835 1889.230 ;
        RECT 355.185 1889.215 355.515 1889.230 ;
        RECT 360.000 1889.080 364.000 1889.230 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 475.250 2768.860 475.570 2768.920 ;
        RECT 603.590 2768.860 603.910 2768.920 ;
        RECT 475.250 2768.720 603.910 2768.860 ;
        RECT 475.250 2768.660 475.570 2768.720 ;
        RECT 603.590 2768.660 603.910 2768.720 ;
        RECT 603.590 2490.060 603.910 2490.120 ;
        RECT 606.810 2490.060 607.130 2490.120 ;
        RECT 1694.250 2490.060 1694.570 2490.120 ;
        RECT 603.590 2489.920 1694.570 2490.060 ;
        RECT 603.590 2489.860 603.910 2489.920 ;
        RECT 606.810 2489.860 607.130 2489.920 ;
        RECT 1694.250 2489.860 1694.570 2489.920 ;
        RECT 604.510 1994.680 604.830 1994.740 ;
        RECT 606.810 1994.680 607.130 1994.740 ;
        RECT 628.430 1994.680 628.750 1994.740 ;
        RECT 604.510 1994.540 628.750 1994.680 ;
        RECT 604.510 1994.480 604.830 1994.540 ;
        RECT 606.810 1994.480 607.130 1994.540 ;
        RECT 628.430 1994.480 628.750 1994.540 ;
        RECT 603.590 592.180 603.910 592.240 ;
        RECT 628.430 592.180 628.750 592.240 ;
        RECT 850.150 592.180 850.470 592.240 ;
        RECT 603.590 592.040 850.470 592.180 ;
        RECT 603.590 591.980 603.910 592.040 ;
        RECT 628.430 591.980 628.750 592.040 ;
        RECT 850.150 591.980 850.470 592.040 ;
        RECT 353.350 22.000 353.670 22.060 ;
        RECT 603.590 22.000 603.910 22.060 ;
        RECT 353.350 21.860 603.910 22.000 ;
        RECT 353.350 21.800 353.670 21.860 ;
        RECT 603.590 21.800 603.910 21.860 ;
      LAYER via ;
        RECT 475.280 2768.660 475.540 2768.920 ;
        RECT 603.620 2768.660 603.880 2768.920 ;
        RECT 603.620 2489.860 603.880 2490.120 ;
        RECT 606.840 2489.860 607.100 2490.120 ;
        RECT 1694.280 2489.860 1694.540 2490.120 ;
        RECT 604.540 1994.480 604.800 1994.740 ;
        RECT 606.840 1994.480 607.100 1994.740 ;
        RECT 628.460 1994.480 628.720 1994.740 ;
        RECT 603.620 591.980 603.880 592.240 ;
        RECT 628.460 591.980 628.720 592.240 ;
        RECT 850.180 591.980 850.440 592.240 ;
        RECT 353.380 21.800 353.640 22.060 ;
        RECT 603.620 21.800 603.880 22.060 ;
      LAYER met2 ;
        RECT 475.280 2768.630 475.540 2768.950 ;
        RECT 603.620 2768.630 603.880 2768.950 ;
        RECT 475.340 2759.520 475.480 2768.630 ;
        RECT 475.170 2759.100 475.480 2759.520 ;
        RECT 475.170 2755.520 475.450 2759.100 ;
        RECT 603.680 2490.150 603.820 2768.630 ;
        RECT 1694.210 2500.000 1694.490 2504.000 ;
        RECT 1694.340 2490.150 1694.480 2500.000 ;
        RECT 603.620 2489.830 603.880 2490.150 ;
        RECT 606.840 2489.830 607.100 2490.150 ;
        RECT 1694.280 2489.830 1694.540 2490.150 ;
        RECT 606.900 1994.770 607.040 2489.830 ;
        RECT 604.540 1994.450 604.800 1994.770 ;
        RECT 606.840 1994.450 607.100 1994.770 ;
        RECT 628.460 1994.450 628.720 1994.770 ;
        RECT 602.970 1981.250 603.250 1981.750 ;
        RECT 604.600 1981.250 604.740 1994.450 ;
        RECT 602.970 1981.110 604.740 1981.250 ;
        RECT 602.970 1977.750 603.250 1981.110 ;
        RECT 628.520 592.270 628.660 1994.450 ;
        RECT 851.790 600.170 852.070 604.000 ;
        RECT 850.240 600.030 852.070 600.170 ;
        RECT 850.240 592.270 850.380 600.030 ;
        RECT 851.790 600.000 852.070 600.030 ;
        RECT 603.620 591.950 603.880 592.270 ;
        RECT 628.460 591.950 628.720 592.270 ;
        RECT 850.180 591.950 850.440 592.270 ;
        RECT 603.680 22.090 603.820 591.950 ;
        RECT 353.380 21.770 353.640 22.090 ;
        RECT 603.620 21.770 603.880 22.090 ;
        RECT 353.440 2.400 353.580 21.770 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 996.890 2917.440 997.210 2917.500 ;
        RECT 1588.450 2917.440 1588.770 2917.500 ;
        RECT 996.890 2917.300 1588.770 2917.440 ;
        RECT 996.890 2917.240 997.210 2917.300 ;
        RECT 1588.450 2917.240 1588.770 2917.300 ;
        RECT 427.410 2749.480 427.730 2749.540 ;
        RECT 432.010 2749.480 432.330 2749.540 ;
        RECT 996.890 2749.480 997.210 2749.540 ;
        RECT 427.410 2749.340 997.210 2749.480 ;
        RECT 427.410 2749.280 427.730 2749.340 ;
        RECT 432.010 2749.280 432.330 2749.340 ;
        RECT 996.890 2749.280 997.210 2749.340 ;
        RECT 358.410 1994.340 358.730 1994.400 ;
        RECT 427.410 1994.340 427.730 1994.400 ;
        RECT 358.410 1994.200 427.730 1994.340 ;
        RECT 358.410 1994.140 358.730 1994.200 ;
        RECT 427.410 1994.140 427.730 1994.200 ;
        RECT 427.410 1993.660 427.730 1993.720 ;
        RECT 451.330 1993.660 451.650 1993.720 ;
        RECT 427.410 1993.520 451.650 1993.660 ;
        RECT 427.410 1993.460 427.730 1993.520 ;
        RECT 451.330 1993.460 451.650 1993.520 ;
        RECT 614.170 589.800 614.490 589.860 ;
        RECT 614.170 589.660 831.980 589.800 ;
        RECT 614.170 589.600 614.490 589.660 ;
        RECT 482.610 589.120 482.930 589.180 ;
        RECT 495.950 589.120 496.270 589.180 ;
        RECT 482.610 588.980 496.270 589.120 ;
        RECT 482.610 588.920 482.930 588.980 ;
        RECT 495.950 588.920 496.270 588.980 ;
        RECT 358.410 588.780 358.730 588.840 ;
        RECT 368.990 588.780 369.310 588.840 ;
        RECT 399.810 588.780 400.130 588.840 ;
        RECT 358.410 588.640 400.130 588.780 ;
        RECT 358.410 588.580 358.730 588.640 ;
        RECT 368.990 588.580 369.310 588.640 ;
        RECT 399.810 588.580 400.130 588.640 ;
        RECT 497.330 588.780 497.650 588.840 ;
        RECT 614.170 588.780 614.490 588.840 ;
        RECT 497.330 588.640 544.940 588.780 ;
        RECT 497.330 588.580 497.650 588.640 ;
        RECT 400.730 588.440 401.050 588.500 ;
        RECT 434.770 588.440 435.090 588.500 ;
        RECT 400.730 588.300 435.090 588.440 ;
        RECT 544.800 588.440 544.940 588.640 ;
        RECT 545.260 588.640 614.490 588.780 ;
        RECT 545.260 588.440 545.400 588.640 ;
        RECT 614.170 588.580 614.490 588.640 ;
        RECT 544.800 588.300 545.400 588.440 ;
        RECT 400.730 588.240 401.050 588.300 ;
        RECT 434.770 588.240 435.090 588.300 ;
        RECT 831.840 588.100 831.980 589.660 ;
        RECT 859.350 588.100 859.670 588.160 ;
        RECT 831.840 587.960 859.670 588.100 ;
        RECT 859.350 587.900 859.670 587.960 ;
        RECT 434.770 587.760 435.090 587.820 ;
        RECT 482.610 587.760 482.930 587.820 ;
        RECT 434.770 587.620 482.930 587.760 ;
        RECT 434.770 587.560 435.090 587.620 ;
        RECT 482.610 587.560 482.930 587.620 ;
        RECT 368.990 16.900 369.310 16.960 ;
        RECT 371.290 16.900 371.610 16.960 ;
        RECT 368.990 16.760 371.610 16.900 ;
        RECT 368.990 16.700 369.310 16.760 ;
        RECT 371.290 16.700 371.610 16.760 ;
      LAYER via ;
        RECT 996.920 2917.240 997.180 2917.500 ;
        RECT 1588.480 2917.240 1588.740 2917.500 ;
        RECT 427.440 2749.280 427.700 2749.540 ;
        RECT 432.040 2749.280 432.300 2749.540 ;
        RECT 996.920 2749.280 997.180 2749.540 ;
        RECT 358.440 1994.140 358.700 1994.400 ;
        RECT 427.440 1994.140 427.700 1994.400 ;
        RECT 427.440 1993.460 427.700 1993.720 ;
        RECT 451.360 1993.460 451.620 1993.720 ;
        RECT 614.200 589.600 614.460 589.860 ;
        RECT 482.640 588.920 482.900 589.180 ;
        RECT 495.980 588.920 496.240 589.180 ;
        RECT 358.440 588.580 358.700 588.840 ;
        RECT 369.020 588.580 369.280 588.840 ;
        RECT 399.840 588.580 400.100 588.840 ;
        RECT 497.360 588.580 497.620 588.840 ;
        RECT 400.760 588.240 401.020 588.500 ;
        RECT 434.800 588.240 435.060 588.500 ;
        RECT 614.200 588.580 614.460 588.840 ;
        RECT 859.380 587.900 859.640 588.160 ;
        RECT 434.800 587.560 435.060 587.820 ;
        RECT 482.640 587.560 482.900 587.820 ;
        RECT 369.020 16.700 369.280 16.960 ;
        RECT 371.320 16.700 371.580 16.960 ;
      LAYER met2 ;
        RECT 996.920 2917.210 997.180 2917.530 ;
        RECT 1588.480 2917.210 1588.740 2917.530 ;
        RECT 427.440 2749.250 427.700 2749.570 ;
        RECT 432.030 2749.395 432.310 2749.765 ;
        RECT 996.980 2749.570 997.120 2917.210 ;
        RECT 1588.540 2900.055 1588.680 2917.210 ;
        RECT 1588.410 2896.055 1588.690 2900.055 ;
        RECT 432.040 2749.250 432.300 2749.395 ;
        RECT 996.920 2749.250 997.180 2749.570 ;
        RECT 427.500 1994.430 427.640 2749.250 ;
        RECT 358.440 1994.110 358.700 1994.430 ;
        RECT 427.440 1994.110 427.700 1994.430 ;
        RECT 358.500 588.870 358.640 1994.110 ;
        RECT 427.500 1993.750 427.640 1994.110 ;
        RECT 427.440 1993.430 427.700 1993.750 ;
        RECT 451.360 1993.430 451.620 1993.750 ;
        RECT 451.420 1981.250 451.560 1993.430 ;
        RECT 453.010 1981.250 453.290 1981.750 ;
        RECT 451.420 1981.110 453.290 1981.250 ;
        RECT 453.010 1977.750 453.290 1981.110 ;
        RECT 860.990 600.170 861.270 604.000 ;
        RECT 859.440 600.030 861.270 600.170 ;
        RECT 614.200 589.570 614.460 589.890 ;
        RECT 482.640 588.890 482.900 589.210 ;
        RECT 495.980 588.890 496.240 589.210 ;
        RECT 358.440 588.550 358.700 588.870 ;
        RECT 369.020 588.550 369.280 588.870 ;
        RECT 399.840 588.610 400.100 588.870 ;
        RECT 399.840 588.550 400.960 588.610 ;
        RECT 369.080 16.990 369.220 588.550 ;
        RECT 399.900 588.530 400.960 588.550 ;
        RECT 399.900 588.470 401.020 588.530 ;
        RECT 400.760 588.210 401.020 588.470 ;
        RECT 434.800 588.210 435.060 588.530 ;
        RECT 434.860 587.850 435.000 588.210 ;
        RECT 482.700 587.850 482.840 588.890 ;
        RECT 496.040 588.610 496.180 588.890 ;
        RECT 614.260 588.870 614.400 589.570 ;
        RECT 497.360 588.610 497.620 588.870 ;
        RECT 496.040 588.550 497.620 588.610 ;
        RECT 614.200 588.550 614.460 588.870 ;
        RECT 496.040 588.470 497.560 588.550 ;
        RECT 859.440 588.190 859.580 600.030 ;
        RECT 860.990 600.000 861.270 600.030 ;
        RECT 859.380 587.870 859.640 588.190 ;
        RECT 434.800 587.530 435.060 587.850 ;
        RECT 482.640 587.530 482.900 587.850 ;
        RECT 369.020 16.670 369.280 16.990 ;
        RECT 371.320 16.670 371.580 16.990 ;
        RECT 371.380 2.400 371.520 16.670 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 432.030 2749.440 432.310 2749.720 ;
      LAYER met3 ;
        RECT 430.000 2752.360 434.000 2752.960 ;
        RECT 431.790 2749.745 432.090 2752.360 ;
        RECT 431.790 2749.430 432.335 2749.745 ;
        RECT 432.005 2749.415 432.335 2749.430 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 503.770 2768.520 504.090 2768.580 ;
        RECT 645.910 2768.520 646.230 2768.580 ;
        RECT 503.770 2768.380 646.230 2768.520 ;
        RECT 503.770 2768.320 504.090 2768.380 ;
        RECT 645.910 2768.320 646.230 2768.380 ;
        RECT 645.910 2484.280 646.230 2484.340 ;
        RECT 1821.210 2484.280 1821.530 2484.340 ;
        RECT 645.910 2484.140 1821.530 2484.280 ;
        RECT 645.910 2484.080 646.230 2484.140 ;
        RECT 1821.210 2484.080 1821.530 2484.140 ;
        RECT 645.910 627.680 646.230 627.940 ;
        RECT 646.000 627.260 646.140 627.680 ;
        RECT 645.910 627.000 646.230 627.260 ;
        RECT 666.150 590.480 666.470 590.540 ;
        RECT 869.470 590.480 869.790 590.540 ;
        RECT 666.150 590.340 869.790 590.480 ;
        RECT 666.150 590.280 666.470 590.340 ;
        RECT 869.470 590.280 869.790 590.340 ;
        RECT 389.230 44.100 389.550 44.160 ;
        RECT 389.230 43.960 630.040 44.100 ;
        RECT 389.230 43.900 389.550 43.960 ;
        RECT 629.900 43.760 630.040 43.960 ;
        RECT 645.910 43.760 646.230 43.820 ;
        RECT 629.900 43.620 646.230 43.760 ;
        RECT 645.910 43.560 646.230 43.620 ;
      LAYER via ;
        RECT 503.800 2768.320 504.060 2768.580 ;
        RECT 645.940 2768.320 646.200 2768.580 ;
        RECT 645.940 2484.080 646.200 2484.340 ;
        RECT 1821.240 2484.080 1821.500 2484.340 ;
        RECT 645.940 627.680 646.200 627.940 ;
        RECT 645.940 627.000 646.200 627.260 ;
        RECT 666.180 590.280 666.440 590.540 ;
        RECT 869.500 590.280 869.760 590.540 ;
        RECT 389.260 43.900 389.520 44.160 ;
        RECT 645.940 43.560 646.200 43.820 ;
      LAYER met2 ;
        RECT 503.800 2768.290 504.060 2768.610 ;
        RECT 645.940 2768.290 646.200 2768.610 ;
        RECT 503.860 2759.520 504.000 2768.290 ;
        RECT 503.690 2759.100 504.000 2759.520 ;
        RECT 503.690 2755.520 503.970 2759.100 ;
        RECT 646.000 2484.370 646.140 2768.290 ;
        RECT 1821.170 2500.000 1821.450 2504.000 ;
        RECT 1821.300 2484.370 1821.440 2500.000 ;
        RECT 645.940 2484.050 646.200 2484.370 ;
        RECT 1821.240 2484.050 1821.500 2484.370 ;
        RECT 646.000 1903.165 646.140 2484.050 ;
        RECT 645.930 1902.795 646.210 1903.165 ;
        RECT 646.000 627.970 646.140 1902.795 ;
        RECT 645.940 627.650 646.200 627.970 ;
        RECT 645.940 626.970 646.200 627.290 ;
        RECT 646.000 590.765 646.140 626.970 ;
        RECT 870.190 600.170 870.470 604.000 ;
        RECT 869.560 600.030 870.470 600.170 ;
        RECT 645.930 590.395 646.210 590.765 ;
        RECT 666.170 590.395 666.450 590.765 ;
        RECT 869.560 590.570 869.700 600.030 ;
        RECT 870.190 600.000 870.470 600.030 ;
        RECT 389.260 43.870 389.520 44.190 ;
        RECT 389.320 2.400 389.460 43.870 ;
        RECT 646.000 43.850 646.140 590.395 ;
        RECT 666.180 590.250 666.440 590.395 ;
        RECT 869.500 590.250 869.760 590.570 ;
        RECT 645.940 43.530 646.200 43.850 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 645.930 1902.840 646.210 1903.120 ;
        RECT 645.930 590.440 646.210 590.720 ;
        RECT 666.170 590.440 666.450 590.720 ;
      LAYER met3 ;
        RECT 627.030 1903.130 631.030 1903.280 ;
        RECT 645.905 1903.130 646.235 1903.145 ;
        RECT 627.030 1902.830 646.235 1903.130 ;
        RECT 627.030 1902.680 631.030 1902.830 ;
        RECT 645.905 1902.815 646.235 1902.830 ;
        RECT 645.905 590.730 646.235 590.745 ;
        RECT 666.145 590.730 666.475 590.745 ;
        RECT 645.905 590.430 666.475 590.730 ;
        RECT 645.905 590.415 646.235 590.430 ;
        RECT 666.145 590.415 666.475 590.430 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 2487.680 419.450 2487.740 ;
        RECT 635.790 2487.680 636.110 2487.740 ;
        RECT 1800.050 2487.680 1800.370 2487.740 ;
        RECT 419.130 2487.540 1800.370 2487.680 ;
        RECT 419.130 2487.480 419.450 2487.540 ;
        RECT 635.790 2487.480 636.110 2487.540 ;
        RECT 1800.050 2487.480 1800.370 2487.540 ;
        RECT 564.030 1689.700 564.350 1689.760 ;
        RECT 565.410 1689.700 565.730 1689.760 ;
        RECT 635.790 1689.700 636.110 1689.760 ;
        RECT 564.030 1689.560 636.110 1689.700 ;
        RECT 564.030 1689.500 564.350 1689.560 ;
        RECT 565.410 1689.500 565.730 1689.560 ;
        RECT 635.790 1689.500 636.110 1689.560 ;
        RECT 565.410 591.160 565.730 591.220 ;
        RECT 877.750 591.160 878.070 591.220 ;
        RECT 565.410 591.020 878.070 591.160 ;
        RECT 565.410 590.960 565.730 591.020 ;
        RECT 877.750 590.960 878.070 591.020 ;
        RECT 548.390 586.740 548.710 586.800 ;
        RECT 565.410 586.740 565.730 586.800 ;
        RECT 548.390 586.600 565.730 586.740 ;
        RECT 548.390 586.540 548.710 586.600 ;
        RECT 565.410 586.540 565.730 586.600 ;
        RECT 407.170 29.140 407.490 29.200 ;
        RECT 548.390 29.140 548.710 29.200 ;
        RECT 407.170 29.000 548.710 29.140 ;
        RECT 407.170 28.940 407.490 29.000 ;
        RECT 548.390 28.940 548.710 29.000 ;
      LAYER via ;
        RECT 419.160 2487.480 419.420 2487.740 ;
        RECT 635.820 2487.480 636.080 2487.740 ;
        RECT 1800.080 2487.480 1800.340 2487.740 ;
        RECT 564.060 1689.500 564.320 1689.760 ;
        RECT 565.440 1689.500 565.700 1689.760 ;
        RECT 635.820 1689.500 636.080 1689.760 ;
        RECT 565.440 590.960 565.700 591.220 ;
        RECT 877.780 590.960 878.040 591.220 ;
        RECT 548.420 586.540 548.680 586.800 ;
        RECT 565.440 586.540 565.700 586.800 ;
        RECT 407.200 28.940 407.460 29.200 ;
        RECT 548.420 28.940 548.680 29.200 ;
      LAYER met2 ;
        RECT 419.150 2643.315 419.430 2643.685 ;
        RECT 419.220 2487.770 419.360 2643.315 ;
        RECT 1800.010 2500.000 1800.290 2504.000 ;
        RECT 1800.140 2487.770 1800.280 2500.000 ;
        RECT 419.160 2487.450 419.420 2487.770 ;
        RECT 635.820 2487.450 636.080 2487.770 ;
        RECT 1800.080 2487.450 1800.340 2487.770 ;
        RECT 562.490 1700.410 562.770 1704.000 ;
        RECT 562.490 1700.270 564.260 1700.410 ;
        RECT 562.490 1700.000 562.770 1700.270 ;
        RECT 564.120 1689.790 564.260 1700.270 ;
        RECT 635.880 1689.790 636.020 2487.450 ;
        RECT 564.060 1689.470 564.320 1689.790 ;
        RECT 565.440 1689.470 565.700 1689.790 ;
        RECT 635.820 1689.470 636.080 1689.790 ;
        RECT 565.500 591.250 565.640 1689.470 ;
        RECT 879.390 600.170 879.670 604.000 ;
        RECT 877.840 600.030 879.670 600.170 ;
        RECT 877.840 591.250 877.980 600.030 ;
        RECT 879.390 600.000 879.670 600.030 ;
        RECT 565.440 590.930 565.700 591.250 ;
        RECT 877.780 590.930 878.040 591.250 ;
        RECT 565.500 586.830 565.640 590.930 ;
        RECT 548.420 586.510 548.680 586.830 ;
        RECT 565.440 586.510 565.700 586.830 ;
        RECT 548.480 29.230 548.620 586.510 ;
        RECT 407.200 28.910 407.460 29.230 ;
        RECT 548.420 28.910 548.680 29.230 ;
        RECT 407.260 2.400 407.400 28.910 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 419.150 2643.360 419.430 2643.640 ;
      LAYER met3 ;
        RECT 430.000 2646.560 434.000 2646.880 ;
        RECT 429.950 2646.280 434.000 2646.560 ;
        RECT 419.125 2643.650 419.455 2643.665 ;
        RECT 429.950 2643.650 430.250 2646.280 ;
        RECT 419.125 2643.350 430.250 2643.650 ;
        RECT 419.125 2643.335 419.455 2643.350 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1682.750 2897.040 1683.070 2897.100 ;
        RECT 1651.100 2896.900 1683.070 2897.040 ;
        RECT 1548.890 2896.500 1549.210 2896.760 ;
        RECT 1549.810 2896.700 1550.130 2896.760 ;
        RECT 1549.810 2896.560 1550.500 2896.700 ;
        RECT 1549.810 2896.500 1550.130 2896.560 ;
        RECT 786.670 2895.340 786.990 2895.400 ;
        RECT 811.970 2895.340 812.290 2895.400 ;
        RECT 786.670 2895.200 812.290 2895.340 ;
        RECT 786.670 2895.140 786.990 2895.200 ;
        RECT 811.970 2895.140 812.290 2895.200 ;
        RECT 883.270 2895.340 883.590 2895.400 ;
        RECT 908.570 2895.340 908.890 2895.400 ;
        RECT 883.270 2895.200 908.890 2895.340 ;
        RECT 883.270 2895.140 883.590 2895.200 ;
        RECT 908.570 2895.140 908.890 2895.200 ;
        RECT 979.870 2895.340 980.190 2895.400 ;
        RECT 1005.170 2895.340 1005.490 2895.400 ;
        RECT 979.870 2895.200 1005.490 2895.340 ;
        RECT 979.870 2895.140 980.190 2895.200 ;
        RECT 1005.170 2895.140 1005.490 2895.200 ;
        RECT 1076.470 2895.340 1076.790 2895.400 ;
        RECT 1101.770 2895.340 1102.090 2895.400 ;
        RECT 1076.470 2895.200 1102.090 2895.340 ;
        RECT 1076.470 2895.140 1076.790 2895.200 ;
        RECT 1101.770 2895.140 1102.090 2895.200 ;
        RECT 1173.070 2895.340 1173.390 2895.400 ;
        RECT 1198.370 2895.340 1198.690 2895.400 ;
        RECT 1173.070 2895.200 1198.690 2895.340 ;
        RECT 1173.070 2895.140 1173.390 2895.200 ;
        RECT 1198.370 2895.140 1198.690 2895.200 ;
        RECT 1269.670 2895.340 1269.990 2895.400 ;
        RECT 1294.970 2895.340 1295.290 2895.400 ;
        RECT 1269.670 2895.200 1295.290 2895.340 ;
        RECT 1269.670 2895.140 1269.990 2895.200 ;
        RECT 1294.970 2895.140 1295.290 2895.200 ;
        RECT 628.430 2894.660 628.750 2894.720 ;
        RECT 689.150 2894.660 689.470 2894.720 ;
        RECT 628.430 2894.520 689.470 2894.660 ;
        RECT 628.430 2894.460 628.750 2894.520 ;
        RECT 689.150 2894.460 689.470 2894.520 ;
        RECT 761.830 2894.660 762.150 2894.720 ;
        RECT 786.210 2894.660 786.530 2894.720 ;
        RECT 761.830 2894.520 786.530 2894.660 ;
        RECT 761.830 2894.460 762.150 2894.520 ;
        RECT 786.210 2894.460 786.530 2894.520 ;
        RECT 858.430 2894.660 858.750 2894.720 ;
        RECT 882.810 2894.660 883.130 2894.720 ;
        RECT 858.430 2894.520 883.130 2894.660 ;
        RECT 858.430 2894.460 858.750 2894.520 ;
        RECT 882.810 2894.460 883.130 2894.520 ;
        RECT 955.030 2894.660 955.350 2894.720 ;
        RECT 979.410 2894.660 979.730 2894.720 ;
        RECT 955.030 2894.520 979.730 2894.660 ;
        RECT 955.030 2894.460 955.350 2894.520 ;
        RECT 979.410 2894.460 979.730 2894.520 ;
        RECT 1051.630 2894.660 1051.950 2894.720 ;
        RECT 1076.010 2894.660 1076.330 2894.720 ;
        RECT 1051.630 2894.520 1076.330 2894.660 ;
        RECT 1051.630 2894.460 1051.950 2894.520 ;
        RECT 1076.010 2894.460 1076.330 2894.520 ;
        RECT 1148.230 2894.660 1148.550 2894.720 ;
        RECT 1172.610 2894.660 1172.930 2894.720 ;
        RECT 1148.230 2894.520 1172.930 2894.660 ;
        RECT 1148.230 2894.460 1148.550 2894.520 ;
        RECT 1172.610 2894.460 1172.930 2894.520 ;
        RECT 1244.830 2894.660 1245.150 2894.720 ;
        RECT 1269.210 2894.660 1269.530 2894.720 ;
        RECT 1244.830 2894.520 1269.530 2894.660 ;
        RECT 1244.830 2894.460 1245.150 2894.520 ;
        RECT 1269.210 2894.460 1269.530 2894.520 ;
        RECT 1341.430 2894.660 1341.750 2894.720 ;
        RECT 1365.810 2894.660 1366.130 2894.720 ;
        RECT 1341.430 2894.520 1366.130 2894.660 ;
        RECT 1341.430 2894.460 1341.750 2894.520 ;
        RECT 1365.810 2894.460 1366.130 2894.520 ;
        RECT 1548.980 2893.640 1549.120 2896.500 ;
        RECT 1550.360 2895.340 1550.500 2896.560 ;
        RECT 1651.100 2895.680 1651.240 2896.900 ;
        RECT 1682.750 2896.840 1683.070 2896.900 ;
        RECT 1645.120 2895.540 1651.240 2895.680 ;
        RECT 1645.120 2895.340 1645.260 2895.540 ;
        RECT 1550.360 2895.200 1645.260 2895.340 ;
        RECT 1520.920 2893.500 1549.120 2893.640 ;
        RECT 690.530 2893.300 690.850 2893.360 ;
        RECT 697.890 2893.300 698.210 2893.360 ;
        RECT 690.530 2893.160 698.210 2893.300 ;
        RECT 690.530 2893.100 690.850 2893.160 ;
        RECT 697.890 2893.100 698.210 2893.160 ;
        RECT 1472.530 2892.960 1472.850 2893.020 ;
        RECT 1520.920 2892.960 1521.060 2893.500 ;
        RECT 1472.530 2892.820 1521.060 2892.960 ;
        RECT 1472.530 2892.760 1472.850 2892.820 ;
        RECT 596.690 2892.620 597.010 2892.680 ;
        RECT 628.430 2892.620 628.750 2892.680 ;
        RECT 596.690 2892.480 628.750 2892.620 ;
        RECT 596.690 2892.420 597.010 2892.480 ;
        RECT 628.430 2892.420 628.750 2892.480 ;
        RECT 689.610 2892.620 689.930 2892.680 ;
        RECT 690.070 2892.620 690.390 2892.680 ;
        RECT 689.610 2892.480 690.390 2892.620 ;
        RECT 689.610 2892.420 689.930 2892.480 ;
        RECT 690.070 2892.420 690.390 2892.480 ;
        RECT 786.210 2892.620 786.530 2892.680 ;
        RECT 786.670 2892.620 786.990 2892.680 ;
        RECT 786.210 2892.480 786.990 2892.620 ;
        RECT 786.210 2892.420 786.530 2892.480 ;
        RECT 786.670 2892.420 786.990 2892.480 ;
        RECT 882.810 2892.620 883.130 2892.680 ;
        RECT 883.270 2892.620 883.590 2892.680 ;
        RECT 882.810 2892.480 883.590 2892.620 ;
        RECT 882.810 2892.420 883.130 2892.480 ;
        RECT 883.270 2892.420 883.590 2892.480 ;
        RECT 979.410 2892.620 979.730 2892.680 ;
        RECT 979.870 2892.620 980.190 2892.680 ;
        RECT 979.410 2892.480 980.190 2892.620 ;
        RECT 979.410 2892.420 979.730 2892.480 ;
        RECT 979.870 2892.420 980.190 2892.480 ;
        RECT 1076.010 2892.620 1076.330 2892.680 ;
        RECT 1076.470 2892.620 1076.790 2892.680 ;
        RECT 1076.010 2892.480 1076.790 2892.620 ;
        RECT 1076.010 2892.420 1076.330 2892.480 ;
        RECT 1076.470 2892.420 1076.790 2892.480 ;
        RECT 1172.610 2892.620 1172.930 2892.680 ;
        RECT 1173.070 2892.620 1173.390 2892.680 ;
        RECT 1172.610 2892.480 1173.390 2892.620 ;
        RECT 1172.610 2892.420 1172.930 2892.480 ;
        RECT 1173.070 2892.420 1173.390 2892.480 ;
        RECT 1269.210 2892.620 1269.530 2892.680 ;
        RECT 1269.670 2892.620 1269.990 2892.680 ;
        RECT 1269.210 2892.480 1269.990 2892.620 ;
        RECT 1269.210 2892.420 1269.530 2892.480 ;
        RECT 1269.670 2892.420 1269.990 2892.480 ;
        RECT 1365.810 2892.620 1366.130 2892.680 ;
        RECT 1365.810 2892.480 1414.340 2892.620 ;
        RECT 1365.810 2892.420 1366.130 2892.480 ;
        RECT 697.890 2892.280 698.210 2892.340 ;
        RECT 761.830 2892.280 762.150 2892.340 ;
        RECT 697.890 2892.140 762.150 2892.280 ;
        RECT 697.890 2892.080 698.210 2892.140 ;
        RECT 761.830 2892.080 762.150 2892.140 ;
        RECT 811.970 2892.280 812.290 2892.340 ;
        RECT 858.430 2892.280 858.750 2892.340 ;
        RECT 811.970 2892.140 858.750 2892.280 ;
        RECT 811.970 2892.080 812.290 2892.140 ;
        RECT 858.430 2892.080 858.750 2892.140 ;
        RECT 908.570 2892.280 908.890 2892.340 ;
        RECT 955.030 2892.280 955.350 2892.340 ;
        RECT 908.570 2892.140 955.350 2892.280 ;
        RECT 908.570 2892.080 908.890 2892.140 ;
        RECT 955.030 2892.080 955.350 2892.140 ;
        RECT 1005.170 2892.280 1005.490 2892.340 ;
        RECT 1051.630 2892.280 1051.950 2892.340 ;
        RECT 1005.170 2892.140 1051.950 2892.280 ;
        RECT 1005.170 2892.080 1005.490 2892.140 ;
        RECT 1051.630 2892.080 1051.950 2892.140 ;
        RECT 1101.770 2892.280 1102.090 2892.340 ;
        RECT 1148.230 2892.280 1148.550 2892.340 ;
        RECT 1101.770 2892.140 1148.550 2892.280 ;
        RECT 1101.770 2892.080 1102.090 2892.140 ;
        RECT 1148.230 2892.080 1148.550 2892.140 ;
        RECT 1198.370 2892.280 1198.690 2892.340 ;
        RECT 1244.830 2892.280 1245.150 2892.340 ;
        RECT 1198.370 2892.140 1245.150 2892.280 ;
        RECT 1198.370 2892.080 1198.690 2892.140 ;
        RECT 1244.830 2892.080 1245.150 2892.140 ;
        RECT 1294.970 2892.280 1295.290 2892.340 ;
        RECT 1341.430 2892.280 1341.750 2892.340 ;
        RECT 1294.970 2892.140 1341.750 2892.280 ;
        RECT 1414.200 2892.280 1414.340 2892.480 ;
        RECT 1472.530 2892.280 1472.850 2892.340 ;
        RECT 1414.200 2892.140 1472.850 2892.280 ;
        RECT 1294.970 2892.080 1295.290 2892.140 ;
        RECT 1341.430 2892.080 1341.750 2892.140 ;
        RECT 1472.530 2892.080 1472.850 2892.140 ;
        RECT 589.790 2649.520 590.110 2649.580 ;
        RECT 596.690 2649.520 597.010 2649.580 ;
        RECT 589.790 2649.380 597.010 2649.520 ;
        RECT 589.790 2649.320 590.110 2649.380 ;
        RECT 596.690 2649.320 597.010 2649.380 ;
        RECT 357.490 1983.800 357.810 1983.860 ;
        RECT 589.790 1983.800 590.110 1983.860 ;
        RECT 631.650 1983.800 631.970 1983.860 ;
        RECT 357.490 1983.660 631.970 1983.800 ;
        RECT 357.490 1983.600 357.810 1983.660 ;
        RECT 589.790 1983.600 590.110 1983.660 ;
        RECT 631.650 1983.600 631.970 1983.660 ;
        RECT 631.650 1924.980 631.970 1925.040 ;
        RECT 651.430 1924.980 651.750 1925.040 ;
        RECT 631.650 1924.840 651.750 1924.980 ;
        RECT 631.650 1924.780 631.970 1924.840 ;
        RECT 651.430 1924.780 651.750 1924.840 ;
        RECT 651.430 1732.540 651.750 1732.600 ;
        RECT 663.850 1732.540 664.170 1732.600 ;
        RECT 651.430 1732.400 664.170 1732.540 ;
        RECT 651.430 1732.340 651.750 1732.400 ;
        RECT 663.850 1732.340 664.170 1732.400 ;
        RECT 663.850 1702.960 664.170 1703.020 ;
        RECT 1918.270 1702.960 1918.590 1703.020 ;
        RECT 663.850 1702.820 1918.590 1702.960 ;
        RECT 663.850 1702.760 664.170 1702.820 ;
        RECT 1918.270 1702.760 1918.590 1702.820 ;
        RECT 663.390 1607.760 663.710 1607.820 ;
        RECT 664.310 1607.760 664.630 1607.820 ;
        RECT 663.390 1607.620 664.630 1607.760 ;
        RECT 663.390 1607.560 663.710 1607.620 ;
        RECT 664.310 1607.560 664.630 1607.620 ;
        RECT 662.010 1593.820 662.330 1593.880 ;
        RECT 664.310 1593.820 664.630 1593.880 ;
        RECT 662.010 1593.680 664.630 1593.820 ;
        RECT 662.010 1593.620 662.330 1593.680 ;
        RECT 664.310 1593.620 664.630 1593.680 ;
        RECT 662.010 1545.880 662.330 1545.940 ;
        RECT 663.850 1545.880 664.170 1545.940 ;
        RECT 662.010 1545.740 664.170 1545.880 ;
        RECT 662.010 1545.680 662.330 1545.740 ;
        RECT 663.850 1545.680 664.170 1545.740 ;
        RECT 663.390 1414.640 663.710 1414.700 ;
        RECT 664.310 1414.640 664.630 1414.700 ;
        RECT 663.390 1414.500 664.630 1414.640 ;
        RECT 663.390 1414.440 663.710 1414.500 ;
        RECT 664.310 1414.440 664.630 1414.500 ;
        RECT 664.310 1052.200 664.630 1052.260 ;
        RECT 667.530 1052.200 667.850 1052.260 ;
        RECT 664.310 1052.060 667.850 1052.200 ;
        RECT 664.310 1052.000 664.630 1052.060 ;
        RECT 667.530 1052.000 667.850 1052.060 ;
        RECT 664.310 926.060 664.630 926.120 ;
        RECT 665.690 926.060 666.010 926.120 ;
        RECT 664.310 925.920 666.010 926.060 ;
        RECT 664.310 925.860 664.630 925.920 ;
        RECT 665.690 925.860 666.010 925.920 ;
        RECT 664.310 675.960 664.630 676.220 ;
        RECT 664.400 675.820 664.540 675.960 ;
        RECT 664.770 675.820 665.090 675.880 ;
        RECT 664.400 675.680 665.090 675.820 ;
        RECT 664.770 675.620 665.090 675.680 ;
        RECT 665.690 497.120 666.010 497.380 ;
        RECT 665.780 496.700 665.920 497.120 ;
        RECT 665.690 496.440 666.010 496.700 ;
        RECT 665.690 338.200 666.010 338.260 ;
        RECT 666.150 338.200 666.470 338.260 ;
        RECT 665.690 338.060 666.470 338.200 ;
        RECT 665.690 338.000 666.010 338.060 ;
        RECT 666.150 338.000 666.470 338.060 ;
        RECT 664.770 289.580 665.090 289.640 ;
        RECT 666.150 289.580 666.470 289.640 ;
        RECT 664.770 289.440 666.470 289.580 ;
        RECT 664.770 289.380 665.090 289.440 ;
        RECT 666.150 289.380 666.470 289.440 ;
        RECT 664.770 193.020 665.090 193.080 ;
        RECT 666.150 193.020 666.470 193.080 ;
        RECT 664.770 192.880 666.470 193.020 ;
        RECT 664.770 192.820 665.090 192.880 ;
        RECT 666.150 192.820 666.470 192.880 ;
        RECT 68.150 45.460 68.470 45.520 ;
        RECT 665.230 45.460 665.550 45.520 ;
        RECT 68.150 45.320 665.550 45.460 ;
        RECT 68.150 45.260 68.470 45.320 ;
        RECT 665.230 45.260 665.550 45.320 ;
      LAYER via ;
        RECT 1548.920 2896.500 1549.180 2896.760 ;
        RECT 1549.840 2896.500 1550.100 2896.760 ;
        RECT 786.700 2895.140 786.960 2895.400 ;
        RECT 812.000 2895.140 812.260 2895.400 ;
        RECT 883.300 2895.140 883.560 2895.400 ;
        RECT 908.600 2895.140 908.860 2895.400 ;
        RECT 979.900 2895.140 980.160 2895.400 ;
        RECT 1005.200 2895.140 1005.460 2895.400 ;
        RECT 1076.500 2895.140 1076.760 2895.400 ;
        RECT 1101.800 2895.140 1102.060 2895.400 ;
        RECT 1173.100 2895.140 1173.360 2895.400 ;
        RECT 1198.400 2895.140 1198.660 2895.400 ;
        RECT 1269.700 2895.140 1269.960 2895.400 ;
        RECT 1295.000 2895.140 1295.260 2895.400 ;
        RECT 628.460 2894.460 628.720 2894.720 ;
        RECT 689.180 2894.460 689.440 2894.720 ;
        RECT 761.860 2894.460 762.120 2894.720 ;
        RECT 786.240 2894.460 786.500 2894.720 ;
        RECT 858.460 2894.460 858.720 2894.720 ;
        RECT 882.840 2894.460 883.100 2894.720 ;
        RECT 955.060 2894.460 955.320 2894.720 ;
        RECT 979.440 2894.460 979.700 2894.720 ;
        RECT 1051.660 2894.460 1051.920 2894.720 ;
        RECT 1076.040 2894.460 1076.300 2894.720 ;
        RECT 1148.260 2894.460 1148.520 2894.720 ;
        RECT 1172.640 2894.460 1172.900 2894.720 ;
        RECT 1244.860 2894.460 1245.120 2894.720 ;
        RECT 1269.240 2894.460 1269.500 2894.720 ;
        RECT 1341.460 2894.460 1341.720 2894.720 ;
        RECT 1365.840 2894.460 1366.100 2894.720 ;
        RECT 1682.780 2896.840 1683.040 2897.100 ;
        RECT 690.560 2893.100 690.820 2893.360 ;
        RECT 697.920 2893.100 698.180 2893.360 ;
        RECT 1472.560 2892.760 1472.820 2893.020 ;
        RECT 596.720 2892.420 596.980 2892.680 ;
        RECT 628.460 2892.420 628.720 2892.680 ;
        RECT 689.640 2892.420 689.900 2892.680 ;
        RECT 690.100 2892.420 690.360 2892.680 ;
        RECT 786.240 2892.420 786.500 2892.680 ;
        RECT 786.700 2892.420 786.960 2892.680 ;
        RECT 882.840 2892.420 883.100 2892.680 ;
        RECT 883.300 2892.420 883.560 2892.680 ;
        RECT 979.440 2892.420 979.700 2892.680 ;
        RECT 979.900 2892.420 980.160 2892.680 ;
        RECT 1076.040 2892.420 1076.300 2892.680 ;
        RECT 1076.500 2892.420 1076.760 2892.680 ;
        RECT 1172.640 2892.420 1172.900 2892.680 ;
        RECT 1173.100 2892.420 1173.360 2892.680 ;
        RECT 1269.240 2892.420 1269.500 2892.680 ;
        RECT 1269.700 2892.420 1269.960 2892.680 ;
        RECT 1365.840 2892.420 1366.100 2892.680 ;
        RECT 697.920 2892.080 698.180 2892.340 ;
        RECT 761.860 2892.080 762.120 2892.340 ;
        RECT 812.000 2892.080 812.260 2892.340 ;
        RECT 858.460 2892.080 858.720 2892.340 ;
        RECT 908.600 2892.080 908.860 2892.340 ;
        RECT 955.060 2892.080 955.320 2892.340 ;
        RECT 1005.200 2892.080 1005.460 2892.340 ;
        RECT 1051.660 2892.080 1051.920 2892.340 ;
        RECT 1101.800 2892.080 1102.060 2892.340 ;
        RECT 1148.260 2892.080 1148.520 2892.340 ;
        RECT 1198.400 2892.080 1198.660 2892.340 ;
        RECT 1244.860 2892.080 1245.120 2892.340 ;
        RECT 1295.000 2892.080 1295.260 2892.340 ;
        RECT 1341.460 2892.080 1341.720 2892.340 ;
        RECT 1472.560 2892.080 1472.820 2892.340 ;
        RECT 589.820 2649.320 590.080 2649.580 ;
        RECT 596.720 2649.320 596.980 2649.580 ;
        RECT 357.520 1983.600 357.780 1983.860 ;
        RECT 589.820 1983.600 590.080 1983.860 ;
        RECT 631.680 1983.600 631.940 1983.860 ;
        RECT 631.680 1924.780 631.940 1925.040 ;
        RECT 651.460 1924.780 651.720 1925.040 ;
        RECT 651.460 1732.340 651.720 1732.600 ;
        RECT 663.880 1732.340 664.140 1732.600 ;
        RECT 663.880 1702.760 664.140 1703.020 ;
        RECT 1918.300 1702.760 1918.560 1703.020 ;
        RECT 663.420 1607.560 663.680 1607.820 ;
        RECT 664.340 1607.560 664.600 1607.820 ;
        RECT 662.040 1593.620 662.300 1593.880 ;
        RECT 664.340 1593.620 664.600 1593.880 ;
        RECT 662.040 1545.680 662.300 1545.940 ;
        RECT 663.880 1545.680 664.140 1545.940 ;
        RECT 663.420 1414.440 663.680 1414.700 ;
        RECT 664.340 1414.440 664.600 1414.700 ;
        RECT 664.340 1052.000 664.600 1052.260 ;
        RECT 667.560 1052.000 667.820 1052.260 ;
        RECT 664.340 925.860 664.600 926.120 ;
        RECT 665.720 925.860 665.980 926.120 ;
        RECT 664.340 675.960 664.600 676.220 ;
        RECT 664.800 675.620 665.060 675.880 ;
        RECT 665.720 497.120 665.980 497.380 ;
        RECT 665.720 496.440 665.980 496.700 ;
        RECT 665.720 338.000 665.980 338.260 ;
        RECT 666.180 338.000 666.440 338.260 ;
        RECT 664.800 289.380 665.060 289.640 ;
        RECT 666.180 289.380 666.440 289.640 ;
        RECT 664.800 192.820 665.060 193.080 ;
        RECT 666.180 192.820 666.440 193.080 ;
        RECT 68.180 45.260 68.440 45.520 ;
        RECT 665.260 45.260 665.520 45.520 ;
      LAYER met2 ;
        RECT 1684.090 2897.210 1684.370 2900.055 ;
        RECT 1682.840 2897.130 1684.370 2897.210 ;
        RECT 1682.780 2897.070 1684.370 2897.130 ;
        RECT 1682.780 2896.810 1683.040 2897.070 ;
        RECT 1548.920 2896.700 1549.180 2896.790 ;
        RECT 1549.840 2896.700 1550.100 2896.790 ;
        RECT 1548.920 2896.560 1550.100 2896.700 ;
        RECT 1548.920 2896.470 1549.180 2896.560 ;
        RECT 1549.840 2896.470 1550.100 2896.560 ;
        RECT 1684.090 2896.055 1684.370 2897.070 ;
        RECT 786.700 2895.110 786.960 2895.430 ;
        RECT 812.000 2895.110 812.260 2895.430 ;
        RECT 883.300 2895.110 883.560 2895.430 ;
        RECT 908.600 2895.110 908.860 2895.430 ;
        RECT 979.900 2895.110 980.160 2895.430 ;
        RECT 1005.200 2895.110 1005.460 2895.430 ;
        RECT 1076.500 2895.110 1076.760 2895.430 ;
        RECT 1101.800 2895.110 1102.060 2895.430 ;
        RECT 1173.100 2895.110 1173.360 2895.430 ;
        RECT 1198.400 2895.110 1198.660 2895.430 ;
        RECT 1269.700 2895.110 1269.960 2895.430 ;
        RECT 1295.000 2895.110 1295.260 2895.430 ;
        RECT 628.460 2894.430 628.720 2894.750 ;
        RECT 689.180 2894.430 689.440 2894.750 ;
        RECT 761.860 2894.430 762.120 2894.750 ;
        RECT 786.240 2894.430 786.500 2894.750 ;
        RECT 628.520 2892.710 628.660 2894.430 ;
        RECT 596.720 2892.390 596.980 2892.710 ;
        RECT 628.460 2892.390 628.720 2892.710 ;
        RECT 689.240 2892.450 689.380 2894.430 ;
        RECT 690.560 2893.070 690.820 2893.390 ;
        RECT 697.920 2893.070 698.180 2893.390 ;
        RECT 689.640 2892.450 689.900 2892.710 ;
        RECT 689.240 2892.390 689.900 2892.450 ;
        RECT 690.100 2892.620 690.360 2892.710 ;
        RECT 690.620 2892.620 690.760 2893.070 ;
        RECT 690.100 2892.480 690.760 2892.620 ;
        RECT 690.100 2892.390 690.360 2892.480 ;
        RECT 596.780 2649.610 596.920 2892.390 ;
        RECT 689.240 2892.310 689.840 2892.390 ;
        RECT 697.980 2892.370 698.120 2893.070 ;
        RECT 761.920 2892.370 762.060 2894.430 ;
        RECT 786.300 2892.710 786.440 2894.430 ;
        RECT 786.760 2892.710 786.900 2895.110 ;
        RECT 786.240 2892.390 786.500 2892.710 ;
        RECT 786.700 2892.390 786.960 2892.710 ;
        RECT 812.060 2892.370 812.200 2895.110 ;
        RECT 858.460 2894.430 858.720 2894.750 ;
        RECT 882.840 2894.430 883.100 2894.750 ;
        RECT 858.520 2892.370 858.660 2894.430 ;
        RECT 882.900 2892.710 883.040 2894.430 ;
        RECT 883.360 2892.710 883.500 2895.110 ;
        RECT 882.840 2892.390 883.100 2892.710 ;
        RECT 883.300 2892.390 883.560 2892.710 ;
        RECT 908.660 2892.370 908.800 2895.110 ;
        RECT 955.060 2894.430 955.320 2894.750 ;
        RECT 979.440 2894.430 979.700 2894.750 ;
        RECT 955.120 2892.370 955.260 2894.430 ;
        RECT 979.500 2892.710 979.640 2894.430 ;
        RECT 979.960 2892.710 980.100 2895.110 ;
        RECT 979.440 2892.390 979.700 2892.710 ;
        RECT 979.900 2892.390 980.160 2892.710 ;
        RECT 1005.260 2892.370 1005.400 2895.110 ;
        RECT 1051.660 2894.430 1051.920 2894.750 ;
        RECT 1076.040 2894.430 1076.300 2894.750 ;
        RECT 1051.720 2892.370 1051.860 2894.430 ;
        RECT 1076.100 2892.710 1076.240 2894.430 ;
        RECT 1076.560 2892.710 1076.700 2895.110 ;
        RECT 1076.040 2892.390 1076.300 2892.710 ;
        RECT 1076.500 2892.390 1076.760 2892.710 ;
        RECT 1101.860 2892.370 1102.000 2895.110 ;
        RECT 1148.260 2894.430 1148.520 2894.750 ;
        RECT 1172.640 2894.430 1172.900 2894.750 ;
        RECT 1148.320 2892.370 1148.460 2894.430 ;
        RECT 1172.700 2892.710 1172.840 2894.430 ;
        RECT 1173.160 2892.710 1173.300 2895.110 ;
        RECT 1172.640 2892.390 1172.900 2892.710 ;
        RECT 1173.100 2892.390 1173.360 2892.710 ;
        RECT 1198.460 2892.370 1198.600 2895.110 ;
        RECT 1244.860 2894.430 1245.120 2894.750 ;
        RECT 1269.240 2894.430 1269.500 2894.750 ;
        RECT 1244.920 2892.370 1245.060 2894.430 ;
        RECT 1269.300 2892.710 1269.440 2894.430 ;
        RECT 1269.760 2892.710 1269.900 2895.110 ;
        RECT 1269.240 2892.390 1269.500 2892.710 ;
        RECT 1269.700 2892.390 1269.960 2892.710 ;
        RECT 1295.060 2892.370 1295.200 2895.110 ;
        RECT 1341.460 2894.430 1341.720 2894.750 ;
        RECT 1365.840 2894.430 1366.100 2894.750 ;
        RECT 1341.520 2892.370 1341.660 2894.430 ;
        RECT 1365.900 2892.710 1366.040 2894.430 ;
        RECT 1472.560 2892.730 1472.820 2893.050 ;
        RECT 1365.840 2892.390 1366.100 2892.710 ;
        RECT 1472.620 2892.370 1472.760 2892.730 ;
        RECT 697.920 2892.050 698.180 2892.370 ;
        RECT 761.860 2892.050 762.120 2892.370 ;
        RECT 812.000 2892.050 812.260 2892.370 ;
        RECT 858.460 2892.050 858.720 2892.370 ;
        RECT 908.600 2892.050 908.860 2892.370 ;
        RECT 955.060 2892.050 955.320 2892.370 ;
        RECT 1005.200 2892.050 1005.460 2892.370 ;
        RECT 1051.660 2892.050 1051.920 2892.370 ;
        RECT 1101.800 2892.050 1102.060 2892.370 ;
        RECT 1148.260 2892.050 1148.520 2892.370 ;
        RECT 1198.400 2892.050 1198.660 2892.370 ;
        RECT 1244.860 2892.050 1245.120 2892.370 ;
        RECT 1295.000 2892.050 1295.260 2892.370 ;
        RECT 1341.460 2892.050 1341.720 2892.370 ;
        RECT 1472.560 2892.050 1472.820 2892.370 ;
        RECT 589.820 2649.290 590.080 2649.610 ;
        RECT 596.720 2649.290 596.980 2649.610 ;
        RECT 589.880 2648.445 590.020 2649.290 ;
        RECT 589.810 2648.075 590.090 2648.445 ;
        RECT 589.880 1983.890 590.020 2648.075 ;
        RECT 357.520 1983.570 357.780 1983.890 ;
        RECT 589.820 1983.570 590.080 1983.890 ;
        RECT 631.680 1983.570 631.940 1983.890 ;
        RECT 357.580 1926.285 357.720 1983.570 ;
        RECT 357.510 1925.915 357.790 1926.285 ;
        RECT 631.740 1925.070 631.880 1983.570 ;
        RECT 631.680 1924.750 631.940 1925.070 ;
        RECT 651.460 1924.750 651.720 1925.070 ;
        RECT 651.520 1732.630 651.660 1924.750 ;
        RECT 1922.850 1750.730 1923.130 1754.000 ;
        RECT 1918.360 1750.590 1923.130 1750.730 ;
        RECT 651.460 1732.310 651.720 1732.630 ;
        RECT 663.880 1732.310 664.140 1732.630 ;
        RECT 663.940 1703.050 664.080 1732.310 ;
        RECT 1918.360 1703.050 1918.500 1750.590 ;
        RECT 1922.850 1750.000 1923.130 1750.590 ;
        RECT 663.880 1702.730 664.140 1703.050 ;
        RECT 1918.300 1702.730 1918.560 1703.050 ;
        RECT 663.940 1607.930 664.080 1702.730 ;
        RECT 663.480 1607.850 664.080 1607.930 ;
        RECT 663.420 1607.790 664.080 1607.850 ;
        RECT 663.420 1607.530 663.680 1607.790 ;
        RECT 664.340 1607.530 664.600 1607.850 ;
        RECT 663.480 1607.375 663.620 1607.530 ;
        RECT 664.400 1593.910 664.540 1607.530 ;
        RECT 662.040 1593.590 662.300 1593.910 ;
        RECT 664.340 1593.590 664.600 1593.910 ;
        RECT 662.100 1545.970 662.240 1593.590 ;
        RECT 662.040 1545.650 662.300 1545.970 ;
        RECT 663.880 1545.650 664.140 1545.970 ;
        RECT 663.940 1511.370 664.080 1545.650 ;
        RECT 663.480 1511.230 664.080 1511.370 ;
        RECT 663.480 1510.690 663.620 1511.230 ;
        RECT 663.480 1510.550 664.080 1510.690 ;
        RECT 663.940 1463.090 664.080 1510.550 ;
        RECT 663.940 1462.950 664.540 1463.090 ;
        RECT 664.400 1414.730 664.540 1462.950 ;
        RECT 663.420 1414.410 663.680 1414.730 ;
        RECT 664.340 1414.410 664.600 1414.730 ;
        RECT 663.480 1414.130 663.620 1414.410 ;
        RECT 663.480 1413.990 664.080 1414.130 ;
        RECT 663.940 1318.250 664.080 1413.990 ;
        RECT 663.480 1318.110 664.080 1318.250 ;
        RECT 663.480 1317.570 663.620 1318.110 ;
        RECT 663.480 1317.430 664.080 1317.570 ;
        RECT 663.940 1269.970 664.080 1317.430 ;
        RECT 663.940 1269.830 664.540 1269.970 ;
        RECT 664.400 1207.525 664.540 1269.830 ;
        RECT 664.330 1207.155 664.610 1207.525 ;
        RECT 667.550 1207.155 667.830 1207.525 ;
        RECT 667.620 1052.290 667.760 1207.155 ;
        RECT 664.340 1051.970 664.600 1052.290 ;
        RECT 667.560 1051.970 667.820 1052.290 ;
        RECT 664.400 980.405 664.540 1051.970 ;
        RECT 664.330 980.035 664.610 980.405 ;
        RECT 664.330 979.355 664.610 979.725 ;
        RECT 664.400 926.150 664.540 979.355 ;
        RECT 664.340 925.830 664.600 926.150 ;
        RECT 665.720 925.830 665.980 926.150 ;
        RECT 665.780 821.285 665.920 925.830 ;
        RECT 664.790 820.915 665.070 821.285 ;
        RECT 665.710 820.915 665.990 821.285 ;
        RECT 664.860 773.685 665.000 820.915 ;
        RECT 664.790 773.315 665.070 773.685 ;
        RECT 664.790 772.890 665.070 773.005 ;
        RECT 664.400 772.750 665.070 772.890 ;
        RECT 664.400 748.410 664.540 772.750 ;
        RECT 664.790 772.635 665.070 772.750 ;
        RECT 664.400 748.270 665.000 748.410 ;
        RECT 664.860 724.440 665.000 748.270 ;
        RECT 664.400 724.300 665.000 724.440 ;
        RECT 664.400 676.250 664.540 724.300 ;
        RECT 664.340 675.930 664.600 676.250 ;
        RECT 664.800 675.590 665.060 675.910 ;
        RECT 664.860 592.805 665.000 675.590 ;
        RECT 705.050 600.170 705.330 604.000 ;
        RECT 703.960 600.030 705.330 600.170 ;
        RECT 703.960 592.805 704.100 600.030 ;
        RECT 705.050 600.000 705.330 600.030 ;
        RECT 664.790 592.435 665.070 592.805 ;
        RECT 703.890 592.435 704.170 592.805 ;
        RECT 664.860 585.890 665.000 592.435 ;
        RECT 664.860 585.750 665.920 585.890 ;
        RECT 665.780 497.410 665.920 585.750 ;
        RECT 665.720 497.090 665.980 497.410 ;
        RECT 665.720 496.410 665.980 496.730 ;
        RECT 665.780 483.210 665.920 496.410 ;
        RECT 665.780 483.070 666.380 483.210 ;
        RECT 666.240 338.290 666.380 483.070 ;
        RECT 665.720 337.970 665.980 338.290 ;
        RECT 666.180 337.970 666.440 338.290 ;
        RECT 665.780 303.690 665.920 337.970 ;
        RECT 665.780 303.550 666.380 303.690 ;
        RECT 666.240 289.670 666.380 303.550 ;
        RECT 664.800 289.350 665.060 289.670 ;
        RECT 666.180 289.350 666.440 289.670 ;
        RECT 664.860 254.730 665.000 289.350 ;
        RECT 664.860 254.590 665.920 254.730 ;
        RECT 665.780 207.130 665.920 254.590 ;
        RECT 665.780 206.990 666.380 207.130 ;
        RECT 666.240 193.110 666.380 206.990 ;
        RECT 664.800 192.790 665.060 193.110 ;
        RECT 666.180 192.790 666.440 193.110 ;
        RECT 664.860 158.170 665.000 192.790 ;
        RECT 664.860 158.030 665.920 158.170 ;
        RECT 665.780 110.570 665.920 158.030 ;
        RECT 665.780 110.430 666.380 110.570 ;
        RECT 666.240 62.290 666.380 110.430 ;
        RECT 665.320 62.150 666.380 62.290 ;
        RECT 665.320 45.550 665.460 62.150 ;
        RECT 68.180 45.230 68.440 45.550 ;
        RECT 665.260 45.230 665.520 45.550 ;
        RECT 68.240 2.400 68.380 45.230 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 589.810 2648.120 590.090 2648.400 ;
        RECT 357.510 1925.960 357.790 1926.240 ;
        RECT 664.330 1207.200 664.610 1207.480 ;
        RECT 667.550 1207.200 667.830 1207.480 ;
        RECT 664.330 980.080 664.610 980.360 ;
        RECT 664.330 979.400 664.610 979.680 ;
        RECT 664.790 820.960 665.070 821.240 ;
        RECT 665.710 820.960 665.990 821.240 ;
        RECT 664.790 773.360 665.070 773.640 ;
        RECT 664.790 772.680 665.070 772.960 ;
        RECT 664.790 592.480 665.070 592.760 ;
        RECT 703.890 592.480 704.170 592.760 ;
      LAYER met3 ;
        RECT 589.785 2648.410 590.115 2648.425 ;
        RECT 578.070 2648.240 590.115 2648.410 ;
        RECT 574.800 2648.110 590.115 2648.240 ;
        RECT 574.800 2647.640 578.800 2648.110 ;
        RECT 589.785 2648.095 590.115 2648.110 ;
        RECT 357.485 1926.250 357.815 1926.265 ;
        RECT 360.000 1926.250 364.000 1926.400 ;
        RECT 357.485 1925.950 364.000 1926.250 ;
        RECT 357.485 1925.935 357.815 1925.950 ;
        RECT 360.000 1925.800 364.000 1925.950 ;
        RECT 664.305 1207.490 664.635 1207.505 ;
        RECT 667.525 1207.490 667.855 1207.505 ;
        RECT 664.305 1207.190 667.855 1207.490 ;
        RECT 664.305 1207.175 664.635 1207.190 ;
        RECT 667.525 1207.175 667.855 1207.190 ;
        RECT 664.305 980.380 664.635 980.385 ;
        RECT 664.305 980.370 664.890 980.380 ;
        RECT 664.080 980.070 664.890 980.370 ;
        RECT 664.305 980.060 664.890 980.070 ;
        RECT 664.305 980.055 664.635 980.060 ;
        RECT 664.305 979.700 664.635 979.705 ;
        RECT 664.305 979.690 664.890 979.700 ;
        RECT 664.080 979.390 664.890 979.690 ;
        RECT 664.305 979.380 664.890 979.390 ;
        RECT 664.305 979.375 664.635 979.380 ;
        RECT 664.765 821.250 665.095 821.265 ;
        RECT 665.685 821.250 666.015 821.265 ;
        RECT 664.765 820.950 666.015 821.250 ;
        RECT 664.765 820.935 665.095 820.950 ;
        RECT 665.685 820.935 666.015 820.950 ;
        RECT 664.765 773.650 665.095 773.665 ;
        RECT 664.765 773.350 665.770 773.650 ;
        RECT 664.765 773.335 665.095 773.350 ;
        RECT 664.765 772.970 665.095 772.985 ;
        RECT 665.470 772.970 665.770 773.350 ;
        RECT 664.765 772.670 665.770 772.970 ;
        RECT 664.765 772.655 665.095 772.670 ;
        RECT 664.765 592.770 665.095 592.785 ;
        RECT 703.865 592.770 704.195 592.785 ;
        RECT 664.765 592.470 704.195 592.770 ;
        RECT 664.765 592.455 665.095 592.470 ;
        RECT 703.865 592.455 704.195 592.470 ;
      LAYER via3 ;
        RECT 664.540 980.060 664.860 980.380 ;
        RECT 664.540 979.380 664.860 979.700 ;
      LAYER met4 ;
        RECT 664.535 980.055 664.865 980.385 ;
        RECT 664.550 979.705 664.850 980.055 ;
        RECT 664.535 979.375 664.865 979.705 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1525.890 2896.500 1526.210 2896.760 ;
        RECT 1579.250 2896.500 1579.570 2896.760 ;
        RECT 1650.090 2896.500 1650.410 2896.760 ;
        RECT 1525.980 2896.360 1526.120 2896.500 ;
        RECT 1525.520 2896.220 1526.120 2896.360 ;
        RECT 1579.340 2896.360 1579.480 2896.500 ;
        RECT 1650.180 2896.360 1650.320 2896.500 ;
        RECT 1579.340 2896.220 1650.320 2896.360 ;
        RECT 1501.050 2894.660 1501.370 2894.720 ;
        RECT 1525.520 2894.660 1525.660 2896.220 ;
        RECT 1501.050 2894.520 1525.660 2894.660 ;
        RECT 1501.050 2894.460 1501.370 2894.520 ;
        RECT 1438.490 2894.320 1438.810 2894.380 ;
        RECT 1449.070 2894.320 1449.390 2894.380 ;
        RECT 1438.490 2894.180 1449.390 2894.320 ;
        RECT 1438.490 2894.120 1438.810 2894.180 ;
        RECT 1449.070 2894.120 1449.390 2894.180 ;
        RECT 1496.910 2893.980 1497.230 2894.040 ;
        RECT 1501.050 2893.980 1501.370 2894.040 ;
        RECT 1496.910 2893.840 1501.370 2893.980 ;
        RECT 1496.910 2893.780 1497.230 2893.840 ;
        RECT 1501.050 2893.780 1501.370 2893.840 ;
        RECT 645.450 2892.960 645.770 2893.020 ;
        RECT 1438.490 2892.960 1438.810 2893.020 ;
        RECT 645.450 2892.820 1438.810 2892.960 ;
        RECT 645.450 2892.760 645.770 2892.820 ;
        RECT 1438.490 2892.760 1438.810 2892.820 ;
        RECT 642.230 2608.040 642.550 2608.100 ;
        RECT 645.450 2608.040 645.770 2608.100 ;
        RECT 642.230 2607.900 645.770 2608.040 ;
        RECT 642.230 2607.840 642.550 2607.900 ;
        RECT 645.450 2607.840 645.770 2607.900 ;
        RECT 586.570 2604.640 586.890 2604.700 ;
        RECT 642.230 2604.640 642.550 2604.700 ;
        RECT 586.570 2604.500 642.550 2604.640 ;
        RECT 586.570 2604.440 586.890 2604.500 ;
        RECT 642.230 2604.440 642.550 2604.500 ;
        RECT 646.370 590.820 646.690 590.880 ;
        RECT 886.950 590.820 887.270 590.880 ;
        RECT 646.370 590.680 887.270 590.820 ;
        RECT 646.370 590.620 646.690 590.680 ;
        RECT 886.950 590.620 887.270 590.680 ;
        RECT 424.650 43.760 424.970 43.820 ;
        RECT 424.650 43.620 629.580 43.760 ;
        RECT 424.650 43.560 424.970 43.620 ;
        RECT 629.440 43.420 629.580 43.620 ;
        RECT 646.370 43.420 646.690 43.480 ;
        RECT 629.440 43.280 646.690 43.420 ;
        RECT 646.370 43.220 646.690 43.280 ;
      LAYER via ;
        RECT 1525.920 2896.500 1526.180 2896.760 ;
        RECT 1579.280 2896.500 1579.540 2896.760 ;
        RECT 1650.120 2896.500 1650.380 2896.760 ;
        RECT 1501.080 2894.460 1501.340 2894.720 ;
        RECT 1438.520 2894.120 1438.780 2894.380 ;
        RECT 1449.100 2894.120 1449.360 2894.380 ;
        RECT 1496.940 2893.780 1497.200 2894.040 ;
        RECT 1501.080 2893.780 1501.340 2894.040 ;
        RECT 645.480 2892.760 645.740 2893.020 ;
        RECT 1438.520 2892.760 1438.780 2893.020 ;
        RECT 642.260 2607.840 642.520 2608.100 ;
        RECT 645.480 2607.840 645.740 2608.100 ;
        RECT 586.600 2604.440 586.860 2604.700 ;
        RECT 642.260 2604.440 642.520 2604.700 ;
        RECT 646.400 590.620 646.660 590.880 ;
        RECT 886.980 590.620 887.240 590.880 ;
        RECT 424.680 43.560 424.940 43.820 ;
        RECT 646.400 43.220 646.660 43.480 ;
      LAYER met2 ;
        RECT 1525.920 2896.645 1526.180 2896.790 ;
        RECT 1579.280 2896.645 1579.540 2896.790 ;
        RECT 1525.910 2896.275 1526.190 2896.645 ;
        RECT 1579.270 2896.275 1579.550 2896.645 ;
        RECT 1650.120 2896.530 1650.380 2896.790 ;
        RECT 1651.890 2896.530 1652.170 2900.055 ;
        RECT 1650.120 2896.470 1652.170 2896.530 ;
        RECT 1650.180 2896.390 1652.170 2896.470 ;
        RECT 1651.890 2896.055 1652.170 2896.390 ;
        RECT 1438.520 2894.090 1438.780 2894.410 ;
        RECT 1449.090 2894.235 1449.370 2894.605 ;
        RECT 1496.930 2894.235 1497.210 2894.605 ;
        RECT 1501.080 2894.430 1501.340 2894.750 ;
        RECT 1449.100 2894.090 1449.360 2894.235 ;
        RECT 1438.580 2893.050 1438.720 2894.090 ;
        RECT 1497.000 2894.070 1497.140 2894.235 ;
        RECT 1501.140 2894.070 1501.280 2894.430 ;
        RECT 1496.940 2893.750 1497.200 2894.070 ;
        RECT 1501.080 2893.750 1501.340 2894.070 ;
        RECT 645.480 2892.730 645.740 2893.050 ;
        RECT 1438.520 2892.730 1438.780 2893.050 ;
        RECT 645.540 2608.130 645.680 2892.730 ;
        RECT 642.260 2607.810 642.520 2608.130 ;
        RECT 645.480 2607.810 645.740 2608.130 ;
        RECT 586.590 2605.235 586.870 2605.605 ;
        RECT 586.660 2604.730 586.800 2605.235 ;
        RECT 642.320 2604.730 642.460 2607.810 ;
        RECT 586.600 2604.410 586.860 2604.730 ;
        RECT 642.260 2604.410 642.520 2604.730 ;
        RECT 642.320 1866.445 642.460 2604.410 ;
        RECT 642.250 1866.075 642.530 1866.445 ;
        RECT 642.320 1863.725 642.460 1866.075 ;
        RECT 642.250 1863.355 642.530 1863.725 ;
        RECT 646.390 1863.355 646.670 1863.725 ;
        RECT 646.460 590.910 646.600 1863.355 ;
        RECT 888.590 600.170 888.870 604.000 ;
        RECT 887.040 600.030 888.870 600.170 ;
        RECT 887.040 590.910 887.180 600.030 ;
        RECT 888.590 600.000 888.870 600.030 ;
        RECT 646.400 590.590 646.660 590.910 ;
        RECT 886.980 590.590 887.240 590.910 ;
        RECT 424.680 43.530 424.940 43.850 ;
        RECT 424.740 2.400 424.880 43.530 ;
        RECT 646.460 43.510 646.600 590.590 ;
        RECT 646.400 43.190 646.660 43.510 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 1525.910 2896.320 1526.190 2896.600 ;
        RECT 1579.270 2896.320 1579.550 2896.600 ;
        RECT 1449.090 2894.280 1449.370 2894.560 ;
        RECT 1496.930 2894.280 1497.210 2894.560 ;
        RECT 586.590 2605.280 586.870 2605.560 ;
        RECT 642.250 1866.120 642.530 1866.400 ;
        RECT 642.250 1863.400 642.530 1863.680 ;
        RECT 646.390 1863.400 646.670 1863.680 ;
      LAYER met3 ;
        RECT 1525.885 2896.610 1526.215 2896.625 ;
        RECT 1579.245 2896.610 1579.575 2896.625 ;
        RECT 1525.885 2896.310 1579.575 2896.610 ;
        RECT 1525.885 2896.295 1526.215 2896.310 ;
        RECT 1579.245 2896.295 1579.575 2896.310 ;
        RECT 1449.065 2894.570 1449.395 2894.585 ;
        RECT 1496.905 2894.570 1497.235 2894.585 ;
        RECT 1449.065 2894.270 1497.235 2894.570 ;
        RECT 1449.065 2894.255 1449.395 2894.270 ;
        RECT 1496.905 2894.255 1497.235 2894.270 ;
        RECT 574.800 2605.570 578.800 2606.080 ;
        RECT 586.565 2605.570 586.895 2605.585 ;
        RECT 574.800 2605.480 586.895 2605.570 ;
        RECT 578.070 2605.270 586.895 2605.480 ;
        RECT 586.565 2605.255 586.895 2605.270 ;
        RECT 627.030 1866.410 631.030 1866.560 ;
        RECT 642.225 1866.410 642.555 1866.425 ;
        RECT 627.030 1866.110 642.555 1866.410 ;
        RECT 627.030 1865.960 631.030 1866.110 ;
        RECT 642.225 1866.095 642.555 1866.110 ;
        RECT 642.225 1863.690 642.555 1863.705 ;
        RECT 646.365 1863.690 646.695 1863.705 ;
        RECT 642.225 1863.390 646.695 1863.690 ;
        RECT 642.225 1863.375 642.555 1863.390 ;
        RECT 646.365 1863.375 646.695 1863.390 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1672.170 2896.500 1672.490 2896.760 ;
        RECT 1672.260 2891.940 1672.400 2896.500 ;
        RECT 1627.640 2891.800 1672.400 2891.940 ;
        RECT 426.950 2891.600 427.270 2891.660 ;
        RECT 627.970 2891.600 628.290 2891.660 ;
        RECT 426.950 2891.460 628.290 2891.600 ;
        RECT 426.950 2891.400 427.270 2891.460 ;
        RECT 627.970 2891.400 628.290 2891.460 ;
        RECT 628.890 2891.600 629.210 2891.660 ;
        RECT 628.890 2891.460 1568.440 2891.600 ;
        RECT 628.890 2891.400 629.210 2891.460 ;
        RECT 1568.300 2890.920 1568.440 2891.460 ;
        RECT 1627.640 2890.920 1627.780 2891.800 ;
        RECT 1568.300 2890.780 1627.780 2890.920 ;
        RECT 351.050 2622.320 351.370 2622.380 ;
        RECT 414.070 2622.320 414.390 2622.380 ;
        RECT 351.050 2622.180 414.390 2622.320 ;
        RECT 351.050 2622.120 351.370 2622.180 ;
        RECT 414.070 2622.120 414.390 2622.180 ;
        RECT 357.950 591.840 358.270 591.900 ;
        RECT 441.670 591.840 441.990 591.900 ;
        RECT 357.950 591.700 441.990 591.840 ;
        RECT 357.950 591.640 358.270 591.700 ;
        RECT 441.670 591.640 441.990 591.700 ;
        RECT 441.670 590.140 441.990 590.200 ;
        RECT 897.070 590.140 897.390 590.200 ;
        RECT 441.670 590.000 897.390 590.140 ;
        RECT 441.670 589.940 441.990 590.000 ;
        RECT 897.070 589.940 897.390 590.000 ;
      LAYER via ;
        RECT 1672.200 2896.500 1672.460 2896.760 ;
        RECT 426.980 2891.400 427.240 2891.660 ;
        RECT 628.000 2891.400 628.260 2891.660 ;
        RECT 628.920 2891.400 629.180 2891.660 ;
        RECT 351.080 2622.120 351.340 2622.380 ;
        RECT 414.100 2622.120 414.360 2622.380 ;
        RECT 357.980 591.640 358.240 591.900 ;
        RECT 441.700 591.640 441.960 591.900 ;
        RECT 441.700 589.940 441.960 590.200 ;
        RECT 897.100 589.940 897.360 590.200 ;
      LAYER met2 ;
        RECT 1672.200 2896.530 1672.460 2896.790 ;
        RECT 1673.050 2896.530 1673.330 2900.055 ;
        RECT 1672.200 2896.470 1673.330 2896.530 ;
        RECT 1672.260 2896.390 1673.330 2896.470 ;
        RECT 1673.050 2896.055 1673.330 2896.390 ;
        RECT 426.980 2891.370 427.240 2891.690 ;
        RECT 628.000 2891.370 628.260 2891.690 ;
        RECT 628.920 2891.370 629.180 2891.690 ;
        RECT 427.040 2628.045 427.180 2891.370 ;
        RECT 628.060 2891.090 628.200 2891.370 ;
        RECT 628.980 2891.090 629.120 2891.370 ;
        RECT 628.060 2890.950 629.120 2891.090 ;
        RECT 426.970 2627.675 427.250 2628.045 ;
        RECT 414.090 2624.275 414.370 2624.645 ;
        RECT 414.160 2622.410 414.300 2624.275 ;
        RECT 351.080 2622.090 351.340 2622.410 ;
        RECT 414.100 2622.090 414.360 2622.410 ;
        RECT 351.140 1741.325 351.280 2622.090 ;
        RECT 351.070 1740.955 351.350 1741.325 ;
        RECT 357.970 1740.955 358.250 1741.325 ;
        RECT 358.040 591.930 358.180 1740.955 ;
        RECT 897.790 600.170 898.070 604.000 ;
        RECT 897.160 600.030 898.070 600.170 ;
        RECT 357.980 591.610 358.240 591.930 ;
        RECT 441.700 591.610 441.960 591.930 ;
        RECT 441.760 590.230 441.900 591.610 ;
        RECT 897.160 590.230 897.300 600.030 ;
        RECT 897.790 600.000 898.070 600.030 ;
        RECT 441.700 589.910 441.960 590.230 ;
        RECT 897.100 589.910 897.360 590.230 ;
        RECT 441.760 17.410 441.900 589.910 ;
        RECT 441.760 17.270 442.820 17.410 ;
        RECT 442.680 2.400 442.820 17.270 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 426.970 2627.720 427.250 2628.000 ;
        RECT 414.090 2624.320 414.370 2624.600 ;
        RECT 351.070 1741.000 351.350 1741.280 ;
        RECT 357.970 1741.000 358.250 1741.280 ;
      LAYER met3 ;
        RECT 426.945 2628.010 427.275 2628.025 ;
        RECT 426.945 2627.710 430.250 2628.010 ;
        RECT 426.945 2627.695 427.275 2627.710 ;
        RECT 429.950 2625.120 430.250 2627.710 ;
        RECT 414.065 2624.610 414.395 2624.625 ;
        RECT 429.950 2624.610 434.000 2625.120 ;
        RECT 414.065 2624.520 434.000 2624.610 ;
        RECT 414.065 2624.310 430.250 2624.520 ;
        RECT 414.065 2624.295 414.395 2624.310 ;
        RECT 351.045 1741.290 351.375 1741.305 ;
        RECT 357.945 1741.290 358.275 1741.305 ;
        RECT 360.000 1741.290 364.000 1741.440 ;
        RECT 351.045 1740.990 364.000 1741.290 ;
        RECT 351.045 1740.975 351.375 1740.990 ;
        RECT 357.945 1740.975 358.275 1740.990 ;
        RECT 360.000 1740.840 364.000 1740.990 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.450 2591.040 461.770 2591.100 ;
        RECT 635.330 2591.040 635.650 2591.100 ;
        RECT 1486.790 2591.040 1487.110 2591.100 ;
        RECT 461.450 2590.900 1487.110 2591.040 ;
        RECT 461.450 2590.840 461.770 2590.900 ;
        RECT 635.330 2590.840 635.650 2590.900 ;
        RECT 1486.790 2590.840 1487.110 2590.900 ;
        RECT 489.510 1690.040 489.830 1690.100 ;
        RECT 635.330 1690.040 635.650 1690.100 ;
        RECT 489.510 1689.900 635.650 1690.040 ;
        RECT 489.510 1689.840 489.830 1689.900 ;
        RECT 635.330 1689.840 635.650 1689.900 ;
        RECT 489.510 592.860 489.830 592.920 ;
        RECT 905.350 592.860 905.670 592.920 ;
        RECT 489.510 592.720 905.670 592.860 ;
        RECT 489.510 592.660 489.830 592.720 ;
        RECT 905.350 592.660 905.670 592.720 ;
        RECT 461.910 586.740 462.230 586.800 ;
        RECT 489.510 586.740 489.830 586.800 ;
        RECT 461.910 586.600 489.830 586.740 ;
        RECT 461.910 586.540 462.230 586.600 ;
        RECT 489.510 586.540 489.830 586.600 ;
        RECT 460.530 2.960 460.850 3.020 ;
        RECT 461.910 2.960 462.230 3.020 ;
        RECT 460.530 2.820 462.230 2.960 ;
        RECT 460.530 2.760 460.850 2.820 ;
        RECT 461.910 2.760 462.230 2.820 ;
      LAYER via ;
        RECT 461.480 2590.840 461.740 2591.100 ;
        RECT 635.360 2590.840 635.620 2591.100 ;
        RECT 1486.820 2590.840 1487.080 2591.100 ;
        RECT 489.540 1689.840 489.800 1690.100 ;
        RECT 635.360 1689.840 635.620 1690.100 ;
        RECT 489.540 592.660 489.800 592.920 ;
        RECT 905.380 592.660 905.640 592.920 ;
        RECT 461.940 586.540 462.200 586.800 ;
        RECT 489.540 586.540 489.800 586.800 ;
        RECT 460.560 2.760 460.820 3.020 ;
        RECT 461.940 2.760 462.200 3.020 ;
      LAYER met2 ;
        RECT 1486.810 2642.635 1487.090 2643.005 ;
        RECT 461.370 2600.660 461.650 2604.000 ;
        RECT 461.370 2600.000 461.680 2600.660 ;
        RECT 461.540 2591.130 461.680 2600.000 ;
        RECT 1486.880 2591.130 1487.020 2642.635 ;
        RECT 461.480 2590.810 461.740 2591.130 ;
        RECT 635.360 2590.810 635.620 2591.130 ;
        RECT 1486.820 2590.810 1487.080 2591.130 ;
        RECT 487.970 1700.410 488.250 1704.000 ;
        RECT 487.970 1700.270 489.740 1700.410 ;
        RECT 487.970 1700.000 488.250 1700.270 ;
        RECT 489.600 1690.130 489.740 1700.270 ;
        RECT 635.420 1690.130 635.560 2590.810 ;
        RECT 489.540 1689.810 489.800 1690.130 ;
        RECT 635.360 1689.810 635.620 1690.130 ;
        RECT 489.600 592.950 489.740 1689.810 ;
        RECT 906.990 600.170 907.270 604.000 ;
        RECT 905.440 600.030 907.270 600.170 ;
        RECT 905.440 592.950 905.580 600.030 ;
        RECT 906.990 600.000 907.270 600.030 ;
        RECT 489.540 592.630 489.800 592.950 ;
        RECT 905.380 592.630 905.640 592.950 ;
        RECT 489.600 586.830 489.740 592.630 ;
        RECT 461.940 586.510 462.200 586.830 ;
        RECT 489.540 586.510 489.800 586.830 ;
        RECT 462.000 3.050 462.140 586.510 ;
        RECT 460.560 2.730 460.820 3.050 ;
        RECT 461.940 2.730 462.200 3.050 ;
        RECT 460.620 2.400 460.760 2.730 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 1486.810 2642.680 1487.090 2642.960 ;
      LAYER met3 ;
        RECT 1500.000 2645.880 1504.000 2646.160 ;
        RECT 1499.910 2645.560 1504.000 2645.880 ;
        RECT 1486.785 2642.970 1487.115 2642.985 ;
        RECT 1499.910 2642.970 1500.210 2645.560 ;
        RECT 1486.785 2642.670 1500.210 2642.970 ;
        RECT 1486.785 2642.655 1487.115 2642.670 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 2917.100 645.310 2917.160 ;
        RECT 1737.490 2917.100 1737.810 2917.160 ;
        RECT 644.990 2916.960 1737.810 2917.100 ;
        RECT 644.990 2916.900 645.310 2916.960 ;
        RECT 1737.490 2916.900 1737.810 2916.960 ;
        RECT 575.530 2769.200 575.850 2769.260 ;
        RECT 642.230 2769.200 642.550 2769.260 ;
        RECT 644.990 2769.200 645.310 2769.260 ;
        RECT 575.530 2769.060 645.310 2769.200 ;
        RECT 575.530 2769.000 575.850 2769.060 ;
        RECT 642.230 2769.000 642.550 2769.060 ;
        RECT 644.990 2769.000 645.310 2769.060 ;
        RECT 642.230 2766.820 642.550 2766.880 ;
        RECT 643.150 2766.820 643.470 2766.880 ;
        RECT 642.230 2766.680 643.470 2766.820 ;
        RECT 642.230 2766.620 642.550 2766.680 ;
        RECT 643.150 2766.620 643.470 2766.680 ;
        RECT 643.150 2719.220 643.470 2719.280 ;
        RECT 642.780 2719.080 643.470 2719.220 ;
        RECT 642.780 2718.600 642.920 2719.080 ;
        RECT 643.150 2719.020 643.470 2719.080 ;
        RECT 642.690 2718.340 643.010 2718.600 ;
        RECT 642.230 2670.600 642.550 2670.660 ;
        RECT 642.230 2670.460 642.920 2670.600 ;
        RECT 642.230 2670.400 642.550 2670.460 ;
        RECT 642.780 2670.320 642.920 2670.460 ;
        RECT 642.690 2670.060 643.010 2670.320 ;
        RECT 642.230 2656.660 642.550 2656.720 ;
        RECT 642.690 2656.660 643.010 2656.720 ;
        RECT 642.230 2656.520 643.010 2656.660 ;
        RECT 642.230 2656.460 642.550 2656.520 ;
        RECT 642.690 2656.460 643.010 2656.520 ;
        RECT 642.230 2622.120 642.550 2622.380 ;
        RECT 642.320 2621.640 642.460 2622.120 ;
        RECT 643.150 2621.640 643.470 2621.700 ;
        RECT 642.320 2621.500 643.470 2621.640 ;
        RECT 643.150 2621.440 643.470 2621.500 ;
        RECT 641.770 2594.780 642.090 2594.840 ;
        RECT 643.150 2594.780 643.470 2594.840 ;
        RECT 641.770 2594.640 643.470 2594.780 ;
        RECT 641.770 2594.580 642.090 2594.640 ;
        RECT 643.150 2594.580 643.470 2594.640 ;
        RECT 641.770 2546.160 642.090 2546.220 ;
        RECT 643.150 2546.160 643.470 2546.220 ;
        RECT 641.770 2546.020 643.470 2546.160 ;
        RECT 641.770 2545.960 642.090 2546.020 ;
        RECT 643.150 2545.960 643.470 2546.020 ;
        RECT 641.770 2497.880 642.090 2497.940 ;
        RECT 643.150 2497.880 643.470 2497.940 ;
        RECT 641.770 2497.740 643.470 2497.880 ;
        RECT 641.770 2497.680 642.090 2497.740 ;
        RECT 643.150 2497.680 643.470 2497.740 ;
        RECT 641.770 2449.260 642.090 2449.320 ;
        RECT 643.150 2449.260 643.470 2449.320 ;
        RECT 641.770 2449.120 643.470 2449.260 ;
        RECT 641.770 2449.060 642.090 2449.120 ;
        RECT 643.150 2449.060 643.470 2449.120 ;
        RECT 641.770 2401.660 642.090 2401.720 ;
        RECT 643.150 2401.660 643.470 2401.720 ;
        RECT 641.770 2401.520 643.470 2401.660 ;
        RECT 641.770 2401.460 642.090 2401.520 ;
        RECT 643.150 2401.460 643.470 2401.520 ;
        RECT 641.770 2159.580 642.090 2159.640 ;
        RECT 643.150 2159.580 643.470 2159.640 ;
        RECT 641.770 2159.440 643.470 2159.580 ;
        RECT 641.770 2159.380 642.090 2159.440 ;
        RECT 643.150 2159.380 643.470 2159.440 ;
        RECT 641.770 2111.980 642.090 2112.040 ;
        RECT 643.150 2111.980 643.470 2112.040 ;
        RECT 641.770 2111.840 643.470 2111.980 ;
        RECT 641.770 2111.780 642.090 2111.840 ;
        RECT 643.150 2111.780 643.470 2111.840 ;
        RECT 641.770 1966.460 642.090 1966.520 ;
        RECT 643.150 1966.460 643.470 1966.520 ;
        RECT 641.770 1966.320 643.470 1966.460 ;
        RECT 641.770 1966.260 642.090 1966.320 ;
        RECT 643.150 1966.260 643.470 1966.320 ;
        RECT 641.770 1918.520 642.090 1918.580 ;
        RECT 643.150 1918.520 643.470 1918.580 ;
        RECT 641.770 1918.380 643.470 1918.520 ;
        RECT 641.770 1918.320 642.090 1918.380 ;
        RECT 643.150 1918.320 643.470 1918.380 ;
        RECT 641.770 1869.900 642.090 1869.960 ;
        RECT 642.690 1869.900 643.010 1869.960 ;
        RECT 641.770 1869.760 643.010 1869.900 ;
        RECT 641.770 1869.700 642.090 1869.760 ;
        RECT 642.690 1869.700 643.010 1869.760 ;
        RECT 642.690 1848.960 643.010 1849.220 ;
        RECT 642.780 1848.820 642.920 1848.960 ;
        RECT 643.150 1848.820 643.470 1848.880 ;
        RECT 642.780 1848.680 643.470 1848.820 ;
        RECT 643.150 1848.620 643.470 1848.680 ;
        RECT 643.610 1739.680 643.930 1739.740 ;
        RECT 643.240 1739.540 643.930 1739.680 ;
        RECT 643.240 1739.060 643.380 1739.540 ;
        RECT 643.610 1739.480 643.930 1739.540 ;
        RECT 643.150 1738.800 643.470 1739.060 ;
        RECT 641.770 1628.500 642.090 1628.560 ;
        RECT 642.230 1628.500 642.550 1628.560 ;
        RECT 641.770 1628.360 642.550 1628.500 ;
        RECT 641.770 1628.300 642.090 1628.360 ;
        RECT 642.230 1628.300 642.550 1628.360 ;
        RECT 643.150 1497.600 643.470 1497.660 ;
        RECT 644.070 1497.600 644.390 1497.660 ;
        RECT 643.150 1497.460 644.390 1497.600 ;
        RECT 643.150 1497.400 643.470 1497.460 ;
        RECT 644.070 1497.400 644.390 1497.460 ;
        RECT 642.230 1452.380 642.550 1452.440 ;
        RECT 643.150 1452.380 643.470 1452.440 ;
        RECT 642.230 1452.240 643.470 1452.380 ;
        RECT 642.230 1452.180 642.550 1452.240 ;
        RECT 643.150 1452.180 643.470 1452.240 ;
        RECT 642.230 1400.700 642.550 1400.760 ;
        RECT 643.150 1400.700 643.470 1400.760 ;
        RECT 642.230 1400.560 643.470 1400.700 ;
        RECT 642.230 1400.500 642.550 1400.560 ;
        RECT 643.150 1400.500 643.470 1400.560 ;
        RECT 642.230 1352.760 642.550 1352.820 ;
        RECT 643.150 1352.760 643.470 1352.820 ;
        RECT 642.230 1352.620 643.470 1352.760 ;
        RECT 642.230 1352.560 642.550 1352.620 ;
        RECT 643.150 1352.560 643.470 1352.620 ;
        RECT 640.390 1304.140 640.710 1304.200 ;
        RECT 642.690 1304.140 643.010 1304.200 ;
        RECT 640.390 1304.000 643.010 1304.140 ;
        RECT 640.390 1303.940 640.710 1304.000 ;
        RECT 642.690 1303.940 643.010 1304.000 ;
        RECT 643.150 1159.300 643.470 1159.360 ;
        RECT 644.070 1159.300 644.390 1159.360 ;
        RECT 643.150 1159.160 644.390 1159.300 ;
        RECT 643.150 1159.100 643.470 1159.160 ;
        RECT 644.070 1159.100 644.390 1159.160 ;
        RECT 642.230 1076.820 642.550 1077.080 ;
        RECT 642.320 1076.400 642.460 1076.820 ;
        RECT 642.230 1076.140 642.550 1076.400 ;
        RECT 642.230 1014.460 642.550 1014.520 ;
        RECT 643.150 1014.460 643.470 1014.520 ;
        RECT 642.230 1014.320 643.470 1014.460 ;
        RECT 642.230 1014.260 642.550 1014.320 ;
        RECT 643.150 1014.260 643.470 1014.320 ;
        RECT 641.770 979.440 642.090 979.500 ;
        RECT 642.690 979.440 643.010 979.500 ;
        RECT 641.770 979.300 643.010 979.440 ;
        RECT 641.770 979.240 642.090 979.300 ;
        RECT 642.690 979.240 643.010 979.300 ;
        RECT 641.770 917.900 642.090 917.960 ;
        RECT 642.690 917.900 643.010 917.960 ;
        RECT 641.770 917.760 643.010 917.900 ;
        RECT 641.770 917.700 642.090 917.760 ;
        RECT 642.690 917.700 643.010 917.760 ;
        RECT 642.690 883.360 643.010 883.620 ;
        RECT 642.780 882.880 642.920 883.360 ;
        RECT 643.150 882.880 643.470 882.940 ;
        RECT 642.780 882.740 643.470 882.880 ;
        RECT 643.150 882.680 643.470 882.740 ;
        RECT 641.770 845.480 642.090 845.540 ;
        RECT 642.690 845.480 643.010 845.540 ;
        RECT 641.770 845.340 643.010 845.480 ;
        RECT 641.770 845.280 642.090 845.340 ;
        RECT 642.690 845.280 643.010 845.340 ;
        RECT 643.150 676.160 643.470 676.220 ;
        RECT 643.610 676.160 643.930 676.220 ;
        RECT 643.150 676.020 643.930 676.160 ;
        RECT 643.150 675.960 643.470 676.020 ;
        RECT 643.610 675.960 643.930 676.020 ;
        RECT 643.610 641.620 643.930 641.880 ;
        RECT 643.150 641.480 643.470 641.540 ;
        RECT 643.700 641.480 643.840 641.620 ;
        RECT 643.150 641.340 643.840 641.480 ;
        RECT 643.150 641.280 643.470 641.340 ;
        RECT 643.610 627.680 643.930 627.940 ;
        RECT 643.700 627.200 643.840 627.680 ;
        RECT 645.450 627.200 645.770 627.260 ;
        RECT 643.700 627.060 645.770 627.200 ;
        RECT 645.450 627.000 645.770 627.060 ;
        RECT 686.390 591.500 686.710 591.560 ;
        RECT 914.550 591.500 914.870 591.560 ;
        RECT 686.390 591.360 914.870 591.500 ;
        RECT 686.390 591.300 686.710 591.360 ;
        RECT 914.550 591.300 914.870 591.360 ;
        RECT 645.450 588.440 645.770 588.500 ;
        RECT 646.830 588.440 647.150 588.500 ;
        RECT 686.390 588.440 686.710 588.500 ;
        RECT 645.450 588.300 686.710 588.440 ;
        RECT 645.450 588.240 645.770 588.300 ;
        RECT 646.830 588.240 647.150 588.300 ;
        RECT 686.390 588.240 686.710 588.300 ;
        RECT 478.470 43.420 478.790 43.480 ;
        RECT 478.470 43.280 628.660 43.420 ;
        RECT 478.470 43.220 478.790 43.280 ;
        RECT 628.520 42.740 628.660 43.280 ;
        RECT 646.830 42.740 647.150 42.800 ;
        RECT 628.520 42.600 647.150 42.740 ;
        RECT 646.830 42.540 647.150 42.600 ;
      LAYER via ;
        RECT 645.020 2916.900 645.280 2917.160 ;
        RECT 1737.520 2916.900 1737.780 2917.160 ;
        RECT 575.560 2769.000 575.820 2769.260 ;
        RECT 642.260 2769.000 642.520 2769.260 ;
        RECT 645.020 2769.000 645.280 2769.260 ;
        RECT 642.260 2766.620 642.520 2766.880 ;
        RECT 643.180 2766.620 643.440 2766.880 ;
        RECT 643.180 2719.020 643.440 2719.280 ;
        RECT 642.720 2718.340 642.980 2718.600 ;
        RECT 642.260 2670.400 642.520 2670.660 ;
        RECT 642.720 2670.060 642.980 2670.320 ;
        RECT 642.260 2656.460 642.520 2656.720 ;
        RECT 642.720 2656.460 642.980 2656.720 ;
        RECT 642.260 2622.120 642.520 2622.380 ;
        RECT 643.180 2621.440 643.440 2621.700 ;
        RECT 641.800 2594.580 642.060 2594.840 ;
        RECT 643.180 2594.580 643.440 2594.840 ;
        RECT 641.800 2545.960 642.060 2546.220 ;
        RECT 643.180 2545.960 643.440 2546.220 ;
        RECT 641.800 2497.680 642.060 2497.940 ;
        RECT 643.180 2497.680 643.440 2497.940 ;
        RECT 641.800 2449.060 642.060 2449.320 ;
        RECT 643.180 2449.060 643.440 2449.320 ;
        RECT 641.800 2401.460 642.060 2401.720 ;
        RECT 643.180 2401.460 643.440 2401.720 ;
        RECT 641.800 2159.380 642.060 2159.640 ;
        RECT 643.180 2159.380 643.440 2159.640 ;
        RECT 641.800 2111.780 642.060 2112.040 ;
        RECT 643.180 2111.780 643.440 2112.040 ;
        RECT 641.800 1966.260 642.060 1966.520 ;
        RECT 643.180 1966.260 643.440 1966.520 ;
        RECT 641.800 1918.320 642.060 1918.580 ;
        RECT 643.180 1918.320 643.440 1918.580 ;
        RECT 641.800 1869.700 642.060 1869.960 ;
        RECT 642.720 1869.700 642.980 1869.960 ;
        RECT 642.720 1848.960 642.980 1849.220 ;
        RECT 643.180 1848.620 643.440 1848.880 ;
        RECT 643.640 1739.480 643.900 1739.740 ;
        RECT 643.180 1738.800 643.440 1739.060 ;
        RECT 641.800 1628.300 642.060 1628.560 ;
        RECT 642.260 1628.300 642.520 1628.560 ;
        RECT 643.180 1497.400 643.440 1497.660 ;
        RECT 644.100 1497.400 644.360 1497.660 ;
        RECT 642.260 1452.180 642.520 1452.440 ;
        RECT 643.180 1452.180 643.440 1452.440 ;
        RECT 642.260 1400.500 642.520 1400.760 ;
        RECT 643.180 1400.500 643.440 1400.760 ;
        RECT 642.260 1352.560 642.520 1352.820 ;
        RECT 643.180 1352.560 643.440 1352.820 ;
        RECT 640.420 1303.940 640.680 1304.200 ;
        RECT 642.720 1303.940 642.980 1304.200 ;
        RECT 643.180 1159.100 643.440 1159.360 ;
        RECT 644.100 1159.100 644.360 1159.360 ;
        RECT 642.260 1076.820 642.520 1077.080 ;
        RECT 642.260 1076.140 642.520 1076.400 ;
        RECT 642.260 1014.260 642.520 1014.520 ;
        RECT 643.180 1014.260 643.440 1014.520 ;
        RECT 641.800 979.240 642.060 979.500 ;
        RECT 642.720 979.240 642.980 979.500 ;
        RECT 641.800 917.700 642.060 917.960 ;
        RECT 642.720 917.700 642.980 917.960 ;
        RECT 642.720 883.360 642.980 883.620 ;
        RECT 643.180 882.680 643.440 882.940 ;
        RECT 641.800 845.280 642.060 845.540 ;
        RECT 642.720 845.280 642.980 845.540 ;
        RECT 643.180 675.960 643.440 676.220 ;
        RECT 643.640 675.960 643.900 676.220 ;
        RECT 643.640 641.620 643.900 641.880 ;
        RECT 643.180 641.280 643.440 641.540 ;
        RECT 643.640 627.680 643.900 627.940 ;
        RECT 645.480 627.000 645.740 627.260 ;
        RECT 686.420 591.300 686.680 591.560 ;
        RECT 914.580 591.300 914.840 591.560 ;
        RECT 645.480 588.240 645.740 588.500 ;
        RECT 646.860 588.240 647.120 588.500 ;
        RECT 686.420 588.240 686.680 588.500 ;
        RECT 478.500 43.220 478.760 43.480 ;
        RECT 646.860 42.540 647.120 42.800 ;
      LAYER met2 ;
        RECT 645.020 2916.870 645.280 2917.190 ;
        RECT 1737.520 2916.870 1737.780 2917.190 ;
        RECT 645.080 2769.290 645.220 2916.870 ;
        RECT 1737.580 2900.055 1737.720 2916.870 ;
        RECT 1737.450 2896.055 1737.730 2900.055 ;
        RECT 575.560 2768.970 575.820 2769.290 ;
        RECT 642.260 2768.970 642.520 2769.290 ;
        RECT 645.020 2768.970 645.280 2769.290 ;
        RECT 575.620 2759.520 575.760 2768.970 ;
        RECT 642.320 2766.910 642.460 2768.970 ;
        RECT 642.260 2766.590 642.520 2766.910 ;
        RECT 643.180 2766.590 643.440 2766.910 ;
        RECT 575.450 2759.100 575.760 2759.520 ;
        RECT 575.450 2755.520 575.730 2759.100 ;
        RECT 643.240 2719.310 643.380 2766.590 ;
        RECT 643.180 2718.990 643.440 2719.310 ;
        RECT 642.720 2718.310 642.980 2718.630 ;
        RECT 642.780 2704.770 642.920 2718.310 ;
        RECT 642.320 2704.630 642.920 2704.770 ;
        RECT 642.320 2670.690 642.460 2704.630 ;
        RECT 642.260 2670.370 642.520 2670.690 ;
        RECT 642.720 2670.030 642.980 2670.350 ;
        RECT 642.780 2656.750 642.920 2670.030 ;
        RECT 642.260 2656.430 642.520 2656.750 ;
        RECT 642.720 2656.430 642.980 2656.750 ;
        RECT 642.320 2622.410 642.460 2656.430 ;
        RECT 642.260 2622.090 642.520 2622.410 ;
        RECT 643.180 2621.410 643.440 2621.730 ;
        RECT 643.240 2594.870 643.380 2621.410 ;
        RECT 641.800 2594.550 642.060 2594.870 ;
        RECT 643.180 2594.550 643.440 2594.870 ;
        RECT 641.860 2546.250 642.000 2594.550 ;
        RECT 641.800 2545.930 642.060 2546.250 ;
        RECT 643.180 2545.930 643.440 2546.250 ;
        RECT 643.240 2497.970 643.380 2545.930 ;
        RECT 641.800 2497.650 642.060 2497.970 ;
        RECT 643.180 2497.650 643.440 2497.970 ;
        RECT 641.860 2449.350 642.000 2497.650 ;
        RECT 641.800 2449.030 642.060 2449.350 ;
        RECT 643.180 2449.030 643.440 2449.350 ;
        RECT 643.240 2401.750 643.380 2449.030 ;
        RECT 641.800 2401.430 642.060 2401.750 ;
        RECT 643.180 2401.430 643.440 2401.750 ;
        RECT 641.860 2159.670 642.000 2401.430 ;
        RECT 641.800 2159.350 642.060 2159.670 ;
        RECT 643.180 2159.350 643.440 2159.670 ;
        RECT 643.240 2112.070 643.380 2159.350 ;
        RECT 641.800 2111.750 642.060 2112.070 ;
        RECT 643.180 2111.750 643.440 2112.070 ;
        RECT 641.860 1966.550 642.000 2111.750 ;
        RECT 641.800 1966.230 642.060 1966.550 ;
        RECT 643.180 1966.230 643.440 1966.550 ;
        RECT 643.240 1918.610 643.380 1966.230 ;
        RECT 641.800 1918.290 642.060 1918.610 ;
        RECT 643.180 1918.290 643.440 1918.610 ;
        RECT 641.860 1869.990 642.000 1918.290 ;
        RECT 641.800 1869.670 642.060 1869.990 ;
        RECT 642.720 1869.670 642.980 1869.990 ;
        RECT 642.780 1849.250 642.920 1869.670 ;
        RECT 642.720 1848.930 642.980 1849.250 ;
        RECT 643.180 1848.590 643.440 1848.910 ;
        RECT 643.240 1793.685 643.380 1848.590 ;
        RECT 643.170 1793.570 643.450 1793.685 ;
        RECT 643.170 1793.430 643.840 1793.570 ;
        RECT 643.170 1793.315 643.450 1793.430 ;
        RECT 643.700 1739.770 643.840 1793.430 ;
        RECT 643.640 1739.450 643.900 1739.770 ;
        RECT 643.180 1738.770 643.440 1739.090 ;
        RECT 643.240 1714.690 643.380 1738.770 ;
        RECT 642.320 1714.550 643.380 1714.690 ;
        RECT 642.320 1690.890 642.460 1714.550 ;
        RECT 642.320 1690.750 642.920 1690.890 ;
        RECT 642.780 1676.725 642.920 1690.750 ;
        RECT 641.790 1676.355 642.070 1676.725 ;
        RECT 642.710 1676.355 642.990 1676.725 ;
        RECT 641.860 1628.590 642.000 1676.355 ;
        RECT 641.800 1628.270 642.060 1628.590 ;
        RECT 642.260 1628.270 642.520 1628.590 ;
        RECT 642.320 1558.970 642.460 1628.270 ;
        RECT 642.320 1558.830 643.380 1558.970 ;
        RECT 643.240 1511.370 643.380 1558.830 ;
        RECT 643.240 1511.230 644.300 1511.370 ;
        RECT 644.160 1497.690 644.300 1511.230 ;
        RECT 643.180 1497.370 643.440 1497.690 ;
        RECT 644.100 1497.370 644.360 1497.690 ;
        RECT 643.240 1452.470 643.380 1497.370 ;
        RECT 642.260 1452.150 642.520 1452.470 ;
        RECT 643.180 1452.150 643.440 1452.470 ;
        RECT 642.320 1414.130 642.460 1452.150 ;
        RECT 642.320 1413.990 643.380 1414.130 ;
        RECT 643.240 1400.790 643.380 1413.990 ;
        RECT 642.260 1400.470 642.520 1400.790 ;
        RECT 643.180 1400.470 643.440 1400.790 ;
        RECT 642.320 1352.850 642.460 1400.470 ;
        RECT 642.260 1352.530 642.520 1352.850 ;
        RECT 643.180 1352.530 643.440 1352.850 ;
        RECT 643.240 1317.570 643.380 1352.530 ;
        RECT 642.780 1317.430 643.380 1317.570 ;
        RECT 642.780 1304.230 642.920 1317.430 ;
        RECT 640.420 1303.910 640.680 1304.230 ;
        RECT 642.720 1303.910 642.980 1304.230 ;
        RECT 640.480 1256.485 640.620 1303.910 ;
        RECT 640.410 1256.115 640.690 1256.485 ;
        RECT 642.250 1256.115 642.530 1256.485 ;
        RECT 642.320 1221.010 642.460 1256.115 ;
        RECT 642.320 1220.870 642.920 1221.010 ;
        RECT 642.780 1207.410 642.920 1220.870 ;
        RECT 642.780 1207.270 644.300 1207.410 ;
        RECT 644.160 1159.390 644.300 1207.270 ;
        RECT 643.180 1159.070 643.440 1159.390 ;
        RECT 644.100 1159.070 644.360 1159.390 ;
        RECT 643.240 1124.450 643.380 1159.070 ;
        RECT 642.780 1124.310 643.380 1124.450 ;
        RECT 642.780 1110.850 642.920 1124.310 ;
        RECT 642.320 1110.710 642.920 1110.850 ;
        RECT 642.320 1077.110 642.460 1110.710 ;
        RECT 642.260 1076.790 642.520 1077.110 ;
        RECT 642.260 1076.110 642.520 1076.430 ;
        RECT 642.320 1062.685 642.460 1076.110 ;
        RECT 642.250 1062.315 642.530 1062.685 ;
        RECT 643.170 1062.315 643.450 1062.685 ;
        RECT 643.240 1014.550 643.380 1062.315 ;
        RECT 642.260 1014.230 642.520 1014.550 ;
        RECT 643.180 1014.230 643.440 1014.550 ;
        RECT 642.320 990.490 642.460 1014.230 ;
        RECT 641.860 990.350 642.460 990.490 ;
        RECT 641.860 979.530 642.000 990.350 ;
        RECT 641.800 979.210 642.060 979.530 ;
        RECT 642.720 979.210 642.980 979.530 ;
        RECT 642.780 966.125 642.920 979.210 ;
        RECT 641.790 965.755 642.070 966.125 ;
        RECT 642.710 965.755 642.990 966.125 ;
        RECT 641.860 917.990 642.000 965.755 ;
        RECT 641.800 917.670 642.060 917.990 ;
        RECT 642.720 917.670 642.980 917.990 ;
        RECT 642.780 883.650 642.920 917.670 ;
        RECT 642.720 883.330 642.980 883.650 ;
        RECT 643.180 882.650 643.440 882.970 ;
        RECT 643.240 869.450 643.380 882.650 ;
        RECT 642.780 869.310 643.380 869.450 ;
        RECT 642.780 845.570 642.920 869.310 ;
        RECT 641.800 845.250 642.060 845.570 ;
        RECT 642.720 845.250 642.980 845.570 ;
        RECT 641.860 821.285 642.000 845.250 ;
        RECT 641.790 820.915 642.070 821.285 ;
        RECT 642.710 820.915 642.990 821.285 ;
        RECT 642.780 774.365 642.920 820.915 ;
        RECT 642.710 773.995 642.990 774.365 ;
        RECT 642.710 772.635 642.990 773.005 ;
        RECT 642.780 676.330 642.920 772.635 ;
        RECT 642.780 676.250 643.380 676.330 ;
        RECT 642.780 676.190 643.440 676.250 ;
        RECT 643.180 675.930 643.440 676.190 ;
        RECT 643.640 675.930 643.900 676.250 ;
        RECT 643.240 675.775 643.380 675.930 ;
        RECT 643.700 641.910 643.840 675.930 ;
        RECT 643.640 641.590 643.900 641.910 ;
        RECT 643.180 641.250 643.440 641.570 ;
        RECT 643.240 628.050 643.380 641.250 ;
        RECT 643.240 627.970 643.840 628.050 ;
        RECT 643.240 627.910 643.900 627.970 ;
        RECT 643.640 627.650 643.900 627.910 ;
        RECT 645.480 626.970 645.740 627.290 ;
        RECT 645.540 588.530 645.680 626.970 ;
        RECT 916.190 600.170 916.470 604.000 ;
        RECT 914.640 600.030 916.470 600.170 ;
        RECT 914.640 591.590 914.780 600.030 ;
        RECT 916.190 600.000 916.470 600.030 ;
        RECT 686.420 591.270 686.680 591.590 ;
        RECT 914.580 591.270 914.840 591.590 ;
        RECT 686.480 588.530 686.620 591.270 ;
        RECT 645.480 588.210 645.740 588.530 ;
        RECT 646.860 588.210 647.120 588.530 ;
        RECT 686.420 588.210 686.680 588.530 ;
        RECT 478.500 43.190 478.760 43.510 ;
        RECT 478.560 2.400 478.700 43.190 ;
        RECT 646.920 42.830 647.060 588.210 ;
        RECT 646.860 42.510 647.120 42.830 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 643.170 1793.360 643.450 1793.640 ;
        RECT 641.790 1676.400 642.070 1676.680 ;
        RECT 642.710 1676.400 642.990 1676.680 ;
        RECT 640.410 1256.160 640.690 1256.440 ;
        RECT 642.250 1256.160 642.530 1256.440 ;
        RECT 642.250 1062.360 642.530 1062.640 ;
        RECT 643.170 1062.360 643.450 1062.640 ;
        RECT 641.790 965.800 642.070 966.080 ;
        RECT 642.710 965.800 642.990 966.080 ;
        RECT 641.790 820.960 642.070 821.240 ;
        RECT 642.710 820.960 642.990 821.240 ;
        RECT 642.710 774.040 642.990 774.320 ;
        RECT 642.710 772.680 642.990 772.960 ;
      LAYER met3 ;
        RECT 643.145 1793.650 643.475 1793.665 ;
        RECT 630.510 1793.350 643.475 1793.650 ;
        RECT 630.510 1791.760 630.810 1793.350 ;
        RECT 643.145 1793.335 643.475 1793.350 ;
        RECT 627.030 1791.160 631.030 1791.760 ;
        RECT 641.765 1676.690 642.095 1676.705 ;
        RECT 642.685 1676.690 643.015 1676.705 ;
        RECT 641.765 1676.390 643.015 1676.690 ;
        RECT 641.765 1676.375 642.095 1676.390 ;
        RECT 642.685 1676.375 643.015 1676.390 ;
        RECT 640.385 1256.450 640.715 1256.465 ;
        RECT 642.225 1256.450 642.555 1256.465 ;
        RECT 640.385 1256.150 642.555 1256.450 ;
        RECT 640.385 1256.135 640.715 1256.150 ;
        RECT 642.225 1256.135 642.555 1256.150 ;
        RECT 642.225 1062.650 642.555 1062.665 ;
        RECT 643.145 1062.650 643.475 1062.665 ;
        RECT 642.225 1062.350 643.475 1062.650 ;
        RECT 642.225 1062.335 642.555 1062.350 ;
        RECT 643.145 1062.335 643.475 1062.350 ;
        RECT 641.765 966.090 642.095 966.105 ;
        RECT 642.685 966.090 643.015 966.105 ;
        RECT 641.765 965.790 643.015 966.090 ;
        RECT 641.765 965.775 642.095 965.790 ;
        RECT 642.685 965.775 643.015 965.790 ;
        RECT 641.765 821.250 642.095 821.265 ;
        RECT 642.685 821.250 643.015 821.265 ;
        RECT 641.765 820.950 643.015 821.250 ;
        RECT 641.765 820.935 642.095 820.950 ;
        RECT 642.685 820.935 643.015 820.950 ;
        RECT 642.685 774.340 643.015 774.345 ;
        RECT 642.430 774.330 643.015 774.340 ;
        RECT 642.230 774.030 643.015 774.330 ;
        RECT 642.430 774.020 643.015 774.030 ;
        RECT 642.685 774.015 643.015 774.020 ;
        RECT 642.685 772.980 643.015 772.985 ;
        RECT 642.430 772.970 643.015 772.980 ;
        RECT 642.430 772.670 643.240 772.970 ;
        RECT 642.430 772.660 643.015 772.670 ;
        RECT 642.685 772.655 643.015 772.660 ;
      LAYER via3 ;
        RECT 642.460 774.020 642.780 774.340 ;
        RECT 642.460 772.660 642.780 772.980 ;
      LAYER met4 ;
        RECT 642.455 774.015 642.785 774.345 ;
        RECT 642.470 772.985 642.770 774.015 ;
        RECT 642.455 772.655 642.785 772.985 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 1687.320 389.550 1687.380 ;
        RECT 496.410 1687.320 496.730 1687.380 ;
        RECT 1649.170 1687.320 1649.490 1687.380 ;
        RECT 389.230 1687.180 1649.490 1687.320 ;
        RECT 389.230 1687.120 389.550 1687.180 ;
        RECT 496.410 1687.120 496.730 1687.180 ;
        RECT 1649.170 1687.120 1649.490 1687.180 ;
        RECT 489.970 37.640 490.290 37.700 ;
        RECT 496.410 37.640 496.730 37.700 ;
        RECT 489.970 37.500 496.730 37.640 ;
        RECT 489.970 37.440 490.290 37.500 ;
        RECT 496.410 37.440 496.730 37.500 ;
      LAYER via ;
        RECT 389.260 1687.120 389.520 1687.380 ;
        RECT 496.440 1687.120 496.700 1687.380 ;
        RECT 1649.200 1687.120 1649.460 1687.380 ;
        RECT 490.000 37.440 490.260 37.700 ;
        RECT 496.440 37.440 496.700 37.700 ;
      LAYER met2 ;
        RECT 1650.970 2500.090 1651.250 2504.000 ;
        RECT 1649.260 2500.000 1651.250 2500.090 ;
        RECT 1649.260 2499.950 1651.170 2500.000 ;
        RECT 387.690 1700.410 387.970 1704.000 ;
        RECT 387.690 1700.270 389.460 1700.410 ;
        RECT 387.690 1700.000 387.970 1700.270 ;
        RECT 389.320 1687.410 389.460 1700.270 ;
        RECT 1649.260 1687.410 1649.400 2499.950 ;
        RECT 389.260 1687.090 389.520 1687.410 ;
        RECT 496.440 1687.090 496.700 1687.410 ;
        RECT 1649.200 1687.090 1649.460 1687.410 ;
        RECT 496.500 589.405 496.640 1687.090 ;
        RECT 925.390 600.170 925.670 604.000 ;
        RECT 924.760 600.030 925.670 600.170 ;
        RECT 924.760 589.405 924.900 600.030 ;
        RECT 925.390 600.000 925.670 600.030 ;
        RECT 489.990 589.035 490.270 589.405 ;
        RECT 496.430 589.035 496.710 589.405 ;
        RECT 924.690 589.035 924.970 589.405 ;
        RECT 490.060 37.730 490.200 589.035 ;
        RECT 490.000 37.410 490.260 37.730 ;
        RECT 496.440 37.410 496.700 37.730 ;
        RECT 496.500 2.400 496.640 37.410 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 489.990 589.080 490.270 589.360 ;
        RECT 496.430 589.080 496.710 589.360 ;
        RECT 924.690 589.080 924.970 589.360 ;
      LAYER met3 ;
        RECT 489.965 589.370 490.295 589.385 ;
        RECT 496.405 589.370 496.735 589.385 ;
        RECT 924.665 589.370 924.995 589.385 ;
        RECT 489.965 589.070 924.995 589.370 ;
        RECT 489.965 589.055 490.295 589.070 ;
        RECT 496.405 589.055 496.735 589.070 ;
        RECT 924.665 589.055 924.995 589.070 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1497.830 2453.000 1498.150 2453.060 ;
        RECT 1502.890 2453.000 1503.210 2453.060 ;
        RECT 1497.830 2452.860 1503.210 2453.000 ;
        RECT 1497.830 2452.800 1498.150 2452.860 ;
        RECT 1502.890 2452.800 1503.210 2452.860 ;
        RECT 364.390 1687.660 364.710 1687.720 ;
        RECT 651.430 1687.660 651.750 1687.720 ;
        RECT 1497.830 1687.660 1498.150 1687.720 ;
        RECT 364.390 1687.520 1498.150 1687.660 ;
        RECT 364.390 1687.460 364.710 1687.520 ;
        RECT 651.430 1687.460 651.750 1687.520 ;
        RECT 1497.830 1687.460 1498.150 1687.520 ;
        RECT 910.870 587.080 911.190 587.140 ;
        RECT 932.490 587.080 932.810 587.140 ;
        RECT 910.870 586.940 932.810 587.080 ;
        RECT 910.870 586.880 911.190 586.940 ;
        RECT 932.490 586.880 932.810 586.940 ;
        RECT 651.430 586.060 651.750 586.120 ;
        RECT 669.370 586.060 669.690 586.120 ;
        RECT 651.430 585.920 669.690 586.060 ;
        RECT 651.430 585.860 651.750 585.920 ;
        RECT 669.370 585.860 669.690 585.920 ;
        RECT 717.210 586.060 717.530 586.120 ;
        RECT 772.410 586.060 772.730 586.120 ;
        RECT 855.670 586.060 855.990 586.120 ;
        RECT 910.870 586.060 911.190 586.120 ;
        RECT 717.210 585.920 772.730 586.060 ;
        RECT 717.210 585.860 717.530 585.920 ;
        RECT 772.410 585.860 772.730 585.920 ;
        RECT 813.900 585.920 855.990 586.060 ;
        RECT 669.370 585.380 669.690 585.440 ;
        RECT 717.210 585.380 717.530 585.440 ;
        RECT 669.370 585.240 717.530 585.380 ;
        RECT 669.370 585.180 669.690 585.240 ;
        RECT 717.210 585.180 717.530 585.240 ;
        RECT 806.910 585.380 807.230 585.440 ;
        RECT 813.900 585.380 814.040 585.920 ;
        RECT 855.670 585.860 855.990 585.920 ;
        RECT 910.500 585.920 911.190 586.060 ;
        RECT 806.910 585.240 814.040 585.380 ;
        RECT 903.510 585.380 903.830 585.440 ;
        RECT 910.500 585.380 910.640 585.920 ;
        RECT 910.870 585.860 911.190 585.920 ;
        RECT 903.510 585.240 910.640 585.380 ;
        RECT 806.910 585.180 807.230 585.240 ;
        RECT 903.510 585.180 903.830 585.240 ;
        RECT 772.410 584.700 772.730 584.760 ;
        RECT 806.910 584.700 807.230 584.760 ;
        RECT 772.410 584.560 807.230 584.700 ;
        RECT 772.410 584.500 772.730 584.560 ;
        RECT 806.910 584.500 807.230 584.560 ;
        RECT 932.490 379.820 932.810 380.080 ;
        RECT 932.580 379.400 932.720 379.820 ;
        RECT 932.490 379.140 932.810 379.400 ;
        RECT 513.890 30.500 514.210 30.560 ;
        RECT 932.490 30.500 932.810 30.560 ;
        RECT 513.890 30.360 932.810 30.500 ;
        RECT 513.890 30.300 514.210 30.360 ;
        RECT 932.490 30.300 932.810 30.360 ;
      LAYER via ;
        RECT 1497.860 2452.800 1498.120 2453.060 ;
        RECT 1502.920 2452.800 1503.180 2453.060 ;
        RECT 364.420 1687.460 364.680 1687.720 ;
        RECT 651.460 1687.460 651.720 1687.720 ;
        RECT 1497.860 1687.460 1498.120 1687.720 ;
        RECT 910.900 586.880 911.160 587.140 ;
        RECT 932.520 586.880 932.780 587.140 ;
        RECT 651.460 585.860 651.720 586.120 ;
        RECT 669.400 585.860 669.660 586.120 ;
        RECT 717.240 585.860 717.500 586.120 ;
        RECT 772.440 585.860 772.700 586.120 ;
        RECT 669.400 585.180 669.660 585.440 ;
        RECT 717.240 585.180 717.500 585.440 ;
        RECT 806.940 585.180 807.200 585.440 ;
        RECT 855.700 585.860 855.960 586.120 ;
        RECT 903.540 585.180 903.800 585.440 ;
        RECT 910.900 585.860 911.160 586.120 ;
        RECT 772.440 584.500 772.700 584.760 ;
        RECT 806.940 584.500 807.200 584.760 ;
        RECT 932.520 379.820 932.780 380.080 ;
        RECT 932.520 379.140 932.780 379.400 ;
        RECT 513.920 30.300 514.180 30.560 ;
        RECT 932.520 30.300 932.780 30.560 ;
      LAYER met2 ;
        RECT 1502.850 2500.000 1503.130 2504.000 ;
        RECT 1502.980 2453.090 1503.120 2500.000 ;
        RECT 1497.860 2452.770 1498.120 2453.090 ;
        RECT 1502.920 2452.770 1503.180 2453.090 ;
        RECT 362.850 1700.410 363.130 1704.000 ;
        RECT 362.850 1700.270 364.620 1700.410 ;
        RECT 362.850 1700.000 363.130 1700.270 ;
        RECT 364.480 1687.750 364.620 1700.270 ;
        RECT 1497.920 1687.750 1498.060 2452.770 ;
        RECT 364.420 1687.430 364.680 1687.750 ;
        RECT 651.460 1687.430 651.720 1687.750 ;
        RECT 1497.860 1687.430 1498.120 1687.750 ;
        RECT 651.520 586.150 651.660 1687.430 ;
        RECT 934.590 600.170 934.870 604.000 ;
        RECT 932.580 600.030 934.870 600.170 ;
        RECT 932.580 587.170 932.720 600.030 ;
        RECT 934.590 600.000 934.870 600.030 ;
        RECT 910.900 586.850 911.160 587.170 ;
        RECT 932.520 586.850 932.780 587.170 ;
        RECT 910.960 586.150 911.100 586.850 ;
        RECT 651.460 585.830 651.720 586.150 ;
        RECT 669.400 585.830 669.660 586.150 ;
        RECT 717.240 585.830 717.500 586.150 ;
        RECT 772.440 585.830 772.700 586.150 ;
        RECT 855.700 586.005 855.960 586.150 ;
        RECT 669.460 585.470 669.600 585.830 ;
        RECT 717.300 585.470 717.440 585.830 ;
        RECT 669.400 585.150 669.660 585.470 ;
        RECT 717.240 585.150 717.500 585.470 ;
        RECT 772.500 584.790 772.640 585.830 ;
        RECT 855.690 585.635 855.970 586.005 ;
        RECT 903.530 585.635 903.810 586.005 ;
        RECT 910.900 585.830 911.160 586.150 ;
        RECT 903.600 585.470 903.740 585.635 ;
        RECT 806.940 585.150 807.200 585.470 ;
        RECT 903.540 585.150 903.800 585.470 ;
        RECT 807.000 584.790 807.140 585.150 ;
        RECT 772.440 584.470 772.700 584.790 ;
        RECT 806.940 584.470 807.200 584.790 ;
        RECT 932.580 380.110 932.720 586.850 ;
        RECT 932.520 379.790 932.780 380.110 ;
        RECT 932.520 379.110 932.780 379.430 ;
        RECT 932.580 30.590 932.720 379.110 ;
        RECT 513.920 30.270 514.180 30.590 ;
        RECT 932.520 30.270 932.780 30.590 ;
        RECT 513.980 2.400 514.120 30.270 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 855.690 585.680 855.970 585.960 ;
        RECT 903.530 585.680 903.810 585.960 ;
      LAYER met3 ;
        RECT 855.665 585.970 855.995 585.985 ;
        RECT 903.505 585.970 903.835 585.985 ;
        RECT 855.665 585.670 903.835 585.970 ;
        RECT 855.665 585.655 855.995 585.670 ;
        RECT 903.505 585.655 903.835 585.670 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 941.690 2039.220 942.010 2039.280 ;
        RECT 1902.630 2039.220 1902.950 2039.280 ;
        RECT 941.690 2039.080 1902.950 2039.220 ;
        RECT 941.690 2039.020 942.010 2039.080 ;
        RECT 1902.630 2039.020 1902.950 2039.080 ;
        RECT 927.890 1780.140 928.210 1780.200 ;
        RECT 941.690 1780.140 942.010 1780.200 ;
        RECT 927.890 1780.000 942.010 1780.140 ;
        RECT 927.890 1779.940 928.210 1780.000 ;
        RECT 941.690 1779.940 942.010 1780.000 ;
        RECT 665.230 843.240 665.550 843.500 ;
        RECT 665.320 842.480 665.460 843.240 ;
        RECT 665.230 842.220 665.550 842.480 ;
        RECT 938.930 598.980 939.250 599.040 ;
        RECT 943.760 598.980 944.080 599.040 ;
        RECT 938.930 598.840 944.080 598.980 ;
        RECT 938.930 598.780 939.250 598.840 ;
        RECT 943.760 598.780 944.080 598.840 ;
        RECT 910.870 591.840 911.190 591.900 ;
        RECT 938.930 591.840 939.250 591.900 ;
        RECT 910.870 591.700 939.250 591.840 ;
        RECT 910.870 591.640 911.190 591.700 ;
        RECT 938.930 591.640 939.250 591.700 ;
        RECT 531.830 29.820 532.150 29.880 ;
        RECT 938.930 29.820 939.250 29.880 ;
        RECT 531.830 29.680 939.250 29.820 ;
        RECT 531.830 29.620 532.150 29.680 ;
        RECT 938.930 29.620 939.250 29.680 ;
      LAYER via ;
        RECT 941.720 2039.020 941.980 2039.280 ;
        RECT 1902.660 2039.020 1902.920 2039.280 ;
        RECT 927.920 1779.940 928.180 1780.200 ;
        RECT 941.720 1779.940 941.980 1780.200 ;
        RECT 665.260 843.240 665.520 843.500 ;
        RECT 665.260 842.220 665.520 842.480 ;
        RECT 938.960 598.780 939.220 599.040 ;
        RECT 943.790 598.780 944.050 599.040 ;
        RECT 910.900 591.640 911.160 591.900 ;
        RECT 938.960 591.640 939.220 591.900 ;
        RECT 531.860 29.620 532.120 29.880 ;
        RECT 938.960 29.620 939.220 29.880 ;
      LAYER met2 ;
        RECT 1902.650 2877.235 1902.930 2877.605 ;
        RECT 1902.720 2039.310 1902.860 2877.235 ;
        RECT 941.720 2038.990 941.980 2039.310 ;
        RECT 1902.660 2038.990 1902.920 2039.310 ;
        RECT 941.780 1780.230 941.920 2038.990 ;
        RECT 927.920 1779.910 928.180 1780.230 ;
        RECT 941.720 1779.910 941.980 1780.230 ;
        RECT 350.610 1777.675 350.890 1778.045 ;
        RECT 350.680 1707.325 350.820 1777.675 ;
        RECT 927.980 1707.325 928.120 1779.910 ;
        RECT 350.610 1706.955 350.890 1707.325 ;
        RECT 671.690 1706.955 671.970 1707.325 ;
        RECT 927.910 1706.955 928.190 1707.325 ;
        RECT 671.760 1000.805 671.900 1706.955 ;
        RECT 671.690 1000.435 671.970 1000.805 ;
        RECT 665.250 924.275 665.530 924.645 ;
        RECT 665.320 843.530 665.460 924.275 ;
        RECT 665.260 843.210 665.520 843.530 ;
        RECT 665.260 842.190 665.520 842.510 ;
        RECT 665.320 588.045 665.460 842.190 ;
        RECT 943.790 600.000 944.070 604.000 ;
        RECT 943.850 599.070 943.990 600.000 ;
        RECT 938.960 598.750 939.220 599.070 ;
        RECT 943.790 598.750 944.050 599.070 ;
        RECT 939.020 591.930 939.160 598.750 ;
        RECT 910.900 591.610 911.160 591.930 ;
        RECT 938.960 591.610 939.220 591.930 ;
        RECT 910.960 590.765 911.100 591.610 ;
        RECT 910.890 590.395 911.170 590.765 ;
        RECT 665.250 587.675 665.530 588.045 ;
        RECT 939.020 29.910 939.160 591.610 ;
        RECT 531.860 29.590 532.120 29.910 ;
        RECT 938.960 29.590 939.220 29.910 ;
        RECT 531.920 2.400 532.060 29.590 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 1902.650 2877.280 1902.930 2877.560 ;
        RECT 350.610 1777.720 350.890 1778.000 ;
        RECT 350.610 1707.000 350.890 1707.280 ;
        RECT 671.690 1707.000 671.970 1707.280 ;
        RECT 927.910 1707.000 928.190 1707.280 ;
        RECT 671.690 1000.480 671.970 1000.760 ;
        RECT 665.250 924.320 665.530 924.600 ;
        RECT 910.890 590.440 911.170 590.720 ;
        RECT 665.250 587.720 665.530 588.000 ;
      LAYER met3 ;
        RECT 1885.335 2879.800 1889.335 2880.080 ;
        RECT 1885.335 2879.480 1889.370 2879.800 ;
        RECT 1889.070 2877.570 1889.370 2879.480 ;
        RECT 1902.625 2877.570 1902.955 2877.585 ;
        RECT 1889.070 2877.270 1902.955 2877.570 ;
        RECT 1902.625 2877.255 1902.955 2877.270 ;
        RECT 350.585 1778.010 350.915 1778.025 ;
        RECT 360.000 1778.010 364.000 1778.160 ;
        RECT 350.585 1777.710 364.000 1778.010 ;
        RECT 350.585 1777.695 350.915 1777.710 ;
        RECT 360.000 1777.560 364.000 1777.710 ;
        RECT 350.585 1707.290 350.915 1707.305 ;
        RECT 671.665 1707.290 671.995 1707.305 ;
        RECT 927.885 1707.290 928.215 1707.305 ;
        RECT 350.585 1706.990 928.215 1707.290 ;
        RECT 350.585 1706.975 350.915 1706.990 ;
        RECT 671.665 1706.975 671.995 1706.990 ;
        RECT 927.885 1706.975 928.215 1706.990 ;
        RECT 665.430 1000.770 665.810 1000.780 ;
        RECT 671.665 1000.770 671.995 1000.785 ;
        RECT 665.430 1000.470 671.995 1000.770 ;
        RECT 665.430 1000.460 665.810 1000.470 ;
        RECT 671.665 1000.455 671.995 1000.470 ;
        RECT 665.225 924.620 665.555 924.625 ;
        RECT 665.225 924.610 665.810 924.620 ;
        RECT 665.000 924.310 665.810 924.610 ;
        RECT 665.225 924.300 665.810 924.310 ;
        RECT 665.225 924.295 665.555 924.300 ;
        RECT 669.110 590.730 669.490 590.740 ;
        RECT 910.865 590.730 911.195 590.745 ;
        RECT 669.110 590.430 772.490 590.730 ;
        RECT 669.110 590.420 669.490 590.430 ;
        RECT 772.190 590.050 772.490 590.430 ;
        RECT 844.870 590.430 911.195 590.730 ;
        RECT 844.870 590.050 845.170 590.430 ;
        RECT 910.865 590.415 911.195 590.430 ;
        RECT 772.190 589.750 845.170 590.050 ;
        RECT 665.225 588.010 665.555 588.025 ;
        RECT 669.110 588.010 669.490 588.020 ;
        RECT 665.225 587.710 669.490 588.010 ;
        RECT 665.225 587.695 665.555 587.710 ;
        RECT 669.110 587.700 669.490 587.710 ;
      LAYER via3 ;
        RECT 665.460 1000.460 665.780 1000.780 ;
        RECT 665.460 924.300 665.780 924.620 ;
        RECT 669.140 590.420 669.460 590.740 ;
        RECT 669.140 587.700 669.460 588.020 ;
      LAYER met4 ;
        RECT 665.455 1000.455 665.785 1000.785 ;
        RECT 665.470 924.625 665.770 1000.455 ;
        RECT 665.455 924.295 665.785 924.625 ;
        RECT 669.135 590.415 669.465 590.745 ;
        RECT 669.150 588.025 669.450 590.415 ;
        RECT 669.135 587.695 669.465 588.025 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 589.790 1688.000 590.110 1688.060 ;
        RECT 640.850 1688.000 641.170 1688.060 ;
        RECT 1486.330 1688.000 1486.650 1688.060 ;
        RECT 589.790 1687.860 1486.650 1688.000 ;
        RECT 589.790 1687.800 590.110 1687.860 ;
        RECT 640.850 1687.800 641.170 1687.860 ;
        RECT 1486.330 1687.800 1486.650 1687.860 ;
        RECT 640.850 590.480 641.170 590.540 ;
        RECT 665.690 590.480 666.010 590.540 ;
        RECT 640.850 590.340 666.010 590.480 ;
        RECT 640.850 590.280 641.170 590.340 ;
        RECT 665.690 590.280 666.010 590.340 ;
        RECT 638.090 588.440 638.410 588.500 ;
        RECT 640.850 588.440 641.170 588.500 ;
        RECT 638.090 588.300 641.170 588.440 ;
        RECT 638.090 588.240 638.410 588.300 ;
        RECT 640.850 588.240 641.170 588.300 ;
        RECT 665.690 586.740 666.010 586.800 ;
        RECT 952.270 586.740 952.590 586.800 ;
        RECT 665.690 586.600 952.590 586.740 ;
        RECT 665.690 586.540 666.010 586.600 ;
        RECT 952.270 586.540 952.590 586.600 ;
        RECT 549.770 36.620 550.090 36.680 ;
        RECT 638.090 36.620 638.410 36.680 ;
        RECT 549.770 36.480 638.410 36.620 ;
        RECT 549.770 36.420 550.090 36.480 ;
        RECT 638.090 36.420 638.410 36.480 ;
      LAYER via ;
        RECT 589.820 1687.800 590.080 1688.060 ;
        RECT 640.880 1687.800 641.140 1688.060 ;
        RECT 1486.360 1687.800 1486.620 1688.060 ;
        RECT 640.880 590.280 641.140 590.540 ;
        RECT 665.720 590.280 665.980 590.540 ;
        RECT 638.120 588.240 638.380 588.500 ;
        RECT 640.880 588.240 641.140 588.500 ;
        RECT 665.720 586.540 665.980 586.800 ;
        RECT 952.300 586.540 952.560 586.800 ;
        RECT 549.800 36.420 550.060 36.680 ;
        RECT 638.120 36.420 638.380 36.680 ;
      LAYER met2 ;
        RECT 1486.350 2705.195 1486.630 2705.565 ;
        RECT 588.250 1700.410 588.530 1704.000 ;
        RECT 588.250 1700.270 590.020 1700.410 ;
        RECT 588.250 1700.000 588.530 1700.270 ;
        RECT 589.880 1688.090 590.020 1700.270 ;
        RECT 1486.420 1688.090 1486.560 2705.195 ;
        RECT 589.820 1687.770 590.080 1688.090 ;
        RECT 640.880 1687.770 641.140 1688.090 ;
        RECT 1486.360 1687.770 1486.620 1688.090 ;
        RECT 640.940 590.570 641.080 1687.770 ;
        RECT 952.990 600.170 953.270 604.000 ;
        RECT 952.360 600.030 953.270 600.170 ;
        RECT 640.880 590.250 641.140 590.570 ;
        RECT 665.720 590.250 665.980 590.570 ;
        RECT 640.940 588.530 641.080 590.250 ;
        RECT 638.120 588.210 638.380 588.530 ;
        RECT 640.880 588.210 641.140 588.530 ;
        RECT 638.180 36.710 638.320 588.210 ;
        RECT 665.780 586.830 665.920 590.250 ;
        RECT 952.360 586.830 952.500 600.030 ;
        RECT 952.990 600.000 953.270 600.030 ;
        RECT 665.720 586.510 665.980 586.830 ;
        RECT 952.300 586.510 952.560 586.830 ;
        RECT 549.800 36.390 550.060 36.710 ;
        RECT 638.120 36.390 638.380 36.710 ;
        RECT 549.860 2.400 550.000 36.390 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 1486.350 2705.240 1486.630 2705.520 ;
      LAYER met3 ;
        RECT 1500.000 2708.440 1504.000 2708.720 ;
        RECT 1499.910 2708.120 1504.000 2708.440 ;
        RECT 1486.325 2705.530 1486.655 2705.545 ;
        RECT 1499.910 2705.530 1500.210 2708.120 ;
        RECT 1486.325 2705.230 1500.210 2705.530 ;
        RECT 1486.325 2705.215 1486.655 2705.230 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 955.490 2532.560 955.810 2532.620 ;
        RECT 1483.570 2532.560 1483.890 2532.620 ;
        RECT 955.490 2532.420 1483.890 2532.560 ;
        RECT 955.490 2532.360 955.810 2532.420 ;
        RECT 1483.570 2532.360 1483.890 2532.420 ;
        RECT 676.270 1714.520 676.590 1714.580 ;
        RECT 955.490 1714.520 955.810 1714.580 ;
        RECT 676.270 1714.380 955.810 1714.520 ;
        RECT 676.270 1714.320 676.590 1714.380 ;
        RECT 955.490 1714.320 955.810 1714.380 ;
        RECT 644.070 1712.480 644.390 1712.540 ;
        RECT 676.270 1712.480 676.590 1712.540 ;
        RECT 644.070 1712.340 676.590 1712.480 ;
        RECT 644.070 1712.280 644.390 1712.340 ;
        RECT 676.270 1712.280 676.590 1712.340 ;
        RECT 667.530 1000.520 667.850 1000.580 ;
        RECT 676.270 1000.520 676.590 1000.580 ;
        RECT 667.530 1000.380 676.590 1000.520 ;
        RECT 667.530 1000.320 667.850 1000.380 ;
        RECT 676.270 1000.320 676.590 1000.380 ;
        RECT 667.530 949.520 667.850 949.580 ;
        RECT 667.160 949.380 667.850 949.520 ;
        RECT 667.160 948.160 667.300 949.380 ;
        RECT 667.530 949.320 667.850 949.380 ;
        RECT 668.910 948.160 669.230 948.220 ;
        RECT 667.160 948.020 669.230 948.160 ;
        RECT 668.910 947.960 669.230 948.020 ;
        RECT 952.730 586.740 953.050 586.800 ;
        RECT 960.550 586.740 960.870 586.800 ;
        RECT 952.730 586.600 960.870 586.740 ;
        RECT 952.730 586.540 953.050 586.600 ;
        RECT 960.550 586.540 960.870 586.600 ;
        RECT 668.910 586.400 669.230 586.460 ;
        RECT 952.820 586.400 952.960 586.540 ;
        RECT 668.910 586.260 952.960 586.400 ;
        RECT 668.910 586.200 669.230 586.260 ;
        RECT 572.310 53.620 572.630 53.680 ;
        RECT 952.730 53.620 953.050 53.680 ;
        RECT 572.310 53.480 953.050 53.620 ;
        RECT 572.310 53.420 572.630 53.480 ;
        RECT 952.730 53.420 953.050 53.480 ;
        RECT 567.710 15.880 568.030 15.940 ;
        RECT 572.310 15.880 572.630 15.940 ;
        RECT 567.710 15.740 572.630 15.880 ;
        RECT 567.710 15.680 568.030 15.740 ;
        RECT 572.310 15.680 572.630 15.740 ;
      LAYER via ;
        RECT 955.520 2532.360 955.780 2532.620 ;
        RECT 1483.600 2532.360 1483.860 2532.620 ;
        RECT 676.300 1714.320 676.560 1714.580 ;
        RECT 955.520 1714.320 955.780 1714.580 ;
        RECT 644.100 1712.280 644.360 1712.540 ;
        RECT 676.300 1712.280 676.560 1712.540 ;
        RECT 667.560 1000.320 667.820 1000.580 ;
        RECT 676.300 1000.320 676.560 1000.580 ;
        RECT 667.560 949.320 667.820 949.580 ;
        RECT 668.940 947.960 669.200 948.220 ;
        RECT 952.760 586.540 953.020 586.800 ;
        RECT 960.580 586.540 960.840 586.800 ;
        RECT 668.940 586.200 669.200 586.460 ;
        RECT 572.340 53.420 572.600 53.680 ;
        RECT 952.760 53.420 953.020 53.680 ;
        RECT 567.740 15.680 568.000 15.940 ;
        RECT 572.340 15.680 572.600 15.940 ;
      LAYER met2 ;
        RECT 955.520 2532.330 955.780 2532.650 ;
        RECT 1483.590 2532.475 1483.870 2532.845 ;
        RECT 1483.600 2532.330 1483.860 2532.475 ;
        RECT 644.090 1717.835 644.370 1718.205 ;
        RECT 644.160 1712.570 644.300 1717.835 ;
        RECT 955.580 1714.610 955.720 2532.330 ;
        RECT 676.300 1714.290 676.560 1714.610 ;
        RECT 955.520 1714.290 955.780 1714.610 ;
        RECT 676.360 1712.570 676.500 1714.290 ;
        RECT 644.100 1712.250 644.360 1712.570 ;
        RECT 676.300 1712.250 676.560 1712.570 ;
        RECT 676.360 1000.610 676.500 1712.250 ;
        RECT 667.560 1000.290 667.820 1000.610 ;
        RECT 676.300 1000.290 676.560 1000.610 ;
        RECT 667.620 949.610 667.760 1000.290 ;
        RECT 667.560 949.290 667.820 949.610 ;
        RECT 668.940 947.930 669.200 948.250 ;
        RECT 669.000 586.490 669.140 947.930 ;
        RECT 962.190 600.170 962.470 604.000 ;
        RECT 960.640 600.030 962.470 600.170 ;
        RECT 960.640 586.830 960.780 600.030 ;
        RECT 962.190 600.000 962.470 600.030 ;
        RECT 952.760 586.510 953.020 586.830 ;
        RECT 960.580 586.510 960.840 586.830 ;
        RECT 668.940 586.170 669.200 586.490 ;
        RECT 952.820 53.710 952.960 586.510 ;
        RECT 572.340 53.390 572.600 53.710 ;
        RECT 952.760 53.390 953.020 53.710 ;
        RECT 572.400 15.970 572.540 53.390 ;
        RECT 567.740 15.650 568.000 15.970 ;
        RECT 572.340 15.650 572.600 15.970 ;
        RECT 567.800 2.400 567.940 15.650 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1483.590 2532.520 1483.870 2532.800 ;
        RECT 644.090 1717.880 644.370 1718.160 ;
      LAYER met3 ;
        RECT 1500.000 2535.720 1504.000 2536.000 ;
        RECT 1499.910 2535.400 1504.000 2535.720 ;
        RECT 1483.565 2532.810 1483.895 2532.825 ;
        RECT 1499.910 2532.810 1500.210 2535.400 ;
        RECT 1483.565 2532.510 1500.210 2532.810 ;
        RECT 1483.565 2532.495 1483.895 2532.510 ;
        RECT 627.030 1718.170 631.030 1718.320 ;
        RECT 644.065 1718.170 644.395 1718.185 ;
        RECT 627.030 1717.870 644.395 1718.170 ;
        RECT 627.030 1717.720 631.030 1717.870 ;
        RECT 644.065 1717.855 644.395 1717.870 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 438.910 1686.980 439.230 1687.040 ;
        RECT 586.110 1686.980 586.430 1687.040 ;
        RECT 1902.170 1686.980 1902.490 1687.040 ;
        RECT 438.910 1686.840 1902.490 1686.980 ;
        RECT 438.910 1686.780 439.230 1686.840 ;
        RECT 586.110 1686.780 586.430 1686.840 ;
        RECT 1902.170 1686.780 1902.490 1686.840 ;
        RECT 579.670 15.880 579.990 15.940 ;
        RECT 585.650 15.880 585.970 15.940 ;
        RECT 579.670 15.740 585.970 15.880 ;
        RECT 579.670 15.680 579.990 15.740 ;
        RECT 585.650 15.680 585.970 15.740 ;
      LAYER via ;
        RECT 438.940 1686.780 439.200 1687.040 ;
        RECT 586.140 1686.780 586.400 1687.040 ;
        RECT 1902.200 1686.780 1902.460 1687.040 ;
        RECT 579.700 15.680 579.960 15.940 ;
        RECT 585.680 15.680 585.940 15.940 ;
      LAYER met2 ;
        RECT 1902.190 2643.315 1902.470 2643.685 ;
        RECT 437.370 1700.410 437.650 1704.000 ;
        RECT 437.370 1700.270 439.140 1700.410 ;
        RECT 437.370 1700.000 437.650 1700.270 ;
        RECT 439.000 1687.070 439.140 1700.270 ;
        RECT 1902.260 1687.070 1902.400 2643.315 ;
        RECT 438.940 1686.750 439.200 1687.070 ;
        RECT 586.140 1686.750 586.400 1687.070 ;
        RECT 1902.200 1686.750 1902.460 1687.070 ;
        RECT 586.200 588.725 586.340 1686.750 ;
        RECT 971.390 600.170 971.670 604.000 ;
        RECT 969.840 600.030 971.670 600.170 ;
        RECT 969.840 588.725 969.980 600.030 ;
        RECT 971.390 600.000 971.670 600.030 ;
        RECT 586.130 588.355 586.410 588.725 ;
        RECT 969.770 588.355 970.050 588.725 ;
        RECT 586.200 586.685 586.340 588.355 ;
        RECT 579.690 586.315 579.970 586.685 ;
        RECT 586.130 586.315 586.410 586.685 ;
        RECT 579.760 15.970 579.900 586.315 ;
        RECT 579.700 15.650 579.960 15.970 ;
        RECT 585.680 15.650 585.940 15.970 ;
        RECT 585.740 2.400 585.880 15.650 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 1902.190 2643.360 1902.470 2643.640 ;
        RECT 586.130 588.400 586.410 588.680 ;
        RECT 969.770 588.400 970.050 588.680 ;
        RECT 579.690 586.360 579.970 586.640 ;
        RECT 586.130 586.360 586.410 586.640 ;
      LAYER met3 ;
        RECT 1885.335 2644.520 1889.335 2644.800 ;
        RECT 1885.335 2644.200 1889.370 2644.520 ;
        RECT 1889.070 2643.650 1889.370 2644.200 ;
        RECT 1902.165 2643.650 1902.495 2643.665 ;
        RECT 1889.070 2643.350 1902.495 2643.650 ;
        RECT 1902.165 2643.335 1902.495 2643.350 ;
        RECT 586.105 588.690 586.435 588.705 ;
        RECT 969.745 588.690 970.075 588.705 ;
        RECT 586.105 588.390 970.075 588.690 ;
        RECT 586.105 588.375 586.435 588.390 ;
        RECT 969.745 588.375 970.075 588.390 ;
        RECT 579.665 586.650 579.995 586.665 ;
        RECT 586.105 586.650 586.435 586.665 ;
        RECT 579.665 586.350 586.435 586.650 ;
        RECT 579.665 586.335 579.995 586.350 ;
        RECT 586.105 586.335 586.435 586.350 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1472.990 2663.800 1473.310 2663.860 ;
        RECT 1486.790 2663.800 1487.110 2663.860 ;
        RECT 1472.990 2663.660 1487.110 2663.800 ;
        RECT 1472.990 2663.600 1473.310 2663.660 ;
        RECT 1486.790 2663.600 1487.110 2663.660 ;
        RECT 1469.770 2608.040 1470.090 2608.100 ;
        RECT 1472.990 2608.040 1473.310 2608.100 ;
        RECT 1469.770 2607.900 1473.310 2608.040 ;
        RECT 1469.770 2607.840 1470.090 2607.900 ;
        RECT 1472.990 2607.840 1473.310 2607.900 ;
        RECT 426.490 2606.340 426.810 2606.400 ;
        RECT 1469.770 2606.340 1470.090 2606.400 ;
        RECT 426.490 2606.200 1470.090 2606.340 ;
        RECT 426.490 2606.140 426.810 2606.200 ;
        RECT 1469.770 2606.140 1470.090 2606.200 ;
        RECT 988.610 2032.760 988.930 2032.820 ;
        RECT 1469.770 2032.760 1470.090 2032.820 ;
        RECT 988.610 2032.620 1470.090 2032.760 ;
        RECT 988.610 2032.560 988.930 2032.620 ;
        RECT 1469.770 2032.560 1470.090 2032.620 ;
        RECT 1469.770 2032.080 1470.090 2032.140 ;
        RECT 1472.990 2032.080 1473.310 2032.140 ;
        RECT 1469.770 2031.940 1473.310 2032.080 ;
        RECT 1469.770 2031.880 1470.090 2031.940 ;
        RECT 1472.990 2031.880 1473.310 2031.940 ;
        RECT 1472.990 1928.380 1473.310 1928.440 ;
        RECT 1941.270 1928.380 1941.590 1928.440 ;
        RECT 1472.990 1928.240 1941.590 1928.380 ;
        RECT 1472.990 1928.180 1473.310 1928.240 ;
        RECT 1941.270 1928.180 1941.590 1928.240 ;
        RECT 644.530 1828.420 644.850 1828.480 ;
        RECT 988.610 1828.420 988.930 1828.480 ;
        RECT 644.530 1828.280 988.930 1828.420 ;
        RECT 644.530 1828.220 644.850 1828.280 ;
        RECT 988.610 1828.220 988.930 1828.280 ;
        RECT 685.930 594.900 686.250 594.960 ;
        RECT 691.450 594.900 691.770 594.960 ;
        RECT 685.930 594.760 691.770 594.900 ;
        RECT 685.930 594.700 686.250 594.760 ;
        RECT 691.450 594.700 691.770 594.760 ;
        RECT 691.450 593.200 691.770 593.260 ;
        RECT 715.370 593.200 715.690 593.260 ;
        RECT 691.450 593.060 715.690 593.200 ;
        RECT 691.450 593.000 691.770 593.060 ;
        RECT 715.370 593.000 715.690 593.060 ;
        RECT 644.530 591.500 644.850 591.560 ;
        RECT 677.190 591.500 677.510 591.560 ;
        RECT 685.930 591.500 686.250 591.560 ;
        RECT 644.530 591.360 686.250 591.500 ;
        RECT 644.530 591.300 644.850 591.360 ;
        RECT 677.190 591.300 677.510 591.360 ;
        RECT 685.930 591.300 686.250 591.360 ;
        RECT 91.610 31.520 91.930 31.580 ;
        RECT 677.190 31.520 677.510 31.580 ;
        RECT 91.610 31.380 677.510 31.520 ;
        RECT 91.610 31.320 91.930 31.380 ;
        RECT 677.190 31.320 677.510 31.380 ;
      LAYER via ;
        RECT 1473.020 2663.600 1473.280 2663.860 ;
        RECT 1486.820 2663.600 1487.080 2663.860 ;
        RECT 1469.800 2607.840 1470.060 2608.100 ;
        RECT 1473.020 2607.840 1473.280 2608.100 ;
        RECT 426.520 2606.140 426.780 2606.400 ;
        RECT 1469.800 2606.140 1470.060 2606.400 ;
        RECT 988.640 2032.560 988.900 2032.820 ;
        RECT 1469.800 2032.560 1470.060 2032.820 ;
        RECT 1469.800 2031.880 1470.060 2032.140 ;
        RECT 1473.020 2031.880 1473.280 2032.140 ;
        RECT 1473.020 1928.180 1473.280 1928.440 ;
        RECT 1941.300 1928.180 1941.560 1928.440 ;
        RECT 644.560 1828.220 644.820 1828.480 ;
        RECT 988.640 1828.220 988.900 1828.480 ;
        RECT 685.960 594.700 686.220 594.960 ;
        RECT 691.480 594.700 691.740 594.960 ;
        RECT 691.480 593.000 691.740 593.260 ;
        RECT 715.400 593.000 715.660 593.260 ;
        RECT 644.560 591.300 644.820 591.560 ;
        RECT 677.220 591.300 677.480 591.560 ;
        RECT 685.960 591.300 686.220 591.560 ;
        RECT 91.640 31.320 91.900 31.580 ;
        RECT 677.220 31.320 677.480 31.580 ;
      LAYER met2 ;
        RECT 1486.810 2864.315 1487.090 2864.685 ;
        RECT 426.510 2665.075 426.790 2665.445 ;
        RECT 426.580 2606.430 426.720 2665.075 ;
        RECT 1486.880 2663.890 1487.020 2864.315 ;
        RECT 1473.020 2663.570 1473.280 2663.890 ;
        RECT 1486.820 2663.570 1487.080 2663.890 ;
        RECT 1473.080 2608.130 1473.220 2663.570 ;
        RECT 1469.800 2607.810 1470.060 2608.130 ;
        RECT 1473.020 2607.810 1473.280 2608.130 ;
        RECT 1469.860 2606.430 1470.000 2607.810 ;
        RECT 426.520 2606.110 426.780 2606.430 ;
        RECT 1469.800 2606.110 1470.060 2606.430 ;
        RECT 1469.860 2032.850 1470.000 2606.110 ;
        RECT 988.640 2032.530 988.900 2032.850 ;
        RECT 1469.800 2032.530 1470.060 2032.850 ;
        RECT 644.550 1829.355 644.830 1829.725 ;
        RECT 644.620 1828.510 644.760 1829.355 ;
        RECT 988.700 1828.510 988.840 2032.530 ;
        RECT 1469.860 2032.170 1470.000 2032.530 ;
        RECT 1469.800 2031.850 1470.060 2032.170 ;
        RECT 1473.020 2031.850 1473.280 2032.170 ;
        RECT 1473.080 1928.470 1473.220 2031.850 ;
        RECT 1473.020 1928.150 1473.280 1928.470 ;
        RECT 1941.300 1928.150 1941.560 1928.470 ;
        RECT 1941.360 1917.095 1941.500 1928.150 ;
        RECT 1941.250 1913.095 1941.530 1917.095 ;
        RECT 644.560 1828.190 644.820 1828.510 ;
        RECT 988.640 1828.190 988.900 1828.510 ;
        RECT 644.620 591.590 644.760 1828.190 ;
        RECT 717.010 600.170 717.290 604.000 ;
        RECT 715.460 600.030 717.290 600.170 ;
        RECT 685.960 594.670 686.220 594.990 ;
        RECT 691.480 594.670 691.740 594.990 ;
        RECT 686.020 591.590 686.160 594.670 ;
        RECT 691.540 593.290 691.680 594.670 ;
        RECT 715.460 593.290 715.600 600.030 ;
        RECT 717.010 600.000 717.290 600.030 ;
        RECT 691.480 592.970 691.740 593.290 ;
        RECT 715.400 592.970 715.660 593.290 ;
        RECT 644.560 591.270 644.820 591.590 ;
        RECT 677.220 591.270 677.480 591.590 ;
        RECT 685.960 591.270 686.220 591.590 ;
        RECT 677.280 31.610 677.420 591.270 ;
        RECT 91.640 31.290 91.900 31.610 ;
        RECT 677.220 31.290 677.480 31.610 ;
        RECT 91.700 2.400 91.840 31.290 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 1486.810 2864.360 1487.090 2864.640 ;
        RECT 426.510 2665.120 426.790 2665.400 ;
        RECT 644.550 1829.400 644.830 1829.680 ;
      LAYER met3 ;
        RECT 1500.000 2864.840 1504.000 2865.120 ;
        RECT 1486.785 2864.650 1487.115 2864.665 ;
        RECT 1499.910 2864.650 1504.000 2864.840 ;
        RECT 1486.785 2864.520 1504.000 2864.650 ;
        RECT 1486.785 2864.350 1500.210 2864.520 ;
        RECT 1486.785 2864.335 1487.115 2864.350 ;
        RECT 430.000 2668.320 434.000 2668.640 ;
        RECT 429.950 2668.040 434.000 2668.320 ;
        RECT 426.485 2665.410 426.815 2665.425 ;
        RECT 429.950 2665.410 430.250 2668.040 ;
        RECT 426.485 2665.110 430.250 2665.410 ;
        RECT 426.485 2665.095 426.815 2665.110 ;
        RECT 627.030 1829.690 631.030 1829.840 ;
        RECT 644.525 1829.690 644.855 1829.705 ;
        RECT 627.030 1829.390 644.855 1829.690 ;
        RECT 627.030 1829.240 631.030 1829.390 ;
        RECT 644.525 1829.375 644.855 1829.390 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 631.190 2918.460 631.510 2918.520 ;
        RECT 1513.930 2918.460 1514.250 2918.520 ;
        RECT 631.190 2918.320 1514.250 2918.460 ;
        RECT 631.190 2918.260 631.510 2918.320 ;
        RECT 1513.930 2918.260 1514.250 2918.320 ;
        RECT 479.390 1988.220 479.710 1988.280 ;
        RECT 631.190 1988.220 631.510 1988.280 ;
        RECT 479.390 1988.080 631.510 1988.220 ;
        RECT 479.390 1988.020 479.710 1988.080 ;
        RECT 631.190 1988.020 631.510 1988.080 ;
        RECT 603.130 43.080 603.450 43.140 ;
        RECT 603.130 42.940 614.400 43.080 ;
        RECT 603.130 42.880 603.450 42.940 ;
        RECT 614.260 42.400 614.400 42.940 ;
        RECT 631.190 42.400 631.510 42.460 ;
        RECT 614.260 42.260 631.510 42.400 ;
        RECT 631.190 42.200 631.510 42.260 ;
      LAYER via ;
        RECT 631.220 2918.260 631.480 2918.520 ;
        RECT 1513.960 2918.260 1514.220 2918.520 ;
        RECT 479.420 1988.020 479.680 1988.280 ;
        RECT 631.220 1988.020 631.480 1988.280 ;
        RECT 603.160 42.880 603.420 43.140 ;
        RECT 631.220 42.200 631.480 42.460 ;
      LAYER met2 ;
        RECT 631.220 2918.230 631.480 2918.550 ;
        RECT 1513.960 2918.230 1514.220 2918.550 ;
        RECT 631.280 1988.310 631.420 2918.230 ;
        RECT 1514.020 2900.055 1514.160 2918.230 ;
        RECT 1513.890 2896.055 1514.170 2900.055 ;
        RECT 479.420 1987.990 479.680 1988.310 ;
        RECT 631.220 1987.990 631.480 1988.310 ;
        RECT 477.850 1981.250 478.130 1981.750 ;
        RECT 479.480 1981.250 479.620 1987.990 ;
        RECT 477.850 1981.110 479.620 1981.250 ;
        RECT 477.850 1977.750 478.130 1981.110 ;
        RECT 631.280 591.445 631.420 1987.990 ;
        RECT 980.590 600.170 980.870 604.000 ;
        RECT 979.960 600.030 980.870 600.170 ;
        RECT 979.960 591.445 980.100 600.030 ;
        RECT 980.590 600.000 980.870 600.030 ;
        RECT 631.210 591.075 631.490 591.445 ;
        RECT 979.890 591.075 980.170 591.445 ;
        RECT 603.160 42.850 603.420 43.170 ;
        RECT 603.220 2.400 603.360 42.850 ;
        RECT 631.280 42.490 631.420 591.075 ;
        RECT 631.220 42.170 631.480 42.490 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 631.210 591.120 631.490 591.400 ;
        RECT 979.890 591.120 980.170 591.400 ;
      LAYER met3 ;
        RECT 631.185 591.410 631.515 591.425 ;
        RECT 979.865 591.410 980.195 591.425 ;
        RECT 631.185 591.110 980.195 591.410 ;
        RECT 631.185 591.095 631.515 591.110 ;
        RECT 979.865 591.095 980.195 591.110 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 624.290 2916.760 624.610 2916.820 ;
        RECT 1620.650 2916.760 1620.970 2916.820 ;
        RECT 624.290 2916.620 1620.970 2916.760 ;
        RECT 624.290 2916.560 624.610 2916.620 ;
        RECT 1620.650 2916.560 1620.970 2916.620 ;
        RECT 403.950 1988.900 404.270 1988.960 ;
        RECT 620.610 1988.900 620.930 1988.960 ;
        RECT 403.950 1988.760 620.930 1988.900 ;
        RECT 403.950 1988.700 404.270 1988.760 ;
        RECT 620.610 1988.700 620.930 1988.760 ;
        RECT 620.610 1987.200 620.930 1987.260 ;
        RECT 624.290 1987.200 624.610 1987.260 ;
        RECT 628.890 1987.200 629.210 1987.260 ;
        RECT 620.610 1987.060 629.210 1987.200 ;
        RECT 620.610 1987.000 620.930 1987.060 ;
        RECT 624.290 1987.000 624.610 1987.060 ;
        RECT 628.890 1987.000 629.210 1987.060 ;
        RECT 621.070 15.200 621.390 15.260 ;
        RECT 627.510 15.200 627.830 15.260 ;
        RECT 621.070 15.060 627.830 15.200 ;
        RECT 621.070 15.000 621.390 15.060 ;
        RECT 627.510 15.000 627.830 15.060 ;
      LAYER via ;
        RECT 624.320 2916.560 624.580 2916.820 ;
        RECT 1620.680 2916.560 1620.940 2916.820 ;
        RECT 403.980 1988.700 404.240 1988.960 ;
        RECT 620.640 1988.700 620.900 1988.960 ;
        RECT 620.640 1987.000 620.900 1987.260 ;
        RECT 624.320 1987.000 624.580 1987.260 ;
        RECT 628.920 1987.000 629.180 1987.260 ;
        RECT 621.100 15.000 621.360 15.260 ;
        RECT 627.540 15.000 627.800 15.260 ;
      LAYER met2 ;
        RECT 624.320 2916.530 624.580 2916.850 ;
        RECT 1620.680 2916.530 1620.940 2916.850 ;
        RECT 403.980 1988.670 404.240 1988.990 ;
        RECT 620.640 1988.670 620.900 1988.990 ;
        RECT 402.410 1981.250 402.690 1981.750 ;
        RECT 404.040 1981.250 404.180 1988.670 ;
        RECT 620.700 1987.290 620.840 1988.670 ;
        RECT 624.380 1987.290 624.520 2916.530 ;
        RECT 1620.740 2900.055 1620.880 2916.530 ;
        RECT 1620.610 2896.055 1620.890 2900.055 ;
        RECT 620.640 1986.970 620.900 1987.290 ;
        RECT 624.320 1986.970 624.580 1987.290 ;
        RECT 628.920 1986.970 629.180 1987.290 ;
        RECT 402.410 1981.110 404.180 1981.250 ;
        RECT 402.410 1977.750 402.690 1981.110 ;
        RECT 628.980 592.125 629.120 1986.970 ;
        RECT 989.790 600.170 990.070 604.000 ;
        RECT 988.240 600.030 990.070 600.170 ;
        RECT 988.240 592.125 988.380 600.030 ;
        RECT 989.790 600.000 990.070 600.030 ;
        RECT 628.910 591.755 629.190 592.125 ;
        RECT 988.170 591.755 988.450 592.125 ;
        RECT 628.980 590.650 629.120 591.755 ;
        RECT 627.600 590.510 629.120 590.650 ;
        RECT 627.600 15.290 627.740 590.510 ;
        RECT 621.100 14.970 621.360 15.290 ;
        RECT 627.540 14.970 627.800 15.290 ;
        RECT 621.160 2.400 621.300 14.970 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 628.910 591.800 629.190 592.080 ;
        RECT 988.170 591.800 988.450 592.080 ;
      LAYER met3 ;
        RECT 628.885 592.090 629.215 592.105 ;
        RECT 988.145 592.090 988.475 592.105 ;
        RECT 628.885 591.790 988.475 592.090 ;
        RECT 628.885 591.775 629.215 591.790 ;
        RECT 988.145 591.775 988.475 591.790 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 2877.660 551.930 2877.720 ;
        RECT 1483.570 2877.660 1483.890 2877.720 ;
        RECT 551.610 2877.520 1483.890 2877.660 ;
        RECT 551.610 2877.460 551.930 2877.520 ;
        RECT 1483.570 2877.460 1483.890 2877.520 ;
        RECT 547.010 2773.960 547.330 2774.020 ;
        RECT 551.610 2773.960 551.930 2774.020 ;
        RECT 579.670 2773.960 579.990 2774.020 ;
        RECT 547.010 2773.820 579.990 2773.960 ;
        RECT 547.010 2773.760 547.330 2773.820 ;
        RECT 551.610 2773.760 551.930 2773.820 ;
        RECT 579.670 2773.760 579.990 2773.820 ;
        RECT 379.110 1990.600 379.430 1990.660 ;
        RECT 579.670 1990.600 579.990 1990.660 ;
        RECT 636.250 1990.600 636.570 1990.660 ;
        RECT 379.110 1990.460 636.570 1990.600 ;
        RECT 379.110 1990.400 379.430 1990.460 ;
        RECT 579.670 1990.400 579.990 1990.460 ;
        RECT 636.250 1990.400 636.570 1990.460 ;
        RECT 636.250 1703.980 636.570 1704.040 ;
        RECT 2021.770 1703.980 2022.090 1704.040 ;
        RECT 636.250 1703.840 2022.090 1703.980 ;
        RECT 636.250 1703.780 636.570 1703.840 ;
        RECT 2021.770 1703.780 2022.090 1703.840 ;
        RECT 551.610 1700.920 551.930 1700.980 ;
        RECT 636.250 1700.920 636.570 1700.980 ;
        RECT 551.610 1700.780 636.570 1700.920 ;
        RECT 551.610 1700.720 551.930 1700.780 ;
        RECT 636.250 1700.720 636.570 1700.780 ;
        RECT 551.610 591.840 551.930 591.900 ;
        RECT 727.790 591.840 728.110 591.900 ;
        RECT 551.610 591.700 728.110 591.840 ;
        RECT 551.610 591.640 551.930 591.700 ;
        RECT 727.790 591.640 728.110 591.700 ;
        RECT 116.910 590.480 117.230 590.540 ;
        RECT 551.610 590.480 551.930 590.540 ;
        RECT 116.910 590.340 551.930 590.480 ;
        RECT 116.910 590.280 117.230 590.340 ;
        RECT 551.610 590.280 551.930 590.340 ;
      LAYER via ;
        RECT 551.640 2877.460 551.900 2877.720 ;
        RECT 1483.600 2877.460 1483.860 2877.720 ;
        RECT 547.040 2773.760 547.300 2774.020 ;
        RECT 551.640 2773.760 551.900 2774.020 ;
        RECT 579.700 2773.760 579.960 2774.020 ;
        RECT 379.140 1990.400 379.400 1990.660 ;
        RECT 579.700 1990.400 579.960 1990.660 ;
        RECT 636.280 1990.400 636.540 1990.660 ;
        RECT 636.280 1703.780 636.540 1704.040 ;
        RECT 2021.800 1703.780 2022.060 1704.040 ;
        RECT 551.640 1700.720 551.900 1700.980 ;
        RECT 636.280 1700.720 636.540 1700.980 ;
        RECT 551.640 591.640 551.900 591.900 ;
        RECT 727.820 591.640 728.080 591.900 ;
        RECT 116.940 590.280 117.200 590.540 ;
        RECT 551.640 590.280 551.900 590.540 ;
      LAYER met2 ;
        RECT 1483.590 2878.595 1483.870 2878.965 ;
        RECT 1483.660 2877.750 1483.800 2878.595 ;
        RECT 551.640 2877.430 551.900 2877.750 ;
        RECT 1483.600 2877.430 1483.860 2877.750 ;
        RECT 551.700 2774.050 551.840 2877.430 ;
        RECT 547.040 2773.730 547.300 2774.050 ;
        RECT 551.640 2773.730 551.900 2774.050 ;
        RECT 579.700 2773.730 579.960 2774.050 ;
        RECT 547.100 2759.520 547.240 2773.730 ;
        RECT 546.930 2759.100 547.240 2759.520 ;
        RECT 546.930 2755.520 547.210 2759.100 ;
        RECT 579.760 1990.690 579.900 2773.730 ;
        RECT 379.140 1990.370 379.400 1990.690 ;
        RECT 579.700 1990.370 579.960 1990.690 ;
        RECT 636.280 1990.370 636.540 1990.690 ;
        RECT 377.570 1981.250 377.850 1981.750 ;
        RECT 379.200 1981.250 379.340 1990.370 ;
        RECT 377.570 1981.110 379.340 1981.250 ;
        RECT 377.570 1977.750 377.850 1981.110 ;
        RECT 636.340 1704.070 636.480 1990.370 ;
        RECT 2025.890 1750.730 2026.170 1754.000 ;
        RECT 2021.860 1750.590 2026.170 1750.730 ;
        RECT 2021.860 1704.070 2022.000 1750.590 ;
        RECT 2025.890 1750.000 2026.170 1750.590 ;
        RECT 636.280 1703.750 636.540 1704.070 ;
        RECT 2021.800 1703.750 2022.060 1704.070 ;
        RECT 636.340 1701.010 636.480 1703.750 ;
        RECT 551.640 1700.690 551.900 1701.010 ;
        RECT 636.280 1700.690 636.540 1701.010 ;
        RECT 551.700 591.930 551.840 1700.690 ;
        RECT 729.430 600.170 729.710 604.000 ;
        RECT 727.880 600.030 729.710 600.170 ;
        RECT 727.880 591.930 728.020 600.030 ;
        RECT 729.430 600.000 729.710 600.030 ;
        RECT 551.640 591.610 551.900 591.930 ;
        RECT 727.820 591.610 728.080 591.930 ;
        RECT 551.700 590.570 551.840 591.610 ;
        RECT 116.940 590.250 117.200 590.570 ;
        RECT 551.640 590.250 551.900 590.570 ;
        RECT 117.000 17.410 117.140 590.250 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 1483.590 2878.640 1483.870 2878.920 ;
      LAYER met3 ;
        RECT 1500.000 2881.160 1504.000 2881.440 ;
        RECT 1499.910 2880.840 1504.000 2881.160 ;
        RECT 1483.565 2878.930 1483.895 2878.945 ;
        RECT 1499.910 2878.930 1500.210 2880.840 ;
        RECT 1483.565 2878.630 1500.210 2878.930 ;
        RECT 1483.565 2878.615 1483.895 2878.630 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 460.530 2769.880 460.850 2769.940 ;
        RECT 576.450 2769.880 576.770 2769.940 ;
        RECT 460.530 2769.740 576.770 2769.880 ;
        RECT 460.530 2769.680 460.850 2769.740 ;
        RECT 576.450 2769.680 576.770 2769.740 ;
        RECT 558.510 2489.380 558.830 2489.440 ;
        RECT 576.450 2489.380 576.770 2489.440 ;
        RECT 1566.370 2489.380 1566.690 2489.440 ;
        RECT 558.510 2489.240 1566.690 2489.380 ;
        RECT 558.510 2489.180 558.830 2489.240 ;
        RECT 576.450 2489.180 576.770 2489.240 ;
        RECT 1566.370 2489.180 1566.690 2489.240 ;
        RECT 554.830 1994.340 555.150 1994.400 ;
        RECT 558.510 1994.340 558.830 1994.400 ;
        RECT 630.270 1994.340 630.590 1994.400 ;
        RECT 554.830 1994.200 630.590 1994.340 ;
        RECT 554.830 1994.140 555.150 1994.200 ;
        RECT 558.510 1994.140 558.830 1994.200 ;
        RECT 630.270 1994.140 630.590 1994.200 ;
        RECT 630.270 1704.320 630.590 1704.380 ;
        RECT 2042.470 1704.320 2042.790 1704.380 ;
        RECT 630.270 1704.180 2042.790 1704.320 ;
        RECT 630.270 1704.120 630.590 1704.180 ;
        RECT 2042.470 1704.120 2042.790 1704.180 ;
        RECT 572.310 1701.260 572.630 1701.320 ;
        RECT 630.270 1701.260 630.590 1701.320 ;
        RECT 572.310 1701.120 630.590 1701.260 ;
        RECT 572.310 1701.060 572.630 1701.120 ;
        RECT 630.270 1701.060 630.590 1701.120 ;
        RECT 144.510 590.820 144.830 590.880 ;
        RECT 572.310 590.820 572.630 590.880 ;
        RECT 144.510 590.680 572.630 590.820 ;
        RECT 144.510 590.620 144.830 590.680 ;
        RECT 572.310 590.620 572.630 590.680 ;
        RECT 572.310 587.080 572.630 587.140 ;
        RECT 740.210 587.080 740.530 587.140 ;
        RECT 572.310 586.940 740.530 587.080 ;
        RECT 572.310 586.880 572.630 586.940 ;
        RECT 740.210 586.880 740.530 586.940 ;
        RECT 139.450 16.900 139.770 16.960 ;
        RECT 144.510 16.900 144.830 16.960 ;
        RECT 139.450 16.760 144.830 16.900 ;
        RECT 139.450 16.700 139.770 16.760 ;
        RECT 144.510 16.700 144.830 16.760 ;
      LAYER via ;
        RECT 460.560 2769.680 460.820 2769.940 ;
        RECT 576.480 2769.680 576.740 2769.940 ;
        RECT 558.540 2489.180 558.800 2489.440 ;
        RECT 576.480 2489.180 576.740 2489.440 ;
        RECT 1566.400 2489.180 1566.660 2489.440 ;
        RECT 554.860 1994.140 555.120 1994.400 ;
        RECT 558.540 1994.140 558.800 1994.400 ;
        RECT 630.300 1994.140 630.560 1994.400 ;
        RECT 630.300 1704.120 630.560 1704.380 ;
        RECT 2042.500 1704.120 2042.760 1704.380 ;
        RECT 572.340 1701.060 572.600 1701.320 ;
        RECT 630.300 1701.060 630.560 1701.320 ;
        RECT 144.540 590.620 144.800 590.880 ;
        RECT 572.340 590.620 572.600 590.880 ;
        RECT 572.340 586.880 572.600 587.140 ;
        RECT 740.240 586.880 740.500 587.140 ;
        RECT 139.480 16.700 139.740 16.960 ;
        RECT 144.540 16.700 144.800 16.960 ;
      LAYER met2 ;
        RECT 460.560 2769.650 460.820 2769.970 ;
        RECT 576.480 2769.650 576.740 2769.970 ;
        RECT 460.620 2759.520 460.760 2769.650 ;
        RECT 460.450 2759.100 460.760 2759.520 ;
        RECT 460.450 2755.520 460.730 2759.100 ;
        RECT 576.540 2489.470 576.680 2769.650 ;
        RECT 1566.330 2500.000 1566.610 2504.000 ;
        RECT 1566.460 2489.470 1566.600 2500.000 ;
        RECT 558.540 2489.150 558.800 2489.470 ;
        RECT 576.480 2489.150 576.740 2489.470 ;
        RECT 1566.400 2489.150 1566.660 2489.470 ;
        RECT 558.600 1994.430 558.740 2489.150 ;
        RECT 554.860 1994.110 555.120 1994.430 ;
        RECT 558.540 1994.110 558.800 1994.430 ;
        RECT 630.300 1994.110 630.560 1994.430 ;
        RECT 553.290 1981.250 553.570 1981.750 ;
        RECT 554.920 1981.250 555.060 1994.110 ;
        RECT 553.290 1981.110 555.060 1981.250 ;
        RECT 553.290 1977.750 553.570 1981.110 ;
        RECT 630.360 1704.410 630.500 1994.110 ;
        RECT 2048.890 1750.730 2049.170 1754.000 ;
        RECT 2042.560 1750.590 2049.170 1750.730 ;
        RECT 2042.560 1704.410 2042.700 1750.590 ;
        RECT 2048.890 1750.000 2049.170 1750.590 ;
        RECT 630.300 1704.090 630.560 1704.410 ;
        RECT 2042.500 1704.090 2042.760 1704.410 ;
        RECT 630.360 1701.350 630.500 1704.090 ;
        RECT 572.340 1701.030 572.600 1701.350 ;
        RECT 630.300 1701.030 630.560 1701.350 ;
        RECT 572.400 590.910 572.540 1701.030 ;
        RECT 741.850 600.170 742.130 604.000 ;
        RECT 740.300 600.030 742.130 600.170 ;
        RECT 144.540 590.590 144.800 590.910 ;
        RECT 572.340 590.590 572.600 590.910 ;
        RECT 144.600 16.990 144.740 590.590 ;
        RECT 572.400 587.170 572.540 590.590 ;
        RECT 740.300 587.170 740.440 600.030 ;
        RECT 741.850 600.000 742.130 600.030 ;
        RECT 572.340 586.850 572.600 587.170 ;
        RECT 740.240 586.850 740.500 587.170 ;
        RECT 139.480 16.670 139.740 16.990 ;
        RECT 144.540 16.670 144.800 16.990 ;
        RECT 139.540 2.400 139.680 16.670 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 590.250 2494.140 590.570 2494.200 ;
        RECT 1510.250 2494.140 1510.570 2494.200 ;
        RECT 590.250 2494.000 1510.570 2494.140 ;
        RECT 590.250 2493.940 590.570 2494.000 ;
        RECT 1510.250 2493.940 1510.570 2494.000 ;
        RECT 1510.250 2463.200 1510.570 2463.260 ;
        RECT 1510.710 2463.200 1511.030 2463.260 ;
        RECT 1510.250 2463.060 1511.030 2463.200 ;
        RECT 1510.250 2463.000 1510.570 2463.060 ;
        RECT 1510.710 2463.000 1511.030 2463.060 ;
        RECT 1509.790 2456.400 1510.110 2456.460 ;
        RECT 1510.710 2456.400 1511.030 2456.460 ;
        RECT 1509.790 2456.260 1511.030 2456.400 ;
        RECT 1509.790 2456.200 1510.110 2456.260 ;
        RECT 1510.710 2456.200 1511.030 2456.260 ;
        RECT 1509.330 2408.460 1509.650 2408.520 ;
        RECT 1509.790 2408.460 1510.110 2408.520 ;
        RECT 1509.330 2408.320 1510.110 2408.460 ;
        RECT 1509.330 2408.260 1509.650 2408.320 ;
        RECT 1509.790 2408.260 1510.110 2408.320 ;
        RECT 1510.250 2345.360 1510.570 2345.620 ;
        RECT 1510.340 2344.940 1510.480 2345.360 ;
        RECT 1510.250 2344.680 1510.570 2344.940 ;
        RECT 1510.250 2242.880 1510.570 2242.940 ;
        RECT 1511.170 2242.880 1511.490 2242.940 ;
        RECT 1510.250 2242.740 1511.490 2242.880 ;
        RECT 1510.250 2242.680 1510.570 2242.740 ;
        RECT 1511.170 2242.680 1511.490 2242.740 ;
        RECT 1509.330 2194.260 1509.650 2194.320 ;
        RECT 1510.250 2194.260 1510.570 2194.320 ;
        RECT 1509.330 2194.120 1510.570 2194.260 ;
        RECT 1509.330 2194.060 1509.650 2194.120 ;
        RECT 1510.250 2194.060 1510.570 2194.120 ;
        RECT 1509.330 2145.980 1509.650 2146.040 ;
        RECT 1510.250 2145.980 1510.570 2146.040 ;
        RECT 1509.330 2145.840 1510.570 2145.980 ;
        RECT 1509.330 2145.780 1509.650 2145.840 ;
        RECT 1510.250 2145.780 1510.570 2145.840 ;
        RECT 1510.710 2139.180 1511.030 2139.240 ;
        RECT 1510.340 2139.040 1511.030 2139.180 ;
        RECT 1510.340 2138.900 1510.480 2139.040 ;
        RECT 1510.710 2138.980 1511.030 2139.040 ;
        RECT 1510.250 2138.640 1510.570 2138.900 ;
        RECT 1510.250 2090.700 1510.570 2090.960 ;
        RECT 1510.340 2090.280 1510.480 2090.700 ;
        RECT 1510.250 2090.020 1510.570 2090.280 ;
        RECT 1508.870 2008.280 1509.190 2008.340 ;
        RECT 1510.250 2008.280 1510.570 2008.340 ;
        RECT 1508.870 2008.140 1510.570 2008.280 ;
        RECT 1508.870 2008.080 1509.190 2008.140 ;
        RECT 1510.250 2008.080 1510.570 2008.140 ;
        RECT 1509.330 1960.000 1509.650 1960.060 ;
        RECT 1510.250 1960.000 1510.570 1960.060 ;
        RECT 1509.330 1959.860 1510.570 1960.000 ;
        RECT 1509.330 1959.800 1509.650 1959.860 ;
        RECT 1510.250 1959.800 1510.570 1959.860 ;
        RECT 1507.490 1907.640 1507.810 1907.700 ;
        RECT 1509.790 1907.640 1510.110 1907.700 ;
        RECT 1904.470 1907.640 1904.790 1907.700 ;
        RECT 1507.490 1907.500 1904.790 1907.640 ;
        RECT 1507.490 1907.440 1507.810 1907.500 ;
        RECT 1509.790 1907.440 1510.110 1907.500 ;
        RECT 1904.470 1907.440 1904.790 1907.500 ;
        RECT 537.810 1690.380 538.130 1690.440 ;
        RECT 1507.490 1690.380 1507.810 1690.440 ;
        RECT 537.810 1690.240 1406.060 1690.380 ;
        RECT 537.810 1690.180 538.130 1690.240 ;
        RECT 1405.920 1690.040 1406.060 1690.240 ;
        RECT 1406.840 1690.240 1507.810 1690.380 ;
        RECT 1406.840 1690.040 1406.980 1690.240 ;
        RECT 1507.490 1690.180 1507.810 1690.240 ;
        RECT 1405.920 1689.900 1406.980 1690.040 ;
        RECT 158.310 591.160 158.630 591.220 ;
        RECT 537.810 591.160 538.130 591.220 ;
        RECT 158.310 591.020 538.130 591.160 ;
        RECT 158.310 590.960 158.630 591.020 ;
        RECT 537.810 590.960 538.130 591.020 ;
        RECT 537.810 589.460 538.130 589.520 ;
        RECT 749.410 589.460 749.730 589.520 ;
        RECT 537.810 589.320 749.730 589.460 ;
        RECT 537.810 589.260 538.130 589.320 ;
        RECT 749.410 589.260 749.730 589.320 ;
      LAYER via ;
        RECT 590.280 2493.940 590.540 2494.200 ;
        RECT 1510.280 2493.940 1510.540 2494.200 ;
        RECT 1510.280 2463.000 1510.540 2463.260 ;
        RECT 1510.740 2463.000 1511.000 2463.260 ;
        RECT 1509.820 2456.200 1510.080 2456.460 ;
        RECT 1510.740 2456.200 1511.000 2456.460 ;
        RECT 1509.360 2408.260 1509.620 2408.520 ;
        RECT 1509.820 2408.260 1510.080 2408.520 ;
        RECT 1510.280 2345.360 1510.540 2345.620 ;
        RECT 1510.280 2344.680 1510.540 2344.940 ;
        RECT 1510.280 2242.680 1510.540 2242.940 ;
        RECT 1511.200 2242.680 1511.460 2242.940 ;
        RECT 1509.360 2194.060 1509.620 2194.320 ;
        RECT 1510.280 2194.060 1510.540 2194.320 ;
        RECT 1509.360 2145.780 1509.620 2146.040 ;
        RECT 1510.280 2145.780 1510.540 2146.040 ;
        RECT 1510.740 2138.980 1511.000 2139.240 ;
        RECT 1510.280 2138.640 1510.540 2138.900 ;
        RECT 1510.280 2090.700 1510.540 2090.960 ;
        RECT 1510.280 2090.020 1510.540 2090.280 ;
        RECT 1508.900 2008.080 1509.160 2008.340 ;
        RECT 1510.280 2008.080 1510.540 2008.340 ;
        RECT 1509.360 1959.800 1509.620 1960.060 ;
        RECT 1510.280 1959.800 1510.540 1960.060 ;
        RECT 1507.520 1907.440 1507.780 1907.700 ;
        RECT 1509.820 1907.440 1510.080 1907.700 ;
        RECT 1904.500 1907.440 1904.760 1907.700 ;
        RECT 537.840 1690.180 538.100 1690.440 ;
        RECT 1507.520 1690.180 1507.780 1690.440 ;
        RECT 158.340 590.960 158.600 591.220 ;
        RECT 537.840 590.960 538.100 591.220 ;
        RECT 537.840 589.260 538.100 589.520 ;
        RECT 749.440 589.260 749.700 589.520 ;
      LAYER met2 ;
        RECT 590.270 2732.395 590.550 2732.765 ;
        RECT 590.340 2494.230 590.480 2732.395 ;
        RECT 1512.970 2500.090 1513.250 2504.000 ;
        RECT 1511.260 2500.000 1513.250 2500.090 ;
        RECT 1511.260 2499.950 1513.170 2500.000 ;
        RECT 1511.260 2499.410 1511.400 2499.950 ;
        RECT 1510.340 2499.270 1511.400 2499.410 ;
        RECT 1510.340 2494.230 1510.480 2499.270 ;
        RECT 590.280 2493.910 590.540 2494.230 ;
        RECT 1510.280 2493.910 1510.540 2494.230 ;
        RECT 1510.340 2463.290 1510.480 2493.910 ;
        RECT 1510.280 2462.970 1510.540 2463.290 ;
        RECT 1510.740 2462.970 1511.000 2463.290 ;
        RECT 1510.800 2456.490 1510.940 2462.970 ;
        RECT 1509.820 2456.170 1510.080 2456.490 ;
        RECT 1510.740 2456.170 1511.000 2456.490 ;
        RECT 1509.880 2408.550 1510.020 2456.170 ;
        RECT 1509.360 2408.230 1509.620 2408.550 ;
        RECT 1509.820 2408.230 1510.080 2408.550 ;
        RECT 1509.420 2366.925 1509.560 2408.230 ;
        RECT 1509.350 2366.555 1509.630 2366.925 ;
        RECT 1510.270 2366.555 1510.550 2366.925 ;
        RECT 1510.340 2345.650 1510.480 2366.555 ;
        RECT 1510.280 2345.330 1510.540 2345.650 ;
        RECT 1510.280 2344.650 1510.540 2344.970 ;
        RECT 1510.340 2311.730 1510.480 2344.650 ;
        RECT 1510.340 2311.590 1511.400 2311.730 ;
        RECT 1511.260 2242.970 1511.400 2311.590 ;
        RECT 1510.280 2242.650 1510.540 2242.970 ;
        RECT 1511.200 2242.650 1511.460 2242.970 ;
        RECT 1510.340 2194.350 1510.480 2242.650 ;
        RECT 1509.360 2194.030 1509.620 2194.350 ;
        RECT 1510.280 2194.030 1510.540 2194.350 ;
        RECT 1509.420 2146.070 1509.560 2194.030 ;
        RECT 1510.340 2146.070 1510.480 2146.225 ;
        RECT 1509.360 2145.750 1509.620 2146.070 ;
        RECT 1510.280 2145.810 1510.540 2146.070 ;
        RECT 1510.280 2145.750 1510.940 2145.810 ;
        RECT 1510.340 2145.670 1510.940 2145.750 ;
        RECT 1510.800 2139.270 1510.940 2145.670 ;
        RECT 1510.740 2138.950 1511.000 2139.270 ;
        RECT 1510.280 2138.610 1510.540 2138.930 ;
        RECT 1510.340 2090.990 1510.480 2138.610 ;
        RECT 1510.280 2090.670 1510.540 2090.990 ;
        RECT 1510.280 2089.990 1510.540 2090.310 ;
        RECT 1510.340 2008.370 1510.480 2089.990 ;
        RECT 1508.900 2008.050 1509.160 2008.370 ;
        RECT 1510.280 2008.050 1510.540 2008.370 ;
        RECT 1508.960 2007.770 1509.100 2008.050 ;
        RECT 1508.960 2007.630 1509.560 2007.770 ;
        RECT 1509.420 1960.090 1509.560 2007.630 ;
        RECT 1509.360 1959.770 1509.620 1960.090 ;
        RECT 1510.280 1959.770 1510.540 1960.090 ;
        RECT 1510.340 1945.890 1510.480 1959.770 ;
        RECT 1509.880 1945.750 1510.480 1945.890 ;
        RECT 1509.880 1907.730 1510.020 1945.750 ;
        RECT 1507.520 1907.410 1507.780 1907.730 ;
        RECT 1509.820 1907.410 1510.080 1907.730 ;
        RECT 1904.500 1907.410 1904.760 1907.730 ;
        RECT 537.650 1700.410 537.930 1704.000 ;
        RECT 537.650 1700.000 538.040 1700.410 ;
        RECT 537.900 1690.470 538.040 1700.000 ;
        RECT 1507.580 1690.470 1507.720 1907.410 ;
        RECT 1904.560 1907.245 1904.700 1907.410 ;
        RECT 1904.490 1906.875 1904.770 1907.245 ;
        RECT 537.840 1690.150 538.100 1690.470 ;
        RECT 1507.520 1690.150 1507.780 1690.470 ;
        RECT 537.900 591.250 538.040 1690.150 ;
        RECT 751.050 600.170 751.330 604.000 ;
        RECT 749.500 600.030 751.330 600.170 ;
        RECT 158.340 590.930 158.600 591.250 ;
        RECT 537.840 590.930 538.100 591.250 ;
        RECT 158.400 3.130 158.540 590.930 ;
        RECT 537.900 589.550 538.040 590.930 ;
        RECT 749.500 589.550 749.640 600.030 ;
        RECT 751.050 600.000 751.330 600.030 ;
        RECT 537.840 589.230 538.100 589.550 ;
        RECT 749.440 589.230 749.700 589.550 ;
        RECT 157.480 2.990 158.540 3.130 ;
        RECT 157.480 2.400 157.620 2.990 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 590.270 2732.440 590.550 2732.720 ;
        RECT 1509.350 2366.600 1509.630 2366.880 ;
        RECT 1510.270 2366.600 1510.550 2366.880 ;
        RECT 1904.490 1906.920 1904.770 1907.200 ;
      LAYER met3 ;
        RECT 574.800 2733.320 578.800 2733.920 ;
        RECT 578.070 2732.730 578.370 2733.320 ;
        RECT 590.245 2732.730 590.575 2732.745 ;
        RECT 578.070 2732.430 590.575 2732.730 ;
        RECT 590.245 2732.415 590.575 2732.430 ;
        RECT 1509.325 2366.890 1509.655 2366.905 ;
        RECT 1510.245 2366.890 1510.575 2366.905 ;
        RECT 1509.325 2366.590 1510.575 2366.890 ;
        RECT 1509.325 2366.575 1509.655 2366.590 ;
        RECT 1510.245 2366.575 1510.575 2366.590 ;
        RECT 1904.465 1907.210 1904.795 1907.225 ;
        RECT 1904.465 1907.040 1920.650 1907.210 ;
        RECT 1904.465 1906.910 1924.000 1907.040 ;
        RECT 1904.465 1906.895 1904.795 1906.910 ;
        RECT 1920.000 1906.440 1924.000 1906.910 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1653.310 2897.720 1653.630 2897.780 ;
        RECT 1675.850 2897.720 1676.170 2897.780 ;
        RECT 1653.310 2897.580 1676.170 2897.720 ;
        RECT 1653.310 2897.520 1653.630 2897.580 ;
        RECT 1675.850 2897.520 1676.170 2897.580 ;
        RECT 1714.950 2897.040 1715.270 2897.100 ;
        RECT 1692.960 2896.900 1715.270 2897.040 ;
        RECT 1653.310 2896.500 1653.630 2896.760 ;
        RECT 1675.850 2896.500 1676.170 2896.760 ;
        RECT 1389.730 2894.660 1390.050 2894.720 ;
        RECT 1472.990 2894.660 1473.310 2894.720 ;
        RECT 1389.730 2894.520 1473.310 2894.660 ;
        RECT 1389.730 2894.460 1390.050 2894.520 ;
        RECT 1472.990 2894.460 1473.310 2894.520 ;
        RECT 693.290 2893.980 693.610 2894.040 ;
        RECT 762.290 2893.980 762.610 2894.040 ;
        RECT 693.290 2893.840 762.610 2893.980 ;
        RECT 693.290 2893.780 693.610 2893.840 ;
        RECT 762.290 2893.780 762.610 2893.840 ;
        RECT 811.510 2893.980 811.830 2894.040 ;
        RECT 858.890 2893.980 859.210 2894.040 ;
        RECT 811.510 2893.840 859.210 2893.980 ;
        RECT 811.510 2893.780 811.830 2893.840 ;
        RECT 858.890 2893.780 859.210 2893.840 ;
        RECT 908.110 2893.980 908.430 2894.040 ;
        RECT 955.490 2893.980 955.810 2894.040 ;
        RECT 908.110 2893.840 955.810 2893.980 ;
        RECT 908.110 2893.780 908.430 2893.840 ;
        RECT 955.490 2893.780 955.810 2893.840 ;
        RECT 1004.710 2893.980 1005.030 2894.040 ;
        RECT 1052.090 2893.980 1052.410 2894.040 ;
        RECT 1004.710 2893.840 1052.410 2893.980 ;
        RECT 1004.710 2893.780 1005.030 2893.840 ;
        RECT 1052.090 2893.780 1052.410 2893.840 ;
        RECT 1101.310 2893.980 1101.630 2894.040 ;
        RECT 1148.690 2893.980 1149.010 2894.040 ;
        RECT 1101.310 2893.840 1149.010 2893.980 ;
        RECT 1101.310 2893.780 1101.630 2893.840 ;
        RECT 1148.690 2893.780 1149.010 2893.840 ;
        RECT 1197.910 2893.980 1198.230 2894.040 ;
        RECT 1245.290 2893.980 1245.610 2894.040 ;
        RECT 1197.910 2893.840 1245.610 2893.980 ;
        RECT 1197.910 2893.780 1198.230 2893.840 ;
        RECT 1245.290 2893.780 1245.610 2893.840 ;
        RECT 1294.510 2893.980 1294.830 2894.040 ;
        RECT 1341.890 2893.980 1342.210 2894.040 ;
        RECT 1653.400 2893.980 1653.540 2896.500 ;
        RECT 1294.510 2893.840 1342.210 2893.980 ;
        RECT 1294.510 2893.780 1294.830 2893.840 ;
        RECT 1341.890 2893.780 1342.210 2893.840 ;
        RECT 1611.080 2893.840 1653.540 2893.980 ;
        RECT 1485.410 2893.640 1485.730 2893.700 ;
        RECT 1500.590 2893.640 1500.910 2893.700 ;
        RECT 1485.410 2893.500 1500.910 2893.640 ;
        RECT 1485.410 2893.440 1485.730 2893.500 ;
        RECT 1500.590 2893.440 1500.910 2893.500 ;
        RECT 1611.080 2893.300 1611.220 2893.840 ;
        RECT 1547.600 2893.160 1611.220 2893.300 ;
        RECT 575.990 2892.960 576.310 2893.020 ;
        RECT 579.670 2892.960 579.990 2893.020 ;
        RECT 575.990 2892.820 579.990 2892.960 ;
        RECT 575.990 2892.760 576.310 2892.820 ;
        RECT 579.670 2892.760 579.990 2892.820 ;
        RECT 1500.590 2892.620 1500.910 2892.680 ;
        RECT 1547.600 2892.620 1547.740 2893.160 ;
        RECT 1500.590 2892.480 1547.740 2892.620 ;
        RECT 1500.590 2892.420 1500.910 2892.480 ;
        RECT 693.290 2892.280 693.610 2892.340 ;
        RECT 640.940 2892.140 693.610 2892.280 ;
        RECT 627.510 2891.940 627.830 2892.000 ;
        RECT 640.940 2891.940 641.080 2892.140 ;
        RECT 693.290 2892.080 693.610 2892.140 ;
        RECT 762.290 2892.280 762.610 2892.340 ;
        RECT 811.510 2892.280 811.830 2892.340 ;
        RECT 762.290 2892.140 811.830 2892.280 ;
        RECT 762.290 2892.080 762.610 2892.140 ;
        RECT 811.510 2892.080 811.830 2892.140 ;
        RECT 858.890 2892.280 859.210 2892.340 ;
        RECT 908.110 2892.280 908.430 2892.340 ;
        RECT 858.890 2892.140 908.430 2892.280 ;
        RECT 858.890 2892.080 859.210 2892.140 ;
        RECT 908.110 2892.080 908.430 2892.140 ;
        RECT 955.490 2892.280 955.810 2892.340 ;
        RECT 1004.710 2892.280 1005.030 2892.340 ;
        RECT 955.490 2892.140 1005.030 2892.280 ;
        RECT 955.490 2892.080 955.810 2892.140 ;
        RECT 1004.710 2892.080 1005.030 2892.140 ;
        RECT 1052.090 2892.280 1052.410 2892.340 ;
        RECT 1101.310 2892.280 1101.630 2892.340 ;
        RECT 1052.090 2892.140 1101.630 2892.280 ;
        RECT 1052.090 2892.080 1052.410 2892.140 ;
        RECT 1101.310 2892.080 1101.630 2892.140 ;
        RECT 1148.690 2892.280 1149.010 2892.340 ;
        RECT 1197.910 2892.280 1198.230 2892.340 ;
        RECT 1148.690 2892.140 1198.230 2892.280 ;
        RECT 1148.690 2892.080 1149.010 2892.140 ;
        RECT 1197.910 2892.080 1198.230 2892.140 ;
        RECT 1245.290 2892.280 1245.610 2892.340 ;
        RECT 1294.510 2892.280 1294.830 2892.340 ;
        RECT 1245.290 2892.140 1294.830 2892.280 ;
        RECT 1245.290 2892.080 1245.610 2892.140 ;
        RECT 1294.510 2892.080 1294.830 2892.140 ;
        RECT 1341.890 2892.280 1342.210 2892.340 ;
        RECT 1389.730 2892.280 1390.050 2892.340 ;
        RECT 1341.890 2892.140 1390.050 2892.280 ;
        RECT 1341.890 2892.080 1342.210 2892.140 ;
        RECT 1389.730 2892.080 1390.050 2892.140 ;
        RECT 1472.990 2892.280 1473.310 2892.340 ;
        RECT 1485.410 2892.280 1485.730 2892.340 ;
        RECT 1472.990 2892.140 1485.730 2892.280 ;
        RECT 1675.940 2892.280 1676.080 2896.500 ;
        RECT 1692.960 2893.300 1693.100 2896.900 ;
        RECT 1714.950 2896.840 1715.270 2896.900 ;
        RECT 1677.320 2893.160 1693.100 2893.300 ;
        RECT 1677.320 2892.280 1677.460 2893.160 ;
        RECT 1675.940 2892.140 1677.460 2892.280 ;
        RECT 1472.990 2892.080 1473.310 2892.140 ;
        RECT 1485.410 2892.080 1485.730 2892.140 ;
        RECT 627.510 2891.800 641.080 2891.940 ;
        RECT 627.510 2891.740 627.830 2891.800 ;
        RECT 547.930 2594.100 548.250 2594.160 ;
        RECT 569.090 2594.100 569.410 2594.160 ;
        RECT 575.990 2594.100 576.310 2594.160 ;
        RECT 547.930 2593.960 576.310 2594.100 ;
        RECT 547.930 2593.900 548.250 2593.960 ;
        RECT 569.090 2593.900 569.410 2593.960 ;
        RECT 575.990 2593.900 576.310 2593.960 ;
        RECT 639.010 2035.820 639.330 2035.880 ;
        RECT 2056.270 2035.820 2056.590 2035.880 ;
        RECT 639.010 2035.680 2056.590 2035.820 ;
        RECT 639.010 2035.620 639.330 2035.680 ;
        RECT 2056.270 2035.620 2056.590 2035.680 ;
        RECT 567.710 1994.000 568.030 1994.060 ;
        RECT 569.090 1994.000 569.410 1994.060 ;
        RECT 634.870 1994.000 635.190 1994.060 ;
        RECT 639.010 1994.000 639.330 1994.060 ;
        RECT 567.710 1993.860 639.330 1994.000 ;
        RECT 567.710 1993.800 568.030 1993.860 ;
        RECT 569.090 1993.800 569.410 1993.860 ;
        RECT 634.870 1993.800 635.190 1993.860 ;
        RECT 639.010 1993.800 639.330 1993.860 ;
        RECT 503.310 1990.940 503.630 1991.000 ;
        RECT 567.710 1990.940 568.030 1991.000 ;
        RECT 503.310 1990.800 568.030 1990.940 ;
        RECT 503.310 1990.740 503.630 1990.800 ;
        RECT 567.710 1990.740 568.030 1990.800 ;
        RECT 575.990 590.480 576.310 590.540 ;
        RECT 634.870 590.480 635.190 590.540 ;
        RECT 575.990 590.340 635.190 590.480 ;
        RECT 575.990 590.280 576.310 590.340 ;
        RECT 634.870 590.280 635.190 590.340 ;
        RECT 174.870 41.380 175.190 41.440 ;
        RECT 575.990 41.380 576.310 41.440 ;
        RECT 174.870 41.240 576.310 41.380 ;
        RECT 174.870 41.180 175.190 41.240 ;
        RECT 575.990 41.180 576.310 41.240 ;
      LAYER via ;
        RECT 1653.340 2897.520 1653.600 2897.780 ;
        RECT 1675.880 2897.520 1676.140 2897.780 ;
        RECT 1653.340 2896.500 1653.600 2896.760 ;
        RECT 1675.880 2896.500 1676.140 2896.760 ;
        RECT 1389.760 2894.460 1390.020 2894.720 ;
        RECT 1473.020 2894.460 1473.280 2894.720 ;
        RECT 693.320 2893.780 693.580 2894.040 ;
        RECT 762.320 2893.780 762.580 2894.040 ;
        RECT 811.540 2893.780 811.800 2894.040 ;
        RECT 858.920 2893.780 859.180 2894.040 ;
        RECT 908.140 2893.780 908.400 2894.040 ;
        RECT 955.520 2893.780 955.780 2894.040 ;
        RECT 1004.740 2893.780 1005.000 2894.040 ;
        RECT 1052.120 2893.780 1052.380 2894.040 ;
        RECT 1101.340 2893.780 1101.600 2894.040 ;
        RECT 1148.720 2893.780 1148.980 2894.040 ;
        RECT 1197.940 2893.780 1198.200 2894.040 ;
        RECT 1245.320 2893.780 1245.580 2894.040 ;
        RECT 1294.540 2893.780 1294.800 2894.040 ;
        RECT 1341.920 2893.780 1342.180 2894.040 ;
        RECT 1485.440 2893.440 1485.700 2893.700 ;
        RECT 1500.620 2893.440 1500.880 2893.700 ;
        RECT 576.020 2892.760 576.280 2893.020 ;
        RECT 579.700 2892.760 579.960 2893.020 ;
        RECT 1500.620 2892.420 1500.880 2892.680 ;
        RECT 627.540 2891.740 627.800 2892.000 ;
        RECT 693.320 2892.080 693.580 2892.340 ;
        RECT 762.320 2892.080 762.580 2892.340 ;
        RECT 811.540 2892.080 811.800 2892.340 ;
        RECT 858.920 2892.080 859.180 2892.340 ;
        RECT 908.140 2892.080 908.400 2892.340 ;
        RECT 955.520 2892.080 955.780 2892.340 ;
        RECT 1004.740 2892.080 1005.000 2892.340 ;
        RECT 1052.120 2892.080 1052.380 2892.340 ;
        RECT 1101.340 2892.080 1101.600 2892.340 ;
        RECT 1148.720 2892.080 1148.980 2892.340 ;
        RECT 1197.940 2892.080 1198.200 2892.340 ;
        RECT 1245.320 2892.080 1245.580 2892.340 ;
        RECT 1294.540 2892.080 1294.800 2892.340 ;
        RECT 1341.920 2892.080 1342.180 2892.340 ;
        RECT 1389.760 2892.080 1390.020 2892.340 ;
        RECT 1473.020 2892.080 1473.280 2892.340 ;
        RECT 1485.440 2892.080 1485.700 2892.340 ;
        RECT 1714.980 2896.840 1715.240 2897.100 ;
        RECT 547.960 2593.900 548.220 2594.160 ;
        RECT 569.120 2593.900 569.380 2594.160 ;
        RECT 576.020 2593.900 576.280 2594.160 ;
        RECT 639.040 2035.620 639.300 2035.880 ;
        RECT 2056.300 2035.620 2056.560 2035.880 ;
        RECT 567.740 1993.800 568.000 1994.060 ;
        RECT 569.120 1993.800 569.380 1994.060 ;
        RECT 634.900 1993.800 635.160 1994.060 ;
        RECT 639.040 1993.800 639.300 1994.060 ;
        RECT 503.340 1990.740 503.600 1991.000 ;
        RECT 567.740 1990.740 568.000 1991.000 ;
        RECT 576.020 590.280 576.280 590.540 ;
        RECT 634.900 590.280 635.160 590.540 ;
        RECT 174.900 41.180 175.160 41.440 ;
        RECT 576.020 41.180 576.280 41.440 ;
      LAYER met2 ;
        RECT 1653.340 2897.490 1653.600 2897.810 ;
        RECT 1675.880 2897.490 1676.140 2897.810 ;
        RECT 1653.400 2896.790 1653.540 2897.490 ;
        RECT 1675.940 2896.790 1676.080 2897.490 ;
        RECT 1716.290 2897.210 1716.570 2900.055 ;
        RECT 1715.040 2897.130 1716.570 2897.210 ;
        RECT 1714.980 2897.070 1716.570 2897.130 ;
        RECT 1714.980 2896.810 1715.240 2897.070 ;
        RECT 1653.340 2896.470 1653.600 2896.790 ;
        RECT 1675.880 2896.470 1676.140 2896.790 ;
        RECT 1716.290 2896.055 1716.570 2897.070 ;
        RECT 1389.760 2894.430 1390.020 2894.750 ;
        RECT 1473.020 2894.430 1473.280 2894.750 ;
        RECT 693.320 2893.750 693.580 2894.070 ;
        RECT 762.320 2893.750 762.580 2894.070 ;
        RECT 811.540 2893.750 811.800 2894.070 ;
        RECT 858.920 2893.750 859.180 2894.070 ;
        RECT 908.140 2893.750 908.400 2894.070 ;
        RECT 955.520 2893.750 955.780 2894.070 ;
        RECT 1004.740 2893.750 1005.000 2894.070 ;
        RECT 1052.120 2893.750 1052.380 2894.070 ;
        RECT 1101.340 2893.750 1101.600 2894.070 ;
        RECT 1148.720 2893.750 1148.980 2894.070 ;
        RECT 1197.940 2893.750 1198.200 2894.070 ;
        RECT 1245.320 2893.750 1245.580 2894.070 ;
        RECT 1294.540 2893.750 1294.800 2894.070 ;
        RECT 1341.920 2893.750 1342.180 2894.070 ;
        RECT 579.760 2893.050 580.360 2893.130 ;
        RECT 576.020 2892.730 576.280 2893.050 ;
        RECT 579.700 2892.990 580.360 2893.050 ;
        RECT 579.700 2892.730 579.960 2892.990 ;
        RECT 547.850 2600.660 548.130 2604.000 ;
        RECT 547.850 2600.000 548.160 2600.660 ;
        RECT 548.020 2594.190 548.160 2600.000 ;
        RECT 576.080 2594.190 576.220 2892.730 ;
        RECT 580.220 2891.885 580.360 2892.990 ;
        RECT 693.380 2892.370 693.520 2893.750 ;
        RECT 762.380 2892.370 762.520 2893.750 ;
        RECT 811.600 2892.370 811.740 2893.750 ;
        RECT 858.980 2892.370 859.120 2893.750 ;
        RECT 908.200 2892.370 908.340 2893.750 ;
        RECT 955.580 2892.370 955.720 2893.750 ;
        RECT 1004.800 2892.370 1004.940 2893.750 ;
        RECT 1052.180 2892.370 1052.320 2893.750 ;
        RECT 1101.400 2892.370 1101.540 2893.750 ;
        RECT 1148.780 2892.370 1148.920 2893.750 ;
        RECT 1198.000 2892.370 1198.140 2893.750 ;
        RECT 1245.380 2892.370 1245.520 2893.750 ;
        RECT 1294.600 2892.370 1294.740 2893.750 ;
        RECT 1341.980 2892.370 1342.120 2893.750 ;
        RECT 1389.820 2892.370 1389.960 2894.430 ;
        RECT 1473.080 2892.370 1473.220 2894.430 ;
        RECT 1485.440 2893.410 1485.700 2893.730 ;
        RECT 1500.620 2893.410 1500.880 2893.730 ;
        RECT 1485.500 2892.370 1485.640 2893.410 ;
        RECT 1500.680 2892.710 1500.820 2893.410 ;
        RECT 1500.620 2892.390 1500.880 2892.710 ;
        RECT 693.320 2892.050 693.580 2892.370 ;
        RECT 762.320 2892.050 762.580 2892.370 ;
        RECT 811.540 2892.050 811.800 2892.370 ;
        RECT 858.920 2892.050 859.180 2892.370 ;
        RECT 908.140 2892.050 908.400 2892.370 ;
        RECT 955.520 2892.050 955.780 2892.370 ;
        RECT 1004.740 2892.050 1005.000 2892.370 ;
        RECT 1052.120 2892.050 1052.380 2892.370 ;
        RECT 1101.340 2892.050 1101.600 2892.370 ;
        RECT 1148.720 2892.050 1148.980 2892.370 ;
        RECT 1197.940 2892.050 1198.200 2892.370 ;
        RECT 1245.320 2892.050 1245.580 2892.370 ;
        RECT 1294.540 2892.050 1294.800 2892.370 ;
        RECT 1341.920 2892.050 1342.180 2892.370 ;
        RECT 1389.760 2892.050 1390.020 2892.370 ;
        RECT 1473.020 2892.050 1473.280 2892.370 ;
        RECT 1485.440 2892.050 1485.700 2892.370 ;
        RECT 627.540 2891.885 627.800 2892.030 ;
        RECT 580.150 2891.515 580.430 2891.885 ;
        RECT 627.530 2891.515 627.810 2891.885 ;
        RECT 547.960 2593.870 548.220 2594.190 ;
        RECT 569.120 2593.870 569.380 2594.190 ;
        RECT 576.020 2593.870 576.280 2594.190 ;
        RECT 569.180 1994.090 569.320 2593.870 ;
        RECT 639.040 2035.590 639.300 2035.910 ;
        RECT 2056.300 2035.590 2056.560 2035.910 ;
        RECT 639.100 1994.090 639.240 2035.590 ;
        RECT 567.740 1993.770 568.000 1994.090 ;
        RECT 569.120 1993.770 569.380 1994.090 ;
        RECT 634.900 1993.770 635.160 1994.090 ;
        RECT 639.040 1993.770 639.300 1994.090 ;
        RECT 567.800 1991.030 567.940 1993.770 ;
        RECT 503.340 1990.710 503.600 1991.030 ;
        RECT 567.740 1990.710 568.000 1991.030 ;
        RECT 502.690 1981.250 502.970 1981.750 ;
        RECT 503.400 1981.250 503.540 1990.710 ;
        RECT 502.690 1981.110 503.540 1981.250 ;
        RECT 502.690 1977.750 502.970 1981.110 ;
        RECT 634.960 593.485 635.100 1993.770 ;
        RECT 2056.360 1917.095 2056.500 2035.590 ;
        RECT 2056.250 1913.095 2056.530 1917.095 ;
        RECT 759.790 600.170 760.070 604.000 ;
        RECT 759.160 600.030 760.070 600.170 ;
        RECT 759.160 593.485 759.300 600.030 ;
        RECT 759.790 600.000 760.070 600.030 ;
        RECT 634.890 593.115 635.170 593.485 ;
        RECT 759.090 593.115 759.370 593.485 ;
        RECT 634.960 590.570 635.100 593.115 ;
        RECT 576.020 590.250 576.280 590.570 ;
        RECT 634.900 590.250 635.160 590.570 ;
        RECT 576.080 41.470 576.220 590.250 ;
        RECT 174.900 41.150 175.160 41.470 ;
        RECT 576.020 41.150 576.280 41.470 ;
        RECT 174.960 2.400 175.100 41.150 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 580.150 2891.560 580.430 2891.840 ;
        RECT 627.530 2891.560 627.810 2891.840 ;
        RECT 634.890 593.160 635.170 593.440 ;
        RECT 759.090 593.160 759.370 593.440 ;
      LAYER met3 ;
        RECT 580.125 2891.850 580.455 2891.865 ;
        RECT 627.505 2891.850 627.835 2891.865 ;
        RECT 580.125 2891.550 627.835 2891.850 ;
        RECT 580.125 2891.535 580.455 2891.550 ;
        RECT 627.505 2891.535 627.835 2891.550 ;
        RECT 634.865 593.450 635.195 593.465 ;
        RECT 759.065 593.450 759.395 593.465 ;
        RECT 634.865 593.150 759.395 593.450 ;
        RECT 634.865 593.135 635.195 593.150 ;
        RECT 759.065 593.135 759.395 593.150 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1673.550 2896.500 1673.870 2896.760 ;
        RECT 1674.470 2896.500 1674.790 2896.760 ;
        RECT 1725.530 2896.500 1725.850 2896.760 ;
        RECT 1673.640 2891.600 1673.780 2896.500 ;
        RECT 1628.560 2891.460 1673.780 2891.600 ;
        RECT 1674.560 2891.600 1674.700 2896.500 ;
        RECT 1693.420 2893.160 1694.940 2893.300 ;
        RECT 1674.560 2891.460 1676.540 2891.600 ;
        RECT 427.870 2891.260 428.190 2891.320 ;
        RECT 427.870 2891.120 1566.600 2891.260 ;
        RECT 427.870 2891.060 428.190 2891.120 ;
        RECT 1566.460 2889.900 1566.600 2891.120 ;
        RECT 1628.560 2890.580 1628.700 2891.460 ;
        RECT 1676.400 2890.920 1676.540 2891.460 ;
        RECT 1693.420 2890.920 1693.560 2893.160 ;
        RECT 1694.800 2892.960 1694.940 2893.160 ;
        RECT 1694.800 2892.820 1696.780 2892.960 ;
        RECT 1696.640 2892.620 1696.780 2892.820 ;
        RECT 1725.620 2892.620 1725.760 2896.500 ;
        RECT 1696.640 2892.480 1725.760 2892.620 ;
        RECT 1676.400 2890.780 1693.560 2890.920 ;
        RECT 1583.480 2890.440 1628.700 2890.580 ;
        RECT 1583.480 2889.900 1583.620 2890.440 ;
        RECT 1566.460 2889.760 1583.620 2889.900 ;
        RECT 996.890 2032.420 997.210 2032.480 ;
        RECT 2014.870 2032.420 2015.190 2032.480 ;
        RECT 996.890 2032.280 2015.190 2032.420 ;
        RECT 996.890 2032.220 997.210 2032.280 ;
        RECT 2014.870 2032.220 2015.190 2032.280 ;
        RECT 419.590 1980.060 419.910 1980.120 ;
        RECT 422.810 1980.060 423.130 1980.120 ;
        RECT 419.590 1979.920 423.130 1980.060 ;
        RECT 419.590 1979.860 419.910 1979.920 ;
        RECT 422.810 1979.860 423.130 1979.920 ;
        RECT 422.810 1978.700 423.130 1978.760 ;
        RECT 422.810 1978.560 496.180 1978.700 ;
        RECT 422.810 1978.500 423.130 1978.560 ;
        RECT 418.670 1978.160 418.990 1978.420 ;
        RECT 496.040 1978.360 496.180 1978.560 ;
        RECT 634.410 1978.360 634.730 1978.420 ;
        RECT 496.040 1978.220 634.730 1978.360 ;
        RECT 634.410 1978.160 634.730 1978.220 ;
        RECT 361.630 1977.680 361.950 1977.740 ;
        RECT 418.760 1977.680 418.900 1978.160 ;
        RECT 361.630 1977.540 418.900 1977.680 ;
        RECT 361.630 1977.480 361.950 1977.540 ;
        RECT 2014.870 1966.460 2015.190 1966.520 ;
        RECT 2019.470 1966.460 2019.790 1966.520 ;
        RECT 2014.870 1966.320 2019.790 1966.460 ;
        RECT 2014.870 1966.260 2015.190 1966.320 ;
        RECT 2019.470 1966.260 2019.790 1966.320 ;
        RECT 634.410 1959.660 634.730 1959.720 ;
        RECT 996.890 1959.660 997.210 1959.720 ;
        RECT 634.410 1959.520 997.210 1959.660 ;
        RECT 634.410 1959.460 634.730 1959.520 ;
        RECT 996.890 1959.460 997.210 1959.520 ;
        RECT 634.410 1931.780 634.730 1931.840 ;
        RECT 651.890 1931.780 652.210 1931.840 ;
        RECT 634.410 1931.640 652.210 1931.780 ;
        RECT 634.410 1931.580 634.730 1931.640 ;
        RECT 651.890 1931.580 652.210 1931.640 ;
        RECT 734.230 591.840 734.550 591.900 ;
        RECT 767.350 591.840 767.670 591.900 ;
        RECT 734.230 591.700 767.670 591.840 ;
        RECT 734.230 591.640 734.550 591.700 ;
        RECT 767.350 591.640 767.670 591.700 ;
        RECT 192.810 51.920 193.130 51.980 ;
        RECT 732.390 51.920 732.710 51.980 ;
        RECT 192.810 51.780 732.710 51.920 ;
        RECT 192.810 51.720 193.130 51.780 ;
        RECT 732.390 51.720 732.710 51.780 ;
      LAYER via ;
        RECT 1673.580 2896.500 1673.840 2896.760 ;
        RECT 1674.500 2896.500 1674.760 2896.760 ;
        RECT 1725.560 2896.500 1725.820 2896.760 ;
        RECT 427.900 2891.060 428.160 2891.320 ;
        RECT 996.920 2032.220 997.180 2032.480 ;
        RECT 2014.900 2032.220 2015.160 2032.480 ;
        RECT 419.620 1979.860 419.880 1980.120 ;
        RECT 422.840 1979.860 423.100 1980.120 ;
        RECT 422.840 1978.500 423.100 1978.760 ;
        RECT 418.700 1978.160 418.960 1978.420 ;
        RECT 634.440 1978.160 634.700 1978.420 ;
        RECT 361.660 1977.480 361.920 1977.740 ;
        RECT 2014.900 1966.260 2015.160 1966.520 ;
        RECT 2019.500 1966.260 2019.760 1966.520 ;
        RECT 634.440 1959.460 634.700 1959.720 ;
        RECT 996.920 1959.460 997.180 1959.720 ;
        RECT 634.440 1931.580 634.700 1931.840 ;
        RECT 651.920 1931.580 652.180 1931.840 ;
        RECT 734.260 591.640 734.520 591.900 ;
        RECT 767.380 591.640 767.640 591.900 ;
        RECT 192.840 51.720 193.100 51.980 ;
        RECT 732.420 51.720 732.680 51.980 ;
      LAYER met2 ;
        RECT 1673.640 2898.430 1674.700 2898.570 ;
        RECT 1673.640 2896.790 1673.780 2898.430 ;
        RECT 1674.560 2896.790 1674.700 2898.430 ;
        RECT 1673.580 2896.470 1673.840 2896.790 ;
        RECT 1674.500 2896.470 1674.760 2896.790 ;
        RECT 1725.560 2896.530 1725.820 2896.790 ;
        RECT 1726.410 2896.530 1726.690 2900.055 ;
        RECT 1725.560 2896.470 1726.690 2896.530 ;
        RECT 1725.620 2896.390 1726.690 2896.470 ;
        RECT 1726.410 2896.055 1726.690 2896.390 ;
        RECT 427.900 2891.030 428.160 2891.350 ;
        RECT 427.960 2688.905 428.100 2891.030 ;
        RECT 427.890 2688.535 428.170 2688.905 ;
        RECT 419.610 2685.475 419.890 2685.845 ;
        RECT 419.680 1980.150 419.820 2685.475 ;
        RECT 996.920 2032.190 997.180 2032.510 ;
        RECT 2014.900 2032.190 2015.160 2032.510 ;
        RECT 419.620 1979.830 419.880 1980.150 ;
        RECT 422.840 1979.830 423.100 1980.150 ;
        RECT 419.680 1978.530 419.820 1979.830 ;
        RECT 422.900 1978.790 423.040 1979.830 ;
        RECT 418.760 1978.450 419.820 1978.530 ;
        RECT 422.840 1978.470 423.100 1978.790 ;
        RECT 418.700 1978.390 419.820 1978.450 ;
        RECT 418.700 1978.130 418.960 1978.390 ;
        RECT 634.440 1978.130 634.700 1978.450 ;
        RECT 361.660 1977.450 361.920 1977.770 ;
        RECT 361.720 1965.045 361.860 1977.450 ;
        RECT 361.650 1964.675 361.930 1965.045 ;
        RECT 634.500 1959.750 634.640 1978.130 ;
        RECT 996.980 1959.750 997.120 2032.190 ;
        RECT 2014.960 1966.550 2015.100 2032.190 ;
        RECT 2014.900 1966.230 2015.160 1966.550 ;
        RECT 2019.500 1966.230 2019.760 1966.550 ;
        RECT 634.440 1959.430 634.700 1959.750 ;
        RECT 996.920 1959.430 997.180 1959.750 ;
        RECT 634.500 1931.870 634.640 1959.430 ;
        RECT 634.440 1931.550 634.700 1931.870 ;
        RECT 651.920 1931.550 652.180 1931.870 ;
        RECT 651.980 590.085 652.120 1931.550 ;
        RECT 2019.560 1916.650 2019.700 1966.230 ;
        RECT 2021.290 1916.650 2021.570 1917.095 ;
        RECT 2019.560 1916.510 2021.570 1916.650 ;
        RECT 2021.290 1913.095 2021.570 1916.510 ;
        RECT 768.990 600.170 769.270 604.000 ;
        RECT 767.440 600.030 769.270 600.170 ;
        RECT 767.440 591.930 767.580 600.030 ;
        RECT 768.990 600.000 769.270 600.030 ;
        RECT 734.260 591.610 734.520 591.930 ;
        RECT 767.380 591.610 767.640 591.930 ;
        RECT 734.320 590.085 734.460 591.610 ;
        RECT 651.910 589.715 652.190 590.085 ;
        RECT 732.410 589.715 732.690 590.085 ;
        RECT 734.250 589.715 734.530 590.085 ;
        RECT 732.480 52.010 732.620 589.715 ;
        RECT 192.840 51.690 193.100 52.010 ;
        RECT 732.420 51.690 732.680 52.010 ;
        RECT 192.900 2.400 193.040 51.690 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 427.890 2688.580 428.170 2688.860 ;
        RECT 419.610 2685.520 419.890 2685.800 ;
        RECT 361.650 1964.720 361.930 1965.000 ;
        RECT 651.910 589.760 652.190 590.040 ;
        RECT 732.410 589.760 732.690 590.040 ;
        RECT 734.250 589.760 734.530 590.040 ;
      LAYER met3 ;
        RECT 427.865 2688.870 428.195 2688.885 ;
        RECT 430.000 2688.870 434.000 2689.040 ;
        RECT 427.865 2688.570 434.000 2688.870 ;
        RECT 427.865 2688.555 428.195 2688.570 ;
        RECT 429.950 2688.440 434.000 2688.570 ;
        RECT 419.585 2685.810 419.915 2685.825 ;
        RECT 429.950 2685.810 430.250 2688.440 ;
        RECT 419.585 2685.510 430.250 2685.810 ;
        RECT 419.585 2685.495 419.915 2685.510 ;
        RECT 361.625 1965.010 361.955 1965.025 ;
        RECT 361.625 1964.695 362.170 1965.010 ;
        RECT 361.870 1963.120 362.170 1964.695 ;
        RECT 360.000 1962.520 364.000 1963.120 ;
        RECT 651.885 590.050 652.215 590.065 ;
        RECT 732.385 590.050 732.715 590.065 ;
        RECT 734.225 590.050 734.555 590.065 ;
        RECT 651.885 589.750 734.555 590.050 ;
        RECT 651.885 589.735 652.215 589.750 ;
        RECT 732.385 589.735 732.715 589.750 ;
        RECT 734.225 589.735 734.555 589.750 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 593.010 2712.080 593.330 2712.140 ;
        RECT 776.090 2712.080 776.410 2712.140 ;
        RECT 593.010 2711.940 776.410 2712.080 ;
        RECT 593.010 2711.880 593.330 2711.940 ;
        RECT 776.090 2711.880 776.410 2711.940 ;
        RECT 776.090 2489.040 776.410 2489.100 ;
        RECT 1598.570 2489.040 1598.890 2489.100 ;
        RECT 776.090 2488.900 1598.890 2489.040 ;
        RECT 776.090 2488.840 776.410 2488.900 ;
        RECT 1598.570 2488.840 1598.890 2488.900 ;
        RECT 776.090 2484.620 776.410 2484.680 ;
        RECT 779.310 2484.620 779.630 2484.680 ;
        RECT 776.090 2484.480 779.630 2484.620 ;
        RECT 776.090 2484.420 776.410 2484.480 ;
        RECT 779.310 2484.420 779.630 2484.480 ;
        RECT 776.090 2038.200 776.410 2038.260 ;
        RECT 779.310 2038.200 779.630 2038.260 ;
        RECT 776.090 2038.060 779.630 2038.200 ;
        RECT 776.090 2038.000 776.410 2038.060 ;
        RECT 779.310 2038.000 779.630 2038.060 ;
        RECT 779.310 2036.160 779.630 2036.220 ;
        RECT 2084.330 2036.160 2084.650 2036.220 ;
        RECT 779.310 2036.020 2084.650 2036.160 ;
        RECT 779.310 2035.960 779.630 2036.020 ;
        RECT 2084.330 2035.960 2084.650 2036.020 ;
        RECT 641.310 1990.600 641.630 1990.660 ;
        RECT 776.090 1990.600 776.410 1990.660 ;
        RECT 641.310 1990.460 776.410 1990.600 ;
        RECT 641.310 1990.400 641.630 1990.460 ;
        RECT 776.090 1990.400 776.410 1990.460 ;
        RECT 429.710 1987.880 430.030 1987.940 ;
        RECT 641.310 1987.880 641.630 1987.940 ;
        RECT 429.710 1987.740 641.630 1987.880 ;
        RECT 429.710 1987.680 430.030 1987.740 ;
        RECT 641.310 1987.680 641.630 1987.740 ;
        RECT 641.310 593.540 641.630 593.600 ;
        RECT 773.330 593.540 773.650 593.600 ;
        RECT 776.550 593.540 776.870 593.600 ;
        RECT 641.310 593.400 776.870 593.540 ;
        RECT 641.310 593.340 641.630 593.400 ;
        RECT 773.330 593.340 773.650 593.400 ;
        RECT 776.550 593.340 776.870 593.400 ;
        RECT 213.510 51.580 213.830 51.640 ;
        RECT 773.330 51.580 773.650 51.640 ;
        RECT 213.510 51.440 773.650 51.580 ;
        RECT 213.510 51.380 213.830 51.440 ;
        RECT 773.330 51.380 773.650 51.440 ;
        RECT 210.750 20.300 211.070 20.360 ;
        RECT 213.510 20.300 213.830 20.360 ;
        RECT 210.750 20.160 213.830 20.300 ;
        RECT 210.750 20.100 211.070 20.160 ;
        RECT 213.510 20.100 213.830 20.160 ;
      LAYER via ;
        RECT 593.040 2711.880 593.300 2712.140 ;
        RECT 776.120 2711.880 776.380 2712.140 ;
        RECT 776.120 2488.840 776.380 2489.100 ;
        RECT 1598.600 2488.840 1598.860 2489.100 ;
        RECT 776.120 2484.420 776.380 2484.680 ;
        RECT 779.340 2484.420 779.600 2484.680 ;
        RECT 776.120 2038.000 776.380 2038.260 ;
        RECT 779.340 2038.000 779.600 2038.260 ;
        RECT 779.340 2035.960 779.600 2036.220 ;
        RECT 2084.360 2035.960 2084.620 2036.220 ;
        RECT 641.340 1990.400 641.600 1990.660 ;
        RECT 776.120 1990.400 776.380 1990.660 ;
        RECT 429.740 1987.680 430.000 1987.940 ;
        RECT 641.340 1987.680 641.600 1987.940 ;
        RECT 641.340 593.340 641.600 593.600 ;
        RECT 773.360 593.340 773.620 593.600 ;
        RECT 776.580 593.340 776.840 593.600 ;
        RECT 213.540 51.380 213.800 51.640 ;
        RECT 773.360 51.380 773.620 51.640 ;
        RECT 210.780 20.100 211.040 20.360 ;
        RECT 213.540 20.100 213.800 20.360 ;
      LAYER met2 ;
        RECT 593.030 2711.995 593.310 2712.365 ;
        RECT 593.040 2711.850 593.300 2711.995 ;
        RECT 776.120 2711.850 776.380 2712.170 ;
        RECT 776.180 2489.130 776.320 2711.850 ;
        RECT 1598.530 2500.000 1598.810 2504.000 ;
        RECT 1598.660 2489.130 1598.800 2500.000 ;
        RECT 776.120 2488.810 776.380 2489.130 ;
        RECT 1598.600 2488.810 1598.860 2489.130 ;
        RECT 776.180 2484.710 776.320 2488.810 ;
        RECT 776.120 2484.390 776.380 2484.710 ;
        RECT 779.340 2484.390 779.600 2484.710 ;
        RECT 779.400 2038.290 779.540 2484.390 ;
        RECT 776.120 2037.970 776.380 2038.290 ;
        RECT 779.340 2037.970 779.600 2038.290 ;
        RECT 776.180 1990.690 776.320 2037.970 ;
        RECT 779.400 2036.250 779.540 2037.970 ;
        RECT 779.340 2035.930 779.600 2036.250 ;
        RECT 2084.360 2035.930 2084.620 2036.250 ;
        RECT 641.340 1990.370 641.600 1990.690 ;
        RECT 776.120 1990.370 776.380 1990.690 ;
        RECT 641.400 1987.970 641.540 1990.370 ;
        RECT 429.740 1987.650 430.000 1987.970 ;
        RECT 641.340 1987.650 641.600 1987.970 ;
        RECT 428.170 1981.250 428.450 1981.750 ;
        RECT 429.800 1981.250 429.940 1987.650 ;
        RECT 428.170 1981.110 429.940 1981.250 ;
        RECT 428.170 1977.750 428.450 1981.110 ;
        RECT 641.400 593.630 641.540 1987.650 ;
        RECT 2084.420 1904.525 2084.560 2035.930 ;
        RECT 2084.350 1904.155 2084.630 1904.525 ;
        RECT 778.190 600.170 778.470 604.000 ;
        RECT 776.640 600.030 778.470 600.170 ;
        RECT 776.640 593.630 776.780 600.030 ;
        RECT 778.190 600.000 778.470 600.030 ;
        RECT 641.340 593.310 641.600 593.630 ;
        RECT 773.360 593.310 773.620 593.630 ;
        RECT 776.580 593.310 776.840 593.630 ;
        RECT 773.420 51.670 773.560 593.310 ;
        RECT 213.540 51.350 213.800 51.670 ;
        RECT 773.360 51.350 773.620 51.670 ;
        RECT 213.600 20.390 213.740 51.350 ;
        RECT 210.780 20.070 211.040 20.390 ;
        RECT 213.540 20.070 213.800 20.390 ;
        RECT 210.840 2.400 210.980 20.070 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 593.030 2712.040 593.310 2712.320 ;
        RECT 2084.350 1904.200 2084.630 1904.480 ;
      LAYER met3 ;
        RECT 593.005 2712.330 593.335 2712.345 ;
        RECT 578.070 2712.160 593.335 2712.330 ;
        RECT 574.800 2712.030 593.335 2712.160 ;
        RECT 574.800 2711.560 578.800 2712.030 ;
        RECT 593.005 2712.015 593.335 2712.030 ;
        RECT 2084.325 1904.490 2084.655 1904.505 ;
        RECT 2075.830 1904.320 2084.655 1904.490 ;
        RECT 2072.375 1904.190 2084.655 1904.320 ;
        RECT 2072.375 1903.720 2076.375 1904.190 ;
        RECT 2084.325 1904.175 2084.655 1904.190 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 489.970 2592.060 490.290 2592.120 ;
        RECT 638.090 2592.060 638.410 2592.120 ;
        RECT 489.970 2591.920 638.410 2592.060 ;
        RECT 489.970 2591.860 490.290 2591.920 ;
        RECT 638.090 2591.860 638.410 2591.920 ;
        RECT 641.310 2489.720 641.630 2489.780 ;
        RECT 1672.170 2489.720 1672.490 2489.780 ;
        RECT 641.310 2489.580 1672.490 2489.720 ;
        RECT 641.310 2489.520 641.630 2489.580 ;
        RECT 1672.170 2489.520 1672.490 2489.580 ;
        RECT 638.090 2488.020 638.410 2488.080 ;
        RECT 641.310 2488.020 641.630 2488.080 ;
        RECT 638.090 2487.880 641.630 2488.020 ;
        RECT 638.090 2487.820 638.410 2487.880 ;
        RECT 641.310 2487.820 641.630 2487.880 ;
        RECT 627.970 1991.280 628.290 1991.340 ;
        RECT 641.310 1991.280 641.630 1991.340 ;
        RECT 690.070 1991.280 690.390 1991.340 ;
        RECT 627.970 1991.140 690.390 1991.280 ;
        RECT 627.970 1991.080 628.290 1991.140 ;
        RECT 641.310 1991.080 641.630 1991.140 ;
        RECT 690.070 1991.080 690.390 1991.140 ;
        RECT 869.470 1702.620 869.790 1702.680 ;
        RECT 834.600 1702.480 869.790 1702.620 ;
        RECT 650.970 1702.280 651.290 1702.340 ;
        RECT 690.070 1702.280 690.390 1702.340 ;
        RECT 772.870 1702.280 773.190 1702.340 ;
        RECT 834.600 1702.280 834.740 1702.480 ;
        RECT 869.470 1702.420 869.790 1702.480 ;
        RECT 1014.000 1702.480 1028.400 1702.620 ;
        RECT 1014.000 1702.340 1014.140 1702.480 ;
        RECT 650.970 1702.140 773.190 1702.280 ;
        RECT 650.970 1702.080 651.290 1702.140 ;
        RECT 690.070 1702.080 690.390 1702.140 ;
        RECT 772.870 1702.080 773.190 1702.140 ;
        RECT 820.800 1702.140 834.740 1702.280 ;
        RECT 917.310 1702.280 917.630 1702.340 ;
        RECT 917.310 1702.140 931.340 1702.280 ;
        RECT 786.670 1701.940 786.990 1702.000 ;
        RECT 820.800 1701.940 820.940 1702.140 ;
        RECT 917.310 1702.080 917.630 1702.140 ;
        RECT 786.670 1701.800 820.940 1701.940 ;
        RECT 931.200 1701.940 931.340 1702.140 ;
        RECT 1013.910 1702.080 1014.230 1702.340 ;
        RECT 1028.260 1702.280 1028.400 1702.480 ;
        RECT 1200.670 1702.420 1200.990 1702.680 ;
        RECT 1296.900 1702.480 1297.500 1702.620 ;
        RECT 1076.010 1702.280 1076.330 1702.340 ;
        RECT 1028.260 1702.140 1076.330 1702.280 ;
        RECT 1076.010 1702.080 1076.330 1702.140 ;
        RECT 1200.210 1702.280 1200.530 1702.340 ;
        RECT 1200.760 1702.280 1200.900 1702.420 ;
        RECT 1200.210 1702.140 1200.900 1702.280 ;
        RECT 1248.510 1702.280 1248.830 1702.340 ;
        RECT 1296.900 1702.280 1297.040 1702.480 ;
        RECT 1297.360 1702.340 1297.500 1702.480 ;
        RECT 1345.110 1702.420 1345.430 1702.680 ;
        RECT 1400.770 1702.620 1401.090 1702.680 ;
        RECT 1393.500 1702.480 1401.090 1702.620 ;
        RECT 1248.510 1702.140 1297.040 1702.280 ;
        RECT 1200.210 1702.080 1200.530 1702.140 ;
        RECT 1248.510 1702.080 1248.830 1702.140 ;
        RECT 1297.270 1702.080 1297.590 1702.340 ;
        RECT 1345.200 1702.280 1345.340 1702.420 ;
        RECT 1345.570 1702.280 1345.890 1702.340 ;
        RECT 1345.200 1702.140 1345.890 1702.280 ;
        RECT 1345.570 1702.080 1345.890 1702.140 ;
        RECT 1366.270 1702.280 1366.590 1702.340 ;
        RECT 1393.500 1702.280 1393.640 1702.480 ;
        RECT 1400.770 1702.420 1401.090 1702.480 ;
        RECT 1704.000 1702.480 1751.980 1702.620 ;
        RECT 1366.270 1702.140 1393.640 1702.280 ;
        RECT 1666.190 1702.280 1666.510 1702.340 ;
        RECT 1704.000 1702.280 1704.140 1702.480 ;
        RECT 1666.190 1702.140 1704.140 1702.280 ;
        RECT 1366.270 1702.080 1366.590 1702.140 ;
        RECT 1666.190 1702.080 1666.510 1702.140 ;
        RECT 966.070 1701.940 966.390 1702.000 ;
        RECT 931.200 1701.800 966.390 1701.940 ;
        RECT 786.670 1701.740 786.990 1701.800 ;
        RECT 966.070 1701.740 966.390 1701.800 ;
        RECT 1124.770 1701.940 1125.090 1702.000 ;
        RECT 1152.370 1701.940 1152.690 1702.000 ;
        RECT 1462.410 1701.940 1462.730 1702.000 ;
        RECT 1594.430 1701.940 1594.750 1702.000 ;
        RECT 1655.610 1701.940 1655.930 1702.000 ;
        RECT 1124.770 1701.800 1152.690 1701.940 ;
        RECT 1124.770 1701.740 1125.090 1701.800 ;
        RECT 1152.370 1701.740 1152.690 1701.800 ;
        RECT 1424.780 1701.800 1462.730 1701.940 ;
        RECT 869.930 1701.600 870.250 1701.660 ;
        RECT 917.310 1701.600 917.630 1701.660 ;
        RECT 869.930 1701.460 917.630 1701.600 ;
        RECT 869.930 1701.400 870.250 1701.460 ;
        RECT 917.310 1701.400 917.630 1701.460 ;
        RECT 1076.930 1701.600 1077.250 1701.660 ;
        RECT 1124.310 1701.600 1124.630 1701.660 ;
        RECT 1076.930 1701.460 1124.630 1701.600 ;
        RECT 1076.930 1701.400 1077.250 1701.460 ;
        RECT 1124.310 1701.400 1124.630 1701.460 ;
        RECT 1400.770 1701.600 1401.090 1701.660 ;
        RECT 1424.780 1701.600 1424.920 1701.800 ;
        RECT 1462.410 1701.740 1462.730 1701.800 ;
        RECT 1521.380 1701.800 1594.200 1701.940 ;
        RECT 1400.770 1701.460 1424.920 1701.600 ;
        RECT 1463.330 1701.600 1463.650 1701.660 ;
        RECT 1521.380 1701.600 1521.520 1701.800 ;
        RECT 1594.060 1701.660 1594.200 1701.800 ;
        RECT 1594.430 1701.800 1655.930 1701.940 ;
        RECT 1594.430 1701.740 1594.750 1701.800 ;
        RECT 1655.610 1701.740 1655.930 1701.800 ;
        RECT 1463.330 1701.460 1521.520 1701.600 ;
        RECT 1400.770 1701.400 1401.090 1701.460 ;
        RECT 1463.330 1701.400 1463.650 1701.460 ;
        RECT 1593.970 1701.400 1594.290 1701.660 ;
        RECT 1751.840 1701.600 1751.980 1702.480 ;
        RECT 1835.100 1702.140 1848.580 1702.280 ;
        RECT 1787.170 1701.940 1787.490 1702.000 ;
        RECT 1786.800 1701.800 1787.490 1701.940 ;
        RECT 1786.800 1701.600 1786.940 1701.800 ;
        RECT 1787.170 1701.740 1787.490 1701.800 ;
        RECT 1811.090 1701.940 1811.410 1702.000 ;
        RECT 1835.100 1701.940 1835.240 1702.140 ;
        RECT 1811.090 1701.800 1835.240 1701.940 ;
        RECT 1848.440 1701.940 1848.580 1702.140 ;
        RECT 1908.610 1701.940 1908.930 1702.000 ;
        RECT 1848.440 1701.800 1908.930 1701.940 ;
        RECT 1811.090 1701.740 1811.410 1701.800 ;
        RECT 1908.610 1701.740 1908.930 1701.800 ;
        RECT 1751.840 1701.460 1786.940 1701.600 ;
        RECT 1655.610 1701.260 1655.930 1701.320 ;
        RECT 1666.190 1701.260 1666.510 1701.320 ;
        RECT 1655.610 1701.120 1666.510 1701.260 ;
        RECT 1655.610 1701.060 1655.930 1701.120 ;
        RECT 1666.190 1701.060 1666.510 1701.120 ;
        RECT 1787.170 1701.260 1787.490 1701.320 ;
        RECT 1811.090 1701.260 1811.410 1701.320 ;
        RECT 1787.170 1701.120 1811.410 1701.260 ;
        RECT 1787.170 1701.060 1787.490 1701.120 ;
        RECT 1811.090 1701.060 1811.410 1701.120 ;
        RECT 650.970 596.940 651.290 597.000 ;
        RECT 696.970 596.940 697.290 597.000 ;
        RECT 650.970 596.800 697.290 596.940 ;
        RECT 650.970 596.740 651.290 596.800 ;
        RECT 696.970 596.740 697.290 596.800 ;
        RECT 733.770 593.200 734.090 593.260 ;
        RECT 786.670 593.200 786.990 593.260 ;
        RECT 733.770 593.060 786.990 593.200 ;
        RECT 733.770 593.000 734.090 593.060 ;
        RECT 786.670 593.000 786.990 593.060 ;
        RECT 693.290 587.760 693.610 587.820 ;
        RECT 696.970 587.760 697.290 587.820 ;
        RECT 733.770 587.760 734.090 587.820 ;
        RECT 693.290 587.620 734.090 587.760 ;
        RECT 693.290 587.560 693.610 587.620 ;
        RECT 696.970 587.560 697.290 587.620 ;
        RECT 733.770 587.560 734.090 587.620 ;
        RECT 228.690 47.840 229.010 47.900 ;
        RECT 693.290 47.840 693.610 47.900 ;
        RECT 228.690 47.700 693.610 47.840 ;
        RECT 228.690 47.640 229.010 47.700 ;
        RECT 693.290 47.640 693.610 47.700 ;
      LAYER via ;
        RECT 490.000 2591.860 490.260 2592.120 ;
        RECT 638.120 2591.860 638.380 2592.120 ;
        RECT 641.340 2489.520 641.600 2489.780 ;
        RECT 1672.200 2489.520 1672.460 2489.780 ;
        RECT 638.120 2487.820 638.380 2488.080 ;
        RECT 641.340 2487.820 641.600 2488.080 ;
        RECT 628.000 1991.080 628.260 1991.340 ;
        RECT 641.340 1991.080 641.600 1991.340 ;
        RECT 690.100 1991.080 690.360 1991.340 ;
        RECT 651.000 1702.080 651.260 1702.340 ;
        RECT 690.100 1702.080 690.360 1702.340 ;
        RECT 772.900 1702.080 773.160 1702.340 ;
        RECT 869.500 1702.420 869.760 1702.680 ;
        RECT 786.700 1701.740 786.960 1702.000 ;
        RECT 917.340 1702.080 917.600 1702.340 ;
        RECT 1013.940 1702.080 1014.200 1702.340 ;
        RECT 1200.700 1702.420 1200.960 1702.680 ;
        RECT 1076.040 1702.080 1076.300 1702.340 ;
        RECT 1200.240 1702.080 1200.500 1702.340 ;
        RECT 1248.540 1702.080 1248.800 1702.340 ;
        RECT 1345.140 1702.420 1345.400 1702.680 ;
        RECT 1297.300 1702.080 1297.560 1702.340 ;
        RECT 1345.600 1702.080 1345.860 1702.340 ;
        RECT 1366.300 1702.080 1366.560 1702.340 ;
        RECT 1400.800 1702.420 1401.060 1702.680 ;
        RECT 1666.220 1702.080 1666.480 1702.340 ;
        RECT 966.100 1701.740 966.360 1702.000 ;
        RECT 1124.800 1701.740 1125.060 1702.000 ;
        RECT 1152.400 1701.740 1152.660 1702.000 ;
        RECT 869.960 1701.400 870.220 1701.660 ;
        RECT 917.340 1701.400 917.600 1701.660 ;
        RECT 1076.960 1701.400 1077.220 1701.660 ;
        RECT 1124.340 1701.400 1124.600 1701.660 ;
        RECT 1400.800 1701.400 1401.060 1701.660 ;
        RECT 1462.440 1701.740 1462.700 1702.000 ;
        RECT 1463.360 1701.400 1463.620 1701.660 ;
        RECT 1594.460 1701.740 1594.720 1702.000 ;
        RECT 1655.640 1701.740 1655.900 1702.000 ;
        RECT 1594.000 1701.400 1594.260 1701.660 ;
        RECT 1787.200 1701.740 1787.460 1702.000 ;
        RECT 1811.120 1701.740 1811.380 1702.000 ;
        RECT 1908.640 1701.740 1908.900 1702.000 ;
        RECT 1655.640 1701.060 1655.900 1701.320 ;
        RECT 1666.220 1701.060 1666.480 1701.320 ;
        RECT 1787.200 1701.060 1787.460 1701.320 ;
        RECT 1811.120 1701.060 1811.380 1701.320 ;
        RECT 651.000 596.740 651.260 597.000 ;
        RECT 697.000 596.740 697.260 597.000 ;
        RECT 733.800 593.000 734.060 593.260 ;
        RECT 786.700 593.000 786.960 593.260 ;
        RECT 693.320 587.560 693.580 587.820 ;
        RECT 697.000 587.560 697.260 587.820 ;
        RECT 733.800 587.560 734.060 587.820 ;
        RECT 228.720 47.640 228.980 47.900 ;
        RECT 693.320 47.640 693.580 47.900 ;
      LAYER met2 ;
        RECT 489.890 2600.660 490.170 2604.000 ;
        RECT 489.890 2600.000 490.200 2600.660 ;
        RECT 490.060 2592.150 490.200 2600.000 ;
        RECT 490.000 2591.830 490.260 2592.150 ;
        RECT 638.120 2591.830 638.380 2592.150 ;
        RECT 638.180 2488.110 638.320 2591.830 ;
        RECT 1672.130 2500.000 1672.410 2504.000 ;
        RECT 1672.260 2489.810 1672.400 2500.000 ;
        RECT 641.340 2489.490 641.600 2489.810 ;
        RECT 1672.200 2489.490 1672.460 2489.810 ;
        RECT 641.400 2488.110 641.540 2489.490 ;
        RECT 638.120 2487.790 638.380 2488.110 ;
        RECT 641.340 2487.790 641.600 2488.110 ;
        RECT 641.400 1991.370 641.540 2487.790 ;
        RECT 628.000 1991.050 628.260 1991.370 ;
        RECT 641.340 1991.050 641.600 1991.370 ;
        RECT 690.100 1991.050 690.360 1991.370 ;
        RECT 628.060 1981.750 628.200 1991.050 ;
        RECT 627.810 1981.110 628.200 1981.750 ;
        RECT 627.810 1977.750 628.090 1981.110 ;
        RECT 690.160 1702.370 690.300 1991.050 ;
        RECT 1908.630 1783.795 1908.910 1784.165 ;
        RECT 869.560 1702.990 870.160 1703.130 ;
        RECT 869.560 1702.710 869.700 1702.990 ;
        RECT 651.000 1702.050 651.260 1702.370 ;
        RECT 690.100 1702.050 690.360 1702.370 ;
        RECT 772.890 1702.195 773.170 1702.565 ;
        RECT 786.690 1702.195 786.970 1702.565 ;
        RECT 869.500 1702.390 869.760 1702.710 ;
        RECT 772.900 1702.050 773.160 1702.195 ;
        RECT 651.060 597.030 651.200 1702.050 ;
        RECT 786.760 1702.030 786.900 1702.195 ;
        RECT 786.700 1701.710 786.960 1702.030 ;
        RECT 870.020 1701.690 870.160 1702.990 ;
        RECT 1344.740 1702.990 1345.340 1703.130 ;
        RECT 1200.700 1702.565 1200.960 1702.710 ;
        RECT 1344.740 1702.565 1344.880 1702.990 ;
        RECT 1345.200 1702.710 1345.340 1702.990 ;
        RECT 917.340 1702.050 917.600 1702.370 ;
        RECT 1013.940 1702.050 1014.200 1702.370 ;
        RECT 1076.040 1702.050 1076.300 1702.370 ;
        RECT 1200.240 1702.050 1200.500 1702.370 ;
        RECT 1200.690 1702.195 1200.970 1702.565 ;
        RECT 1248.530 1702.195 1248.810 1702.565 ;
        RECT 1297.290 1702.195 1297.570 1702.565 ;
        RECT 1344.670 1702.195 1344.950 1702.565 ;
        RECT 1345.140 1702.390 1345.400 1702.710 ;
        RECT 1345.590 1702.195 1345.870 1702.565 ;
        RECT 1366.290 1702.195 1366.570 1702.565 ;
        RECT 1400.800 1702.390 1401.060 1702.710 ;
        RECT 1248.540 1702.050 1248.800 1702.195 ;
        RECT 1297.300 1702.050 1297.560 1702.195 ;
        RECT 1345.600 1702.050 1345.860 1702.195 ;
        RECT 1366.300 1702.050 1366.560 1702.195 ;
        RECT 917.400 1701.690 917.540 1702.050 ;
        RECT 966.100 1701.885 966.360 1702.030 ;
        RECT 1014.000 1701.885 1014.140 1702.050 ;
        RECT 869.960 1701.370 870.220 1701.690 ;
        RECT 917.340 1701.370 917.600 1701.690 ;
        RECT 966.090 1701.515 966.370 1701.885 ;
        RECT 1013.930 1701.515 1014.210 1701.885 ;
        RECT 1076.100 1701.770 1076.240 1702.050 ;
        RECT 1124.800 1701.770 1125.060 1702.030 ;
        RECT 1152.400 1701.885 1152.660 1702.030 ;
        RECT 1200.300 1701.885 1200.440 1702.050 ;
        RECT 1076.100 1701.690 1077.160 1701.770 ;
        RECT 1124.400 1701.710 1125.060 1701.770 ;
        RECT 1124.400 1701.690 1125.000 1701.710 ;
        RECT 1076.100 1701.630 1077.220 1701.690 ;
        RECT 1076.960 1701.370 1077.220 1701.630 ;
        RECT 1124.340 1701.630 1125.000 1701.690 ;
        RECT 1124.340 1701.370 1124.600 1701.630 ;
        RECT 1152.390 1701.515 1152.670 1701.885 ;
        RECT 1200.230 1701.515 1200.510 1701.885 ;
        RECT 1400.860 1701.690 1401.000 1702.390 ;
        RECT 1666.220 1702.050 1666.480 1702.370 ;
        RECT 1462.440 1701.770 1462.700 1702.030 ;
        RECT 1594.460 1701.770 1594.720 1702.030 ;
        RECT 1462.440 1701.710 1463.560 1701.770 ;
        RECT 1462.500 1701.690 1463.560 1701.710 ;
        RECT 1594.060 1701.710 1594.720 1701.770 ;
        RECT 1655.640 1701.710 1655.900 1702.030 ;
        RECT 1594.060 1701.690 1594.660 1701.710 ;
        RECT 1400.800 1701.370 1401.060 1701.690 ;
        RECT 1462.500 1701.630 1463.620 1701.690 ;
        RECT 1463.360 1701.370 1463.620 1701.630 ;
        RECT 1594.000 1701.630 1594.660 1701.690 ;
        RECT 1594.000 1701.370 1594.260 1701.630 ;
        RECT 1655.700 1701.350 1655.840 1701.710 ;
        RECT 1666.280 1701.350 1666.420 1702.050 ;
        RECT 1908.700 1702.030 1908.840 1783.795 ;
        RECT 1787.200 1701.710 1787.460 1702.030 ;
        RECT 1811.120 1701.710 1811.380 1702.030 ;
        RECT 1908.640 1701.710 1908.900 1702.030 ;
        RECT 1787.260 1701.350 1787.400 1701.710 ;
        RECT 1811.180 1701.350 1811.320 1701.710 ;
        RECT 1655.640 1701.030 1655.900 1701.350 ;
        RECT 1666.220 1701.030 1666.480 1701.350 ;
        RECT 1787.200 1701.030 1787.460 1701.350 ;
        RECT 1811.120 1701.030 1811.380 1701.350 ;
        RECT 787.390 600.170 787.670 604.000 ;
        RECT 786.760 600.030 787.670 600.170 ;
        RECT 651.000 596.710 651.260 597.030 ;
        RECT 697.000 596.710 697.260 597.030 ;
        RECT 697.060 587.850 697.200 596.710 ;
        RECT 786.760 593.290 786.900 600.030 ;
        RECT 787.390 600.000 787.670 600.030 ;
        RECT 733.800 592.970 734.060 593.290 ;
        RECT 786.700 592.970 786.960 593.290 ;
        RECT 733.860 587.850 734.000 592.970 ;
        RECT 693.320 587.530 693.580 587.850 ;
        RECT 697.000 587.530 697.260 587.850 ;
        RECT 733.800 587.530 734.060 587.850 ;
        RECT 693.380 47.930 693.520 587.530 ;
        RECT 228.720 47.610 228.980 47.930 ;
        RECT 693.320 47.610 693.580 47.930 ;
        RECT 228.780 2.400 228.920 47.610 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 1908.630 1783.840 1908.910 1784.120 ;
        RECT 772.890 1702.240 773.170 1702.520 ;
        RECT 786.690 1702.240 786.970 1702.520 ;
        RECT 1200.690 1702.240 1200.970 1702.520 ;
        RECT 1248.530 1702.240 1248.810 1702.520 ;
        RECT 1297.290 1702.240 1297.570 1702.520 ;
        RECT 1344.670 1702.240 1344.950 1702.520 ;
        RECT 1345.590 1702.240 1345.870 1702.520 ;
        RECT 1366.290 1702.240 1366.570 1702.520 ;
        RECT 966.090 1701.560 966.370 1701.840 ;
        RECT 1013.930 1701.560 1014.210 1701.840 ;
        RECT 1152.390 1701.560 1152.670 1701.840 ;
        RECT 1200.230 1701.560 1200.510 1701.840 ;
      LAYER met3 ;
        RECT 1920.000 1786.760 1924.000 1787.360 ;
        RECT 1908.605 1784.130 1908.935 1784.145 ;
        RECT 1920.350 1784.130 1920.650 1786.760 ;
        RECT 1908.605 1783.830 1920.650 1784.130 ;
        RECT 1908.605 1783.815 1908.935 1783.830 ;
        RECT 772.865 1702.530 773.195 1702.545 ;
        RECT 786.665 1702.530 786.995 1702.545 ;
        RECT 772.865 1702.230 786.995 1702.530 ;
        RECT 772.865 1702.215 773.195 1702.230 ;
        RECT 786.665 1702.215 786.995 1702.230 ;
        RECT 1200.665 1702.530 1200.995 1702.545 ;
        RECT 1248.505 1702.530 1248.835 1702.545 ;
        RECT 1200.665 1702.230 1248.835 1702.530 ;
        RECT 1200.665 1702.215 1200.995 1702.230 ;
        RECT 1248.505 1702.215 1248.835 1702.230 ;
        RECT 1297.265 1702.530 1297.595 1702.545 ;
        RECT 1344.645 1702.530 1344.975 1702.545 ;
        RECT 1297.265 1702.230 1344.975 1702.530 ;
        RECT 1297.265 1702.215 1297.595 1702.230 ;
        RECT 1344.645 1702.215 1344.975 1702.230 ;
        RECT 1345.565 1702.530 1345.895 1702.545 ;
        RECT 1366.265 1702.530 1366.595 1702.545 ;
        RECT 1345.565 1702.230 1366.595 1702.530 ;
        RECT 1345.565 1702.215 1345.895 1702.230 ;
        RECT 1366.265 1702.215 1366.595 1702.230 ;
        RECT 966.065 1701.850 966.395 1701.865 ;
        RECT 1013.905 1701.850 1014.235 1701.865 ;
        RECT 966.065 1701.550 1014.235 1701.850 ;
        RECT 966.065 1701.535 966.395 1701.550 ;
        RECT 1013.905 1701.535 1014.235 1701.550 ;
        RECT 1152.365 1701.850 1152.695 1701.865 ;
        RECT 1200.205 1701.850 1200.535 1701.865 ;
        RECT 1152.365 1701.550 1200.535 1701.850 ;
        RECT 1152.365 1701.535 1152.695 1701.550 ;
        RECT 1200.205 1701.535 1200.535 1701.550 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 690.530 497.120 690.850 497.380 ;
        RECT 690.620 496.700 690.760 497.120 ;
        RECT 690.530 496.440 690.850 496.700 ;
        RECT 690.530 355.540 690.850 355.600 ;
        RECT 691.450 355.540 691.770 355.600 ;
        RECT 690.530 355.400 691.770 355.540 ;
        RECT 690.530 355.340 690.850 355.400 ;
        RECT 691.450 355.340 691.770 355.400 ;
        RECT 690.530 331.400 690.850 331.460 ;
        RECT 691.450 331.400 691.770 331.460 ;
        RECT 690.530 331.260 691.770 331.400 ;
        RECT 690.530 331.200 690.850 331.260 ;
        RECT 691.450 331.200 691.770 331.260 ;
        RECT 690.530 159.360 690.850 159.420 ;
        RECT 691.450 159.360 691.770 159.420 ;
        RECT 690.530 159.220 691.770 159.360 ;
        RECT 690.530 159.160 690.850 159.220 ;
        RECT 691.450 159.160 691.770 159.220 ;
        RECT 690.530 131.480 690.850 131.540 ;
        RECT 691.450 131.480 691.770 131.540 ;
        RECT 690.530 131.340 691.770 131.480 ;
        RECT 690.530 131.280 690.850 131.340 ;
        RECT 691.450 131.280 691.770 131.340 ;
        RECT 690.070 34.580 690.390 34.640 ;
        RECT 690.990 34.580 691.310 34.640 ;
        RECT 690.070 34.440 691.310 34.580 ;
        RECT 690.070 34.380 690.390 34.440 ;
        RECT 690.990 34.380 691.310 34.440 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 690.070 17.580 690.390 17.640 ;
        RECT 50.210 17.440 690.390 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 690.070 17.380 690.390 17.440 ;
      LAYER via ;
        RECT 690.560 497.120 690.820 497.380 ;
        RECT 690.560 496.440 690.820 496.700 ;
        RECT 690.560 355.340 690.820 355.600 ;
        RECT 691.480 355.340 691.740 355.600 ;
        RECT 690.560 331.200 690.820 331.460 ;
        RECT 691.480 331.200 691.740 331.460 ;
        RECT 690.560 159.160 690.820 159.420 ;
        RECT 691.480 159.160 691.740 159.420 ;
        RECT 690.560 131.280 690.820 131.540 ;
        RECT 691.480 131.280 691.740 131.540 ;
        RECT 690.100 34.380 690.360 34.640 ;
        RECT 691.020 34.380 691.280 34.640 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 690.100 17.380 690.360 17.640 ;
      LAYER met2 ;
        RECT 695.850 600.170 696.130 604.000 ;
        RECT 693.380 600.030 696.130 600.170 ;
        RECT 693.380 588.440 693.520 600.030 ;
        RECT 695.850 600.000 696.130 600.030 ;
        RECT 690.620 588.300 693.520 588.440 ;
        RECT 690.620 497.410 690.760 588.300 ;
        RECT 690.560 497.090 690.820 497.410 ;
        RECT 690.560 496.410 690.820 496.730 ;
        RECT 690.620 355.630 690.760 496.410 ;
        RECT 690.560 355.310 690.820 355.630 ;
        RECT 691.480 355.310 691.740 355.630 ;
        RECT 691.540 331.490 691.680 355.310 ;
        RECT 690.560 331.170 690.820 331.490 ;
        RECT 691.480 331.170 691.740 331.490 ;
        RECT 690.620 159.450 690.760 331.170 ;
        RECT 690.560 159.130 690.820 159.450 ;
        RECT 691.480 159.130 691.740 159.450 ;
        RECT 691.540 131.570 691.680 159.130 ;
        RECT 690.560 131.250 690.820 131.570 ;
        RECT 691.480 131.250 691.740 131.570 ;
        RECT 690.620 74.530 690.760 131.250 ;
        RECT 690.620 74.390 691.220 74.530 ;
        RECT 691.080 34.670 691.220 74.390 ;
        RECT 690.100 34.350 690.360 34.670 ;
        RECT 691.020 34.350 691.280 34.670 ;
        RECT 690.160 17.670 690.300 34.350 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 690.100 17.350 690.360 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 795.410 545.260 795.730 545.320 ;
        RECT 795.040 545.120 795.730 545.260 ;
        RECT 795.040 544.980 795.180 545.120 ;
        RECT 795.410 545.060 795.730 545.120 ;
        RECT 794.950 544.720 795.270 544.980 ;
        RECT 795.410 283.260 795.730 283.520 ;
        RECT 795.500 283.120 795.640 283.260 ;
        RECT 795.870 283.120 796.190 283.180 ;
        RECT 795.500 282.980 796.190 283.120 ;
        RECT 795.870 282.920 796.190 282.980 ;
        RECT 795.410 241.440 795.730 241.700 ;
        RECT 795.500 241.300 795.640 241.440 ;
        RECT 795.870 241.300 796.190 241.360 ;
        RECT 795.500 241.160 796.190 241.300 ;
        RECT 795.870 241.100 796.190 241.160 ;
        RECT 794.950 234.840 795.270 234.900 ;
        RECT 795.870 234.840 796.190 234.900 ;
        RECT 794.950 234.700 796.190 234.840 ;
        RECT 794.950 234.640 795.270 234.700 ;
        RECT 795.870 234.640 796.190 234.700 ;
        RECT 793.570 186.220 793.890 186.280 ;
        RECT 794.950 186.220 795.270 186.280 ;
        RECT 793.570 186.080 795.270 186.220 ;
        RECT 793.570 186.020 793.890 186.080 ;
        RECT 794.950 186.020 795.270 186.080 ;
        RECT 793.570 138.280 793.890 138.340 ;
        RECT 794.950 138.280 795.270 138.340 ;
        RECT 793.570 138.140 795.270 138.280 ;
        RECT 793.570 138.080 793.890 138.140 ;
        RECT 794.950 138.080 795.270 138.140 ;
        RECT 793.570 89.320 793.890 89.380 ;
        RECT 794.950 89.320 795.270 89.380 ;
        RECT 793.570 89.180 795.270 89.320 ;
        RECT 793.570 89.120 793.890 89.180 ;
        RECT 794.950 89.120 795.270 89.180 ;
        RECT 252.610 32.880 252.930 32.940 ;
        RECT 793.570 32.880 793.890 32.940 ;
        RECT 252.610 32.740 793.890 32.880 ;
        RECT 252.610 32.680 252.930 32.740 ;
        RECT 793.570 32.680 793.890 32.740 ;
      LAYER via ;
        RECT 795.440 545.060 795.700 545.320 ;
        RECT 794.980 544.720 795.240 544.980 ;
        RECT 795.440 283.260 795.700 283.520 ;
        RECT 795.900 282.920 796.160 283.180 ;
        RECT 795.440 241.440 795.700 241.700 ;
        RECT 795.900 241.100 796.160 241.360 ;
        RECT 794.980 234.640 795.240 234.900 ;
        RECT 795.900 234.640 796.160 234.900 ;
        RECT 793.600 186.020 793.860 186.280 ;
        RECT 794.980 186.020 795.240 186.280 ;
        RECT 793.600 138.080 793.860 138.340 ;
        RECT 794.980 138.080 795.240 138.340 ;
        RECT 793.600 89.120 793.860 89.380 ;
        RECT 794.980 89.120 795.240 89.380 ;
        RECT 252.640 32.680 252.900 32.940 ;
        RECT 793.600 32.680 793.860 32.940 ;
      LAYER met2 ;
        RECT 799.810 600.850 800.090 604.000 ;
        RECT 797.340 600.710 800.090 600.850 ;
        RECT 797.340 596.770 797.480 600.710 ;
        RECT 799.810 600.000 800.090 600.710 ;
        RECT 795.500 596.630 797.480 596.770 ;
        RECT 795.500 545.350 795.640 596.630 ;
        RECT 795.440 545.030 795.700 545.350 ;
        RECT 794.980 544.690 795.240 545.010 ;
        RECT 795.040 434.930 795.180 544.690 ;
        RECT 795.040 434.790 795.640 434.930 ;
        RECT 795.500 400.930 795.640 434.790 ;
        RECT 795.500 400.790 796.100 400.930 ;
        RECT 795.960 400.250 796.100 400.790 ;
        RECT 795.040 400.110 796.100 400.250 ;
        RECT 795.040 362.170 795.180 400.110 ;
        RECT 795.040 362.030 795.640 362.170 ;
        RECT 795.500 283.550 795.640 362.030 ;
        RECT 795.440 283.230 795.700 283.550 ;
        RECT 795.900 282.890 796.160 283.210 ;
        RECT 795.960 282.610 796.100 282.890 ;
        RECT 795.500 282.470 796.100 282.610 ;
        RECT 795.500 241.730 795.640 282.470 ;
        RECT 795.440 241.410 795.700 241.730 ;
        RECT 795.900 241.070 796.160 241.390 ;
        RECT 795.960 234.930 796.100 241.070 ;
        RECT 794.980 234.610 795.240 234.930 ;
        RECT 795.900 234.610 796.160 234.930 ;
        RECT 795.040 186.310 795.180 234.610 ;
        RECT 793.600 185.990 793.860 186.310 ;
        RECT 794.980 185.990 795.240 186.310 ;
        RECT 793.660 138.370 793.800 185.990 ;
        RECT 793.600 138.050 793.860 138.370 ;
        RECT 794.980 138.050 795.240 138.370 ;
        RECT 795.040 89.410 795.180 138.050 ;
        RECT 793.600 89.090 793.860 89.410 ;
        RECT 794.980 89.090 795.240 89.410 ;
        RECT 793.660 32.970 793.800 89.090 ;
        RECT 252.640 32.650 252.900 32.970 ;
        RECT 793.600 32.650 793.860 32.970 ;
        RECT 252.700 2.400 252.840 32.650 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 33.220 270.410 33.280 ;
        RECT 807.370 33.220 807.690 33.280 ;
        RECT 270.090 33.080 807.690 33.220 ;
        RECT 270.090 33.020 270.410 33.080 ;
        RECT 807.370 33.020 807.690 33.080 ;
      LAYER via ;
        RECT 270.120 33.020 270.380 33.280 ;
        RECT 807.400 33.020 807.660 33.280 ;
      LAYER met2 ;
        RECT 809.010 600.170 809.290 604.000 ;
        RECT 807.460 600.030 809.290 600.170 ;
        RECT 807.460 33.310 807.600 600.030 ;
        RECT 809.010 600.000 809.290 600.030 ;
        RECT 270.120 32.990 270.380 33.310 ;
        RECT 807.400 32.990 807.660 33.310 ;
        RECT 270.180 2.400 270.320 32.990 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 814.730 497.120 815.050 497.380 ;
        RECT 814.820 496.700 814.960 497.120 ;
        RECT 814.730 496.440 815.050 496.700 ;
        RECT 814.730 355.540 815.050 355.600 ;
        RECT 815.650 355.540 815.970 355.600 ;
        RECT 814.730 355.400 815.970 355.540 ;
        RECT 814.730 355.340 815.050 355.400 ;
        RECT 815.650 355.340 815.970 355.400 ;
        RECT 814.730 331.400 815.050 331.460 ;
        RECT 815.650 331.400 815.970 331.460 ;
        RECT 814.730 331.260 815.970 331.400 ;
        RECT 814.730 331.200 815.050 331.260 ;
        RECT 815.650 331.200 815.970 331.260 ;
        RECT 814.730 282.780 815.050 282.840 ;
        RECT 815.650 282.780 815.970 282.840 ;
        RECT 814.730 282.640 815.970 282.780 ;
        RECT 814.730 282.580 815.050 282.640 ;
        RECT 815.650 282.580 815.970 282.640 ;
        RECT 814.730 234.840 815.050 234.900 ;
        RECT 815.650 234.840 815.970 234.900 ;
        RECT 814.730 234.700 815.970 234.840 ;
        RECT 814.730 234.640 815.050 234.700 ;
        RECT 815.650 234.640 815.970 234.700 ;
        RECT 814.730 96.800 815.050 96.860 ;
        RECT 814.730 96.660 815.420 96.800 ;
        RECT 814.730 96.600 815.050 96.660 ;
        RECT 815.280 96.520 815.420 96.660 ;
        RECT 815.190 96.260 815.510 96.520 ;
        RECT 815.190 90.000 815.510 90.060 ;
        RECT 815.650 90.000 815.970 90.060 ;
        RECT 815.190 89.860 815.970 90.000 ;
        RECT 815.190 89.800 815.510 89.860 ;
        RECT 815.650 89.800 815.970 89.860 ;
        RECT 814.270 48.520 814.590 48.580 ;
        RECT 815.650 48.520 815.970 48.580 ;
        RECT 814.270 48.380 815.970 48.520 ;
        RECT 814.270 48.320 814.590 48.380 ;
        RECT 815.650 48.320 815.970 48.380 ;
        RECT 288.030 33.560 288.350 33.620 ;
        RECT 814.270 33.560 814.590 33.620 ;
        RECT 288.030 33.420 814.590 33.560 ;
        RECT 288.030 33.360 288.350 33.420 ;
        RECT 814.270 33.360 814.590 33.420 ;
      LAYER via ;
        RECT 814.760 497.120 815.020 497.380 ;
        RECT 814.760 496.440 815.020 496.700 ;
        RECT 814.760 355.340 815.020 355.600 ;
        RECT 815.680 355.340 815.940 355.600 ;
        RECT 814.760 331.200 815.020 331.460 ;
        RECT 815.680 331.200 815.940 331.460 ;
        RECT 814.760 282.580 815.020 282.840 ;
        RECT 815.680 282.580 815.940 282.840 ;
        RECT 814.760 234.640 815.020 234.900 ;
        RECT 815.680 234.640 815.940 234.900 ;
        RECT 814.760 96.600 815.020 96.860 ;
        RECT 815.220 96.260 815.480 96.520 ;
        RECT 815.220 89.800 815.480 90.060 ;
        RECT 815.680 89.800 815.940 90.060 ;
        RECT 814.300 48.320 814.560 48.580 ;
        RECT 815.680 48.320 815.940 48.580 ;
        RECT 288.060 33.360 288.320 33.620 ;
        RECT 814.300 33.360 814.560 33.620 ;
      LAYER met2 ;
        RECT 818.210 600.850 818.490 604.000 ;
        RECT 815.740 600.710 818.490 600.850 ;
        RECT 815.740 596.770 815.880 600.710 ;
        RECT 818.210 600.000 818.490 600.710 ;
        RECT 814.820 596.630 815.880 596.770 ;
        RECT 814.820 497.410 814.960 596.630 ;
        RECT 814.760 497.090 815.020 497.410 ;
        RECT 814.760 496.410 815.020 496.730 ;
        RECT 814.820 355.630 814.960 496.410 ;
        RECT 814.760 355.310 815.020 355.630 ;
        RECT 815.680 355.310 815.940 355.630 ;
        RECT 815.740 331.490 815.880 355.310 ;
        RECT 814.760 331.170 815.020 331.490 ;
        RECT 815.680 331.170 815.940 331.490 ;
        RECT 814.820 282.870 814.960 331.170 ;
        RECT 814.760 282.550 815.020 282.870 ;
        RECT 815.680 282.550 815.940 282.870 ;
        RECT 815.740 234.930 815.880 282.550 ;
        RECT 814.760 234.610 815.020 234.930 ;
        RECT 815.680 234.610 815.940 234.930 ;
        RECT 814.820 96.890 814.960 234.610 ;
        RECT 814.760 96.570 815.020 96.890 ;
        RECT 815.220 96.230 815.480 96.550 ;
        RECT 815.280 90.090 815.420 96.230 ;
        RECT 815.220 89.770 815.480 90.090 ;
        RECT 815.680 89.770 815.940 90.090 ;
        RECT 815.740 48.610 815.880 89.770 ;
        RECT 814.300 48.290 814.560 48.610 ;
        RECT 815.680 48.290 815.940 48.610 ;
        RECT 814.360 33.650 814.500 48.290 ;
        RECT 288.060 33.330 288.320 33.650 ;
        RECT 814.300 33.330 814.560 33.650 ;
        RECT 288.120 2.400 288.260 33.330 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 822.550 410.620 822.870 410.680 ;
        RECT 822.550 410.480 823.240 410.620 ;
        RECT 822.550 410.420 822.870 410.480 ;
        RECT 823.100 410.340 823.240 410.480 ;
        RECT 823.010 410.080 823.330 410.340 ;
        RECT 822.550 324.260 822.870 324.320 ;
        RECT 823.930 324.260 824.250 324.320 ;
        RECT 822.550 324.120 824.250 324.260 ;
        RECT 822.550 324.060 822.870 324.120 ;
        RECT 823.930 324.060 824.250 324.120 ;
        RECT 823.010 234.840 823.330 234.900 ;
        RECT 823.930 234.840 824.250 234.900 ;
        RECT 823.010 234.700 824.250 234.840 ;
        RECT 823.010 234.640 823.330 234.700 ;
        RECT 823.930 234.640 824.250 234.700 ;
        RECT 305.970 33.900 306.290 33.960 ;
        RECT 822.550 33.900 822.870 33.960 ;
        RECT 305.970 33.760 822.870 33.900 ;
        RECT 305.970 33.700 306.290 33.760 ;
        RECT 822.550 33.700 822.870 33.760 ;
      LAYER via ;
        RECT 822.580 410.420 822.840 410.680 ;
        RECT 823.040 410.080 823.300 410.340 ;
        RECT 822.580 324.060 822.840 324.320 ;
        RECT 823.960 324.060 824.220 324.320 ;
        RECT 823.040 234.640 823.300 234.900 ;
        RECT 823.960 234.640 824.220 234.900 ;
        RECT 306.000 33.700 306.260 33.960 ;
        RECT 822.580 33.700 822.840 33.960 ;
      LAYER met2 ;
        RECT 827.410 600.850 827.690 604.000 ;
        RECT 824.940 600.710 827.690 600.850 ;
        RECT 824.940 596.770 825.080 600.710 ;
        RECT 827.410 600.000 827.690 600.710 ;
        RECT 823.100 596.630 825.080 596.770 ;
        RECT 823.100 569.400 823.240 596.630 ;
        RECT 822.640 569.260 823.240 569.400 ;
        RECT 822.640 410.710 822.780 569.260 ;
        RECT 822.580 410.390 822.840 410.710 ;
        RECT 823.040 410.050 823.300 410.370 ;
        RECT 823.100 386.650 823.240 410.050 ;
        RECT 822.640 386.510 823.240 386.650 ;
        RECT 822.640 385.970 822.780 386.510 ;
        RECT 822.640 385.830 823.240 385.970 ;
        RECT 823.100 331.570 823.240 385.830 ;
        RECT 822.640 331.430 823.240 331.570 ;
        RECT 822.640 324.350 822.780 331.430 ;
        RECT 822.580 324.030 822.840 324.350 ;
        RECT 823.960 324.030 824.220 324.350 ;
        RECT 824.020 234.930 824.160 324.030 ;
        RECT 823.040 234.610 823.300 234.930 ;
        RECT 823.960 234.610 824.220 234.930 ;
        RECT 823.100 146.045 823.240 234.610 ;
        RECT 823.030 145.675 823.310 146.045 ;
        RECT 822.570 144.995 822.850 145.365 ;
        RECT 822.640 144.740 822.780 144.995 ;
        RECT 822.640 144.600 823.240 144.740 ;
        RECT 823.100 120.770 823.240 144.600 ;
        RECT 822.640 120.630 823.240 120.770 ;
        RECT 822.640 33.990 822.780 120.630 ;
        RECT 306.000 33.670 306.260 33.990 ;
        RECT 822.580 33.670 822.840 33.990 ;
        RECT 306.060 2.400 306.200 33.670 ;
        RECT 305.850 -4.800 306.410 2.400 ;
      LAYER via2 ;
        RECT 823.030 145.720 823.310 146.000 ;
        RECT 822.570 145.040 822.850 145.320 ;
      LAYER met3 ;
        RECT 823.005 146.010 823.335 146.025 ;
        RECT 821.870 145.710 823.335 146.010 ;
        RECT 821.870 145.330 822.170 145.710 ;
        RECT 823.005 145.695 823.335 145.710 ;
        RECT 822.545 145.330 822.875 145.345 ;
        RECT 821.870 145.030 822.875 145.330 ;
        RECT 822.545 145.015 822.875 145.030 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 52.260 324.230 52.320 ;
        RECT 835.430 52.260 835.750 52.320 ;
        RECT 323.910 52.120 835.750 52.260 ;
        RECT 323.910 52.060 324.230 52.120 ;
        RECT 835.430 52.060 835.750 52.120 ;
      LAYER via ;
        RECT 323.940 52.060 324.200 52.320 ;
        RECT 835.460 52.060 835.720 52.320 ;
      LAYER met2 ;
        RECT 836.610 600.170 836.890 604.000 ;
        RECT 835.520 600.030 836.890 600.170 ;
        RECT 835.520 52.350 835.660 600.030 ;
        RECT 836.610 600.000 836.890 600.030 ;
        RECT 323.940 52.030 324.200 52.350 ;
        RECT 835.460 52.030 835.720 52.350 ;
        RECT 324.000 2.400 324.140 52.030 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 842.330 579.600 842.650 579.660 ;
        RECT 842.790 579.600 843.110 579.660 ;
        RECT 842.330 579.460 843.110 579.600 ;
        RECT 842.330 579.400 842.650 579.460 ;
        RECT 842.790 579.400 843.110 579.460 ;
        RECT 842.790 545.260 843.110 545.320 ;
        RECT 842.420 545.120 843.110 545.260 ;
        RECT 842.420 544.980 842.560 545.120 ;
        RECT 842.790 545.060 843.110 545.120 ;
        RECT 842.330 544.720 842.650 544.980 ;
        RECT 841.870 496.980 842.190 497.040 ;
        RECT 842.790 496.980 843.110 497.040 ;
        RECT 841.870 496.840 843.110 496.980 ;
        RECT 841.870 496.780 842.190 496.840 ;
        RECT 842.790 496.780 843.110 496.840 ;
        RECT 841.870 483.040 842.190 483.100 ;
        RECT 842.790 483.040 843.110 483.100 ;
        RECT 841.870 482.900 843.110 483.040 ;
        RECT 841.870 482.840 842.190 482.900 ;
        RECT 842.790 482.840 843.110 482.900 ;
        RECT 842.330 234.840 842.650 234.900 ;
        RECT 842.790 234.840 843.110 234.900 ;
        RECT 842.330 234.700 843.110 234.840 ;
        RECT 842.330 234.640 842.650 234.700 ;
        RECT 842.790 234.640 843.110 234.700 ;
        RECT 841.870 193.020 842.190 193.080 ;
        RECT 842.790 193.020 843.110 193.080 ;
        RECT 841.870 192.880 843.110 193.020 ;
        RECT 841.870 192.820 842.190 192.880 ;
        RECT 842.790 192.820 843.110 192.880 ;
        RECT 842.330 144.740 842.650 144.800 ;
        RECT 843.250 144.740 843.570 144.800 ;
        RECT 842.330 144.600 843.570 144.740 ;
        RECT 842.330 144.540 842.650 144.600 ;
        RECT 843.250 144.540 843.570 144.600 ;
        RECT 840.950 96.460 841.270 96.520 ;
        RECT 841.870 96.460 842.190 96.520 ;
        RECT 840.950 96.320 842.190 96.460 ;
        RECT 840.950 96.260 841.270 96.320 ;
        RECT 841.870 96.260 842.190 96.320 ;
        RECT 840.950 48.520 841.270 48.580 ;
        RECT 842.330 48.520 842.650 48.580 ;
        RECT 840.950 48.380 842.650 48.520 ;
        RECT 840.950 48.320 841.270 48.380 ;
        RECT 842.330 48.320 842.650 48.380 ;
        RECT 341.390 39.680 341.710 39.740 ;
        RECT 842.330 39.680 842.650 39.740 ;
        RECT 341.390 39.540 842.650 39.680 ;
        RECT 341.390 39.480 341.710 39.540 ;
        RECT 842.330 39.480 842.650 39.540 ;
      LAYER via ;
        RECT 842.360 579.400 842.620 579.660 ;
        RECT 842.820 579.400 843.080 579.660 ;
        RECT 842.820 545.060 843.080 545.320 ;
        RECT 842.360 544.720 842.620 544.980 ;
        RECT 841.900 496.780 842.160 497.040 ;
        RECT 842.820 496.780 843.080 497.040 ;
        RECT 841.900 482.840 842.160 483.100 ;
        RECT 842.820 482.840 843.080 483.100 ;
        RECT 842.360 234.640 842.620 234.900 ;
        RECT 842.820 234.640 843.080 234.900 ;
        RECT 841.900 192.820 842.160 193.080 ;
        RECT 842.820 192.820 843.080 193.080 ;
        RECT 842.360 144.540 842.620 144.800 ;
        RECT 843.280 144.540 843.540 144.800 ;
        RECT 840.980 96.260 841.240 96.520 ;
        RECT 841.900 96.260 842.160 96.520 ;
        RECT 840.980 48.320 841.240 48.580 ;
        RECT 842.360 48.320 842.620 48.580 ;
        RECT 341.420 39.480 341.680 39.740 ;
        RECT 842.360 39.480 842.620 39.740 ;
      LAYER met2 ;
        RECT 845.810 600.170 846.090 604.000 ;
        RECT 844.260 600.030 846.090 600.170 ;
        RECT 844.260 596.770 844.400 600.030 ;
        RECT 845.810 600.000 846.090 600.030 ;
        RECT 842.420 596.630 844.400 596.770 ;
        RECT 842.420 579.690 842.560 596.630 ;
        RECT 842.360 579.370 842.620 579.690 ;
        RECT 842.820 579.370 843.080 579.690 ;
        RECT 842.880 545.350 843.020 579.370 ;
        RECT 842.820 545.030 843.080 545.350 ;
        RECT 842.360 544.690 842.620 545.010 ;
        RECT 842.420 531.490 842.560 544.690 ;
        RECT 842.420 531.350 843.020 531.490 ;
        RECT 841.960 497.070 842.100 497.225 ;
        RECT 842.880 497.070 843.020 531.350 ;
        RECT 841.900 496.810 842.160 497.070 ;
        RECT 842.820 496.810 843.080 497.070 ;
        RECT 841.900 496.750 843.080 496.810 ;
        RECT 841.960 496.670 843.020 496.750 ;
        RECT 842.880 483.130 843.020 496.670 ;
        RECT 841.900 482.810 842.160 483.130 ;
        RECT 842.820 482.810 843.080 483.130 ;
        RECT 841.960 447.170 842.100 482.810 ;
        RECT 841.960 447.030 843.020 447.170 ;
        RECT 842.880 351.290 843.020 447.030 ;
        RECT 842.420 351.150 843.020 351.290 ;
        RECT 842.420 303.690 842.560 351.150 ;
        RECT 842.420 303.550 843.020 303.690 ;
        RECT 842.880 234.930 843.020 303.550 ;
        RECT 842.360 234.610 842.620 234.930 ;
        RECT 842.820 234.610 843.080 234.930 ;
        RECT 842.420 207.130 842.560 234.610 ;
        RECT 842.420 206.990 843.020 207.130 ;
        RECT 842.880 193.110 843.020 206.990 ;
        RECT 841.900 192.790 842.160 193.110 ;
        RECT 842.820 192.790 843.080 193.110 ;
        RECT 841.960 145.250 842.100 192.790 ;
        RECT 841.960 145.110 842.560 145.250 ;
        RECT 842.420 144.830 842.560 145.110 ;
        RECT 842.360 144.510 842.620 144.830 ;
        RECT 843.280 144.510 843.540 144.830 ;
        RECT 843.340 96.970 843.480 144.510 ;
        RECT 841.960 96.830 843.480 96.970 ;
        RECT 841.960 96.550 842.100 96.830 ;
        RECT 840.980 96.230 841.240 96.550 ;
        RECT 841.900 96.230 842.160 96.550 ;
        RECT 841.040 48.610 841.180 96.230 ;
        RECT 840.980 48.290 841.240 48.610 ;
        RECT 842.360 48.290 842.620 48.610 ;
        RECT 842.420 39.770 842.560 48.290 ;
        RECT 341.420 39.450 341.680 39.770 ;
        RECT 842.360 39.450 842.620 39.770 ;
        RECT 341.480 2.400 341.620 39.450 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 849.230 569.400 849.550 569.460 ;
        RECT 853.370 569.400 853.690 569.460 ;
        RECT 849.230 569.260 853.690 569.400 ;
        RECT 849.230 569.200 849.550 569.260 ;
        RECT 853.370 569.200 853.690 569.260 ;
        RECT 364.850 52.600 365.170 52.660 ;
        RECT 849.230 52.600 849.550 52.660 ;
        RECT 364.850 52.460 849.550 52.600 ;
        RECT 364.850 52.400 365.170 52.460 ;
        RECT 849.230 52.400 849.550 52.460 ;
        RECT 359.330 16.900 359.650 16.960 ;
        RECT 364.850 16.900 365.170 16.960 ;
        RECT 359.330 16.760 365.170 16.900 ;
        RECT 359.330 16.700 359.650 16.760 ;
        RECT 364.850 16.700 365.170 16.760 ;
      LAYER via ;
        RECT 849.260 569.200 849.520 569.460 ;
        RECT 853.400 569.200 853.660 569.460 ;
        RECT 364.880 52.400 365.140 52.660 ;
        RECT 849.260 52.400 849.520 52.660 ;
        RECT 359.360 16.700 359.620 16.960 ;
        RECT 364.880 16.700 365.140 16.960 ;
      LAYER met2 ;
        RECT 855.010 600.170 855.290 604.000 ;
        RECT 853.460 600.030 855.290 600.170 ;
        RECT 853.460 569.490 853.600 600.030 ;
        RECT 855.010 600.000 855.290 600.030 ;
        RECT 849.260 569.170 849.520 569.490 ;
        RECT 853.400 569.170 853.660 569.490 ;
        RECT 849.320 52.690 849.460 569.170 ;
        RECT 364.880 52.370 365.140 52.690 ;
        RECT 849.260 52.370 849.520 52.690 ;
        RECT 364.940 16.990 365.080 52.370 ;
        RECT 359.360 16.670 359.620 16.990 ;
        RECT 364.880 16.670 365.140 16.990 ;
        RECT 359.420 2.400 359.560 16.670 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 377.270 40.020 377.590 40.080 ;
        RECT 863.030 40.020 863.350 40.080 ;
        RECT 377.270 39.880 863.350 40.020 ;
        RECT 377.270 39.820 377.590 39.880 ;
        RECT 863.030 39.820 863.350 39.880 ;
      LAYER via ;
        RECT 377.300 39.820 377.560 40.080 ;
        RECT 863.060 39.820 863.320 40.080 ;
      LAYER met2 ;
        RECT 864.210 600.170 864.490 604.000 ;
        RECT 863.120 600.030 864.490 600.170 ;
        RECT 863.120 40.110 863.260 600.030 ;
        RECT 864.210 600.000 864.490 600.030 ;
        RECT 377.300 39.790 377.560 40.110 ;
        RECT 863.060 39.790 863.320 40.110 ;
        RECT 377.360 2.400 377.500 39.790 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 869.010 493.580 869.330 493.640 ;
        RECT 869.930 493.580 870.250 493.640 ;
        RECT 869.010 493.440 870.250 493.580 ;
        RECT 869.010 493.380 869.330 493.440 ;
        RECT 869.930 493.380 870.250 493.440 ;
        RECT 869.010 469.440 869.330 469.500 ;
        RECT 869.930 469.440 870.250 469.500 ;
        RECT 869.010 469.300 870.250 469.440 ;
        RECT 869.010 469.240 869.330 469.300 ;
        RECT 869.930 469.240 870.250 469.300 ;
        RECT 869.010 420.820 869.330 420.880 ;
        RECT 869.930 420.820 870.250 420.880 ;
        RECT 869.010 420.680 870.250 420.820 ;
        RECT 869.010 420.620 869.330 420.680 ;
        RECT 869.930 420.620 870.250 420.680 ;
        RECT 869.010 372.880 869.330 372.940 ;
        RECT 869.470 372.880 869.790 372.940 ;
        RECT 869.010 372.740 869.790 372.880 ;
        RECT 869.010 372.680 869.330 372.740 ;
        RECT 869.470 372.680 869.790 372.740 ;
        RECT 869.010 324.260 869.330 324.320 ;
        RECT 869.930 324.260 870.250 324.320 ;
        RECT 869.010 324.120 870.250 324.260 ;
        RECT 869.010 324.060 869.330 324.120 ;
        RECT 869.930 324.060 870.250 324.120 ;
        RECT 869.010 276.320 869.330 276.380 ;
        RECT 870.390 276.320 870.710 276.380 ;
        RECT 869.010 276.180 870.710 276.320 ;
        RECT 869.010 276.120 869.330 276.180 ;
        RECT 870.390 276.120 870.710 276.180 ;
        RECT 869.470 234.840 869.790 234.900 ;
        RECT 870.390 234.840 870.710 234.900 ;
        RECT 869.470 234.700 870.710 234.840 ;
        RECT 869.470 234.640 869.790 234.700 ;
        RECT 870.390 234.640 870.710 234.700 ;
        RECT 868.550 227.700 868.870 227.760 ;
        RECT 869.470 227.700 869.790 227.760 ;
        RECT 868.550 227.560 869.790 227.700 ;
        RECT 868.550 227.500 868.870 227.560 ;
        RECT 869.470 227.500 869.790 227.560 ;
        RECT 868.550 179.760 868.870 179.820 ;
        RECT 869.930 179.760 870.250 179.820 ;
        RECT 868.550 179.620 870.250 179.760 ;
        RECT 868.550 179.560 868.870 179.620 ;
        RECT 869.930 179.560 870.250 179.620 ;
        RECT 869.930 144.540 870.250 144.800 ;
        RECT 870.020 144.120 870.160 144.540 ;
        RECT 869.930 143.860 870.250 144.120 ;
        RECT 869.930 96.460 870.250 96.520 ;
        RECT 870.850 96.460 871.170 96.520 ;
        RECT 869.930 96.320 871.170 96.460 ;
        RECT 869.930 96.260 870.250 96.320 ;
        RECT 870.850 96.260 871.170 96.320 ;
        RECT 399.810 52.940 400.130 53.000 ;
        RECT 870.850 52.940 871.170 53.000 ;
        RECT 399.810 52.800 871.170 52.940 ;
        RECT 399.810 52.740 400.130 52.800 ;
        RECT 870.850 52.740 871.170 52.800 ;
        RECT 395.210 15.200 395.530 15.260 ;
        RECT 399.810 15.200 400.130 15.260 ;
        RECT 395.210 15.060 400.130 15.200 ;
        RECT 395.210 15.000 395.530 15.060 ;
        RECT 399.810 15.000 400.130 15.060 ;
      LAYER via ;
        RECT 869.040 493.380 869.300 493.640 ;
        RECT 869.960 493.380 870.220 493.640 ;
        RECT 869.040 469.240 869.300 469.500 ;
        RECT 869.960 469.240 870.220 469.500 ;
        RECT 869.040 420.620 869.300 420.880 ;
        RECT 869.960 420.620 870.220 420.880 ;
        RECT 869.040 372.680 869.300 372.940 ;
        RECT 869.500 372.680 869.760 372.940 ;
        RECT 869.040 324.060 869.300 324.320 ;
        RECT 869.960 324.060 870.220 324.320 ;
        RECT 869.040 276.120 869.300 276.380 ;
        RECT 870.420 276.120 870.680 276.380 ;
        RECT 869.500 234.640 869.760 234.900 ;
        RECT 870.420 234.640 870.680 234.900 ;
        RECT 868.580 227.500 868.840 227.760 ;
        RECT 869.500 227.500 869.760 227.760 ;
        RECT 868.580 179.560 868.840 179.820 ;
        RECT 869.960 179.560 870.220 179.820 ;
        RECT 869.960 144.540 870.220 144.800 ;
        RECT 869.960 143.860 870.220 144.120 ;
        RECT 869.960 96.260 870.220 96.520 ;
        RECT 870.880 96.260 871.140 96.520 ;
        RECT 399.840 52.740 400.100 53.000 ;
        RECT 870.880 52.740 871.140 53.000 ;
        RECT 395.240 15.000 395.500 15.260 ;
        RECT 399.840 15.000 400.100 15.260 ;
      LAYER met2 ;
        RECT 873.410 600.170 873.690 604.000 ;
        RECT 871.860 600.030 873.690 600.170 ;
        RECT 871.860 596.770 872.000 600.030 ;
        RECT 873.410 600.000 873.690 600.030 ;
        RECT 870.020 596.630 872.000 596.770 ;
        RECT 870.020 493.670 870.160 596.630 ;
        RECT 869.040 493.350 869.300 493.670 ;
        RECT 869.960 493.350 870.220 493.670 ;
        RECT 869.100 469.530 869.240 493.350 ;
        RECT 869.040 469.210 869.300 469.530 ;
        RECT 869.960 469.210 870.220 469.530 ;
        RECT 870.020 420.910 870.160 469.210 ;
        RECT 869.040 420.590 869.300 420.910 ;
        RECT 869.960 420.590 870.220 420.910 ;
        RECT 869.100 372.970 869.240 420.590 ;
        RECT 869.040 372.650 869.300 372.970 ;
        RECT 869.500 372.650 869.760 372.970 ;
        RECT 869.560 331.570 869.700 372.650 ;
        RECT 869.560 331.430 870.160 331.570 ;
        RECT 870.020 324.350 870.160 331.430 ;
        RECT 869.040 324.030 869.300 324.350 ;
        RECT 869.960 324.030 870.220 324.350 ;
        RECT 869.100 276.410 869.240 324.030 ;
        RECT 869.040 276.090 869.300 276.410 ;
        RECT 870.420 276.090 870.680 276.410 ;
        RECT 870.480 234.930 870.620 276.090 ;
        RECT 869.500 234.610 869.760 234.930 ;
        RECT 870.420 234.610 870.680 234.930 ;
        RECT 869.560 227.790 869.700 234.610 ;
        RECT 868.580 227.470 868.840 227.790 ;
        RECT 869.500 227.470 869.760 227.790 ;
        RECT 868.640 179.850 868.780 227.470 ;
        RECT 868.580 179.530 868.840 179.850 ;
        RECT 869.960 179.530 870.220 179.850 ;
        RECT 870.020 144.830 870.160 179.530 ;
        RECT 869.960 144.510 870.220 144.830 ;
        RECT 869.960 143.830 870.220 144.150 ;
        RECT 870.020 96.550 870.160 143.830 ;
        RECT 869.960 96.230 870.220 96.550 ;
        RECT 870.880 96.230 871.140 96.550 ;
        RECT 870.940 53.030 871.080 96.230 ;
        RECT 399.840 52.710 400.100 53.030 ;
        RECT 870.880 52.710 871.140 53.030 ;
        RECT 399.900 15.290 400.040 52.710 ;
        RECT 395.240 14.970 395.500 15.290 ;
        RECT 399.840 14.970 400.100 15.290 ;
        RECT 395.300 2.400 395.440 14.970 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 876.830 558.860 877.150 558.920 ;
        RECT 880.970 558.860 881.290 558.920 ;
        RECT 876.830 558.720 881.290 558.860 ;
        RECT 876.830 558.660 877.150 558.720 ;
        RECT 880.970 558.660 881.290 558.720 ;
        RECT 413.150 40.360 413.470 40.420 ;
        RECT 876.830 40.360 877.150 40.420 ;
        RECT 413.150 40.220 877.150 40.360 ;
        RECT 413.150 40.160 413.470 40.220 ;
        RECT 876.830 40.160 877.150 40.220 ;
      LAYER via ;
        RECT 876.860 558.660 877.120 558.920 ;
        RECT 881.000 558.660 881.260 558.920 ;
        RECT 413.180 40.160 413.440 40.420 ;
        RECT 876.860 40.160 877.120 40.420 ;
      LAYER met2 ;
        RECT 882.610 600.170 882.890 604.000 ;
        RECT 881.060 600.030 882.890 600.170 ;
        RECT 881.060 558.950 881.200 600.030 ;
        RECT 882.610 600.000 882.890 600.030 ;
        RECT 876.860 558.630 877.120 558.950 ;
        RECT 881.000 558.630 881.260 558.950 ;
        RECT 876.920 40.450 877.060 558.630 ;
        RECT 413.180 40.130 413.440 40.450 ;
        RECT 876.860 40.130 877.120 40.450 ;
        RECT 413.240 2.400 413.380 40.130 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 703.870 531.320 704.190 531.380 ;
        RECT 704.790 531.320 705.110 531.380 ;
        RECT 703.870 531.180 705.110 531.320 ;
        RECT 703.870 531.120 704.190 531.180 ;
        RECT 704.790 531.120 705.110 531.180 ;
        RECT 704.790 524.180 705.110 524.240 ;
        RECT 705.710 524.180 706.030 524.240 ;
        RECT 704.790 524.040 706.030 524.180 ;
        RECT 704.790 523.980 705.110 524.040 ;
        RECT 705.710 523.980 706.030 524.040 ;
        RECT 704.330 435.100 704.650 435.160 ;
        RECT 704.790 435.100 705.110 435.160 ;
        RECT 704.330 434.960 705.110 435.100 ;
        RECT 704.330 434.900 704.650 434.960 ;
        RECT 704.790 434.900 705.110 434.960 ;
        RECT 704.330 96.260 704.650 96.520 ;
        RECT 704.420 96.120 704.560 96.260 ;
        RECT 704.790 96.120 705.110 96.180 ;
        RECT 704.420 95.980 705.110 96.120 ;
        RECT 704.790 95.920 705.110 95.980 ;
        RECT 74.130 18.260 74.450 18.320 ;
        RECT 704.790 18.260 705.110 18.320 ;
        RECT 74.130 18.120 705.110 18.260 ;
        RECT 74.130 18.060 74.450 18.120 ;
        RECT 704.790 18.060 705.110 18.120 ;
      LAYER via ;
        RECT 703.900 531.120 704.160 531.380 ;
        RECT 704.820 531.120 705.080 531.380 ;
        RECT 704.820 523.980 705.080 524.240 ;
        RECT 705.740 523.980 706.000 524.240 ;
        RECT 704.360 434.900 704.620 435.160 ;
        RECT 704.820 434.900 705.080 435.160 ;
        RECT 704.360 96.260 704.620 96.520 ;
        RECT 704.820 95.920 705.080 96.180 ;
        RECT 74.160 18.060 74.420 18.320 ;
        RECT 704.820 18.060 705.080 18.320 ;
      LAYER met2 ;
        RECT 707.810 600.170 708.090 604.000 ;
        RECT 706.260 600.030 708.090 600.170 ;
        RECT 706.260 596.770 706.400 600.030 ;
        RECT 707.810 600.000 708.090 600.030 ;
        RECT 704.420 596.630 706.400 596.770 ;
        RECT 704.420 532.285 704.560 596.630 ;
        RECT 704.350 531.915 704.630 532.285 ;
        RECT 703.890 531.235 704.170 531.605 ;
        RECT 703.900 531.090 704.160 531.235 ;
        RECT 704.820 531.090 705.080 531.410 ;
        RECT 704.880 524.270 705.020 531.090 ;
        RECT 704.820 523.950 705.080 524.270 ;
        RECT 705.740 523.950 706.000 524.270 ;
        RECT 705.800 481.850 705.940 523.950 ;
        RECT 704.880 481.710 705.940 481.850 ;
        RECT 704.880 435.190 705.020 481.710 ;
        RECT 704.360 434.870 704.620 435.190 ;
        RECT 704.820 434.870 705.080 435.190 ;
        RECT 704.420 331.570 704.560 434.870 ;
        RECT 703.960 331.430 704.560 331.570 ;
        RECT 703.960 304.485 704.100 331.430 ;
        RECT 703.890 304.115 704.170 304.485 ;
        RECT 703.890 276.235 704.170 276.605 ;
        RECT 703.960 220.730 704.100 276.235 ;
        RECT 703.960 220.590 704.560 220.730 ;
        RECT 704.420 207.245 704.560 220.590 ;
        RECT 704.350 206.875 704.630 207.245 ;
        RECT 703.890 206.195 704.170 206.565 ;
        RECT 703.960 158.850 704.100 206.195 ;
        RECT 703.960 158.710 704.560 158.850 ;
        RECT 704.420 96.550 704.560 158.710 ;
        RECT 704.360 96.230 704.620 96.550 ;
        RECT 704.820 95.890 705.080 96.210 ;
        RECT 704.880 18.350 705.020 95.890 ;
        RECT 74.160 18.030 74.420 18.350 ;
        RECT 704.820 18.030 705.080 18.350 ;
        RECT 74.220 2.400 74.360 18.030 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 704.350 531.960 704.630 532.240 ;
        RECT 703.890 531.280 704.170 531.560 ;
        RECT 703.890 304.160 704.170 304.440 ;
        RECT 703.890 276.280 704.170 276.560 ;
        RECT 704.350 206.920 704.630 207.200 ;
        RECT 703.890 206.240 704.170 206.520 ;
      LAYER met3 ;
        RECT 704.325 532.250 704.655 532.265 ;
        RECT 704.110 531.935 704.655 532.250 ;
        RECT 704.110 531.585 704.410 531.935 ;
        RECT 703.865 531.270 704.410 531.585 ;
        RECT 703.865 531.255 704.195 531.270 ;
        RECT 703.865 304.460 704.195 304.465 ;
        RECT 703.865 304.450 704.450 304.460 ;
        RECT 703.865 304.150 704.650 304.450 ;
        RECT 703.865 304.140 704.450 304.150 ;
        RECT 703.865 304.135 704.195 304.140 ;
        RECT 703.865 276.580 704.195 276.585 ;
        RECT 703.865 276.570 704.450 276.580 ;
        RECT 703.865 276.270 704.650 276.570 ;
        RECT 703.865 276.260 704.450 276.270 ;
        RECT 703.865 276.255 704.195 276.260 ;
        RECT 704.325 207.210 704.655 207.225 ;
        RECT 704.110 206.895 704.655 207.210 ;
        RECT 704.110 206.545 704.410 206.895 ;
        RECT 703.865 206.230 704.410 206.545 ;
        RECT 703.865 206.215 704.195 206.230 ;
      LAYER via3 ;
        RECT 704.100 304.140 704.420 304.460 ;
        RECT 704.100 276.260 704.420 276.580 ;
      LAYER met4 ;
        RECT 704.095 304.135 704.425 304.465 ;
        RECT 704.110 276.585 704.410 304.135 ;
        RECT 704.095 276.255 704.425 276.585 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.310 53.280 434.630 53.340 ;
        RECT 890.630 53.280 890.950 53.340 ;
        RECT 434.310 53.140 890.950 53.280 ;
        RECT 434.310 53.080 434.630 53.140 ;
        RECT 890.630 53.080 890.950 53.140 ;
        RECT 430.630 16.900 430.950 16.960 ;
        RECT 434.310 16.900 434.630 16.960 ;
        RECT 430.630 16.760 434.630 16.900 ;
        RECT 430.630 16.700 430.950 16.760 ;
        RECT 434.310 16.700 434.630 16.760 ;
      LAYER via ;
        RECT 434.340 53.080 434.600 53.340 ;
        RECT 890.660 53.080 890.920 53.340 ;
        RECT 430.660 16.700 430.920 16.960 ;
        RECT 434.340 16.700 434.600 16.960 ;
      LAYER met2 ;
        RECT 891.810 600.170 892.090 604.000 ;
        RECT 890.720 600.030 892.090 600.170 ;
        RECT 890.720 53.370 890.860 600.030 ;
        RECT 891.810 600.000 892.090 600.030 ;
        RECT 434.340 53.050 434.600 53.370 ;
        RECT 890.660 53.050 890.920 53.370 ;
        RECT 434.400 16.990 434.540 53.050 ;
        RECT 430.660 16.670 430.920 16.990 ;
        RECT 434.340 16.670 434.600 16.990 ;
        RECT 430.720 2.400 430.860 16.670 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 897.990 572.800 898.310 572.860 ;
        RECT 899.830 572.800 900.150 572.860 ;
        RECT 897.990 572.660 900.150 572.800 ;
        RECT 897.990 572.600 898.310 572.660 ;
        RECT 899.830 572.600 900.150 572.660 ;
        RECT 897.990 545.400 898.310 545.660 ;
        RECT 898.080 544.980 898.220 545.400 ;
        RECT 897.990 544.720 898.310 544.980 ;
        RECT 897.990 517.380 898.310 517.440 ;
        RECT 898.450 517.380 898.770 517.440 ;
        RECT 897.990 517.240 898.770 517.380 ;
        RECT 897.990 517.180 898.310 517.240 ;
        RECT 898.450 517.180 898.770 517.240 ;
        RECT 897.990 496.980 898.310 497.040 ;
        RECT 897.990 496.840 898.680 496.980 ;
        RECT 897.990 496.780 898.310 496.840 ;
        RECT 898.540 496.700 898.680 496.840 ;
        RECT 898.450 496.440 898.770 496.700 ;
        RECT 897.990 338.340 898.310 338.600 ;
        RECT 898.080 337.520 898.220 338.340 ;
        RECT 898.450 337.520 898.770 337.580 ;
        RECT 898.080 337.380 898.770 337.520 ;
        RECT 898.450 337.320 898.770 337.380 ;
        RECT 897.530 282.780 897.850 282.840 ;
        RECT 897.990 282.780 898.310 282.840 ;
        RECT 897.530 282.640 898.310 282.780 ;
        RECT 897.530 282.580 897.850 282.640 ;
        RECT 897.990 282.580 898.310 282.640 ;
        RECT 897.530 234.840 897.850 234.900 ;
        RECT 898.450 234.840 898.770 234.900 ;
        RECT 897.530 234.700 898.770 234.840 ;
        RECT 897.530 234.640 897.850 234.700 ;
        RECT 898.450 234.640 898.770 234.700 ;
        RECT 897.070 227.700 897.390 227.760 ;
        RECT 898.450 227.700 898.770 227.760 ;
        RECT 897.070 227.560 898.770 227.700 ;
        RECT 897.070 227.500 897.390 227.560 ;
        RECT 898.450 227.500 898.770 227.560 ;
        RECT 897.070 179.760 897.390 179.820 ;
        RECT 897.990 179.760 898.310 179.820 ;
        RECT 897.070 179.620 898.310 179.760 ;
        RECT 897.070 179.560 897.390 179.620 ;
        RECT 897.990 179.560 898.310 179.620 ;
        RECT 897.990 144.740 898.310 144.800 ;
        RECT 898.450 144.740 898.770 144.800 ;
        RECT 897.990 144.600 898.770 144.740 ;
        RECT 897.990 144.540 898.310 144.600 ;
        RECT 898.450 144.540 898.770 144.600 ;
        RECT 448.570 40.700 448.890 40.760 ;
        RECT 897.990 40.700 898.310 40.760 ;
        RECT 448.570 40.560 898.310 40.700 ;
        RECT 448.570 40.500 448.890 40.560 ;
        RECT 897.990 40.500 898.310 40.560 ;
      LAYER via ;
        RECT 898.020 572.600 898.280 572.860 ;
        RECT 899.860 572.600 900.120 572.860 ;
        RECT 898.020 545.400 898.280 545.660 ;
        RECT 898.020 544.720 898.280 544.980 ;
        RECT 898.020 517.180 898.280 517.440 ;
        RECT 898.480 517.180 898.740 517.440 ;
        RECT 898.020 496.780 898.280 497.040 ;
        RECT 898.480 496.440 898.740 496.700 ;
        RECT 898.020 338.340 898.280 338.600 ;
        RECT 898.480 337.320 898.740 337.580 ;
        RECT 897.560 282.580 897.820 282.840 ;
        RECT 898.020 282.580 898.280 282.840 ;
        RECT 897.560 234.640 897.820 234.900 ;
        RECT 898.480 234.640 898.740 234.900 ;
        RECT 897.100 227.500 897.360 227.760 ;
        RECT 898.480 227.500 898.740 227.760 ;
        RECT 897.100 179.560 897.360 179.820 ;
        RECT 898.020 179.560 898.280 179.820 ;
        RECT 898.020 144.540 898.280 144.800 ;
        RECT 898.480 144.540 898.740 144.800 ;
        RECT 448.600 40.500 448.860 40.760 ;
        RECT 898.020 40.500 898.280 40.760 ;
      LAYER met2 ;
        RECT 901.010 600.170 901.290 604.000 ;
        RECT 899.920 600.030 901.290 600.170 ;
        RECT 899.920 572.890 900.060 600.030 ;
        RECT 901.010 600.000 901.290 600.030 ;
        RECT 898.020 572.570 898.280 572.890 ;
        RECT 899.860 572.570 900.120 572.890 ;
        RECT 898.080 545.690 898.220 572.570 ;
        RECT 898.020 545.370 898.280 545.690 ;
        RECT 898.020 544.690 898.280 545.010 ;
        RECT 898.080 524.690 898.220 544.690 ;
        RECT 898.080 524.550 898.680 524.690 ;
        RECT 898.540 517.470 898.680 524.550 ;
        RECT 898.020 517.150 898.280 517.470 ;
        RECT 898.480 517.150 898.740 517.470 ;
        RECT 898.080 497.070 898.220 517.150 ;
        RECT 898.020 496.750 898.280 497.070 ;
        RECT 898.480 496.410 898.740 496.730 ;
        RECT 898.540 386.650 898.680 496.410 ;
        RECT 898.080 386.510 898.680 386.650 ;
        RECT 898.080 338.630 898.220 386.510 ;
        RECT 898.020 338.310 898.280 338.630 ;
        RECT 898.480 337.290 898.740 337.610 ;
        RECT 898.540 303.690 898.680 337.290 ;
        RECT 898.080 303.550 898.680 303.690 ;
        RECT 898.080 282.870 898.220 303.550 ;
        RECT 897.560 282.550 897.820 282.870 ;
        RECT 898.020 282.550 898.280 282.870 ;
        RECT 897.620 234.930 897.760 282.550 ;
        RECT 897.560 234.610 897.820 234.930 ;
        RECT 898.480 234.610 898.740 234.930 ;
        RECT 898.540 227.790 898.680 234.610 ;
        RECT 897.100 227.470 897.360 227.790 ;
        RECT 898.480 227.470 898.740 227.790 ;
        RECT 897.160 179.850 897.300 227.470 ;
        RECT 897.100 179.530 897.360 179.850 ;
        RECT 898.020 179.530 898.280 179.850 ;
        RECT 898.080 144.830 898.220 179.530 ;
        RECT 898.020 144.510 898.280 144.830 ;
        RECT 898.480 144.510 898.740 144.830 ;
        RECT 898.540 110.060 898.680 144.510 ;
        RECT 898.080 109.920 898.680 110.060 ;
        RECT 898.080 40.790 898.220 109.920 ;
        RECT 448.600 40.470 448.860 40.790 ;
        RECT 898.020 40.470 898.280 40.790 ;
        RECT 448.660 2.400 448.800 40.470 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 904.890 483.040 905.210 483.100 ;
        RECT 905.810 483.040 906.130 483.100 ;
        RECT 904.890 482.900 906.130 483.040 ;
        RECT 904.890 482.840 905.210 482.900 ;
        RECT 905.810 482.840 906.130 482.900 ;
        RECT 904.890 448.360 905.210 448.420 ;
        RECT 905.810 448.360 906.130 448.420 ;
        RECT 904.890 448.220 906.130 448.360 ;
        RECT 904.890 448.160 905.210 448.220 ;
        RECT 905.810 448.160 906.130 448.220 ;
        RECT 905.350 338.340 905.670 338.600 ;
        RECT 905.440 337.520 905.580 338.340 ;
        RECT 905.810 337.520 906.130 337.580 ;
        RECT 905.440 337.380 906.130 337.520 ;
        RECT 905.810 337.320 906.130 337.380 ;
        RECT 905.350 289.580 905.670 289.640 ;
        RECT 905.810 289.580 906.130 289.640 ;
        RECT 905.350 289.440 906.130 289.580 ;
        RECT 905.350 289.380 905.670 289.440 ;
        RECT 905.810 289.380 906.130 289.440 ;
        RECT 904.890 282.780 905.210 282.840 ;
        RECT 905.350 282.780 905.670 282.840 ;
        RECT 904.890 282.640 905.670 282.780 ;
        RECT 904.890 282.580 905.210 282.640 ;
        RECT 905.350 282.580 905.670 282.640 ;
        RECT 904.890 234.840 905.210 234.900 ;
        RECT 905.810 234.840 906.130 234.900 ;
        RECT 904.890 234.700 906.130 234.840 ;
        RECT 904.890 234.640 905.210 234.700 ;
        RECT 905.810 234.640 906.130 234.700 ;
        RECT 903.510 137.940 903.830 138.000 ;
        RECT 905.810 137.940 906.130 138.000 ;
        RECT 903.510 137.800 906.130 137.940 ;
        RECT 903.510 137.740 903.830 137.800 ;
        RECT 905.810 137.740 906.130 137.800 ;
        RECT 903.510 90.000 903.830 90.060 ;
        RECT 905.350 90.000 905.670 90.060 ;
        RECT 903.510 89.860 905.670 90.000 ;
        RECT 903.510 89.800 903.830 89.860 ;
        RECT 905.350 89.800 905.670 89.860 ;
        RECT 466.510 16.900 466.830 16.960 ;
        RECT 871.310 16.900 871.630 16.960 ;
        RECT 466.510 16.760 871.630 16.900 ;
        RECT 466.510 16.700 466.830 16.760 ;
        RECT 871.310 16.700 871.630 16.760 ;
      LAYER via ;
        RECT 904.920 482.840 905.180 483.100 ;
        RECT 905.840 482.840 906.100 483.100 ;
        RECT 904.920 448.160 905.180 448.420 ;
        RECT 905.840 448.160 906.100 448.420 ;
        RECT 905.380 338.340 905.640 338.600 ;
        RECT 905.840 337.320 906.100 337.580 ;
        RECT 905.380 289.380 905.640 289.640 ;
        RECT 905.840 289.380 906.100 289.640 ;
        RECT 904.920 282.580 905.180 282.840 ;
        RECT 905.380 282.580 905.640 282.840 ;
        RECT 904.920 234.640 905.180 234.900 ;
        RECT 905.840 234.640 906.100 234.900 ;
        RECT 903.540 137.740 903.800 138.000 ;
        RECT 905.840 137.740 906.100 138.000 ;
        RECT 903.540 89.800 903.800 90.060 ;
        RECT 905.380 89.800 905.640 90.060 ;
        RECT 466.540 16.700 466.800 16.960 ;
        RECT 871.340 16.700 871.600 16.960 ;
      LAYER met2 ;
        RECT 910.210 600.850 910.490 604.000 ;
        RECT 907.740 600.710 910.490 600.850 ;
        RECT 907.740 596.770 907.880 600.710 ;
        RECT 910.210 600.000 910.490 600.710 ;
        RECT 905.900 596.630 907.880 596.770 ;
        RECT 905.900 569.400 906.040 596.630 ;
        RECT 905.440 569.260 906.040 569.400 ;
        RECT 905.440 545.090 905.580 569.260 ;
        RECT 905.440 544.950 906.040 545.090 ;
        RECT 905.900 483.130 906.040 544.950 ;
        RECT 904.920 482.810 905.180 483.130 ;
        RECT 905.840 482.810 906.100 483.130 ;
        RECT 904.980 448.450 905.120 482.810 ;
        RECT 904.920 448.130 905.180 448.450 ;
        RECT 905.840 448.130 906.100 448.450 ;
        RECT 905.900 409.770 906.040 448.130 ;
        RECT 905.440 409.630 906.040 409.770 ;
        RECT 905.440 338.630 905.580 409.630 ;
        RECT 905.380 338.310 905.640 338.630 ;
        RECT 905.840 337.290 906.100 337.610 ;
        RECT 905.900 289.670 906.040 337.290 ;
        RECT 905.380 289.350 905.640 289.670 ;
        RECT 905.840 289.350 906.100 289.670 ;
        RECT 905.440 282.870 905.580 289.350 ;
        RECT 904.920 282.550 905.180 282.870 ;
        RECT 905.380 282.550 905.640 282.870 ;
        RECT 904.980 234.930 905.120 282.550 ;
        RECT 904.920 234.610 905.180 234.930 ;
        RECT 905.840 234.610 906.100 234.930 ;
        RECT 905.900 207.810 906.040 234.610 ;
        RECT 905.900 207.670 906.500 207.810 ;
        RECT 906.360 179.930 906.500 207.670 ;
        RECT 905.900 179.790 906.500 179.930 ;
        RECT 905.900 138.030 906.040 179.790 ;
        RECT 903.540 137.710 903.800 138.030 ;
        RECT 905.840 137.710 906.100 138.030 ;
        RECT 903.600 90.090 903.740 137.710 ;
        RECT 903.540 89.770 903.800 90.090 ;
        RECT 905.380 89.770 905.640 90.090 ;
        RECT 905.440 48.125 905.580 89.770 ;
        RECT 871.330 47.755 871.610 48.125 ;
        RECT 905.370 47.755 905.650 48.125 ;
        RECT 871.400 16.990 871.540 47.755 ;
        RECT 466.540 16.670 466.800 16.990 ;
        RECT 871.340 16.670 871.600 16.990 ;
        RECT 466.600 2.400 466.740 16.670 ;
        RECT 466.390 -4.800 466.950 2.400 ;
      LAYER via2 ;
        RECT 871.330 47.800 871.610 48.080 ;
        RECT 905.370 47.800 905.650 48.080 ;
      LAYER met3 ;
        RECT 871.305 48.090 871.635 48.105 ;
        RECT 905.345 48.090 905.675 48.105 ;
        RECT 871.305 47.790 905.675 48.090 ;
        RECT 871.305 47.775 871.635 47.790 ;
        RECT 905.345 47.775 905.675 47.790 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 41.040 484.770 41.100 ;
        RECT 917.770 41.040 918.090 41.100 ;
        RECT 484.450 40.900 918.090 41.040 ;
        RECT 484.450 40.840 484.770 40.900 ;
        RECT 917.770 40.840 918.090 40.900 ;
      LAYER via ;
        RECT 484.480 40.840 484.740 41.100 ;
        RECT 917.800 40.840 918.060 41.100 ;
      LAYER met2 ;
        RECT 919.410 600.170 919.690 604.000 ;
        RECT 917.860 600.030 919.690 600.170 ;
        RECT 917.860 41.130 918.000 600.030 ;
        RECT 919.410 600.000 919.690 600.030 ;
        RECT 484.480 40.810 484.740 41.130 ;
        RECT 917.800 40.810 918.060 41.130 ;
        RECT 484.540 2.400 484.680 40.810 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 925.130 572.460 925.450 572.520 ;
        RECT 925.590 572.460 925.910 572.520 ;
        RECT 925.130 572.320 925.910 572.460 ;
        RECT 925.130 572.260 925.450 572.320 ;
        RECT 925.590 572.260 925.910 572.320 ;
        RECT 925.130 449.040 925.450 449.100 ;
        RECT 924.760 448.900 925.450 449.040 ;
        RECT 924.760 448.420 924.900 448.900 ;
        RECT 925.130 448.840 925.450 448.900 ;
        RECT 924.670 448.160 924.990 448.420 ;
        RECT 923.750 434.760 924.070 434.820 ;
        RECT 924.670 434.760 924.990 434.820 ;
        RECT 923.750 434.620 924.990 434.760 ;
        RECT 923.750 434.560 924.070 434.620 ;
        RECT 924.670 434.560 924.990 434.620 ;
        RECT 923.750 386.480 924.070 386.540 ;
        RECT 925.130 386.480 925.450 386.540 ;
        RECT 923.750 386.340 925.450 386.480 ;
        RECT 923.750 386.280 924.070 386.340 ;
        RECT 925.130 386.280 925.450 386.340 ;
        RECT 923.750 355.540 924.070 355.600 ;
        RECT 925.130 355.540 925.450 355.600 ;
        RECT 923.750 355.400 925.450 355.540 ;
        RECT 923.750 355.340 924.070 355.400 ;
        RECT 925.130 355.340 925.450 355.400 ;
        RECT 923.750 283.120 924.070 283.180 ;
        RECT 924.670 283.120 924.990 283.180 ;
        RECT 923.750 282.980 924.990 283.120 ;
        RECT 923.750 282.920 924.070 282.980 ;
        RECT 924.670 282.920 924.990 282.980 ;
        RECT 924.670 193.020 924.990 193.080 ;
        RECT 925.130 193.020 925.450 193.080 ;
        RECT 924.670 192.880 925.450 193.020 ;
        RECT 924.670 192.820 924.990 192.880 ;
        RECT 925.130 192.820 925.450 192.880 ;
        RECT 921.450 48.180 921.770 48.240 ;
        RECT 925.130 48.180 925.450 48.240 ;
        RECT 921.450 48.040 925.450 48.180 ;
        RECT 921.450 47.980 921.770 48.040 ;
        RECT 925.130 47.980 925.450 48.040 ;
        RECT 502.390 16.560 502.710 16.620 ;
        RECT 921.450 16.560 921.770 16.620 ;
        RECT 502.390 16.420 921.770 16.560 ;
        RECT 502.390 16.360 502.710 16.420 ;
        RECT 921.450 16.360 921.770 16.420 ;
      LAYER via ;
        RECT 925.160 572.260 925.420 572.520 ;
        RECT 925.620 572.260 925.880 572.520 ;
        RECT 925.160 448.840 925.420 449.100 ;
        RECT 924.700 448.160 924.960 448.420 ;
        RECT 923.780 434.560 924.040 434.820 ;
        RECT 924.700 434.560 924.960 434.820 ;
        RECT 923.780 386.280 924.040 386.540 ;
        RECT 925.160 386.280 925.420 386.540 ;
        RECT 923.780 355.340 924.040 355.600 ;
        RECT 925.160 355.340 925.420 355.600 ;
        RECT 923.780 282.920 924.040 283.180 ;
        RECT 924.700 282.920 924.960 283.180 ;
        RECT 924.700 192.820 924.960 193.080 ;
        RECT 925.160 192.820 925.420 193.080 ;
        RECT 921.480 47.980 921.740 48.240 ;
        RECT 925.160 47.980 925.420 48.240 ;
        RECT 502.420 16.360 502.680 16.620 ;
        RECT 921.480 16.360 921.740 16.620 ;
      LAYER met2 ;
        RECT 928.610 600.170 928.890 604.000 ;
        RECT 927.060 600.030 928.890 600.170 ;
        RECT 927.060 596.770 927.200 600.030 ;
        RECT 928.610 600.000 928.890 600.030 ;
        RECT 925.220 596.630 927.200 596.770 ;
        RECT 925.220 572.550 925.360 596.630 ;
        RECT 925.160 572.230 925.420 572.550 ;
        RECT 925.620 572.230 925.880 572.550 ;
        RECT 925.680 495.450 925.820 572.230 ;
        RECT 925.220 495.310 925.820 495.450 ;
        RECT 925.220 449.130 925.360 495.310 ;
        RECT 925.160 448.810 925.420 449.130 ;
        RECT 924.700 448.130 924.960 448.450 ;
        RECT 924.760 434.850 924.900 448.130 ;
        RECT 923.780 434.530 924.040 434.850 ;
        RECT 924.700 434.530 924.960 434.850 ;
        RECT 923.840 386.570 923.980 434.530 ;
        RECT 923.780 386.250 924.040 386.570 ;
        RECT 925.160 386.250 925.420 386.570 ;
        RECT 925.220 355.630 925.360 386.250 ;
        RECT 923.780 355.310 924.040 355.630 ;
        RECT 925.160 355.310 925.420 355.630 ;
        RECT 923.840 283.210 923.980 355.310 ;
        RECT 923.780 282.890 924.040 283.210 ;
        RECT 924.700 282.890 924.960 283.210 ;
        RECT 924.760 217.330 924.900 282.890 ;
        RECT 924.760 217.190 925.360 217.330 ;
        RECT 925.220 193.110 925.360 217.190 ;
        RECT 924.700 192.790 924.960 193.110 ;
        RECT 925.160 192.790 925.420 193.110 ;
        RECT 924.760 144.570 924.900 192.790 ;
        RECT 924.760 144.430 925.360 144.570 ;
        RECT 925.220 48.270 925.360 144.430 ;
        RECT 921.480 47.950 921.740 48.270 ;
        RECT 925.160 47.950 925.420 48.270 ;
        RECT 921.540 16.650 921.680 47.950 ;
        RECT 502.420 16.330 502.680 16.650 ;
        RECT 921.480 16.330 921.740 16.650 ;
        RECT 502.480 2.400 502.620 16.330 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 931.570 569.400 931.890 569.460 ;
        RECT 935.710 569.400 936.030 569.460 ;
        RECT 931.570 569.260 936.030 569.400 ;
        RECT 931.570 569.200 931.890 569.260 ;
        RECT 935.710 569.200 936.030 569.260 ;
        RECT 931.570 379.820 931.890 380.080 ;
        RECT 931.660 379.400 931.800 379.820 ;
        RECT 931.570 379.140 931.890 379.400 ;
        RECT 519.870 16.220 520.190 16.280 ;
        RECT 931.570 16.220 931.890 16.280 ;
        RECT 519.870 16.080 931.890 16.220 ;
        RECT 519.870 16.020 520.190 16.080 ;
        RECT 931.570 16.020 931.890 16.080 ;
      LAYER via ;
        RECT 931.600 569.200 931.860 569.460 ;
        RECT 935.740 569.200 936.000 569.460 ;
        RECT 931.600 379.820 931.860 380.080 ;
        RECT 931.600 379.140 931.860 379.400 ;
        RECT 519.900 16.020 520.160 16.280 ;
        RECT 931.600 16.020 931.860 16.280 ;
      LAYER met2 ;
        RECT 937.350 600.170 937.630 604.000 ;
        RECT 935.800 600.030 937.630 600.170 ;
        RECT 935.800 569.490 935.940 600.030 ;
        RECT 937.350 600.000 937.630 600.030 ;
        RECT 931.600 569.170 931.860 569.490 ;
        RECT 935.740 569.170 936.000 569.490 ;
        RECT 931.660 380.110 931.800 569.170 ;
        RECT 931.600 379.790 931.860 380.110 ;
        RECT 931.600 379.110 931.860 379.430 ;
        RECT 931.660 16.310 931.800 379.110 ;
        RECT 519.900 15.990 520.160 16.310 ;
        RECT 931.600 15.990 931.860 16.310 ;
        RECT 519.960 2.400 520.100 15.990 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 838.650 589.120 838.970 589.180 ;
        RECT 945.370 589.120 945.690 589.180 ;
        RECT 838.650 588.980 945.690 589.120 ;
        RECT 838.650 588.920 838.970 588.980 ;
        RECT 945.370 588.920 945.690 588.980 ;
        RECT 838.190 15.880 838.510 15.940 ;
        RECT 589.880 15.740 838.510 15.880 ;
        RECT 537.810 15.540 538.130 15.600 ;
        RECT 589.880 15.540 590.020 15.740 ;
        RECT 838.190 15.680 838.510 15.740 ;
        RECT 537.810 15.400 590.020 15.540 ;
        RECT 537.810 15.340 538.130 15.400 ;
      LAYER via ;
        RECT 838.680 588.920 838.940 589.180 ;
        RECT 945.400 588.920 945.660 589.180 ;
        RECT 537.840 15.340 538.100 15.600 ;
        RECT 838.220 15.680 838.480 15.940 ;
      LAYER met2 ;
        RECT 946.550 600.170 946.830 604.000 ;
        RECT 945.460 600.030 946.830 600.170 ;
        RECT 945.460 589.210 945.600 600.030 ;
        RECT 946.550 600.000 946.830 600.030 ;
        RECT 838.680 588.890 838.940 589.210 ;
        RECT 945.400 588.890 945.660 589.210 ;
        RECT 838.740 566.850 838.880 588.890 ;
        RECT 838.280 566.710 838.880 566.850 ;
        RECT 838.280 15.970 838.420 566.710 ;
        RECT 838.220 15.650 838.480 15.970 ;
        RECT 537.840 15.310 538.100 15.630 ;
        RECT 537.900 2.400 538.040 15.310 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 953.650 545.600 953.970 545.660 ;
        RECT 953.280 545.460 953.970 545.600 ;
        RECT 953.280 544.980 953.420 545.460 ;
        RECT 953.650 545.400 953.970 545.460 ;
        RECT 953.190 544.720 953.510 544.980 ;
        RECT 953.190 482.700 953.510 482.760 ;
        RECT 953.650 482.700 953.970 482.760 ;
        RECT 953.190 482.560 953.970 482.700 ;
        RECT 953.190 482.500 953.510 482.560 ;
        RECT 953.650 482.500 953.970 482.560 ;
        RECT 953.190 158.680 953.510 158.740 ;
        RECT 954.110 158.680 954.430 158.740 ;
        RECT 953.190 158.540 954.430 158.680 ;
        RECT 953.190 158.480 953.510 158.540 ;
        RECT 954.110 158.480 954.430 158.540 ;
        RECT 555.750 37.640 556.070 37.700 ;
        RECT 953.190 37.640 953.510 37.700 ;
        RECT 555.750 37.500 953.510 37.640 ;
        RECT 555.750 37.440 556.070 37.500 ;
        RECT 953.190 37.440 953.510 37.500 ;
      LAYER via ;
        RECT 953.680 545.400 953.940 545.660 ;
        RECT 953.220 544.720 953.480 544.980 ;
        RECT 953.220 482.500 953.480 482.760 ;
        RECT 953.680 482.500 953.940 482.760 ;
        RECT 953.220 158.480 953.480 158.740 ;
        RECT 954.140 158.480 954.400 158.740 ;
        RECT 555.780 37.440 556.040 37.700 ;
        RECT 953.220 37.440 953.480 37.700 ;
      LAYER met2 ;
        RECT 955.750 600.170 956.030 604.000 ;
        RECT 953.740 600.030 956.030 600.170 ;
        RECT 953.740 545.690 953.880 600.030 ;
        RECT 955.750 600.000 956.030 600.030 ;
        RECT 953.680 545.370 953.940 545.690 ;
        RECT 953.220 544.690 953.480 545.010 ;
        RECT 953.280 482.790 953.420 544.690 ;
        RECT 953.220 482.470 953.480 482.790 ;
        RECT 953.680 482.470 953.940 482.790 ;
        RECT 953.740 400.930 953.880 482.470 ;
        RECT 953.280 400.790 953.880 400.930 ;
        RECT 953.280 158.770 953.420 400.790 ;
        RECT 953.220 158.450 953.480 158.770 ;
        RECT 954.140 158.450 954.400 158.770 ;
        RECT 954.200 109.890 954.340 158.450 ;
        RECT 953.740 109.750 954.340 109.890 ;
        RECT 953.740 62.290 953.880 109.750 ;
        RECT 953.280 62.150 953.880 62.290 ;
        RECT 953.280 37.730 953.420 62.150 ;
        RECT 555.780 37.410 556.040 37.730 ;
        RECT 953.220 37.410 953.480 37.730 ;
        RECT 555.840 2.400 555.980 37.410 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 845.090 588.440 845.410 588.500 ;
        RECT 963.310 588.440 963.630 588.500 ;
        RECT 845.090 588.300 963.630 588.440 ;
        RECT 845.090 588.240 845.410 588.300 ;
        RECT 963.310 588.240 963.630 588.300 ;
        RECT 845.090 15.540 845.410 15.600 ;
        RECT 590.800 15.400 845.410 15.540 ;
        RECT 573.690 15.200 574.010 15.260 ;
        RECT 590.800 15.200 590.940 15.400 ;
        RECT 845.090 15.340 845.410 15.400 ;
        RECT 573.690 15.060 590.940 15.200 ;
        RECT 573.690 15.000 574.010 15.060 ;
      LAYER via ;
        RECT 845.120 588.240 845.380 588.500 ;
        RECT 963.340 588.240 963.600 588.500 ;
        RECT 573.720 15.000 573.980 15.260 ;
        RECT 845.120 15.340 845.380 15.600 ;
      LAYER met2 ;
        RECT 964.950 600.170 965.230 604.000 ;
        RECT 963.400 600.030 965.230 600.170 ;
        RECT 963.400 588.530 963.540 600.030 ;
        RECT 964.950 600.000 965.230 600.030 ;
        RECT 845.120 588.210 845.380 588.530 ;
        RECT 963.340 588.210 963.600 588.530 ;
        RECT 845.180 15.630 845.320 588.210 ;
        RECT 845.120 15.310 845.380 15.630 ;
        RECT 573.720 14.970 573.980 15.290 ;
        RECT 573.780 2.400 573.920 14.970 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 591.170 41.380 591.490 41.440 ;
        RECT 973.430 41.380 973.750 41.440 ;
        RECT 591.170 41.240 973.750 41.380 ;
        RECT 591.170 41.180 591.490 41.240 ;
        RECT 973.430 41.180 973.750 41.240 ;
      LAYER via ;
        RECT 591.200 41.180 591.460 41.440 ;
        RECT 973.460 41.180 973.720 41.440 ;
      LAYER met2 ;
        RECT 974.150 600.170 974.430 604.000 ;
        RECT 973.520 600.030 974.430 600.170 ;
        RECT 973.520 41.470 973.660 600.030 ;
        RECT 974.150 600.000 974.430 600.030 ;
        RECT 591.200 41.150 591.460 41.470 ;
        RECT 973.460 41.150 973.720 41.470 ;
        RECT 591.260 2.400 591.400 41.150 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 18.600 97.910 18.660 ;
        RECT 717.670 18.600 717.990 18.660 ;
        RECT 97.590 18.460 717.990 18.600 ;
        RECT 97.590 18.400 97.910 18.460 ;
        RECT 717.670 18.400 717.990 18.460 ;
      LAYER via ;
        RECT 97.620 18.400 97.880 18.660 ;
        RECT 717.700 18.400 717.960 18.660 ;
      LAYER met2 ;
        RECT 720.230 600.170 720.510 604.000 ;
        RECT 717.760 600.030 720.510 600.170 ;
        RECT 717.760 18.690 717.900 600.030 ;
        RECT 720.230 600.000 720.510 600.030 ;
        RECT 97.620 18.370 97.880 18.690 ;
        RECT 717.700 18.370 717.960 18.690 ;
        RECT 97.680 2.400 97.820 18.370 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 980.330 545.400 980.650 545.660 ;
        RECT 980.420 544.980 980.560 545.400 ;
        RECT 980.330 544.720 980.650 544.980 ;
        RECT 980.790 400.900 981.110 401.160 ;
        RECT 980.880 400.480 981.020 400.900 ;
        RECT 980.790 400.220 981.110 400.480 ;
        RECT 980.330 255.040 980.650 255.300 ;
        RECT 980.420 254.900 980.560 255.040 ;
        RECT 980.790 254.900 981.110 254.960 ;
        RECT 980.420 254.760 981.110 254.900 ;
        RECT 980.790 254.700 981.110 254.760 ;
        RECT 609.110 37.300 609.430 37.360 ;
        RECT 979.870 37.300 980.190 37.360 ;
        RECT 609.110 37.160 980.190 37.300 ;
        RECT 609.110 37.100 609.430 37.160 ;
        RECT 979.870 37.100 980.190 37.160 ;
      LAYER via ;
        RECT 980.360 545.400 980.620 545.660 ;
        RECT 980.360 544.720 980.620 544.980 ;
        RECT 980.820 400.900 981.080 401.160 ;
        RECT 980.820 400.220 981.080 400.480 ;
        RECT 980.360 255.040 980.620 255.300 ;
        RECT 980.820 254.700 981.080 254.960 ;
        RECT 609.140 37.100 609.400 37.360 ;
        RECT 979.900 37.100 980.160 37.360 ;
      LAYER met2 ;
        RECT 983.350 600.170 983.630 604.000 ;
        RECT 981.340 600.030 983.630 600.170 ;
        RECT 981.340 596.770 981.480 600.030 ;
        RECT 983.350 600.000 983.630 600.030 ;
        RECT 980.420 596.630 981.480 596.770 ;
        RECT 980.420 545.690 980.560 596.630 ;
        RECT 980.360 545.370 980.620 545.690 ;
        RECT 980.360 544.690 980.620 545.010 ;
        RECT 980.420 531.490 980.560 544.690 ;
        RECT 980.420 531.350 981.020 531.490 ;
        RECT 980.880 401.190 981.020 531.350 ;
        RECT 980.820 400.870 981.080 401.190 ;
        RECT 980.820 400.190 981.080 400.510 ;
        RECT 980.880 399.570 981.020 400.190 ;
        RECT 980.420 399.430 981.020 399.570 ;
        RECT 980.420 351.970 980.560 399.430 ;
        RECT 980.420 351.830 981.020 351.970 ;
        RECT 980.880 304.370 981.020 351.830 ;
        RECT 980.420 304.230 981.020 304.370 ;
        RECT 980.420 303.690 980.560 304.230 ;
        RECT 979.960 303.550 980.560 303.690 ;
        RECT 979.960 303.010 980.100 303.550 ;
        RECT 979.960 302.870 980.560 303.010 ;
        RECT 980.420 255.330 980.560 302.870 ;
        RECT 980.360 255.010 980.620 255.330 ;
        RECT 980.820 254.670 981.080 254.990 ;
        RECT 980.880 62.970 981.020 254.670 ;
        RECT 980.420 62.830 981.020 62.970 ;
        RECT 980.420 62.290 980.560 62.830 ;
        RECT 979.960 62.150 980.560 62.290 ;
        RECT 979.960 37.390 980.100 62.150 ;
        RECT 609.140 37.070 609.400 37.390 ;
        RECT 979.900 37.070 980.160 37.390 ;
        RECT 609.200 2.400 609.340 37.070 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 851.990 593.200 852.310 593.260 ;
        RECT 990.910 593.200 991.230 593.260 ;
        RECT 851.990 593.060 991.230 593.200 ;
        RECT 851.990 593.000 852.310 593.060 ;
        RECT 990.910 593.000 991.230 593.060 ;
        RECT 627.050 20.640 627.370 20.700 ;
        RECT 851.990 20.640 852.310 20.700 ;
        RECT 627.050 20.500 852.310 20.640 ;
        RECT 627.050 20.440 627.370 20.500 ;
        RECT 851.990 20.440 852.310 20.500 ;
      LAYER via ;
        RECT 852.020 593.000 852.280 593.260 ;
        RECT 990.940 593.000 991.200 593.260 ;
        RECT 627.080 20.440 627.340 20.700 ;
        RECT 852.020 20.440 852.280 20.700 ;
      LAYER met2 ;
        RECT 992.550 600.170 992.830 604.000 ;
        RECT 991.000 600.030 992.830 600.170 ;
        RECT 991.000 593.290 991.140 600.030 ;
        RECT 992.550 600.000 992.830 600.030 ;
        RECT 852.020 592.970 852.280 593.290 ;
        RECT 990.940 592.970 991.200 593.290 ;
        RECT 852.080 20.730 852.220 592.970 ;
        RECT 627.080 20.410 627.340 20.730 ;
        RECT 852.020 20.410 852.280 20.730 ;
        RECT 627.140 2.400 627.280 20.410 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 19.280 121.830 19.340 ;
        RECT 731.470 19.280 731.790 19.340 ;
        RECT 121.510 19.140 731.790 19.280 ;
        RECT 121.510 19.080 121.830 19.140 ;
        RECT 731.470 19.080 731.790 19.140 ;
      LAYER via ;
        RECT 121.540 19.080 121.800 19.340 ;
        RECT 731.500 19.080 731.760 19.340 ;
      LAYER met2 ;
        RECT 732.650 600.170 732.930 604.000 ;
        RECT 731.560 600.030 732.930 600.170 ;
        RECT 731.560 19.370 731.700 600.030 ;
        RECT 732.650 600.000 732.930 600.030 ;
        RECT 121.540 19.050 121.800 19.370 ;
        RECT 731.500 19.050 731.760 19.370 ;
        RECT 121.600 2.400 121.740 19.050 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 739.750 572.800 740.070 572.860 ;
        RECT 742.970 572.800 743.290 572.860 ;
        RECT 739.750 572.660 743.290 572.800 ;
        RECT 739.750 572.600 740.070 572.660 ;
        RECT 742.970 572.600 743.290 572.660 ;
        RECT 739.750 572.120 740.070 572.180 ;
        RECT 741.130 572.120 741.450 572.180 ;
        RECT 739.750 571.980 741.450 572.120 ;
        RECT 739.750 571.920 740.070 571.980 ;
        RECT 741.130 571.920 741.450 571.980 ;
        RECT 740.210 524.180 740.530 524.240 ;
        RECT 741.130 524.180 741.450 524.240 ;
        RECT 740.210 524.040 741.450 524.180 ;
        RECT 740.210 523.980 740.530 524.040 ;
        RECT 741.130 523.980 741.450 524.040 ;
        RECT 740.210 476.240 740.530 476.300 ;
        RECT 741.130 476.240 741.450 476.300 ;
        RECT 740.210 476.100 741.450 476.240 ;
        RECT 740.210 476.040 740.530 476.100 ;
        RECT 741.130 476.040 741.450 476.100 ;
        RECT 739.290 435.100 739.610 435.160 ;
        RECT 740.210 435.100 740.530 435.160 ;
        RECT 739.290 434.960 740.530 435.100 ;
        RECT 739.290 434.900 739.610 434.960 ;
        RECT 740.210 434.900 740.530 434.960 ;
        RECT 145.430 19.620 145.750 19.680 ;
        RECT 739.750 19.620 740.070 19.680 ;
        RECT 145.430 19.480 740.070 19.620 ;
        RECT 145.430 19.420 145.750 19.480 ;
        RECT 739.750 19.420 740.070 19.480 ;
      LAYER via ;
        RECT 739.780 572.600 740.040 572.860 ;
        RECT 743.000 572.600 743.260 572.860 ;
        RECT 739.780 571.920 740.040 572.180 ;
        RECT 741.160 571.920 741.420 572.180 ;
        RECT 740.240 523.980 740.500 524.240 ;
        RECT 741.160 523.980 741.420 524.240 ;
        RECT 740.240 476.040 740.500 476.300 ;
        RECT 741.160 476.040 741.420 476.300 ;
        RECT 739.320 434.900 739.580 435.160 ;
        RECT 740.240 434.900 740.500 435.160 ;
        RECT 145.460 19.420 145.720 19.680 ;
        RECT 739.780 19.420 740.040 19.680 ;
      LAYER met2 ;
        RECT 744.610 600.170 744.890 604.000 ;
        RECT 743.060 600.030 744.890 600.170 ;
        RECT 743.060 572.890 743.200 600.030 ;
        RECT 744.610 600.000 744.890 600.030 ;
        RECT 739.780 572.570 740.040 572.890 ;
        RECT 743.000 572.570 743.260 572.890 ;
        RECT 739.840 572.210 739.980 572.570 ;
        RECT 739.780 571.890 740.040 572.210 ;
        RECT 741.160 571.890 741.420 572.210 ;
        RECT 741.220 524.805 741.360 571.890 ;
        RECT 740.230 524.435 740.510 524.805 ;
        RECT 741.150 524.435 741.430 524.805 ;
        RECT 740.300 524.270 740.440 524.435 ;
        RECT 740.240 523.950 740.500 524.270 ;
        RECT 741.160 523.950 741.420 524.270 ;
        RECT 741.220 476.330 741.360 523.950 ;
        RECT 740.240 476.010 740.500 476.330 ;
        RECT 741.160 476.010 741.420 476.330 ;
        RECT 740.300 435.190 740.440 476.010 ;
        RECT 739.320 434.870 739.580 435.190 ;
        RECT 740.240 434.870 740.500 435.190 ;
        RECT 739.380 144.570 739.520 434.870 ;
        RECT 739.380 144.430 739.980 144.570 ;
        RECT 739.840 19.710 739.980 144.430 ;
        RECT 145.460 19.390 145.720 19.710 ;
        RECT 739.780 19.390 740.040 19.710 ;
        RECT 145.520 2.400 145.660 19.390 ;
        RECT 145.310 -4.800 145.870 2.400 ;
      LAYER via2 ;
        RECT 740.230 524.480 740.510 524.760 ;
        RECT 741.150 524.480 741.430 524.760 ;
      LAYER met3 ;
        RECT 740.205 524.770 740.535 524.785 ;
        RECT 741.125 524.770 741.455 524.785 ;
        RECT 740.205 524.470 741.455 524.770 ;
        RECT 740.205 524.455 740.535 524.470 ;
        RECT 741.125 524.455 741.455 524.470 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 31.180 163.690 31.240 ;
        RECT 420.970 31.180 421.290 31.240 ;
        RECT 163.370 31.040 421.290 31.180 ;
        RECT 163.370 30.980 163.690 31.040 ;
        RECT 420.970 30.980 421.290 31.040 ;
        RECT 517.110 31.180 517.430 31.240 ;
        RECT 565.870 31.180 566.190 31.240 ;
        RECT 517.110 31.040 566.190 31.180 ;
        RECT 517.110 30.980 517.430 31.040 ;
        RECT 565.870 30.980 566.190 31.040 ;
        RECT 613.710 31.180 614.030 31.240 ;
        RECT 641.770 31.180 642.090 31.240 ;
        RECT 613.710 31.040 642.090 31.180 ;
        RECT 613.710 30.980 614.030 31.040 ;
        RECT 641.770 30.980 642.090 31.040 ;
        RECT 676.730 30.840 677.050 30.900 ;
        RECT 751.710 30.840 752.030 30.900 ;
        RECT 676.730 30.700 752.030 30.840 ;
        RECT 676.730 30.640 677.050 30.700 ;
        RECT 751.710 30.640 752.030 30.700 ;
        RECT 420.970 30.160 421.290 30.220 ;
        RECT 517.110 30.160 517.430 30.220 ;
        RECT 420.970 30.020 517.430 30.160 ;
        RECT 420.970 29.960 421.290 30.020 ;
        RECT 517.110 29.960 517.430 30.020 ;
        RECT 565.870 28.120 566.190 28.180 ;
        RECT 613.710 28.120 614.030 28.180 ;
        RECT 565.870 27.980 614.030 28.120 ;
        RECT 565.870 27.920 566.190 27.980 ;
        RECT 613.710 27.920 614.030 27.980 ;
        RECT 641.770 27.780 642.090 27.840 ;
        RECT 676.730 27.780 677.050 27.840 ;
        RECT 641.770 27.640 677.050 27.780 ;
        RECT 641.770 27.580 642.090 27.640 ;
        RECT 676.730 27.580 677.050 27.640 ;
      LAYER via ;
        RECT 163.400 30.980 163.660 31.240 ;
        RECT 421.000 30.980 421.260 31.240 ;
        RECT 517.140 30.980 517.400 31.240 ;
        RECT 565.900 30.980 566.160 31.240 ;
        RECT 613.740 30.980 614.000 31.240 ;
        RECT 641.800 30.980 642.060 31.240 ;
        RECT 676.760 30.640 677.020 30.900 ;
        RECT 751.740 30.640 752.000 30.900 ;
        RECT 421.000 29.960 421.260 30.220 ;
        RECT 517.140 29.960 517.400 30.220 ;
        RECT 565.900 27.920 566.160 28.180 ;
        RECT 613.740 27.920 614.000 28.180 ;
        RECT 641.800 27.580 642.060 27.840 ;
        RECT 676.760 27.580 677.020 27.840 ;
      LAYER met2 ;
        RECT 753.810 600.170 754.090 604.000 ;
        RECT 752.260 600.030 754.090 600.170 ;
        RECT 752.260 31.690 752.400 600.030 ;
        RECT 753.810 600.000 754.090 600.030 ;
        RECT 751.800 31.550 752.400 31.690 ;
        RECT 163.400 30.950 163.660 31.270 ;
        RECT 421.000 30.950 421.260 31.270 ;
        RECT 517.140 30.950 517.400 31.270 ;
        RECT 565.900 30.950 566.160 31.270 ;
        RECT 613.740 30.950 614.000 31.270 ;
        RECT 641.800 30.950 642.060 31.270 ;
        RECT 163.460 2.400 163.600 30.950 ;
        RECT 421.060 30.250 421.200 30.950 ;
        RECT 517.200 30.250 517.340 30.950 ;
        RECT 421.000 29.930 421.260 30.250 ;
        RECT 517.140 29.930 517.400 30.250 ;
        RECT 565.960 28.210 566.100 30.950 ;
        RECT 613.800 28.210 613.940 30.950 ;
        RECT 565.900 27.890 566.160 28.210 ;
        RECT 613.740 27.890 614.000 28.210 ;
        RECT 641.860 27.870 642.000 30.950 ;
        RECT 751.800 30.930 751.940 31.550 ;
        RECT 676.760 30.610 677.020 30.930 ;
        RECT 751.740 30.610 752.000 30.930 ;
        RECT 676.820 27.870 676.960 30.610 ;
        RECT 641.800 27.550 642.060 27.870 ;
        RECT 676.760 27.550 677.020 27.870 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 760.450 524.180 760.770 524.240 ;
        RECT 760.910 524.180 761.230 524.240 ;
        RECT 760.450 524.040 761.230 524.180 ;
        RECT 760.450 523.980 760.770 524.040 ;
        RECT 760.910 523.980 761.230 524.040 ;
        RECT 759.070 476.240 759.390 476.300 ;
        RECT 760.450 476.240 760.770 476.300 ;
        RECT 759.070 476.100 760.770 476.240 ;
        RECT 759.070 476.040 759.390 476.100 ;
        RECT 760.450 476.040 760.770 476.100 ;
        RECT 759.070 434.760 759.390 434.820 ;
        RECT 759.530 434.760 759.850 434.820 ;
        RECT 759.070 434.620 759.850 434.760 ;
        RECT 759.070 434.560 759.390 434.620 ;
        RECT 759.530 434.560 759.850 434.620 ;
        RECT 759.070 144.740 759.390 144.800 ;
        RECT 759.530 144.740 759.850 144.800 ;
        RECT 759.070 144.600 759.850 144.740 ;
        RECT 759.070 144.540 759.390 144.600 ;
        RECT 759.530 144.540 759.850 144.600 ;
        RECT 180.850 19.960 181.170 20.020 ;
        RECT 759.530 19.960 759.850 20.020 ;
        RECT 180.850 19.820 759.850 19.960 ;
        RECT 180.850 19.760 181.170 19.820 ;
        RECT 759.530 19.760 759.850 19.820 ;
      LAYER via ;
        RECT 760.480 523.980 760.740 524.240 ;
        RECT 760.940 523.980 761.200 524.240 ;
        RECT 759.100 476.040 759.360 476.300 ;
        RECT 760.480 476.040 760.740 476.300 ;
        RECT 759.100 434.560 759.360 434.820 ;
        RECT 759.560 434.560 759.820 434.820 ;
        RECT 759.100 144.540 759.360 144.800 ;
        RECT 759.560 144.540 759.820 144.800 ;
        RECT 180.880 19.760 181.140 20.020 ;
        RECT 759.560 19.760 759.820 20.020 ;
      LAYER met2 ;
        RECT 763.010 600.170 763.290 604.000 ;
        RECT 762.380 600.030 763.290 600.170 ;
        RECT 762.380 579.885 762.520 600.030 ;
        RECT 763.010 600.000 763.290 600.030 ;
        RECT 760.930 579.515 761.210 579.885 ;
        RECT 762.310 579.515 762.590 579.885 ;
        RECT 761.000 524.270 761.140 579.515 ;
        RECT 760.480 523.950 760.740 524.270 ;
        RECT 760.940 523.950 761.200 524.270 ;
        RECT 760.540 476.330 760.680 523.950 ;
        RECT 759.100 476.010 759.360 476.330 ;
        RECT 760.480 476.010 760.740 476.330 ;
        RECT 759.160 434.930 759.300 476.010 ;
        RECT 759.160 434.850 759.760 434.930 ;
        RECT 759.100 434.790 759.820 434.850 ;
        RECT 759.100 434.530 759.360 434.790 ;
        RECT 759.560 434.530 759.820 434.790 ;
        RECT 759.160 144.830 759.300 434.530 ;
        RECT 759.100 144.510 759.360 144.830 ;
        RECT 759.560 144.510 759.820 144.830 ;
        RECT 759.620 20.050 759.760 144.510 ;
        RECT 180.880 19.730 181.140 20.050 ;
        RECT 759.560 19.730 759.820 20.050 ;
        RECT 180.940 2.400 181.080 19.730 ;
        RECT 180.730 -4.800 181.290 2.400 ;
      LAYER via2 ;
        RECT 760.930 579.560 761.210 579.840 ;
        RECT 762.310 579.560 762.590 579.840 ;
      LAYER met3 ;
        RECT 760.905 579.850 761.235 579.865 ;
        RECT 762.285 579.850 762.615 579.865 ;
        RECT 760.905 579.550 762.615 579.850 ;
        RECT 760.905 579.535 761.235 579.550 ;
        RECT 762.285 579.535 762.615 579.550 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 766.430 549.000 766.750 549.060 ;
        RECT 770.570 549.000 770.890 549.060 ;
        RECT 766.430 548.860 770.890 549.000 ;
        RECT 766.430 548.800 766.750 548.860 ;
        RECT 770.570 548.800 770.890 548.860 ;
        RECT 198.790 31.860 199.110 31.920 ;
        RECT 766.430 31.860 766.750 31.920 ;
        RECT 198.790 31.720 766.750 31.860 ;
        RECT 198.790 31.660 199.110 31.720 ;
        RECT 766.430 31.660 766.750 31.720 ;
      LAYER via ;
        RECT 766.460 548.800 766.720 549.060 ;
        RECT 770.600 548.800 770.860 549.060 ;
        RECT 198.820 31.660 199.080 31.920 ;
        RECT 766.460 31.660 766.720 31.920 ;
      LAYER met2 ;
        RECT 772.210 600.170 772.490 604.000 ;
        RECT 770.660 600.030 772.490 600.170 ;
        RECT 770.660 549.090 770.800 600.030 ;
        RECT 772.210 600.000 772.490 600.030 ;
        RECT 766.460 548.770 766.720 549.090 ;
        RECT 770.600 548.770 770.860 549.090 ;
        RECT 766.520 31.950 766.660 548.770 ;
        RECT 198.820 31.630 199.080 31.950 ;
        RECT 766.460 31.630 766.720 31.950 ;
        RECT 198.880 2.400 199.020 31.630 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 20.300 217.050 20.360 ;
        RECT 779.770 20.300 780.090 20.360 ;
        RECT 216.730 20.160 780.090 20.300 ;
        RECT 216.730 20.100 217.050 20.160 ;
        RECT 779.770 20.100 780.090 20.160 ;
      LAYER via ;
        RECT 216.760 20.100 217.020 20.360 ;
        RECT 779.800 20.100 780.060 20.360 ;
      LAYER met2 ;
        RECT 781.410 600.170 781.690 604.000 ;
        RECT 779.860 600.030 781.690 600.170 ;
        RECT 779.860 20.390 780.000 600.030 ;
        RECT 781.410 600.000 781.690 600.030 ;
        RECT 216.760 20.070 217.020 20.390 ;
        RECT 779.800 20.070 780.060 20.390 ;
        RECT 216.820 2.400 216.960 20.070 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 787.130 572.800 787.450 572.860 ;
        RECT 788.970 572.800 789.290 572.860 ;
        RECT 787.130 572.660 789.290 572.800 ;
        RECT 787.130 572.600 787.450 572.660 ;
        RECT 788.970 572.600 789.290 572.660 ;
        RECT 786.670 193.360 786.990 193.420 ;
        RECT 787.130 193.360 787.450 193.420 ;
        RECT 786.670 193.220 787.450 193.360 ;
        RECT 786.670 193.160 786.990 193.220 ;
        RECT 787.130 193.160 787.450 193.220 ;
        RECT 786.670 144.740 786.990 144.800 ;
        RECT 787.130 144.740 787.450 144.800 ;
        RECT 786.670 144.600 787.450 144.740 ;
        RECT 786.670 144.540 786.990 144.600 ;
        RECT 787.130 144.540 787.450 144.600 ;
        RECT 786.670 96.800 786.990 96.860 ;
        RECT 787.130 96.800 787.450 96.860 ;
        RECT 786.670 96.660 787.450 96.800 ;
        RECT 786.670 96.600 786.990 96.660 ;
        RECT 787.130 96.600 787.450 96.660 ;
        RECT 234.670 32.540 234.990 32.600 ;
        RECT 786.670 32.540 786.990 32.600 ;
        RECT 234.670 32.400 786.990 32.540 ;
        RECT 234.670 32.340 234.990 32.400 ;
        RECT 786.670 32.340 786.990 32.400 ;
      LAYER via ;
        RECT 787.160 572.600 787.420 572.860 ;
        RECT 789.000 572.600 789.260 572.860 ;
        RECT 786.700 193.160 786.960 193.420 ;
        RECT 787.160 193.160 787.420 193.420 ;
        RECT 786.700 144.540 786.960 144.800 ;
        RECT 787.160 144.540 787.420 144.800 ;
        RECT 786.700 96.600 786.960 96.860 ;
        RECT 787.160 96.600 787.420 96.860 ;
        RECT 234.700 32.340 234.960 32.600 ;
        RECT 786.700 32.340 786.960 32.600 ;
      LAYER met2 ;
        RECT 790.610 600.170 790.890 604.000 ;
        RECT 789.060 600.030 790.890 600.170 ;
        RECT 789.060 572.890 789.200 600.030 ;
        RECT 790.610 600.000 790.890 600.030 ;
        RECT 787.160 572.570 787.420 572.890 ;
        RECT 789.000 572.570 789.260 572.890 ;
        RECT 787.220 265.610 787.360 572.570 ;
        RECT 786.760 265.470 787.360 265.610 ;
        RECT 786.760 193.450 786.900 265.470 ;
        RECT 786.700 193.130 786.960 193.450 ;
        RECT 787.160 193.130 787.420 193.450 ;
        RECT 787.220 144.830 787.360 193.130 ;
        RECT 786.700 144.510 786.960 144.830 ;
        RECT 787.160 144.510 787.420 144.830 ;
        RECT 786.760 96.890 786.900 144.510 ;
        RECT 786.700 96.570 786.960 96.890 ;
        RECT 787.160 96.570 787.420 96.890 ;
        RECT 787.220 62.970 787.360 96.570 ;
        RECT 787.220 62.830 787.820 62.970 ;
        RECT 787.680 61.610 787.820 62.830 ;
        RECT 786.760 61.470 787.820 61.610 ;
        RECT 786.760 32.630 786.900 61.470 ;
        RECT 234.700 32.310 234.960 32.630 ;
        RECT 786.700 32.310 786.960 32.630 ;
        RECT 234.760 2.400 234.900 32.310 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 56.190 17.240 56.510 17.300 ;
        RECT 697.890 17.240 698.210 17.300 ;
        RECT 56.190 17.100 698.210 17.240 ;
        RECT 56.190 17.040 56.510 17.100 ;
        RECT 697.890 17.040 698.210 17.100 ;
      LAYER via ;
        RECT 56.220 17.040 56.480 17.300 ;
        RECT 697.920 17.040 698.180 17.300 ;
      LAYER met2 ;
        RECT 698.610 600.170 698.890 604.000 ;
        RECT 697.980 600.030 698.890 600.170 ;
        RECT 697.980 17.330 698.120 600.030 ;
        RECT 698.610 600.000 698.890 600.030 ;
        RECT 56.220 17.010 56.480 17.330 ;
        RECT 697.920 17.010 698.180 17.330 ;
        RECT 56.280 2.400 56.420 17.010 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 80.110 17.920 80.430 17.980 ;
        RECT 711.690 17.920 712.010 17.980 ;
        RECT 80.110 17.780 712.010 17.920 ;
        RECT 80.110 17.720 80.430 17.780 ;
        RECT 711.690 17.720 712.010 17.780 ;
      LAYER via ;
        RECT 80.140 17.720 80.400 17.980 ;
        RECT 711.720 17.720 711.980 17.980 ;
      LAYER met2 ;
        RECT 711.030 600.170 711.310 604.000 ;
        RECT 711.030 600.030 711.920 600.170 ;
        RECT 711.030 600.000 711.310 600.030 ;
        RECT 711.780 18.010 711.920 600.030 ;
        RECT 80.140 17.690 80.400 18.010 ;
        RECT 711.720 17.690 711.980 18.010 ;
        RECT 80.200 2.400 80.340 17.690 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 718.130 596.940 718.450 597.000 ;
        RECT 721.810 596.940 722.130 597.000 ;
        RECT 718.130 596.800 722.130 596.940 ;
        RECT 718.130 596.740 718.450 596.800 ;
        RECT 721.810 596.740 722.130 596.800 ;
        RECT 718.130 579.600 718.450 579.660 ;
        RECT 718.590 579.600 718.910 579.660 ;
        RECT 718.130 579.460 718.910 579.600 ;
        RECT 718.130 579.400 718.450 579.460 ;
        RECT 718.590 579.400 718.910 579.460 ;
        RECT 718.130 531.660 718.450 531.720 ;
        RECT 718.590 531.660 718.910 531.720 ;
        RECT 718.130 531.520 718.910 531.660 ;
        RECT 718.130 531.460 718.450 531.520 ;
        RECT 718.590 531.460 718.910 531.520 ;
        RECT 718.130 524.180 718.450 524.240 ;
        RECT 719.510 524.180 719.830 524.240 ;
        RECT 718.130 524.040 719.830 524.180 ;
        RECT 718.130 523.980 718.450 524.040 ;
        RECT 719.510 523.980 719.830 524.040 ;
        RECT 718.130 435.100 718.450 435.160 ;
        RECT 719.510 435.100 719.830 435.160 ;
        RECT 718.130 434.960 719.830 435.100 ;
        RECT 718.130 434.900 718.450 434.960 ;
        RECT 719.510 434.900 719.830 434.960 ;
        RECT 718.130 427.620 718.450 427.680 ;
        RECT 719.050 427.620 719.370 427.680 ;
        RECT 718.130 427.480 719.370 427.620 ;
        RECT 718.130 427.420 718.450 427.480 ;
        RECT 719.050 427.420 719.370 427.480 ;
        RECT 718.130 379.680 718.450 379.740 ;
        RECT 719.050 379.680 719.370 379.740 ;
        RECT 718.130 379.540 719.370 379.680 ;
        RECT 718.130 379.480 718.450 379.540 ;
        RECT 719.050 379.480 719.370 379.540 ;
        RECT 718.130 331.060 718.450 331.120 ;
        RECT 719.050 331.060 719.370 331.120 ;
        RECT 718.130 330.920 719.370 331.060 ;
        RECT 718.130 330.860 718.450 330.920 ;
        RECT 719.050 330.860 719.370 330.920 ;
        RECT 718.130 283.120 718.450 283.180 ;
        RECT 719.050 283.120 719.370 283.180 ;
        RECT 718.130 282.980 719.370 283.120 ;
        RECT 718.130 282.920 718.450 282.980 ;
        RECT 719.050 282.920 719.370 282.980 ;
        RECT 719.050 172.620 719.370 172.680 ;
        RECT 719.970 172.620 720.290 172.680 ;
        RECT 719.050 172.480 720.290 172.620 ;
        RECT 719.050 172.420 719.370 172.480 ;
        RECT 719.970 172.420 720.290 172.480 ;
        RECT 718.590 96.800 718.910 96.860 ;
        RECT 719.050 96.800 719.370 96.860 ;
        RECT 718.590 96.660 719.370 96.800 ;
        RECT 718.590 96.600 718.910 96.660 ;
        RECT 719.050 96.600 719.370 96.660 ;
        RECT 103.570 18.940 103.890 19.000 ;
        RECT 718.590 18.940 718.910 19.000 ;
        RECT 103.570 18.800 718.910 18.940 ;
        RECT 103.570 18.740 103.890 18.800 ;
        RECT 718.590 18.740 718.910 18.800 ;
      LAYER via ;
        RECT 718.160 596.740 718.420 597.000 ;
        RECT 721.840 596.740 722.100 597.000 ;
        RECT 718.160 579.400 718.420 579.660 ;
        RECT 718.620 579.400 718.880 579.660 ;
        RECT 718.160 531.460 718.420 531.720 ;
        RECT 718.620 531.460 718.880 531.720 ;
        RECT 718.160 523.980 718.420 524.240 ;
        RECT 719.540 523.980 719.800 524.240 ;
        RECT 718.160 434.900 718.420 435.160 ;
        RECT 719.540 434.900 719.800 435.160 ;
        RECT 718.160 427.420 718.420 427.680 ;
        RECT 719.080 427.420 719.340 427.680 ;
        RECT 718.160 379.480 718.420 379.740 ;
        RECT 719.080 379.480 719.340 379.740 ;
        RECT 718.160 330.860 718.420 331.120 ;
        RECT 719.080 330.860 719.340 331.120 ;
        RECT 718.160 282.920 718.420 283.180 ;
        RECT 719.080 282.920 719.340 283.180 ;
        RECT 719.080 172.420 719.340 172.680 ;
        RECT 720.000 172.420 720.260 172.680 ;
        RECT 718.620 96.600 718.880 96.860 ;
        RECT 719.080 96.600 719.340 96.860 ;
        RECT 103.600 18.740 103.860 19.000 ;
        RECT 718.620 18.740 718.880 19.000 ;
      LAYER met2 ;
        RECT 723.450 600.170 723.730 604.000 ;
        RECT 721.900 600.030 723.730 600.170 ;
        RECT 721.900 597.030 722.040 600.030 ;
        RECT 723.450 600.000 723.730 600.030 ;
        RECT 718.160 596.710 718.420 597.030 ;
        RECT 721.840 596.710 722.100 597.030 ;
        RECT 718.220 579.690 718.360 596.710 ;
        RECT 718.160 579.370 718.420 579.690 ;
        RECT 718.620 579.370 718.880 579.690 ;
        RECT 718.680 531.750 718.820 579.370 ;
        RECT 718.160 531.430 718.420 531.750 ;
        RECT 718.620 531.430 718.880 531.750 ;
        RECT 718.220 524.270 718.360 531.430 ;
        RECT 718.160 523.950 718.420 524.270 ;
        RECT 719.540 523.950 719.800 524.270 ;
        RECT 719.600 435.190 719.740 523.950 ;
        RECT 718.160 434.870 718.420 435.190 ;
        RECT 719.540 434.870 719.800 435.190 ;
        RECT 718.220 427.710 718.360 434.870 ;
        RECT 718.160 427.390 718.420 427.710 ;
        RECT 719.080 427.390 719.340 427.710 ;
        RECT 719.140 379.770 719.280 427.390 ;
        RECT 718.160 379.450 718.420 379.770 ;
        RECT 719.080 379.450 719.340 379.770 ;
        RECT 718.220 331.150 718.360 379.450 ;
        RECT 718.160 330.830 718.420 331.150 ;
        RECT 719.080 330.830 719.340 331.150 ;
        RECT 719.140 283.210 719.280 330.830 ;
        RECT 718.160 282.890 718.420 283.210 ;
        RECT 719.080 282.890 719.340 283.210 ;
        RECT 718.220 282.610 718.360 282.890 ;
        RECT 718.220 282.470 718.820 282.610 ;
        RECT 718.680 220.845 718.820 282.470 ;
        RECT 718.610 220.475 718.890 220.845 ;
        RECT 719.990 220.475 720.270 220.845 ;
        RECT 720.060 172.710 720.200 220.475 ;
        RECT 719.080 172.390 719.340 172.710 ;
        RECT 720.000 172.390 720.260 172.710 ;
        RECT 719.140 96.890 719.280 172.390 ;
        RECT 718.620 96.570 718.880 96.890 ;
        RECT 719.080 96.570 719.340 96.890 ;
        RECT 718.680 19.030 718.820 96.570 ;
        RECT 103.600 18.710 103.860 19.030 ;
        RECT 718.620 18.710 718.880 19.030 ;
        RECT 103.660 2.400 103.800 18.710 ;
        RECT 103.450 -4.800 104.010 2.400 ;
      LAYER via2 ;
        RECT 718.610 220.520 718.890 220.800 ;
        RECT 719.990 220.520 720.270 220.800 ;
      LAYER met3 ;
        RECT 718.585 220.810 718.915 220.825 ;
        RECT 719.965 220.810 720.295 220.825 ;
        RECT 718.585 220.510 720.295 220.810 ;
        RECT 718.585 220.495 718.915 220.510 ;
        RECT 719.965 220.495 720.295 220.510 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 604.050 22.000 604.370 22.060 ;
        RECT 731.930 22.000 732.250 22.060 ;
        RECT 604.050 21.860 732.250 22.000 ;
        RECT 604.050 21.800 604.370 21.860 ;
        RECT 731.930 21.800 732.250 21.860 ;
        RECT 127.490 20.640 127.810 20.700 ;
        RECT 604.050 20.640 604.370 20.700 ;
        RECT 127.490 20.500 604.370 20.640 ;
        RECT 127.490 20.440 127.810 20.500 ;
        RECT 604.050 20.440 604.370 20.500 ;
      LAYER via ;
        RECT 604.080 21.800 604.340 22.060 ;
        RECT 731.960 21.800 732.220 22.060 ;
        RECT 127.520 20.440 127.780 20.700 ;
        RECT 604.080 20.440 604.340 20.700 ;
      LAYER met2 ;
        RECT 735.410 600.170 735.690 604.000 ;
        RECT 733.400 600.030 735.690 600.170 ;
        RECT 733.400 590.650 733.540 600.030 ;
        RECT 735.410 600.000 735.690 600.030 ;
        RECT 732.020 590.510 733.540 590.650 ;
        RECT 732.020 22.090 732.160 590.510 ;
        RECT 604.080 21.770 604.340 22.090 ;
        RECT 731.960 21.770 732.220 22.090 ;
        RECT 604.140 20.730 604.280 21.770 ;
        RECT 127.520 20.410 127.780 20.730 ;
        RECT 604.080 20.410 604.340 20.730 ;
        RECT 127.580 2.400 127.720 20.410 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 44.780 26.610 44.840 ;
        RECT 684.090 44.780 684.410 44.840 ;
        RECT 26.290 44.640 684.410 44.780 ;
        RECT 26.290 44.580 26.610 44.640 ;
        RECT 684.090 44.580 684.410 44.640 ;
      LAYER via ;
        RECT 26.320 44.580 26.580 44.840 ;
        RECT 684.120 44.580 684.380 44.840 ;
      LAYER met2 ;
        RECT 683.430 600.170 683.710 604.000 ;
        RECT 683.430 600.030 684.320 600.170 ;
        RECT 683.430 600.000 683.710 600.030 ;
        RECT 684.180 44.870 684.320 600.030 ;
        RECT 26.320 44.550 26.580 44.870 ;
        RECT 684.120 44.550 684.380 44.870 ;
        RECT 26.380 2.400 26.520 44.550 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 683.630 569.400 683.950 569.460 ;
        RECT 685.010 569.400 685.330 569.460 ;
        RECT 683.630 569.260 685.330 569.400 ;
        RECT 683.630 569.200 683.950 569.260 ;
        RECT 685.010 569.200 685.330 569.260 ;
        RECT 32.270 45.120 32.590 45.180 ;
        RECT 683.630 45.120 683.950 45.180 ;
        RECT 32.270 44.980 683.950 45.120 ;
        RECT 32.270 44.920 32.590 44.980 ;
        RECT 683.630 44.920 683.950 44.980 ;
      LAYER via ;
        RECT 683.660 569.200 683.920 569.460 ;
        RECT 685.040 569.200 685.300 569.460 ;
        RECT 32.300 44.920 32.560 45.180 ;
        RECT 683.660 44.920 683.920 45.180 ;
      LAYER met2 ;
        RECT 686.650 600.170 686.930 604.000 ;
        RECT 685.100 600.030 686.930 600.170 ;
        RECT 685.100 569.490 685.240 600.030 ;
        RECT 686.650 600.000 686.930 600.030 ;
        RECT 683.660 569.170 683.920 569.490 ;
        RECT 685.040 569.170 685.300 569.490 ;
        RECT 683.720 45.210 683.860 569.170 ;
        RECT 32.300 44.890 32.560 45.210 ;
        RECT 683.660 44.890 683.920 45.210 ;
        RECT 32.360 2.400 32.500 44.890 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 1982.750 367.020 3529.000 ;
        RECT 544.020 2760.520 547.020 3529.000 ;
        RECT 457.645 2610.640 459.245 2747.120 ;
        RECT 544.020 1982.750 547.020 2599.000 ;
        RECT 381.040 1710.640 382.640 1969.520 ;
        RECT 364.020 -9.320 367.020 1699.000 ;
        RECT 544.020 -9.320 547.020 1699.000 ;
        RECT 724.020 1001.000 727.020 3529.000 ;
        RECT 904.020 1001.000 907.020 3529.000 ;
        RECT 1084.020 2801.000 1087.020 3529.000 ;
        RECT 1019.545 2610.640 1021.145 2787.920 ;
        RECT 1084.020 2045.110 1087.020 2599.000 ;
        RECT 1264.020 2045.110 1267.020 3529.000 ;
        RECT 1021.040 1710.640 1022.640 2032.080 ;
        RECT 1084.020 1001.000 1087.020 1699.000 ;
        RECT 1264.020 1001.000 1267.020 1699.000 ;
        RECT 1444.020 1001.000 1447.020 3529.000 ;
        RECT 1624.020 2901.055 1627.020 3529.000 ;
        RECT 1804.020 2901.055 1807.020 3529.000 ;
        RECT 1521.040 2510.640 1522.640 2889.200 ;
        RECT 1624.020 1001.000 1627.020 2499.000 ;
        RECT 1804.020 1001.000 1807.020 2499.000 ;
        RECT 1984.020 1918.095 1987.020 3529.000 ;
        RECT 1948.870 1760.640 1950.470 1905.280 ;
        RECT 1984.020 1001.000 1987.020 1749.000 ;
        RECT 2164.020 1001.000 2167.020 3529.000 ;
        RECT 2344.020 1938.745 2347.020 3529.000 ;
        RECT 2524.020 2774.820 2527.020 3529.000 ;
        RECT 2427.190 2610.640 2428.790 2760.720 ;
        RECT 2524.020 1938.745 2527.020 2599.000 ;
        RECT 2321.040 1710.640 2322.640 1926.000 ;
        RECT 691.040 610.640 692.640 989.200 ;
        RECT 724.020 -9.320 727.020 599.000 ;
        RECT 904.020 -9.320 907.020 599.000 ;
        RECT 1084.020 -9.320 1087.020 599.000 ;
        RECT 1264.020 -9.320 1267.020 599.000 ;
        RECT 1444.020 -9.320 1447.020 599.000 ;
        RECT 1624.020 -9.320 1627.020 599.000 ;
        RECT 1804.020 -9.320 1807.020 599.000 ;
        RECT 1984.020 -9.320 1987.020 599.000 ;
        RECT 2164.020 -9.320 2167.020 599.000 ;
        RECT 2344.020 -9.320 2347.020 1699.000 ;
        RECT 2524.020 -9.320 2527.020 1699.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 457.855 2711.090 459.035 2712.270 ;
        RECT 457.855 2709.490 459.035 2710.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 381.250 1811.090 382.430 1812.270 ;
        RECT 381.250 1809.490 382.430 1810.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 1019.755 2711.090 1020.935 2712.270 ;
        RECT 1019.755 2709.490 1020.935 2710.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1521.250 2711.090 1522.430 2712.270 ;
        RECT 1521.250 2709.490 1522.430 2710.670 ;
        RECT 1521.250 2531.090 1522.430 2532.270 ;
        RECT 1521.250 2529.490 1522.430 2530.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 1021.250 1991.090 1022.430 1992.270 ;
        RECT 1021.250 1989.490 1022.430 1990.670 ;
        RECT 1021.250 1811.090 1022.430 1812.270 ;
        RECT 1021.250 1809.490 1022.430 1810.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1949.080 1811.090 1950.260 1812.270 ;
        RECT 1949.080 1809.490 1950.260 1810.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2427.400 2711.090 2428.580 2712.270 ;
        RECT 2427.400 2709.490 2428.580 2710.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 2321.250 1811.090 2322.430 1812.270 ;
        RECT 2321.250 1809.490 2322.430 1810.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 691.250 911.090 692.430 912.270 ;
        RECT 691.250 909.490 692.430 910.670 ;
        RECT 691.250 731.090 692.430 732.270 ;
        RECT 691.250 729.490 692.430 730.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 457.645 2712.380 459.245 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1019.545 2712.380 1021.145 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1521.040 2712.380 1522.640 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2427.190 2712.380 2428.790 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 457.645 2709.370 459.245 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1019.545 2709.370 1021.145 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1521.040 2709.370 1522.640 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2427.190 2709.370 2428.790 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1521.040 2532.380 1522.640 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1521.040 2529.370 1522.640 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1021.040 1992.380 1022.640 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1021.040 1989.370 1022.640 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 381.040 1812.380 382.640 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1021.040 1812.380 1022.640 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1948.870 1812.380 1950.470 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2321.040 1812.380 2322.640 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 381.040 1809.370 382.640 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1021.040 1809.370 1022.640 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1948.870 1809.370 1950.470 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2321.040 1809.370 2322.640 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 691.040 912.380 692.640 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 691.040 909.370 692.640 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 691.040 732.380 692.640 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 691.040 729.370 692.640 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 2760.520 457.020 3529.000 ;
        RECT 480.565 2610.640 482.165 2747.120 ;
        RECT 454.020 1982.750 457.020 2599.000 ;
        RECT 457.840 1710.640 459.440 1969.520 ;
        RECT 454.020 -9.320 457.020 1699.000 ;
        RECT 634.020 -9.320 637.020 3529.000 ;
        RECT 814.020 1001.000 817.020 3529.000 ;
        RECT 994.020 1001.000 997.020 3529.000 ;
        RECT 1034.375 2610.640 1035.975 2787.920 ;
        RECT 1174.020 2045.110 1177.020 3529.000 ;
        RECT 1097.840 1710.640 1099.440 2032.080 ;
        RECT 1174.020 1001.000 1177.020 1699.000 ;
        RECT 1354.020 1001.000 1357.020 3529.000 ;
        RECT 1534.020 2901.055 1537.020 3529.000 ;
        RECT 1714.020 2901.055 1717.020 3529.000 ;
        RECT 1597.840 2510.640 1599.440 2889.200 ;
        RECT 1534.020 1001.000 1537.020 2499.000 ;
        RECT 1714.020 1001.000 1717.020 2499.000 ;
        RECT 1894.020 1001.000 1897.020 3529.000 ;
        RECT 2074.020 1918.095 2077.020 3529.000 ;
        RECT 1973.020 1760.640 1974.620 1905.280 ;
        RECT 2074.020 1001.000 2077.020 1749.000 ;
        RECT 767.840 610.640 769.440 989.200 ;
        RECT 814.020 -9.320 817.020 599.000 ;
        RECT 994.020 -9.320 997.020 599.000 ;
        RECT 1174.020 -9.320 1177.020 599.000 ;
        RECT 1354.020 -9.320 1357.020 599.000 ;
        RECT 1534.020 -9.320 1537.020 599.000 ;
        RECT 1714.020 -9.320 1717.020 599.000 ;
        RECT 1894.020 -9.320 1897.020 599.000 ;
        RECT 2074.020 -9.320 2077.020 599.000 ;
        RECT 2254.020 -9.320 2257.020 3529.000 ;
        RECT 2434.020 2774.820 2437.020 3529.000 ;
        RECT 2452.490 2610.640 2454.090 2760.720 ;
        RECT 2434.020 1938.745 2437.020 2599.000 ;
        RECT 2397.840 1710.640 2399.440 1926.000 ;
        RECT 2434.020 -9.320 2437.020 1699.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 480.775 2621.090 481.955 2622.270 ;
        RECT 480.775 2619.490 481.955 2620.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 458.050 1901.090 459.230 1902.270 ;
        RECT 458.050 1899.490 459.230 1900.670 ;
        RECT 458.050 1721.090 459.230 1722.270 ;
        RECT 458.050 1719.490 459.230 1720.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 1034.585 2621.090 1035.765 2622.270 ;
        RECT 1034.585 2619.490 1035.765 2620.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1598.050 2801.090 1599.230 2802.270 ;
        RECT 1598.050 2799.490 1599.230 2800.670 ;
        RECT 1598.050 2621.090 1599.230 2622.270 ;
        RECT 1598.050 2619.490 1599.230 2620.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 1098.050 1901.090 1099.230 1902.270 ;
        RECT 1098.050 1899.490 1099.230 1900.670 ;
        RECT 1098.050 1721.090 1099.230 1722.270 ;
        RECT 1098.050 1719.490 1099.230 1720.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2452.700 2621.090 2453.880 2622.270 ;
        RECT 2452.700 2619.490 2453.880 2620.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1973.230 1901.090 1974.410 1902.270 ;
        RECT 1973.230 1899.490 1974.410 1900.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2398.050 1901.090 2399.230 1902.270 ;
        RECT 2398.050 1899.490 2399.230 1900.670 ;
        RECT 2398.050 1721.090 2399.230 1722.270 ;
        RECT 2398.050 1719.490 2399.230 1720.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 768.050 821.090 769.230 822.270 ;
        RECT 768.050 819.490 769.230 820.670 ;
        RECT 768.050 641.090 769.230 642.270 ;
        RECT 768.050 639.490 769.230 640.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1597.840 2802.380 1599.440 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1597.840 2799.370 1599.440 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 480.565 2622.380 482.165 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1034.375 2622.380 1035.975 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1597.840 2622.380 1599.440 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2452.490 2622.380 2454.090 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 480.565 2619.370 482.165 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1034.375 2619.370 1035.975 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1597.840 2619.370 1599.440 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2452.490 2619.370 2454.090 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 457.840 1902.380 459.440 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1097.840 1902.380 1099.440 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 1973.020 1902.380 1974.620 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2397.840 1902.380 2399.440 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 457.840 1899.370 459.440 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1097.840 1899.370 1099.440 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 1973.020 1899.370 1974.620 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2397.840 1899.370 2399.440 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 457.840 1722.380 459.440 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1097.840 1722.380 1099.440 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2397.840 1722.380 2399.440 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 457.840 1719.370 459.440 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1097.840 1719.370 1099.440 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2397.840 1719.370 2399.440 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 767.840 822.380 769.440 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 767.840 819.370 769.440 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 767.840 642.380 769.440 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 767.840 639.370 769.440 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 382.020 1982.750 385.020 3538.400 ;
        RECT 562.020 2760.520 565.020 3538.400 ;
        RECT 562.020 1982.750 565.020 2599.000 ;
        RECT 382.020 -18.720 385.020 1699.000 ;
        RECT 562.020 -18.720 565.020 1699.000 ;
        RECT 742.020 1001.000 745.020 3538.400 ;
        RECT 922.020 1001.000 925.020 3538.400 ;
        RECT 1102.020 2045.110 1105.020 3538.400 ;
        RECT 1282.020 2045.110 1285.020 3538.400 ;
        RECT 1102.020 1001.000 1105.020 1699.000 ;
        RECT 1282.020 1001.000 1285.020 1699.000 ;
        RECT 1462.020 1001.000 1465.020 3538.400 ;
        RECT 1642.020 2901.055 1645.020 3538.400 ;
        RECT 1822.020 2901.055 1825.020 3538.400 ;
        RECT 1642.020 1001.000 1645.020 2499.000 ;
        RECT 1822.020 1001.000 1825.020 2499.000 ;
        RECT 2002.020 1918.095 2005.020 3538.400 ;
        RECT 2002.020 1001.000 2005.020 1749.000 ;
        RECT 742.020 -18.720 745.020 599.000 ;
        RECT 922.020 -18.720 925.020 599.000 ;
        RECT 1102.020 -18.720 1105.020 599.000 ;
        RECT 1282.020 -18.720 1285.020 599.000 ;
        RECT 1462.020 -18.720 1465.020 599.000 ;
        RECT 1642.020 -18.720 1645.020 599.000 ;
        RECT 1822.020 -18.720 1825.020 599.000 ;
        RECT 2002.020 -18.720 2005.020 599.000 ;
        RECT 2182.020 -18.720 2185.020 3538.400 ;
        RECT 2362.020 1938.745 2365.020 3538.400 ;
        RECT 2542.020 2774.820 2545.020 3538.400 ;
        RECT 2362.020 -18.720 2365.020 1699.000 ;
        RECT 2542.020 -18.720 2545.020 2599.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 292.020 -18.720 295.020 3538.400 ;
        RECT 472.020 2760.520 475.020 3538.400 ;
        RECT 472.020 1982.750 475.020 2599.000 ;
        RECT 472.020 -18.720 475.020 1699.000 ;
        RECT 652.020 -18.720 655.020 3538.400 ;
        RECT 832.020 1001.000 835.020 3538.400 ;
        RECT 1012.020 2801.000 1015.020 3538.400 ;
        RECT 1012.020 2045.110 1015.020 2599.000 ;
        RECT 1192.020 2045.110 1195.020 3538.400 ;
        RECT 1012.020 1001.000 1015.020 1699.000 ;
        RECT 1192.020 1001.000 1195.020 1699.000 ;
        RECT 1372.020 1001.000 1375.020 3538.400 ;
        RECT 1552.020 2901.055 1555.020 3538.400 ;
        RECT 1732.020 2901.055 1735.020 3538.400 ;
        RECT 1552.020 1001.000 1555.020 2499.000 ;
        RECT 1732.020 1001.000 1735.020 2499.000 ;
        RECT 1912.020 1001.000 1915.020 3538.400 ;
        RECT 2092.020 1001.000 2095.020 3538.400 ;
        RECT 832.020 -18.720 835.020 599.000 ;
        RECT 1012.020 -18.720 1015.020 599.000 ;
        RECT 1192.020 -18.720 1195.020 599.000 ;
        RECT 1372.020 -18.720 1375.020 599.000 ;
        RECT 1552.020 -18.720 1555.020 599.000 ;
        RECT 1732.020 -18.720 1735.020 599.000 ;
        RECT 1912.020 -18.720 1915.020 599.000 ;
        RECT 2092.020 -18.720 2095.020 599.000 ;
        RECT 2272.020 -18.720 2275.020 3538.400 ;
        RECT 2452.020 2774.820 2455.020 3538.400 ;
        RECT 2452.020 1938.745 2455.020 2599.000 ;
        RECT 2452.020 -18.720 2455.020 1699.000 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 400.020 1982.750 403.020 3547.800 ;
        RECT 580.020 1982.750 583.020 3547.800 ;
        RECT 400.020 -28.120 403.020 1699.000 ;
        RECT 580.020 -28.120 583.020 1699.000 ;
        RECT 760.020 1001.000 763.020 3547.800 ;
        RECT 940.020 1001.000 943.020 3547.800 ;
        RECT 1120.020 2045.110 1123.020 3547.800 ;
        RECT 1300.020 2045.110 1303.020 3547.800 ;
        RECT 1120.020 1001.000 1123.020 1699.000 ;
        RECT 1300.020 1001.000 1303.020 1699.000 ;
        RECT 1480.020 1001.000 1483.020 3547.800 ;
        RECT 1660.020 2901.055 1663.020 3547.800 ;
        RECT 1840.020 2901.055 1843.020 3547.800 ;
        RECT 1660.020 1001.000 1663.020 2499.000 ;
        RECT 1840.020 1001.000 1843.020 2499.000 ;
        RECT 2020.020 1918.095 2023.020 3547.800 ;
        RECT 2020.020 1001.000 2023.020 1749.000 ;
        RECT 760.020 -28.120 763.020 599.000 ;
        RECT 940.020 -28.120 943.020 599.000 ;
        RECT 1120.020 -28.120 1123.020 599.000 ;
        RECT 1300.020 -28.120 1303.020 599.000 ;
        RECT 1480.020 -28.120 1483.020 599.000 ;
        RECT 1660.020 -28.120 1663.020 599.000 ;
        RECT 1840.020 -28.120 1843.020 599.000 ;
        RECT 2020.020 -28.120 2023.020 599.000 ;
        RECT 2200.020 -28.120 2203.020 3547.800 ;
        RECT 2380.020 1938.745 2383.020 3547.800 ;
        RECT 2380.020 -28.120 2383.020 1699.000 ;
        RECT 2560.020 -28.120 2563.020 3547.800 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 310.020 -28.120 313.020 3547.800 ;
        RECT 490.020 2760.520 493.020 3547.800 ;
        RECT 490.020 1982.750 493.020 2599.000 ;
        RECT 490.020 -28.120 493.020 1699.000 ;
        RECT 670.020 1001.000 673.020 3547.800 ;
        RECT 850.020 1001.000 853.020 3547.800 ;
        RECT 1030.020 2801.000 1033.020 3547.800 ;
        RECT 1030.020 2045.110 1033.020 2599.000 ;
        RECT 1210.020 2045.110 1213.020 3547.800 ;
        RECT 1030.020 1001.000 1033.020 1699.000 ;
        RECT 1210.020 1001.000 1213.020 1699.000 ;
        RECT 1390.020 1001.000 1393.020 3547.800 ;
        RECT 1570.020 2901.055 1573.020 3547.800 ;
        RECT 1750.020 2901.055 1753.020 3547.800 ;
        RECT 1570.020 1001.000 1573.020 2499.000 ;
        RECT 1750.020 1001.000 1753.020 2499.000 ;
        RECT 1930.020 1918.095 1933.020 3547.800 ;
        RECT 1930.020 1001.000 1933.020 1749.000 ;
        RECT 2110.020 1001.000 2113.020 3547.800 ;
        RECT 670.020 -28.120 673.020 599.000 ;
        RECT 850.020 -28.120 853.020 599.000 ;
        RECT 1030.020 -28.120 1033.020 599.000 ;
        RECT 1210.020 -28.120 1213.020 599.000 ;
        RECT 1390.020 -28.120 1393.020 599.000 ;
        RECT 1570.020 -28.120 1573.020 599.000 ;
        RECT 1750.020 -28.120 1753.020 599.000 ;
        RECT 1930.020 -28.120 1933.020 599.000 ;
        RECT 2110.020 -28.120 2113.020 599.000 ;
        RECT 2290.020 -28.120 2293.020 3547.800 ;
        RECT 2470.020 2774.820 2473.020 3547.800 ;
        RECT 2470.020 1938.745 2473.020 2599.000 ;
        RECT 2470.020 -28.120 2473.020 1699.000 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 418.020 1982.750 421.020 3557.200 ;
        RECT 598.020 1982.750 601.020 3557.200 ;
        RECT 418.020 -37.520 421.020 1699.000 ;
        RECT 598.020 -37.520 601.020 1699.000 ;
        RECT 778.020 1001.000 781.020 3557.200 ;
        RECT 958.020 1001.000 961.020 3557.200 ;
        RECT 1138.020 2045.110 1141.020 3557.200 ;
        RECT 1318.020 2045.110 1321.020 3557.200 ;
        RECT 1498.020 2901.055 1501.020 3557.200 ;
        RECT 1678.020 2901.055 1681.020 3557.200 ;
        RECT 1858.020 2901.055 1861.020 3557.200 ;
        RECT 1138.020 1001.000 1141.020 1699.000 ;
        RECT 1318.020 1001.000 1321.020 1699.000 ;
        RECT 1498.020 1001.000 1501.020 2499.000 ;
        RECT 1678.020 1001.000 1681.020 2499.000 ;
        RECT 1858.020 1001.000 1861.020 2499.000 ;
        RECT 2038.020 1918.095 2041.020 3557.200 ;
        RECT 2038.020 1001.000 2041.020 1749.000 ;
        RECT 778.020 -37.520 781.020 599.000 ;
        RECT 958.020 -37.520 961.020 599.000 ;
        RECT 1138.020 -37.520 1141.020 599.000 ;
        RECT 1318.020 -37.520 1321.020 599.000 ;
        RECT 1498.020 -37.520 1501.020 599.000 ;
        RECT 1678.020 -37.520 1681.020 599.000 ;
        RECT 1858.020 -37.520 1861.020 599.000 ;
        RECT 2038.020 -37.520 2041.020 599.000 ;
        RECT 2218.020 -37.520 2221.020 3557.200 ;
        RECT 2398.020 2774.820 2401.020 3557.200 ;
        RECT 2398.020 1938.745 2401.020 2599.000 ;
        RECT 2398.020 -37.520 2401.020 1699.000 ;
        RECT 2578.020 -37.520 2581.020 3557.200 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 328.020 -37.520 331.020 3557.200 ;
        RECT 508.020 2760.520 511.020 3557.200 ;
        RECT 508.020 1982.750 511.020 2599.000 ;
        RECT 508.020 -37.520 511.020 1699.000 ;
        RECT 688.020 1001.000 691.020 3557.200 ;
        RECT 868.020 1001.000 871.020 3557.200 ;
        RECT 1048.020 2801.000 1051.020 3557.200 ;
        RECT 1048.020 2045.110 1051.020 2599.000 ;
        RECT 1228.020 2045.110 1231.020 3557.200 ;
        RECT 1048.020 1001.000 1051.020 1699.000 ;
        RECT 1228.020 1001.000 1231.020 1699.000 ;
        RECT 1408.020 1001.000 1411.020 3557.200 ;
        RECT 1588.020 2901.055 1591.020 3557.200 ;
        RECT 1768.020 2901.055 1771.020 3557.200 ;
        RECT 1588.020 1001.000 1591.020 2499.000 ;
        RECT 1768.020 1001.000 1771.020 2499.000 ;
        RECT 1948.020 1918.095 1951.020 3557.200 ;
        RECT 1948.020 1001.000 1951.020 1749.000 ;
        RECT 2128.020 1001.000 2131.020 3557.200 ;
        RECT 2308.020 1938.745 2311.020 3557.200 ;
        RECT 2488.020 2774.820 2491.020 3557.200 ;
        RECT 2488.020 1938.745 2491.020 2599.000 ;
        RECT 688.020 -37.520 691.020 599.000 ;
        RECT 868.020 -37.520 871.020 599.000 ;
        RECT 1048.020 -37.520 1051.020 599.000 ;
        RECT 1228.020 -37.520 1231.020 599.000 ;
        RECT 1408.020 -37.520 1411.020 599.000 ;
        RECT 1588.020 -37.520 1591.020 599.000 ;
        RECT 1768.020 -37.520 1771.020 599.000 ;
        RECT 1948.020 -37.520 1951.020 599.000 ;
        RECT 2128.020 -37.520 2131.020 599.000 ;
        RECT 2308.020 -37.520 2311.020 1699.000 ;
        RECT 2488.020 -37.520 2491.020 1699.000 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 435.520 2610.795 573.060 2746.965 ;
        RECT 1005.520 2610.795 1094.300 2787.765 ;
        RECT 1505.520 2510.795 1883.640 2889.045 ;
        RECT 2402.690 2610.795 2554.490 2760.565 ;
        RECT 365.520 1710.795 625.420 1969.365 ;
        RECT 1005.520 1710.795 1327.520 2031.925 ;
        RECT 1925.520 1760.795 2070.420 1905.125 ;
        RECT 2305.520 1710.795 2521.260 1925.845 ;
        RECT 675.520 610.795 2164.080 998.055 ;
      LAYER met1 ;
        RECT 1352.010 2918.120 1352.330 2918.180 ;
        RECT 1535.090 2918.120 1535.410 2918.180 ;
        RECT 1352.010 2917.980 1535.410 2918.120 ;
        RECT 1352.010 2917.920 1352.330 2917.980 ;
        RECT 1535.090 2917.920 1535.410 2917.980 ;
        RECT 1414.110 2917.780 1414.430 2917.840 ;
        RECT 1567.290 2917.780 1567.610 2917.840 ;
        RECT 1414.110 2917.640 1567.610 2917.780 ;
        RECT 1414.110 2917.580 1414.430 2917.640 ;
        RECT 1567.290 2917.580 1567.610 2917.640 ;
        RECT 1448.610 2916.080 1448.930 2916.140 ;
        RECT 1641.810 2916.080 1642.130 2916.140 ;
        RECT 1448.610 2915.940 1642.130 2916.080 ;
        RECT 1448.610 2915.880 1448.930 2915.940 ;
        RECT 1641.810 2915.880 1642.130 2915.940 ;
        RECT 1379.610 2915.740 1379.930 2915.800 ;
        RECT 1598.570 2915.740 1598.890 2915.800 ;
        RECT 1379.610 2915.600 1598.890 2915.740 ;
        RECT 1379.610 2915.540 1379.930 2915.600 ;
        RECT 1598.570 2915.540 1598.890 2915.600 ;
        RECT 1405.830 2915.400 1406.150 2915.460 ;
        RECT 1630.770 2915.400 1631.090 2915.460 ;
        RECT 1405.830 2915.260 1631.090 2915.400 ;
        RECT 1405.830 2915.200 1406.150 2915.260 ;
        RECT 1630.770 2915.200 1631.090 2915.260 ;
        RECT 1469.310 2915.060 1469.630 2915.120 ;
        RECT 1694.250 2915.060 1694.570 2915.120 ;
        RECT 1469.310 2914.920 1694.570 2915.060 ;
        RECT 1469.310 2914.860 1469.630 2914.920 ;
        RECT 1694.250 2914.860 1694.570 2914.920 ;
        RECT 1501.970 2914.720 1502.290 2914.780 ;
        RECT 1768.770 2914.720 1769.090 2914.780 ;
        RECT 1501.970 2914.580 1769.090 2914.720 ;
        RECT 1501.970 2914.520 1502.290 2914.580 ;
        RECT 1768.770 2914.520 1769.090 2914.580 ;
        RECT 1502.430 2914.380 1502.750 2914.440 ;
        RECT 1779.810 2914.380 1780.130 2914.440 ;
        RECT 1502.430 2914.240 1780.130 2914.380 ;
        RECT 1502.430 2914.180 1502.750 2914.240 ;
        RECT 1779.810 2914.180 1780.130 2914.240 ;
        RECT 1455.510 2914.040 1455.830 2914.100 ;
        RECT 1758.650 2914.040 1758.970 2914.100 ;
        RECT 1455.510 2913.900 1758.970 2914.040 ;
        RECT 1455.510 2913.840 1455.830 2913.900 ;
        RECT 1758.650 2913.840 1758.970 2913.900 ;
        RECT 1372.710 2913.700 1373.030 2913.760 ;
        RECT 1843.290 2913.700 1843.610 2913.760 ;
        RECT 1372.710 2913.560 1843.610 2913.700 ;
        RECT 1372.710 2913.500 1373.030 2913.560 ;
        RECT 1843.290 2913.500 1843.610 2913.560 ;
        RECT 1494.610 2913.360 1494.930 2913.420 ;
        RECT 1705.290 2913.360 1705.610 2913.420 ;
        RECT 1494.610 2913.220 1705.610 2913.360 ;
        RECT 1494.610 2913.160 1494.930 2913.220 ;
        RECT 1705.290 2913.160 1705.610 2913.220 ;
        RECT 1789.930 2913.360 1790.250 2913.420 ;
        RECT 1895.270 2913.360 1895.590 2913.420 ;
        RECT 1789.930 2913.220 1895.590 2913.360 ;
        RECT 1789.930 2913.160 1790.250 2913.220 ;
        RECT 1895.270 2913.160 1895.590 2913.220 ;
        RECT 1501.510 2913.020 1501.830 2913.080 ;
        RECT 1812.010 2913.020 1812.330 2913.080 ;
        RECT 1501.510 2912.880 1812.330 2913.020 ;
        RECT 1501.510 2912.820 1501.830 2912.880 ;
        RECT 1812.010 2912.820 1812.330 2912.880 ;
        RECT 1833.170 2913.020 1833.490 2913.080 ;
        RECT 1887.910 2913.020 1888.230 2913.080 ;
        RECT 1833.170 2912.880 1888.230 2913.020 ;
        RECT 1833.170 2912.820 1833.490 2912.880 ;
        RECT 1887.910 2912.820 1888.230 2912.880 ;
        RECT 1496.450 2912.680 1496.770 2912.740 ;
        RECT 1662.970 2912.680 1663.290 2912.740 ;
        RECT 1496.450 2912.540 1663.290 2912.680 ;
        RECT 1496.450 2912.480 1496.770 2912.540 ;
        RECT 1662.970 2912.480 1663.290 2912.540 ;
        RECT 1854.330 2912.680 1854.650 2912.740 ;
        RECT 1886.530 2912.680 1886.850 2912.740 ;
        RECT 1854.330 2912.540 1886.850 2912.680 ;
        RECT 1854.330 2912.480 1854.650 2912.540 ;
        RECT 1886.530 2912.480 1886.850 2912.540 ;
        RECT 1493.690 2912.340 1494.010 2912.400 ;
        RECT 1609.610 2912.340 1609.930 2912.400 ;
        RECT 1493.690 2912.200 1609.930 2912.340 ;
        RECT 1493.690 2912.140 1494.010 2912.200 ;
        RECT 1609.610 2912.140 1609.930 2912.200 ;
        RECT 1864.450 2912.340 1864.770 2912.400 ;
        RECT 1887.450 2912.340 1887.770 2912.400 ;
        RECT 1864.450 2912.200 1887.770 2912.340 ;
        RECT 1864.450 2912.140 1864.770 2912.200 ;
        RECT 1887.450 2912.140 1887.770 2912.200 ;
        RECT 1494.150 2912.000 1494.470 2912.060 ;
        RECT 1546.130 2912.000 1546.450 2912.060 ;
        RECT 1494.150 2911.860 1546.450 2912.000 ;
        RECT 1494.150 2911.800 1494.470 2911.860 ;
        RECT 1546.130 2911.800 1546.450 2911.860 ;
        RECT 1495.990 2898.400 1496.310 2898.460 ;
        RECT 1524.050 2898.400 1524.370 2898.460 ;
        RECT 1495.990 2898.260 1524.370 2898.400 ;
        RECT 1495.990 2898.200 1496.310 2898.260 ;
        RECT 1524.050 2898.200 1524.370 2898.260 ;
        RECT 1652.850 2897.380 1653.170 2897.440 ;
        RECT 1693.330 2897.380 1693.650 2897.440 ;
        RECT 1652.850 2897.240 1693.650 2897.380 ;
        RECT 1652.850 2897.180 1653.170 2897.240 ;
        RECT 1693.330 2897.180 1693.650 2897.240 ;
        RECT 1534.720 2896.900 1549.580 2897.040 ;
        RECT 1497.370 2896.700 1497.690 2896.760 ;
        RECT 1503.350 2896.700 1503.670 2896.760 ;
        RECT 1497.370 2896.560 1503.670 2896.700 ;
        RECT 1497.370 2896.500 1497.690 2896.560 ;
        RECT 1503.350 2896.500 1503.670 2896.560 ;
        RECT 1490.010 2894.320 1490.330 2894.380 ;
        RECT 1490.010 2894.180 1521.520 2894.320 ;
        RECT 1490.010 2894.120 1490.330 2894.180 ;
        RECT 1521.380 2893.980 1521.520 2894.180 ;
        RECT 1534.720 2893.980 1534.860 2896.900 ;
        RECT 1549.440 2895.680 1549.580 2896.900 ;
        RECT 1715.960 2896.900 1727.600 2897.040 ;
        RECT 1652.850 2896.500 1653.170 2896.760 ;
        RECT 1693.330 2896.500 1693.650 2896.760 ;
        RECT 1549.440 2895.540 1550.040 2895.680 ;
        RECT 1549.900 2895.000 1550.040 2895.540 ;
        RECT 1549.440 2894.860 1550.040 2895.000 ;
        RECT 1549.440 2894.320 1549.580 2894.860 ;
        RECT 1611.080 2894.520 1635.140 2894.660 ;
        RECT 1611.080 2894.320 1611.220 2894.520 ;
        RECT 1549.440 2894.180 1587.300 2894.320 ;
        RECT 1521.380 2893.840 1534.860 2893.980 ;
        RECT 1587.160 2893.980 1587.300 2894.180 ;
        RECT 1609.700 2894.180 1611.220 2894.320 ;
        RECT 1635.000 2894.320 1635.140 2894.520 ;
        RECT 1652.940 2894.320 1653.080 2896.500 ;
        RECT 1693.420 2896.360 1693.560 2896.500 ;
        RECT 1693.420 2896.220 1695.400 2896.360 ;
        RECT 1695.260 2895.000 1695.400 2896.220 ;
        RECT 1715.960 2895.000 1716.100 2896.900 ;
        RECT 1695.260 2894.860 1716.100 2895.000 ;
        RECT 1635.000 2894.180 1653.080 2894.320 ;
        RECT 1609.700 2893.980 1609.840 2894.180 ;
        RECT 1587.160 2893.840 1609.840 2893.980 ;
        RECT 1727.460 2893.640 1727.600 2896.900 ;
        RECT 1801.890 2896.500 1802.210 2896.760 ;
        RECT 1876.870 2896.700 1877.190 2896.760 ;
        RECT 1894.810 2896.700 1895.130 2896.760 ;
        RECT 1876.870 2896.560 1895.130 2896.700 ;
        RECT 1876.870 2896.500 1877.190 2896.560 ;
        RECT 1894.810 2896.500 1895.130 2896.560 ;
        RECT 1801.980 2894.660 1802.120 2896.500 ;
        RECT 1801.060 2894.520 1802.120 2894.660 ;
        RECT 1801.060 2894.320 1801.200 2894.520 ;
        RECT 1800.600 2894.180 1801.200 2894.320 ;
        RECT 1800.600 2893.980 1800.740 2894.180 ;
        RECT 1752.760 2893.840 1800.740 2893.980 ;
        RECT 1752.760 2893.640 1752.900 2893.840 ;
        RECT 1727.460 2893.500 1752.900 2893.640 ;
        RECT 1406.290 2863.520 1406.610 2863.780 ;
        RECT 1406.380 2863.100 1406.520 2863.520 ;
        RECT 1406.290 2862.840 1406.610 2863.100 ;
        RECT 1358.910 2849.780 1359.230 2849.840 ;
        RECT 1483.570 2849.780 1483.890 2849.840 ;
        RECT 1358.910 2849.640 1483.890 2849.780 ;
        RECT 1358.910 2849.580 1359.230 2849.640 ;
        RECT 1483.570 2849.580 1483.890 2849.640 ;
        RECT 1405.370 2849.100 1405.690 2849.160 ;
        RECT 1406.290 2849.100 1406.610 2849.160 ;
        RECT 1405.370 2848.960 1406.610 2849.100 ;
        RECT 1405.370 2848.900 1405.690 2848.960 ;
        RECT 1406.290 2848.900 1406.610 2848.960 ;
        RECT 1000.570 2810.680 1000.890 2810.740 ;
        RECT 1048.410 2810.680 1048.730 2810.740 ;
        RECT 1000.570 2810.540 1048.730 2810.680 ;
        RECT 1000.570 2810.480 1000.890 2810.540 ;
        RECT 1048.410 2810.480 1048.730 2810.540 ;
        RECT 978.950 2810.340 979.270 2810.400 ;
        RECT 1073.710 2810.340 1074.030 2810.400 ;
        RECT 978.950 2810.200 1074.030 2810.340 ;
        RECT 978.950 2810.140 979.270 2810.200 ;
        RECT 1073.710 2810.140 1074.030 2810.200 ;
        RECT 978.490 2810.000 978.810 2810.060 ;
        RECT 1027.710 2810.000 1028.030 2810.060 ;
        RECT 978.490 2809.860 1028.030 2810.000 ;
        RECT 978.490 2809.800 978.810 2809.860 ;
        RECT 1027.710 2809.800 1028.030 2809.860 ;
        RECT 986.310 2809.660 986.630 2809.720 ;
        RECT 1043.350 2809.660 1043.670 2809.720 ;
        RECT 986.310 2809.520 1043.670 2809.660 ;
        RECT 986.310 2809.460 986.630 2809.520 ;
        RECT 1043.350 2809.460 1043.670 2809.520 ;
        RECT 979.410 2809.320 979.730 2809.380 ;
        RECT 1058.070 2809.320 1058.390 2809.380 ;
        RECT 979.410 2809.180 1058.390 2809.320 ;
        RECT 979.410 2809.120 979.730 2809.180 ;
        RECT 1058.070 2809.120 1058.390 2809.180 ;
        RECT 985.850 2808.980 986.170 2809.040 ;
        RECT 1000.570 2808.980 1000.890 2809.040 ;
        RECT 985.850 2808.840 1000.890 2808.980 ;
        RECT 985.850 2808.780 986.170 2808.840 ;
        RECT 1000.570 2808.780 1000.890 2808.840 ;
        RECT 1048.410 2808.640 1048.730 2808.700 ;
        RECT 1089.350 2808.640 1089.670 2808.700 ;
        RECT 1048.410 2808.500 1089.670 2808.640 ;
        RECT 1048.410 2808.440 1048.730 2808.500 ;
        RECT 1089.350 2808.440 1089.670 2808.500 ;
        RECT 1405.370 2801.500 1405.690 2801.560 ;
        RECT 1406.290 2801.500 1406.610 2801.560 ;
        RECT 1405.370 2801.360 1406.610 2801.500 ;
        RECT 1405.370 2801.300 1405.690 2801.360 ;
        RECT 1406.290 2801.300 1406.610 2801.360 ;
        RECT 985.390 2801.160 985.710 2801.220 ;
        RECT 1010.230 2801.160 1010.550 2801.220 ;
        RECT 985.390 2801.020 1010.550 2801.160 ;
        RECT 985.390 2800.960 985.710 2801.020 ;
        RECT 1010.230 2800.960 1010.550 2801.020 ;
        RECT 445.810 2769.540 446.130 2769.600 ;
        RECT 782.990 2769.540 783.310 2769.600 ;
        RECT 445.810 2769.400 783.310 2769.540 ;
        RECT 445.810 2769.340 446.130 2769.400 ;
        RECT 782.990 2769.340 783.310 2769.400 ;
        RECT 532.290 2768.180 532.610 2768.240 ;
        RECT 686.390 2768.180 686.710 2768.240 ;
        RECT 532.290 2768.040 686.710 2768.180 ;
        RECT 532.290 2767.980 532.610 2768.040 ;
        RECT 686.390 2767.980 686.710 2768.040 ;
        RECT 518.490 2767.840 518.810 2767.900 ;
        RECT 707.090 2767.840 707.410 2767.900 ;
        RECT 518.490 2767.700 707.410 2767.840 ;
        RECT 518.490 2767.640 518.810 2767.700 ;
        RECT 707.090 2767.640 707.410 2767.700 ;
        RECT 489.050 2767.500 489.370 2767.560 ;
        RECT 755.390 2767.500 755.710 2767.560 ;
        RECT 489.050 2767.360 755.710 2767.500 ;
        RECT 489.050 2767.300 489.370 2767.360 ;
        RECT 755.390 2767.300 755.710 2767.360 ;
      LAYER met1 ;
        RECT 432.830 2606.500 575.750 2747.120 ;
      LAYER met1 ;
        RECT 588.870 2684.200 589.190 2684.260 ;
        RECT 700.190 2684.200 700.510 2684.260 ;
        RECT 588.870 2684.060 700.510 2684.200 ;
        RECT 588.870 2684.000 589.190 2684.060 ;
        RECT 700.190 2684.000 700.510 2684.060 ;
        RECT 588.870 2663.800 589.190 2663.860 ;
        RECT 769.190 2663.800 769.510 2663.860 ;
        RECT 588.870 2663.660 769.510 2663.800 ;
        RECT 588.870 2663.600 589.190 2663.660 ;
        RECT 769.190 2663.600 769.510 2663.660 ;
      LAYER met1 ;
        RECT 1002.830 2610.640 1095.150 2787.920 ;
      LAYER met1 ;
        RECT 1365.810 2781.100 1366.130 2781.160 ;
        RECT 1489.090 2781.100 1489.410 2781.160 ;
        RECT 1365.810 2780.960 1489.410 2781.100 ;
        RECT 1365.810 2780.900 1366.130 2780.960 ;
        RECT 1489.090 2780.900 1489.410 2780.960 ;
        RECT 1406.290 2767.160 1406.610 2767.220 ;
        RECT 1406.290 2767.020 1406.980 2767.160 ;
        RECT 1406.290 2766.960 1406.610 2767.020 ;
        RECT 1406.840 2766.880 1406.980 2767.020 ;
        RECT 1406.750 2766.620 1407.070 2766.880 ;
        RECT 1357.530 2753.220 1357.850 2753.280 ;
        RECT 1358.910 2753.220 1359.230 2753.280 ;
        RECT 1357.530 2753.080 1359.230 2753.220 ;
        RECT 1357.530 2753.020 1357.850 2753.080 ;
        RECT 1358.910 2753.020 1359.230 2753.080 ;
        RECT 1406.290 2753.220 1406.610 2753.280 ;
        RECT 1406.750 2753.220 1407.070 2753.280 ;
        RECT 1406.290 2753.080 1407.070 2753.220 ;
        RECT 1406.290 2753.020 1406.610 2753.080 ;
        RECT 1406.750 2753.020 1407.070 2753.080 ;
        RECT 1405.370 2752.540 1405.690 2752.600 ;
        RECT 1406.290 2752.540 1406.610 2752.600 ;
        RECT 1405.370 2752.400 1406.610 2752.540 ;
        RECT 1405.370 2752.340 1405.690 2752.400 ;
        RECT 1406.290 2752.340 1406.610 2752.400 ;
        RECT 1357.530 2729.080 1357.850 2729.140 ;
        RECT 1358.910 2729.080 1359.230 2729.140 ;
        RECT 1357.530 2728.940 1359.230 2729.080 ;
        RECT 1357.530 2728.880 1357.850 2728.940 ;
        RECT 1358.910 2728.880 1359.230 2728.940 ;
        RECT 1357.530 2704.940 1357.850 2705.000 ;
        RECT 1357.990 2704.940 1358.310 2705.000 ;
        RECT 1357.530 2704.800 1358.310 2704.940 ;
        RECT 1357.530 2704.740 1357.850 2704.800 ;
        RECT 1357.990 2704.740 1358.310 2704.800 ;
        RECT 1405.370 2704.940 1405.690 2705.000 ;
        RECT 1406.290 2704.940 1406.610 2705.000 ;
        RECT 1405.370 2704.800 1406.610 2704.940 ;
        RECT 1405.370 2704.740 1405.690 2704.800 ;
        RECT 1406.290 2704.740 1406.610 2704.800 ;
        RECT 1434.810 2691.340 1435.130 2691.400 ;
        RECT 1488.170 2691.340 1488.490 2691.400 ;
        RECT 1434.810 2691.200 1488.490 2691.340 ;
        RECT 1434.810 2691.140 1435.130 2691.200 ;
        RECT 1488.170 2691.140 1488.490 2691.200 ;
        RECT 1406.290 2670.400 1406.610 2670.660 ;
        RECT 1406.380 2670.260 1406.520 2670.400 ;
        RECT 1406.750 2670.260 1407.070 2670.320 ;
        RECT 1406.380 2670.120 1407.070 2670.260 ;
        RECT 1406.750 2670.060 1407.070 2670.120 ;
        RECT 1358.910 2656.660 1359.230 2656.720 ;
        RECT 1359.830 2656.660 1360.150 2656.720 ;
        RECT 1358.910 2656.520 1360.150 2656.660 ;
        RECT 1358.910 2656.460 1359.230 2656.520 ;
        RECT 1359.830 2656.460 1360.150 2656.520 ;
        RECT 1406.290 2656.660 1406.610 2656.720 ;
        RECT 1406.750 2656.660 1407.070 2656.720 ;
        RECT 1406.290 2656.520 1407.070 2656.660 ;
        RECT 1406.290 2656.460 1406.610 2656.520 ;
        RECT 1406.750 2656.460 1407.070 2656.520 ;
        RECT 1358.910 2622.460 1359.230 2622.720 ;
        RECT 1406.290 2622.460 1406.610 2622.720 ;
        RECT 1359.000 2622.040 1359.140 2622.460 ;
        RECT 1406.380 2622.040 1406.520 2622.460 ;
        RECT 1358.910 2621.780 1359.230 2622.040 ;
        RECT 1406.290 2621.780 1406.610 2622.040 ;
        RECT 1400.310 2608.380 1400.630 2608.440 ;
        RECT 1487.710 2608.380 1488.030 2608.440 ;
        RECT 1400.310 2608.240 1488.030 2608.380 ;
        RECT 1400.310 2608.180 1400.630 2608.240 ;
        RECT 1487.710 2608.180 1488.030 2608.240 ;
        RECT 998.730 2605.660 999.050 2605.720 ;
        RECT 1111.890 2605.660 1112.210 2605.720 ;
        RECT 998.730 2605.520 1112.210 2605.660 ;
        RECT 998.730 2605.460 999.050 2605.520 ;
        RECT 1111.890 2605.460 1112.210 2605.520 ;
        RECT 999.190 2605.320 999.510 2605.380 ;
        RECT 1112.810 2605.320 1113.130 2605.380 ;
        RECT 999.190 2605.180 1113.130 2605.320 ;
        RECT 999.190 2605.120 999.510 2605.180 ;
        RECT 1112.810 2605.120 1113.130 2605.180 ;
        RECT 982.170 2604.980 982.490 2605.040 ;
        RECT 1112.350 2604.980 1112.670 2605.040 ;
        RECT 982.170 2604.840 1112.670 2604.980 ;
        RECT 982.170 2604.780 982.490 2604.840 ;
        RECT 1112.350 2604.780 1112.670 2604.840 ;
        RECT 975.270 2604.640 975.590 2604.700 ;
        RECT 1113.270 2604.640 1113.590 2604.700 ;
        RECT 975.270 2604.500 1113.590 2604.640 ;
        RECT 975.270 2604.440 975.590 2604.500 ;
        RECT 1113.270 2604.440 1113.590 2604.500 ;
        RECT 1393.410 2594.780 1393.730 2594.840 ;
        RECT 1487.250 2594.780 1487.570 2594.840 ;
        RECT 1393.410 2594.640 1487.570 2594.780 ;
        RECT 1393.410 2594.580 1393.730 2594.640 ;
        RECT 1487.250 2594.580 1487.570 2594.640 ;
        RECT 533.210 2591.720 533.530 2591.780 ;
        RECT 720.890 2591.720 721.210 2591.780 ;
        RECT 533.210 2591.580 721.210 2591.720 ;
        RECT 533.210 2591.520 533.530 2591.580 ;
        RECT 720.890 2591.520 721.210 2591.580 ;
        RECT 504.690 2591.380 505.010 2591.440 ;
        RECT 762.290 2591.380 762.610 2591.440 ;
        RECT 504.690 2591.240 762.610 2591.380 ;
        RECT 504.690 2591.180 505.010 2591.240 ;
        RECT 762.290 2591.180 762.610 2591.240 ;
        RECT 981.710 2591.380 982.030 2591.440 ;
        RECT 1094.870 2591.380 1095.190 2591.440 ;
        RECT 981.710 2591.240 1095.190 2591.380 ;
        RECT 981.710 2591.180 982.030 2591.240 ;
        RECT 1094.870 2591.180 1095.190 2591.240 ;
        RECT 1028.170 2587.640 1028.490 2587.700 ;
        RECT 1033.230 2587.640 1033.550 2587.700 ;
        RECT 1028.170 2587.500 1033.550 2587.640 ;
        RECT 1028.170 2587.440 1028.490 2587.500 ;
        RECT 1033.230 2587.440 1033.550 2587.500 ;
        RECT 1413.650 2580.840 1413.970 2580.900 ;
        RECT 1487.250 2580.840 1487.570 2580.900 ;
        RECT 1413.650 2580.700 1487.570 2580.840 ;
        RECT 1413.650 2580.640 1413.970 2580.700 ;
        RECT 1487.250 2580.640 1487.570 2580.700 ;
        RECT 1358.910 2574.040 1359.230 2574.100 ;
        RECT 1358.540 2573.900 1359.230 2574.040 ;
        RECT 1358.540 2573.760 1358.680 2573.900 ;
        RECT 1358.910 2573.840 1359.230 2573.900 ;
        RECT 1406.290 2573.840 1406.610 2574.100 ;
        RECT 1358.450 2573.500 1358.770 2573.760 ;
        RECT 1406.380 2573.700 1406.520 2573.840 ;
        RECT 1406.750 2573.700 1407.070 2573.760 ;
        RECT 1406.380 2573.560 1407.070 2573.700 ;
        RECT 1406.750 2573.500 1407.070 2573.560 ;
        RECT 1358.450 2560.100 1358.770 2560.160 ;
        RECT 1358.910 2560.100 1359.230 2560.160 ;
        RECT 1358.450 2559.960 1359.230 2560.100 ;
        RECT 1358.450 2559.900 1358.770 2559.960 ;
        RECT 1358.910 2559.900 1359.230 2559.960 ;
        RECT 1406.290 2560.100 1406.610 2560.160 ;
        RECT 1406.750 2560.100 1407.070 2560.160 ;
        RECT 1406.290 2559.960 1407.070 2560.100 ;
        RECT 1406.290 2559.900 1406.610 2559.960 ;
        RECT 1406.750 2559.900 1407.070 2559.960 ;
        RECT 1405.370 2559.420 1405.690 2559.480 ;
        RECT 1406.290 2559.420 1406.610 2559.480 ;
        RECT 1405.370 2559.280 1406.610 2559.420 ;
        RECT 1405.370 2559.220 1405.690 2559.280 ;
        RECT 1406.290 2559.220 1406.610 2559.280 ;
        RECT 1468.850 2546.500 1469.170 2546.560 ;
        RECT 1483.570 2546.500 1483.890 2546.560 ;
        RECT 1468.850 2546.360 1483.890 2546.500 ;
        RECT 1468.850 2546.300 1469.170 2546.360 ;
        RECT 1483.570 2546.300 1483.890 2546.360 ;
        RECT 1357.530 2535.960 1357.850 2536.020 ;
        RECT 1358.910 2535.960 1359.230 2536.020 ;
        RECT 1357.530 2535.820 1359.230 2535.960 ;
        RECT 1357.530 2535.760 1357.850 2535.820 ;
        RECT 1358.910 2535.760 1359.230 2535.820 ;
        RECT 1485.870 2525.420 1486.190 2525.480 ;
        RECT 1490.010 2525.420 1490.330 2525.480 ;
        RECT 1485.870 2525.280 1490.330 2525.420 ;
        RECT 1485.870 2525.220 1486.190 2525.280 ;
        RECT 1490.010 2525.220 1490.330 2525.280 ;
        RECT 1357.530 2511.820 1357.850 2511.880 ;
        RECT 1357.990 2511.820 1358.310 2511.880 ;
        RECT 1357.530 2511.680 1358.310 2511.820 ;
        RECT 1357.530 2511.620 1357.850 2511.680 ;
        RECT 1357.990 2511.620 1358.310 2511.680 ;
        RECT 1405.370 2511.820 1405.690 2511.880 ;
        RECT 1406.290 2511.820 1406.610 2511.880 ;
        RECT 1405.370 2511.680 1406.610 2511.820 ;
        RECT 1405.370 2511.620 1405.690 2511.680 ;
        RECT 1406.290 2511.620 1406.610 2511.680 ;
      LAYER met1 ;
        RECT 1502.830 2510.640 1885.870 2889.200 ;
      LAYER met1 ;
        RECT 2093.990 2781.440 2094.310 2781.500 ;
        RECT 2556.290 2781.440 2556.610 2781.500 ;
        RECT 2093.990 2781.300 2556.610 2781.440 ;
        RECT 2093.990 2781.240 2094.310 2781.300 ;
        RECT 2556.290 2781.240 2556.610 2781.300 ;
        RECT 1893.890 2781.100 1894.210 2781.160 ;
        RECT 2421.970 2781.100 2422.290 2781.160 ;
        RECT 1893.890 2780.960 2422.290 2781.100 ;
        RECT 1893.890 2780.900 1894.210 2780.960 ;
        RECT 2421.970 2780.900 2422.290 2780.960 ;
      LAYER met1 ;
        RECT 2400.000 2610.640 2556.720 2760.720 ;
      LAYER met1 ;
        RECT 2528.690 2587.640 2529.010 2587.700 ;
        RECT 2534.210 2587.640 2534.530 2587.700 ;
        RECT 2528.690 2587.500 2534.530 2587.640 ;
        RECT 2528.690 2587.440 2529.010 2587.500 ;
        RECT 2534.210 2587.440 2534.530 2587.500 ;
        RECT 1494.150 2497.200 1494.470 2497.260 ;
        RECT 1512.090 2497.200 1512.410 2497.260 ;
        RECT 1494.150 2497.060 1512.410 2497.200 ;
        RECT 1494.150 2497.000 1494.470 2497.060 ;
        RECT 1512.090 2497.000 1512.410 2497.060 ;
        RECT 1621.110 2495.500 1621.430 2495.560 ;
        RECT 1895.270 2495.500 1895.590 2495.560 ;
        RECT 1621.110 2495.360 1895.590 2495.500 ;
        RECT 1621.110 2495.300 1621.430 2495.360 ;
        RECT 1895.270 2495.300 1895.590 2495.360 ;
        RECT 1494.610 2495.160 1494.930 2495.220 ;
        RECT 1552.570 2495.160 1552.890 2495.220 ;
        RECT 1494.610 2495.020 1552.890 2495.160 ;
        RECT 1494.610 2494.960 1494.930 2495.020 ;
        RECT 1552.570 2494.960 1552.890 2495.020 ;
        RECT 1607.310 2495.160 1607.630 2495.220 ;
        RECT 1894.810 2495.160 1895.130 2495.220 ;
        RECT 1607.310 2495.020 1895.130 2495.160 ;
        RECT 1607.310 2494.960 1607.630 2495.020 ;
        RECT 1894.810 2494.960 1895.130 2495.020 ;
        RECT 1501.510 2494.820 1501.830 2494.880 ;
        RECT 1559.470 2494.820 1559.790 2494.880 ;
        RECT 1501.510 2494.680 1559.790 2494.820 ;
        RECT 1501.510 2494.620 1501.830 2494.680 ;
        RECT 1559.470 2494.620 1559.790 2494.680 ;
        RECT 1586.610 2494.820 1586.930 2494.880 ;
        RECT 1887.910 2494.820 1888.230 2494.880 ;
        RECT 1586.610 2494.680 1888.230 2494.820 ;
        RECT 1586.610 2494.620 1586.930 2494.680 ;
        RECT 1887.910 2494.620 1888.230 2494.680 ;
        RECT 1545.210 2494.480 1545.530 2494.540 ;
        RECT 1887.450 2494.480 1887.770 2494.540 ;
        RECT 1545.210 2494.340 1887.770 2494.480 ;
        RECT 1545.210 2494.280 1545.530 2494.340 ;
        RECT 1887.450 2494.280 1887.770 2494.340 ;
        RECT 1876.410 2494.140 1876.730 2494.200 ;
        RECT 2394.370 2494.140 2394.690 2494.200 ;
        RECT 1876.410 2494.000 2394.690 2494.140 ;
        RECT 1876.410 2493.940 1876.730 2494.000 ;
        RECT 2394.370 2493.940 2394.690 2494.000 ;
        RECT 1679.990 2489.720 1680.310 2489.780 ;
        RECT 1746.690 2489.720 1747.010 2489.780 ;
        RECT 1679.990 2489.580 1747.010 2489.720 ;
        RECT 1679.990 2489.520 1680.310 2489.580 ;
        RECT 1746.690 2489.520 1747.010 2489.580 ;
        RECT 1593.510 2489.380 1593.830 2489.440 ;
        RECT 1778.890 2489.380 1779.210 2489.440 ;
        RECT 1593.510 2489.240 1779.210 2489.380 ;
        RECT 1593.510 2489.180 1593.830 2489.240 ;
        RECT 1778.890 2489.180 1779.210 2489.240 ;
        RECT 1600.410 2489.040 1600.730 2489.100 ;
        RECT 1789.930 2489.040 1790.250 2489.100 ;
        RECT 1600.410 2488.900 1790.250 2489.040 ;
        RECT 1600.410 2488.840 1600.730 2488.900 ;
        RECT 1789.930 2488.840 1790.250 2488.900 ;
        RECT 1421.010 2488.700 1421.330 2488.760 ;
        RECT 1842.370 2488.700 1842.690 2488.760 ;
        RECT 1421.010 2488.560 1842.690 2488.700 ;
        RECT 1421.010 2488.500 1421.330 2488.560 ;
        RECT 1842.370 2488.500 1842.690 2488.560 ;
        RECT 1455.050 2488.360 1455.370 2488.420 ;
        RECT 1885.610 2488.360 1885.930 2488.420 ;
        RECT 1455.050 2488.220 1885.930 2488.360 ;
        RECT 1455.050 2488.160 1455.370 2488.220 ;
        RECT 1885.610 2488.160 1885.930 2488.220 ;
        RECT 1405.370 2488.020 1405.690 2488.080 ;
        RECT 1406.290 2488.020 1406.610 2488.080 ;
        RECT 1405.370 2487.880 1406.610 2488.020 ;
        RECT 1405.370 2487.820 1405.690 2487.880 ;
        RECT 1406.290 2487.820 1406.610 2487.880 ;
        RECT 1420.550 2488.020 1420.870 2488.080 ;
        RECT 1874.570 2488.020 1874.890 2488.080 ;
        RECT 1420.550 2487.880 1874.890 2488.020 ;
        RECT 1420.550 2487.820 1420.870 2487.880 ;
        RECT 1874.570 2487.820 1874.890 2487.880 ;
        RECT 1448.150 2487.000 1448.470 2487.060 ;
        RECT 1832.250 2487.000 1832.570 2487.060 ;
        RECT 1448.150 2486.860 1832.570 2487.000 ;
        RECT 1448.150 2486.800 1448.470 2486.860 ;
        RECT 1832.250 2486.800 1832.570 2486.860 ;
        RECT 1427.910 2486.660 1428.230 2486.720 ;
        RECT 1725.530 2486.660 1725.850 2486.720 ;
        RECT 1427.910 2486.520 1725.850 2486.660 ;
        RECT 1427.910 2486.460 1428.230 2486.520 ;
        RECT 1725.530 2486.460 1725.850 2486.520 ;
        RECT 1461.950 2486.320 1462.270 2486.380 ;
        RECT 1757.730 2486.320 1758.050 2486.380 ;
        RECT 1461.950 2486.180 1758.050 2486.320 ;
        RECT 1461.950 2486.120 1462.270 2486.180 ;
        RECT 1757.730 2486.120 1758.050 2486.180 ;
        RECT 1379.150 2485.980 1379.470 2486.040 ;
        RECT 1534.170 2485.980 1534.490 2486.040 ;
        RECT 1379.150 2485.840 1534.490 2485.980 ;
        RECT 1379.150 2485.780 1379.470 2485.840 ;
        RECT 1534.170 2485.780 1534.490 2485.840 ;
        RECT 1535.090 2485.980 1535.410 2486.040 ;
        RECT 1811.090 2485.980 1811.410 2486.040 ;
        RECT 1535.090 2485.840 1811.410 2485.980 ;
        RECT 1535.090 2485.780 1535.410 2485.840 ;
        RECT 1811.090 2485.780 1811.410 2485.840 ;
        RECT 1386.510 2485.640 1386.830 2485.700 ;
        RECT 1587.530 2485.640 1587.850 2485.700 ;
        RECT 1386.510 2485.500 1587.850 2485.640 ;
        RECT 1386.510 2485.440 1386.830 2485.500 ;
        RECT 1587.530 2485.440 1587.850 2485.500 ;
        RECT 1673.090 2485.640 1673.410 2485.700 ;
        RECT 1715.410 2485.640 1715.730 2485.700 ;
        RECT 1673.090 2485.500 1715.730 2485.640 ;
        RECT 1673.090 2485.440 1673.410 2485.500 ;
        RECT 1715.410 2485.440 1715.730 2485.500 ;
        RECT 1441.250 2485.300 1441.570 2485.360 ;
        RECT 1608.690 2485.300 1609.010 2485.360 ;
        RECT 1441.250 2485.160 1609.010 2485.300 ;
        RECT 1441.250 2485.100 1441.570 2485.160 ;
        RECT 1608.690 2485.100 1609.010 2485.160 ;
        RECT 1537.850 2484.960 1538.170 2485.020 ;
        RECT 1575.110 2484.960 1575.430 2485.020 ;
        RECT 1537.850 2484.820 1575.430 2484.960 ;
        RECT 1537.850 2484.760 1538.170 2484.820 ;
        RECT 1575.110 2484.760 1575.430 2484.820 ;
        RECT 1576.490 2484.960 1576.810 2485.020 ;
        RECT 1619.730 2484.960 1620.050 2485.020 ;
        RECT 1576.490 2484.820 1620.050 2484.960 ;
        RECT 1576.490 2484.760 1576.810 2484.820 ;
        RECT 1619.730 2484.760 1620.050 2484.820 ;
        RECT 1524.050 2484.620 1524.370 2484.680 ;
        RECT 1546.590 2484.620 1546.910 2484.680 ;
        RECT 1524.050 2484.480 1546.910 2484.620 ;
        RECT 1524.050 2484.420 1524.370 2484.480 ;
        RECT 1546.590 2484.420 1546.910 2484.480 ;
        RECT 1624.790 2484.620 1625.110 2484.680 ;
        RECT 1640.890 2484.620 1641.210 2484.680 ;
        RECT 1624.790 2484.480 1641.210 2484.620 ;
        RECT 1624.790 2484.420 1625.110 2484.480 ;
        RECT 1640.890 2484.420 1641.210 2484.480 ;
        RECT 1659.290 2484.620 1659.610 2484.680 ;
        RECT 1683.210 2484.620 1683.530 2484.680 ;
        RECT 1659.290 2484.480 1683.530 2484.620 ;
        RECT 1659.290 2484.420 1659.610 2484.480 ;
        RECT 1683.210 2484.420 1683.530 2484.480 ;
        RECT 1485.870 2477.480 1486.190 2477.540 ;
        RECT 1490.010 2477.480 1490.330 2477.540 ;
        RECT 1485.870 2477.340 1490.330 2477.480 ;
        RECT 1485.870 2477.280 1486.190 2477.340 ;
        RECT 1490.010 2477.280 1490.330 2477.340 ;
        RECT 1544.290 2463.880 1544.610 2463.940 ;
        RECT 1545.210 2463.880 1545.530 2463.940 ;
        RECT 1544.290 2463.740 1545.530 2463.880 ;
        RECT 1544.290 2463.680 1544.610 2463.740 ;
        RECT 1545.210 2463.680 1545.530 2463.740 ;
        RECT 1357.530 2439.060 1357.850 2439.120 ;
        RECT 1358.910 2439.060 1359.230 2439.120 ;
        RECT 1357.530 2438.920 1359.230 2439.060 ;
        RECT 1357.530 2438.860 1357.850 2438.920 ;
        RECT 1358.910 2438.860 1359.230 2438.920 ;
        RECT 1406.290 2429.340 1406.610 2429.600 ;
        RECT 1406.380 2428.920 1406.520 2429.340 ;
        RECT 1406.290 2428.660 1406.610 2428.920 ;
        RECT 1357.530 2415.600 1357.850 2415.660 ;
        RECT 1358.450 2415.600 1358.770 2415.660 ;
        RECT 1357.530 2415.460 1358.770 2415.600 ;
        RECT 1357.530 2415.400 1357.850 2415.460 ;
        RECT 1358.450 2415.400 1358.770 2415.460 ;
        RECT 1358.450 2414.920 1358.770 2414.980 ;
        RECT 1358.910 2414.920 1359.230 2414.980 ;
        RECT 1358.450 2414.780 1359.230 2414.920 ;
        RECT 1358.450 2414.720 1358.770 2414.780 ;
        RECT 1358.910 2414.720 1359.230 2414.780 ;
        RECT 1543.830 2408.120 1544.150 2408.180 ;
        RECT 1544.290 2408.120 1544.610 2408.180 ;
        RECT 1543.830 2407.980 1544.610 2408.120 ;
        RECT 1543.830 2407.920 1544.150 2407.980 ;
        RECT 1544.290 2407.920 1544.610 2407.980 ;
        RECT 1358.910 2380.580 1359.230 2380.640 ;
        RECT 1358.540 2380.440 1359.230 2380.580 ;
        RECT 1358.540 2380.300 1358.680 2380.440 ;
        RECT 1358.910 2380.380 1359.230 2380.440 ;
        RECT 1406.290 2380.580 1406.610 2380.640 ;
        RECT 1406.750 2380.580 1407.070 2380.640 ;
        RECT 1406.290 2380.440 1407.070 2380.580 ;
        RECT 1406.290 2380.380 1406.610 2380.440 ;
        RECT 1406.750 2380.380 1407.070 2380.440 ;
        RECT 1358.450 2380.040 1358.770 2380.300 ;
        RECT 1406.290 2366.980 1406.610 2367.040 ;
        RECT 1406.750 2366.980 1407.070 2367.040 ;
        RECT 1406.290 2366.840 1407.070 2366.980 ;
        RECT 1406.290 2366.780 1406.610 2366.840 ;
        RECT 1406.750 2366.780 1407.070 2366.840 ;
        RECT 1544.290 2366.780 1544.610 2367.040 ;
        RECT 1543.830 2366.640 1544.150 2366.700 ;
        RECT 1544.380 2366.640 1544.520 2366.780 ;
        RECT 1543.830 2366.500 1544.520 2366.640 ;
        RECT 1543.830 2366.440 1544.150 2366.500 ;
        RECT 1357.530 2342.500 1357.850 2342.560 ;
        RECT 1358.910 2342.500 1359.230 2342.560 ;
        RECT 1357.530 2342.360 1359.230 2342.500 ;
        RECT 1357.530 2342.300 1357.850 2342.360 ;
        RECT 1358.910 2342.300 1359.230 2342.360 ;
        RECT 1406.290 2332.440 1406.610 2332.700 ;
        RECT 1406.380 2332.020 1406.520 2332.440 ;
        RECT 1406.290 2331.760 1406.610 2332.020 ;
        RECT 1357.530 2319.040 1357.850 2319.100 ;
        RECT 1358.450 2319.040 1358.770 2319.100 ;
        RECT 1357.530 2318.900 1358.770 2319.040 ;
        RECT 1357.530 2318.840 1357.850 2318.900 ;
        RECT 1358.450 2318.840 1358.770 2318.900 ;
        RECT 1358.450 2318.360 1358.770 2318.420 ;
        RECT 1358.910 2318.360 1359.230 2318.420 ;
        RECT 1358.450 2318.220 1359.230 2318.360 ;
        RECT 1358.450 2318.160 1358.770 2318.220 ;
        RECT 1358.910 2318.160 1359.230 2318.220 ;
        RECT 1534.170 2318.360 1534.490 2318.420 ;
        RECT 1535.090 2318.360 1535.410 2318.420 ;
        RECT 1534.170 2318.220 1535.410 2318.360 ;
        RECT 1534.170 2318.160 1534.490 2318.220 ;
        RECT 1535.090 2318.160 1535.410 2318.220 ;
        RECT 1405.370 2294.220 1405.690 2294.280 ;
        RECT 1406.290 2294.220 1406.610 2294.280 ;
        RECT 1405.370 2294.080 1406.610 2294.220 ;
        RECT 1405.370 2294.020 1405.690 2294.080 ;
        RECT 1406.290 2294.020 1406.610 2294.080 ;
        RECT 1358.910 2284.020 1359.230 2284.080 ;
        RECT 1358.540 2283.880 1359.230 2284.020 ;
        RECT 1358.540 2283.740 1358.680 2283.880 ;
        RECT 1358.910 2283.820 1359.230 2283.880 ;
        RECT 1358.450 2283.480 1358.770 2283.740 ;
        RECT 1357.530 2245.940 1357.850 2246.000 ;
        RECT 1358.910 2245.940 1359.230 2246.000 ;
        RECT 1357.530 2245.800 1359.230 2245.940 ;
        RECT 1357.530 2245.740 1357.850 2245.800 ;
        RECT 1358.910 2245.740 1359.230 2245.800 ;
        RECT 1406.290 2235.880 1406.610 2236.140 ;
        RECT 1406.380 2235.460 1406.520 2235.880 ;
        RECT 1406.290 2235.200 1406.610 2235.460 ;
        RECT 1357.530 2222.480 1357.850 2222.540 ;
        RECT 1358.450 2222.480 1358.770 2222.540 ;
        RECT 1357.530 2222.340 1358.770 2222.480 ;
        RECT 1357.530 2222.280 1357.850 2222.340 ;
        RECT 1358.450 2222.280 1358.770 2222.340 ;
        RECT 1358.450 2221.800 1358.770 2221.860 ;
        RECT 1358.910 2221.800 1359.230 2221.860 ;
        RECT 1358.450 2221.660 1359.230 2221.800 ;
        RECT 1358.450 2221.600 1358.770 2221.660 ;
        RECT 1358.910 2221.600 1359.230 2221.660 ;
        RECT 1534.170 2221.800 1534.490 2221.860 ;
        RECT 1535.090 2221.800 1535.410 2221.860 ;
        RECT 1534.170 2221.660 1535.410 2221.800 ;
        RECT 1534.170 2221.600 1534.490 2221.660 ;
        RECT 1535.090 2221.600 1535.410 2221.660 ;
        RECT 1543.830 2215.000 1544.150 2215.060 ;
        RECT 1544.290 2215.000 1544.610 2215.060 ;
        RECT 1543.830 2214.860 1544.610 2215.000 ;
        RECT 1543.830 2214.800 1544.150 2214.860 ;
        RECT 1544.290 2214.800 1544.610 2214.860 ;
        RECT 1405.370 2197.660 1405.690 2197.720 ;
        RECT 1406.290 2197.660 1406.610 2197.720 ;
        RECT 1405.370 2197.520 1406.610 2197.660 ;
        RECT 1405.370 2197.460 1405.690 2197.520 ;
        RECT 1406.290 2197.460 1406.610 2197.520 ;
        RECT 1358.910 2187.460 1359.230 2187.520 ;
        RECT 1358.540 2187.320 1359.230 2187.460 ;
        RECT 1358.540 2187.180 1358.680 2187.320 ;
        RECT 1358.910 2187.260 1359.230 2187.320 ;
        RECT 1358.450 2186.920 1358.770 2187.180 ;
        RECT 1534.170 2173.860 1534.490 2173.920 ;
        RECT 1535.090 2173.860 1535.410 2173.920 ;
        RECT 1534.170 2173.720 1535.410 2173.860 ;
        RECT 1534.170 2173.660 1534.490 2173.720 ;
        RECT 1535.090 2173.660 1535.410 2173.720 ;
        RECT 1357.530 2149.380 1357.850 2149.440 ;
        RECT 1358.910 2149.380 1359.230 2149.440 ;
        RECT 1357.530 2149.240 1359.230 2149.380 ;
        RECT 1357.530 2149.180 1357.850 2149.240 ;
        RECT 1358.910 2149.180 1359.230 2149.240 ;
        RECT 1406.290 2139.320 1406.610 2139.580 ;
        RECT 1406.380 2138.900 1406.520 2139.320 ;
        RECT 1406.290 2138.640 1406.610 2138.900 ;
        RECT 1357.530 2125.920 1357.850 2125.980 ;
        RECT 1358.450 2125.920 1358.770 2125.980 ;
        RECT 1357.530 2125.780 1358.770 2125.920 ;
        RECT 1357.530 2125.720 1357.850 2125.780 ;
        RECT 1358.450 2125.720 1358.770 2125.780 ;
        RECT 1358.450 2125.240 1358.770 2125.300 ;
        RECT 1358.910 2125.240 1359.230 2125.300 ;
        RECT 1358.450 2125.100 1359.230 2125.240 ;
        RECT 1358.450 2125.040 1358.770 2125.100 ;
        RECT 1358.910 2125.040 1359.230 2125.100 ;
        RECT 1543.830 2118.440 1544.150 2118.500 ;
        RECT 1544.290 2118.440 1544.610 2118.500 ;
        RECT 1543.830 2118.300 1544.610 2118.440 ;
        RECT 1543.830 2118.240 1544.150 2118.300 ;
        RECT 1544.290 2118.240 1544.610 2118.300 ;
        RECT 1406.290 2118.100 1406.610 2118.160 ;
        RECT 1407.670 2118.100 1407.990 2118.160 ;
        RECT 1406.290 2117.960 1407.990 2118.100 ;
        RECT 1406.290 2117.900 1406.610 2117.960 ;
        RECT 1407.670 2117.900 1407.990 2117.960 ;
        RECT 1408.130 2069.820 1408.450 2069.880 ;
        RECT 1409.050 2069.820 1409.370 2069.880 ;
        RECT 1408.130 2069.680 1409.370 2069.820 ;
        RECT 1408.130 2069.620 1408.450 2069.680 ;
        RECT 1409.050 2069.620 1409.370 2069.680 ;
        RECT 1272.890 2055.540 1273.210 2055.600 ;
        RECT 1347.870 2055.540 1348.190 2055.600 ;
        RECT 1272.890 2055.400 1348.190 2055.540 ;
        RECT 1272.890 2055.340 1273.210 2055.400 ;
        RECT 1347.870 2055.340 1348.190 2055.400 ;
        RECT 1273.350 2055.200 1273.670 2055.260 ;
        RECT 1331.770 2055.200 1332.090 2055.260 ;
        RECT 1273.350 2055.060 1332.090 2055.200 ;
        RECT 1273.350 2055.000 1273.670 2055.060 ;
        RECT 1331.770 2055.000 1332.090 2055.060 ;
        RECT 1293.590 2054.860 1293.910 2054.920 ;
        RECT 1334.990 2054.860 1335.310 2054.920 ;
        RECT 1293.590 2054.720 1335.310 2054.860 ;
        RECT 1293.590 2054.660 1293.910 2054.720 ;
        RECT 1334.990 2054.660 1335.310 2054.720 ;
        RECT 1130.750 2054.520 1131.070 2054.580 ;
        RECT 1353.850 2054.520 1354.170 2054.580 ;
        RECT 1130.750 2054.380 1354.170 2054.520 ;
        RECT 1130.750 2054.320 1131.070 2054.380 ;
        RECT 1353.850 2054.320 1354.170 2054.380 ;
        RECT 1116.950 2054.180 1117.270 2054.240 ;
        RECT 1332.690 2054.180 1333.010 2054.240 ;
        RECT 1116.950 2054.040 1333.010 2054.180 ;
        RECT 1116.950 2053.980 1117.270 2054.040 ;
        RECT 1332.690 2053.980 1333.010 2054.040 ;
        RECT 1230.110 2053.840 1230.430 2053.900 ;
        RECT 1353.390 2053.840 1353.710 2053.900 ;
        RECT 1230.110 2053.700 1353.710 2053.840 ;
        RECT 1230.110 2053.640 1230.430 2053.700 ;
        RECT 1353.390 2053.640 1353.710 2053.700 ;
        RECT 1059.910 2053.500 1060.230 2053.560 ;
        RECT 1293.590 2053.500 1293.910 2053.560 ;
        RECT 1059.910 2053.360 1293.910 2053.500 ;
        RECT 1059.910 2053.300 1060.230 2053.360 ;
        RECT 1293.590 2053.300 1293.910 2053.360 ;
        RECT 1294.050 2053.500 1294.370 2053.560 ;
        RECT 1333.610 2053.500 1333.930 2053.560 ;
        RECT 1294.050 2053.360 1333.930 2053.500 ;
        RECT 1294.050 2053.300 1294.370 2053.360 ;
        RECT 1333.610 2053.300 1333.930 2053.360 ;
        RECT 1031.390 2053.160 1031.710 2053.220 ;
        RECT 1352.470 2053.160 1352.790 2053.220 ;
        RECT 1031.390 2053.020 1352.790 2053.160 ;
        RECT 1031.390 2052.960 1031.710 2053.020 ;
        RECT 1352.470 2052.960 1352.790 2053.020 ;
        RECT 1016.670 2052.820 1016.990 2052.880 ;
        RECT 1272.890 2052.820 1273.210 2052.880 ;
        RECT 1016.670 2052.680 1273.210 2052.820 ;
        RECT 1016.670 2052.620 1016.990 2052.680 ;
        RECT 1272.890 2052.620 1273.210 2052.680 ;
        RECT 1286.230 2052.820 1286.550 2052.880 ;
        RECT 1346.030 2052.820 1346.350 2052.880 ;
        RECT 1286.230 2052.680 1346.350 2052.820 ;
        RECT 1286.230 2052.620 1286.550 2052.680 ;
        RECT 1346.030 2052.620 1346.350 2052.680 ;
        RECT 1201.590 2052.480 1201.910 2052.540 ;
        RECT 1332.230 2052.480 1332.550 2052.540 ;
        RECT 1201.590 2052.340 1332.550 2052.480 ;
        RECT 1201.590 2052.280 1201.910 2052.340 ;
        RECT 1332.230 2052.280 1332.550 2052.340 ;
        RECT 1187.790 2052.140 1188.110 2052.200 ;
        RECT 1294.050 2052.140 1294.370 2052.200 ;
        RECT 1187.790 2052.000 1294.370 2052.140 ;
        RECT 1187.790 2051.940 1188.110 2052.000 ;
        RECT 1294.050 2051.940 1294.370 2052.000 ;
        RECT 1301.870 2052.140 1302.190 2052.200 ;
        RECT 1336.370 2052.140 1336.690 2052.200 ;
        RECT 1301.870 2052.000 1336.690 2052.140 ;
        RECT 1301.870 2051.940 1302.190 2052.000 ;
        RECT 1336.370 2051.940 1336.690 2052.000 ;
        RECT 1173.070 2051.800 1173.390 2051.860 ;
        RECT 1286.230 2051.800 1286.550 2051.860 ;
        RECT 1173.070 2051.660 1286.550 2051.800 ;
        RECT 1173.070 2051.600 1173.390 2051.660 ;
        RECT 1286.230 2051.600 1286.550 2051.660 ;
        RECT 1286.690 2051.800 1287.010 2051.860 ;
        RECT 1346.490 2051.800 1346.810 2051.860 ;
        RECT 1286.690 2051.660 1346.810 2051.800 ;
        RECT 1286.690 2051.600 1287.010 2051.660 ;
        RECT 1346.490 2051.600 1346.810 2051.660 ;
        RECT 1159.270 2051.460 1159.590 2051.520 ;
        RECT 1354.310 2051.460 1354.630 2051.520 ;
        RECT 1159.270 2051.320 1354.630 2051.460 ;
        RECT 1159.270 2051.260 1159.590 2051.320 ;
        RECT 1354.310 2051.260 1354.630 2051.320 ;
        RECT 1144.550 2051.120 1144.870 2051.180 ;
        RECT 1352.930 2051.120 1353.250 2051.180 ;
        RECT 1144.550 2050.980 1353.250 2051.120 ;
        RECT 1144.550 2050.920 1144.870 2050.980 ;
        RECT 1352.930 2050.920 1353.250 2050.980 ;
        RECT 1000.110 2050.780 1000.430 2050.840 ;
        RECT 1088.430 2050.780 1088.750 2050.840 ;
        RECT 1000.110 2050.640 1088.750 2050.780 ;
        RECT 1000.110 2050.580 1000.430 2050.640 ;
        RECT 1088.430 2050.580 1088.750 2050.640 ;
        RECT 1258.630 2050.780 1258.950 2050.840 ;
        RECT 1286.690 2050.780 1287.010 2050.840 ;
        RECT 1258.630 2050.640 1287.010 2050.780 ;
        RECT 1258.630 2050.580 1258.950 2050.640 ;
        RECT 1286.690 2050.580 1287.010 2050.640 ;
        RECT 1287.150 2050.780 1287.470 2050.840 ;
        RECT 1346.950 2050.780 1347.270 2050.840 ;
        RECT 1287.150 2050.640 1347.270 2050.780 ;
        RECT 1287.150 2050.580 1287.470 2050.640 ;
        RECT 1346.950 2050.580 1347.270 2050.640 ;
        RECT 977.570 2050.440 977.890 2050.500 ;
        RECT 1102.230 2050.440 1102.550 2050.500 ;
        RECT 1347.410 2050.440 1347.730 2050.500 ;
        RECT 977.570 2050.300 1102.550 2050.440 ;
        RECT 977.570 2050.240 977.890 2050.300 ;
        RECT 1102.230 2050.240 1102.550 2050.300 ;
        RECT 1293.220 2050.300 1347.730 2050.440 ;
        RECT 978.030 2050.100 978.350 2050.160 ;
        RECT 1073.710 2050.100 1074.030 2050.160 ;
        RECT 978.030 2049.960 1074.030 2050.100 ;
        RECT 978.030 2049.900 978.350 2049.960 ;
        RECT 1073.710 2049.900 1074.030 2049.960 ;
        RECT 1244.830 2050.100 1245.150 2050.160 ;
        RECT 1293.220 2050.100 1293.360 2050.300 ;
        RECT 1347.410 2050.240 1347.730 2050.300 ;
        RECT 1333.150 2050.100 1333.470 2050.160 ;
        RECT 1244.830 2049.960 1293.360 2050.100 ;
        RECT 1293.680 2049.960 1333.470 2050.100 ;
        RECT 1244.830 2049.900 1245.150 2049.960 ;
        RECT 999.650 2049.760 999.970 2049.820 ;
        RECT 1045.190 2049.760 1045.510 2049.820 ;
        RECT 999.650 2049.620 1045.510 2049.760 ;
        RECT 999.650 2049.560 999.970 2049.620 ;
        RECT 1045.190 2049.560 1045.510 2049.620 ;
        RECT 1216.310 2049.760 1216.630 2049.820 ;
        RECT 1293.680 2049.760 1293.820 2049.960 ;
        RECT 1333.150 2049.900 1333.470 2049.960 ;
        RECT 1216.310 2049.620 1293.820 2049.760 ;
        RECT 1315.670 2049.760 1315.990 2049.820 ;
        RECT 1336.830 2049.760 1337.150 2049.820 ;
        RECT 1315.670 2049.620 1337.150 2049.760 ;
        RECT 1216.310 2049.560 1216.630 2049.620 ;
        RECT 1315.670 2049.560 1315.990 2049.620 ;
        RECT 1336.830 2049.560 1337.150 2049.620 ;
        RECT 984.930 2049.420 985.250 2049.480 ;
        RECT 1002.870 2049.420 1003.190 2049.480 ;
        RECT 984.930 2049.280 1003.190 2049.420 ;
        RECT 984.930 2049.220 985.250 2049.280 ;
        RECT 1002.870 2049.220 1003.190 2049.280 ;
        RECT 1329.470 2049.420 1329.790 2049.480 ;
        RECT 1343.730 2049.420 1344.050 2049.480 ;
        RECT 1329.470 2049.280 1344.050 2049.420 ;
        RECT 1329.470 2049.220 1329.790 2049.280 ;
        RECT 1343.730 2049.220 1344.050 2049.280 ;
        RECT 984.010 2048.400 984.330 2048.460 ;
        RECT 1014.370 2048.400 1014.690 2048.460 ;
        RECT 984.010 2048.260 1014.690 2048.400 ;
        RECT 984.010 2048.200 984.330 2048.260 ;
        RECT 1014.370 2048.200 1014.690 2048.260 ;
        RECT 984.470 2048.060 984.790 2048.120 ;
        RECT 1028.170 2048.060 1028.490 2048.120 ;
        RECT 984.470 2047.920 1028.490 2048.060 ;
        RECT 984.470 2047.860 984.790 2047.920 ;
        RECT 1028.170 2047.860 1028.490 2047.920 ;
        RECT 977.110 2047.720 977.430 2047.780 ;
        RECT 1048.870 2047.720 1049.190 2047.780 ;
        RECT 977.110 2047.580 1049.190 2047.720 ;
        RECT 977.110 2047.520 977.430 2047.580 ;
        RECT 1048.870 2047.520 1049.190 2047.580 ;
        RECT 975.730 2047.380 976.050 2047.440 ;
        RECT 1062.670 2047.380 1062.990 2047.440 ;
        RECT 975.730 2047.240 1062.990 2047.380 ;
        RECT 975.730 2047.180 976.050 2047.240 ;
        RECT 1062.670 2047.180 1062.990 2047.240 ;
        RECT 983.090 2047.040 983.410 2047.100 ;
        RECT 1076.470 2047.040 1076.790 2047.100 ;
        RECT 983.090 2046.900 1076.790 2047.040 ;
        RECT 983.090 2046.840 983.410 2046.900 ;
        RECT 1076.470 2046.840 1076.790 2046.900 ;
        RECT 983.550 2046.700 983.870 2046.760 ;
        RECT 1097.170 2046.700 1097.490 2046.760 ;
        RECT 983.550 2046.560 1097.490 2046.700 ;
        RECT 983.550 2046.500 983.870 2046.560 ;
        RECT 1097.170 2046.500 1097.490 2046.560 ;
        RECT 976.650 2046.360 976.970 2046.420 ;
        RECT 1097.630 2046.360 1097.950 2046.420 ;
        RECT 976.650 2046.220 1097.950 2046.360 ;
        RECT 976.650 2046.160 976.970 2046.220 ;
        RECT 1097.630 2046.160 1097.950 2046.220 ;
        RECT 982.630 2046.020 982.950 2046.080 ;
        RECT 1110.970 2046.020 1111.290 2046.080 ;
        RECT 982.630 2045.880 1111.290 2046.020 ;
        RECT 982.630 2045.820 982.950 2045.880 ;
        RECT 1110.970 2045.820 1111.290 2045.880 ;
        RECT 976.190 2045.680 976.510 2045.740 ;
        RECT 1111.430 2045.680 1111.750 2045.740 ;
        RECT 976.190 2045.540 1111.750 2045.680 ;
        RECT 976.190 2045.480 976.510 2045.540 ;
        RECT 1111.430 2045.480 1111.750 2045.540 ;
        RECT 1357.990 2042.620 1358.310 2042.680 ;
        RECT 1359.830 2042.620 1360.150 2042.680 ;
        RECT 1357.990 2042.480 1360.150 2042.620 ;
        RECT 1357.990 2042.420 1358.310 2042.480 ;
        RECT 1359.830 2042.420 1360.150 2042.480 ;
        RECT 529.990 1988.560 530.310 1988.620 ;
        RECT 650.510 1988.560 650.830 1988.620 ;
        RECT 529.990 1988.420 650.830 1988.560 ;
        RECT 529.990 1988.360 530.310 1988.420 ;
        RECT 650.510 1988.360 650.830 1988.420 ;
        RECT 579.210 1987.540 579.530 1987.600 ;
        RECT 638.090 1987.540 638.410 1987.600 ;
        RECT 579.210 1987.400 638.410 1987.540 ;
        RECT 579.210 1987.340 579.530 1987.400 ;
        RECT 638.090 1987.340 638.410 1987.400 ;
        RECT 420.510 1978.700 420.830 1978.760 ;
        RECT 419.680 1978.560 420.830 1978.700 ;
        RECT 419.680 1977.680 419.820 1978.560 ;
        RECT 420.510 1978.500 420.830 1978.560 ;
        RECT 420.050 1978.160 420.370 1978.420 ;
        RECT 420.140 1978.020 420.280 1978.160 ;
        RECT 843.250 1978.020 843.570 1978.080 ;
        RECT 420.140 1977.880 843.570 1978.020 ;
        RECT 843.250 1977.820 843.570 1977.880 ;
        RECT 897.530 1977.680 897.850 1977.740 ;
        RECT 419.680 1977.540 897.850 1977.680 ;
        RECT 897.530 1977.480 897.850 1977.540 ;
      LAYER met1 ;
        RECT 362.830 1704.460 628.110 1977.400 ;
      LAYER met1 ;
        RECT 998.270 1713.840 998.590 1713.900 ;
        RECT 1001.030 1713.840 1001.350 1713.900 ;
        RECT 998.270 1713.700 1001.350 1713.840 ;
        RECT 998.270 1713.640 998.590 1713.700 ;
        RECT 1001.030 1713.640 1001.350 1713.700 ;
      LAYER met1 ;
        RECT 1002.830 1710.640 1329.750 2032.080 ;
      LAYER met1 ;
        RECT 1543.830 2021.880 1544.150 2021.940 ;
        RECT 1544.290 2021.880 1544.610 2021.940 ;
        RECT 1543.830 2021.740 1544.610 2021.880 ;
        RECT 1543.830 2021.680 1544.150 2021.740 ;
        RECT 1544.290 2021.680 1544.610 2021.740 ;
        RECT 1357.990 1994.000 1358.310 1994.060 ;
        RECT 1358.910 1994.000 1359.230 1994.060 ;
        RECT 1357.990 1993.860 1359.230 1994.000 ;
        RECT 1357.990 1993.800 1358.310 1993.860 ;
        RECT 1358.910 1993.800 1359.230 1993.860 ;
        RECT 1542.910 1972.920 1543.230 1972.980 ;
        RECT 1544.290 1972.920 1544.610 1972.980 ;
        RECT 1542.910 1972.780 1544.610 1972.920 ;
        RECT 1542.910 1972.720 1543.230 1972.780 ;
        RECT 1544.290 1972.720 1544.610 1972.780 ;
        RECT 2294.090 1947.080 2294.410 1947.140 ;
        RECT 2379.190 1947.080 2379.510 1947.140 ;
        RECT 2294.090 1946.940 2379.510 1947.080 ;
        RECT 2294.090 1946.880 2294.410 1946.940 ;
        RECT 2379.190 1946.880 2379.510 1946.940 ;
        RECT 2083.410 1946.740 2083.730 1946.800 ;
        RECT 2321.230 1946.740 2321.550 1946.800 ;
        RECT 2083.410 1946.600 2321.550 1946.740 ;
        RECT 2083.410 1946.540 2083.730 1946.600 ;
        RECT 2321.230 1946.540 2321.550 1946.600 ;
        RECT 2090.310 1946.400 2090.630 1946.460 ;
        RECT 2437.150 1946.400 2437.470 1946.460 ;
        RECT 2090.310 1946.260 2437.470 1946.400 ;
        RECT 2090.310 1946.200 2090.630 1946.260 ;
        RECT 2437.150 1946.200 2437.470 1946.260 ;
        RECT 2082.950 1946.060 2083.270 1946.120 ;
        RECT 2495.110 1946.060 2495.430 1946.120 ;
        RECT 2082.950 1945.920 2495.430 1946.060 ;
        RECT 2082.950 1945.860 2083.270 1945.920 ;
        RECT 2495.110 1945.860 2495.430 1945.920 ;
        RECT 1357.530 1945.720 1357.850 1945.780 ;
        RECT 1357.990 1945.720 1358.310 1945.780 ;
        RECT 1357.530 1945.580 1358.310 1945.720 ;
        RECT 1357.530 1945.520 1357.850 1945.580 ;
        RECT 1357.990 1945.520 1358.310 1945.580 ;
        RECT 1485.870 1945.720 1486.190 1945.780 ;
        RECT 1490.010 1945.720 1490.330 1945.780 ;
        RECT 1485.870 1945.580 1490.330 1945.720 ;
        RECT 1485.870 1945.520 1486.190 1945.580 ;
        RECT 1490.010 1945.520 1490.330 1945.580 ;
        RECT 1406.750 1931.780 1407.070 1931.840 ;
        RECT 1407.670 1931.780 1407.990 1931.840 ;
        RECT 1406.750 1931.640 1407.990 1931.780 ;
        RECT 1406.750 1931.580 1407.070 1931.640 ;
        RECT 1407.670 1931.580 1407.990 1931.640 ;
        RECT 1534.170 1931.780 1534.490 1931.840 ;
        RECT 1535.090 1931.780 1535.410 1931.840 ;
        RECT 1534.170 1931.640 1535.410 1931.780 ;
        RECT 1534.170 1931.580 1534.490 1931.640 ;
        RECT 1535.090 1931.580 1535.410 1931.640 ;
        RECT 1724.610 1928.720 1724.930 1928.780 ;
        RECT 2044.310 1928.720 2044.630 1928.780 ;
        RECT 1724.610 1928.580 2044.630 1928.720 ;
        RECT 1724.610 1928.520 1724.930 1928.580 ;
        RECT 2044.310 1928.520 2044.630 1928.580 ;
        RECT 1828.110 1928.040 1828.430 1928.100 ;
        RECT 1964.270 1928.040 1964.590 1928.100 ;
        RECT 1828.110 1927.900 1964.590 1928.040 ;
        RECT 1828.110 1927.840 1828.430 1927.900 ;
        RECT 1964.270 1927.840 1964.590 1927.900 ;
        RECT 1745.310 1927.700 1745.630 1927.760 ;
        RECT 1929.310 1927.700 1929.630 1927.760 ;
        RECT 1745.310 1927.560 1929.630 1927.700 ;
        RECT 1745.310 1927.500 1745.630 1927.560 ;
        RECT 1929.310 1927.500 1929.630 1927.560 ;
        RECT 1779.350 1927.360 1779.670 1927.420 ;
        RECT 1998.310 1927.360 1998.630 1927.420 ;
        RECT 1779.350 1927.220 1998.630 1927.360 ;
        RECT 1779.350 1927.160 1779.670 1927.220 ;
        RECT 1998.310 1927.160 1998.630 1927.220 ;
        RECT 1766.010 1927.020 1766.330 1927.080 ;
        RECT 2010.270 1927.020 2010.590 1927.080 ;
        RECT 1766.010 1926.880 2010.590 1927.020 ;
        RECT 1766.010 1926.820 1766.330 1926.880 ;
        RECT 2010.270 1926.820 2010.590 1926.880 ;
        RECT 1786.710 1926.680 1787.030 1926.740 ;
        RECT 2033.270 1926.680 2033.590 1926.740 ;
        RECT 1786.710 1926.540 2033.590 1926.680 ;
        RECT 1786.710 1926.480 1787.030 1926.540 ;
        RECT 2033.270 1926.480 2033.590 1926.540 ;
        RECT 1738.410 1926.340 1738.730 1926.400 ;
        RECT 1987.270 1926.340 1987.590 1926.400 ;
        RECT 1738.410 1926.200 1987.590 1926.340 ;
        RECT 1738.410 1926.140 1738.730 1926.200 ;
        RECT 1987.270 1926.140 1987.590 1926.200 ;
        RECT 1717.710 1926.000 1718.030 1926.060 ;
        RECT 1975.310 1926.000 1975.630 1926.060 ;
        RECT 1717.710 1925.860 1975.630 1926.000 ;
        RECT 1717.710 1925.800 1718.030 1925.860 ;
        RECT 1975.310 1925.800 1975.630 1925.860 ;
        RECT 1779.810 1925.660 1780.130 1925.720 ;
        RECT 2067.310 1925.660 2067.630 1925.720 ;
        RECT 1779.810 1925.520 2067.630 1925.660 ;
        RECT 1779.810 1925.460 1780.130 1925.520 ;
        RECT 2067.310 1925.460 2067.630 1925.520 ;
        RECT 1835.010 1925.320 1835.330 1925.380 ;
        RECT 1952.310 1925.320 1952.630 1925.380 ;
        RECT 1835.010 1925.180 1952.630 1925.320 ;
        RECT 1835.010 1925.120 1835.330 1925.180 ;
        RECT 1952.310 1925.120 1952.630 1925.180 ;
        RECT 1357.530 1921.240 1357.850 1921.300 ;
        RECT 1358.450 1921.240 1358.770 1921.300 ;
        RECT 1357.530 1921.100 1358.770 1921.240 ;
        RECT 1357.530 1921.040 1357.850 1921.100 ;
        RECT 1358.450 1921.040 1358.770 1921.100 ;
        RECT 1485.870 1897.780 1486.190 1897.840 ;
        RECT 1490.010 1897.780 1490.330 1897.840 ;
        RECT 1485.870 1897.640 1490.330 1897.780 ;
        RECT 1485.870 1897.580 1486.190 1897.640 ;
        RECT 1490.010 1897.580 1490.330 1897.640 ;
        RECT 1358.450 1897.440 1358.770 1897.500 ;
        RECT 1358.910 1897.440 1359.230 1897.500 ;
        RECT 1358.450 1897.300 1359.230 1897.440 ;
        RECT 1358.450 1897.240 1358.770 1897.300 ;
        RECT 1358.910 1897.240 1359.230 1897.300 ;
        RECT 1405.830 1884.180 1406.150 1884.240 ;
        RECT 1407.670 1884.180 1407.990 1884.240 ;
        RECT 1405.830 1884.040 1407.990 1884.180 ;
        RECT 1405.830 1883.980 1406.150 1884.040 ;
        RECT 1407.670 1883.980 1407.990 1884.040 ;
        RECT 1534.170 1883.840 1534.490 1883.900 ;
        RECT 1535.090 1883.840 1535.410 1883.900 ;
        RECT 1534.170 1883.700 1535.410 1883.840 ;
        RECT 1534.170 1883.640 1534.490 1883.700 ;
        RECT 1535.090 1883.640 1535.410 1883.700 ;
        RECT 1542.910 1883.840 1543.230 1883.900 ;
        RECT 1543.370 1883.840 1543.690 1883.900 ;
        RECT 1542.910 1883.700 1543.690 1883.840 ;
        RECT 1542.910 1883.640 1543.230 1883.700 ;
        RECT 1543.370 1883.640 1543.690 1883.700 ;
        RECT 1759.110 1883.840 1759.430 1883.900 ;
        RECT 1904.470 1883.840 1904.790 1883.900 ;
        RECT 1759.110 1883.700 1904.790 1883.840 ;
        RECT 1759.110 1883.640 1759.430 1883.700 ;
        RECT 1904.470 1883.640 1904.790 1883.700 ;
        RECT 1405.370 1883.500 1405.690 1883.560 ;
        RECT 1405.830 1883.500 1406.150 1883.560 ;
        RECT 1405.370 1883.360 1406.150 1883.500 ;
        RECT 1405.370 1883.300 1405.690 1883.360 ;
        RECT 1405.830 1883.300 1406.150 1883.360 ;
        RECT 1821.210 1870.240 1821.530 1870.300 ;
        RECT 1904.470 1870.240 1904.790 1870.300 ;
        RECT 1821.210 1870.100 1904.790 1870.240 ;
        RECT 1821.210 1870.040 1821.530 1870.100 ;
        RECT 1904.470 1870.040 1904.790 1870.100 ;
        RECT 1737.950 1849.500 1738.270 1849.560 ;
        RECT 1904.470 1849.500 1904.790 1849.560 ;
        RECT 1737.950 1849.360 1904.790 1849.500 ;
        RECT 1737.950 1849.300 1738.270 1849.360 ;
        RECT 1904.470 1849.300 1904.790 1849.360 ;
        RECT 1405.370 1835.900 1405.690 1835.960 ;
        RECT 1406.750 1835.900 1407.070 1835.960 ;
        RECT 1405.370 1835.760 1407.070 1835.900 ;
        RECT 1405.370 1835.700 1405.690 1835.760 ;
        RECT 1406.750 1835.700 1407.070 1835.760 ;
        RECT 1405.370 1835.220 1405.690 1835.280 ;
        RECT 1406.750 1835.220 1407.070 1835.280 ;
        RECT 1405.370 1835.080 1407.070 1835.220 ;
        RECT 1405.370 1835.020 1405.690 1835.080 ;
        RECT 1406.750 1835.020 1407.070 1835.080 ;
        RECT 1534.170 1835.220 1534.490 1835.280 ;
        RECT 1535.090 1835.220 1535.410 1835.280 ;
        RECT 1534.170 1835.080 1535.410 1835.220 ;
        RECT 1534.170 1835.020 1534.490 1835.080 ;
        RECT 1535.090 1835.020 1535.410 1835.080 ;
        RECT 1543.370 1829.100 1543.690 1829.160 ;
        RECT 1544.290 1829.100 1544.610 1829.160 ;
        RECT 1543.370 1828.960 1544.610 1829.100 ;
        RECT 1543.370 1828.900 1543.690 1828.960 ;
        RECT 1544.290 1828.900 1544.610 1828.960 ;
        RECT 1543.370 1828.420 1543.690 1828.480 ;
        RECT 1544.290 1828.420 1544.610 1828.480 ;
        RECT 1543.370 1828.280 1544.610 1828.420 ;
        RECT 1543.370 1828.220 1543.690 1828.280 ;
        RECT 1544.290 1828.220 1544.610 1828.280 ;
        RECT 1669.410 1814.820 1669.730 1814.880 ;
        RECT 1904.470 1814.820 1904.790 1814.880 ;
        RECT 1669.410 1814.680 1904.790 1814.820 ;
        RECT 1669.410 1814.620 1669.730 1814.680 ;
        RECT 1904.470 1814.620 1904.790 1814.680 ;
        RECT 1358.450 1801.220 1358.770 1801.280 ;
        RECT 1358.910 1801.220 1359.230 1801.280 ;
        RECT 1358.450 1801.080 1359.230 1801.220 ;
        RECT 1358.450 1801.020 1358.770 1801.080 ;
        RECT 1358.910 1801.020 1359.230 1801.080 ;
        RECT 1405.370 1787.620 1405.690 1787.680 ;
        RECT 1405.830 1787.620 1406.150 1787.680 ;
        RECT 1405.370 1787.480 1406.150 1787.620 ;
        RECT 1405.370 1787.420 1405.690 1787.480 ;
        RECT 1405.830 1787.420 1406.150 1787.480 ;
        RECT 1534.170 1787.280 1534.490 1787.340 ;
        RECT 1535.090 1787.280 1535.410 1787.340 ;
        RECT 1534.170 1787.140 1535.410 1787.280 ;
        RECT 1534.170 1787.080 1534.490 1787.140 ;
        RECT 1535.090 1787.080 1535.410 1787.140 ;
        RECT 1543.370 1787.280 1543.690 1787.340 ;
        RECT 1543.370 1787.140 1544.520 1787.280 ;
        RECT 1543.370 1787.080 1543.690 1787.140 ;
        RECT 1544.380 1787.000 1544.520 1787.140 ;
        RECT 1405.370 1786.940 1405.690 1787.000 ;
        RECT 1405.830 1786.940 1406.150 1787.000 ;
        RECT 1405.370 1786.800 1406.150 1786.940 ;
        RECT 1405.370 1786.740 1405.690 1786.800 ;
        RECT 1405.830 1786.740 1406.150 1786.800 ;
        RECT 1544.290 1786.740 1544.610 1787.000 ;
        RECT 1772.910 1766.540 1773.230 1766.600 ;
        RECT 1904.470 1766.540 1904.790 1766.600 ;
        RECT 1772.910 1766.400 1904.790 1766.540 ;
        RECT 1772.910 1766.340 1773.230 1766.400 ;
        RECT 1904.470 1766.340 1904.790 1766.400 ;
      LAYER met1 ;
        RECT 1922.830 1760.240 2072.190 1905.280 ;
      LAYER met1 ;
        RECT 2073.290 1870.240 2073.610 1870.300 ;
        RECT 2283.970 1870.240 2284.290 1870.300 ;
        RECT 2073.290 1870.100 2284.290 1870.240 ;
        RECT 2073.290 1870.040 2073.610 1870.100 ;
        RECT 2283.970 1870.040 2284.290 1870.100 ;
        RECT 1405.370 1739.340 1405.690 1739.400 ;
        RECT 1406.750 1739.340 1407.070 1739.400 ;
        RECT 1405.370 1739.200 1407.070 1739.340 ;
        RECT 1405.370 1739.140 1405.690 1739.200 ;
        RECT 1406.750 1739.140 1407.070 1739.200 ;
        RECT 1405.370 1738.660 1405.690 1738.720 ;
        RECT 1406.750 1738.660 1407.070 1738.720 ;
        RECT 1405.370 1738.520 1407.070 1738.660 ;
        RECT 1405.370 1738.460 1405.690 1738.520 ;
        RECT 1406.750 1738.460 1407.070 1738.520 ;
        RECT 1534.170 1738.660 1534.490 1738.720 ;
        RECT 1534.630 1738.660 1534.950 1738.720 ;
        RECT 1534.170 1738.520 1534.950 1738.660 ;
        RECT 1534.170 1738.460 1534.490 1738.520 ;
        RECT 1534.630 1738.460 1534.950 1738.520 ;
        RECT 1827.650 1738.660 1827.970 1738.720 ;
        RECT 1933.910 1738.660 1934.230 1738.720 ;
        RECT 1827.650 1738.520 1934.230 1738.660 ;
        RECT 1827.650 1738.460 1827.970 1738.520 ;
        RECT 1933.910 1738.460 1934.230 1738.520 ;
        RECT 1800.510 1738.320 1800.830 1738.380 ;
        RECT 1956.910 1738.320 1957.230 1738.380 ;
        RECT 1800.510 1738.180 1957.230 1738.320 ;
        RECT 1800.510 1738.120 1800.830 1738.180 ;
        RECT 1956.910 1738.120 1957.230 1738.180 ;
        RECT 1793.610 1737.980 1793.930 1738.040 ;
        RECT 1967.950 1737.980 1968.270 1738.040 ;
        RECT 1793.610 1737.840 1968.270 1737.980 ;
        RECT 1793.610 1737.780 1793.930 1737.840 ;
        RECT 1967.950 1737.780 1968.270 1737.840 ;
        RECT 1814.310 1737.640 1814.630 1737.700 ;
        RECT 1990.950 1737.640 1991.270 1737.700 ;
        RECT 1814.310 1737.500 1991.270 1737.640 ;
        RECT 1814.310 1737.440 1814.630 1737.500 ;
        RECT 1990.950 1737.440 1991.270 1737.500 ;
        RECT 1813.850 1737.300 1814.170 1737.360 ;
        RECT 2013.950 1737.300 2014.270 1737.360 ;
        RECT 1813.850 1737.160 2014.270 1737.300 ;
        RECT 1813.850 1737.100 1814.170 1737.160 ;
        RECT 2013.950 1737.100 2014.270 1737.160 ;
        RECT 1752.670 1736.960 1752.990 1737.020 ;
        RECT 1979.910 1736.960 1980.230 1737.020 ;
        RECT 1752.670 1736.820 1980.230 1736.960 ;
        RECT 1752.670 1736.760 1752.990 1736.820 ;
        RECT 1979.910 1736.760 1980.230 1736.820 ;
        RECT 1710.810 1736.620 1711.130 1736.680 ;
        RECT 1944.950 1736.620 1945.270 1736.680 ;
        RECT 1710.810 1736.480 1945.270 1736.620 ;
        RECT 1710.810 1736.420 1711.130 1736.480 ;
        RECT 1944.950 1736.420 1945.270 1736.480 ;
        RECT 1807.410 1736.280 1807.730 1736.340 ;
        RECT 2036.950 1736.280 2037.270 1736.340 ;
        RECT 1807.410 1736.140 2037.270 1736.280 ;
        RECT 1807.410 1736.080 1807.730 1736.140 ;
        RECT 2036.950 1736.080 2037.270 1736.140 ;
        RECT 1772.450 1735.940 1772.770 1736.000 ;
        RECT 2002.910 1735.940 2003.230 1736.000 ;
        RECT 1772.450 1735.800 2003.230 1735.940 ;
        RECT 1772.450 1735.740 1772.770 1735.800 ;
        RECT 2002.910 1735.740 2003.230 1735.800 ;
        RECT 1806.950 1735.600 1807.270 1735.660 ;
        RECT 2071.910 1735.600 2072.230 1735.660 ;
        RECT 1806.950 1735.460 2072.230 1735.600 ;
        RECT 1806.950 1735.400 1807.270 1735.460 ;
        RECT 2071.910 1735.400 2072.230 1735.460 ;
        RECT 1372.250 1735.260 1372.570 1735.320 ;
        RECT 1553.030 1735.260 1553.350 1735.320 ;
        RECT 1372.250 1735.120 1553.350 1735.260 ;
        RECT 1372.250 1735.060 1372.570 1735.120 ;
        RECT 1553.030 1735.060 1553.350 1735.120 ;
        RECT 1668.950 1735.260 1669.270 1735.320 ;
        RECT 2059.950 1735.260 2060.270 1735.320 ;
        RECT 1668.950 1735.120 2060.270 1735.260 ;
        RECT 1668.950 1735.060 1669.270 1735.120 ;
        RECT 2059.950 1735.060 2060.270 1735.120 ;
        RECT 1543.370 1732.200 1543.690 1732.260 ;
        RECT 1543.830 1732.200 1544.150 1732.260 ;
        RECT 1543.370 1732.060 1544.150 1732.200 ;
        RECT 1543.370 1732.000 1543.690 1732.060 ;
        RECT 1543.830 1732.000 1544.150 1732.060 ;
      LAYER met1 ;
        RECT 2302.830 1710.640 2521.260 1926.000 ;
      LAYER met1 ;
        RECT 2519.030 1710.100 2519.350 1710.160 ;
        RECT 2520.870 1710.100 2521.190 1710.160 ;
        RECT 2519.030 1709.960 2521.190 1710.100 ;
        RECT 2519.030 1709.900 2519.350 1709.960 ;
        RECT 2520.870 1709.900 2521.190 1709.960 ;
        RECT 2523.630 1704.320 2523.950 1704.380 ;
        RECT 2520.500 1704.180 2523.950 1704.320 ;
        RECT 2519.490 1703.980 2519.810 1704.040 ;
        RECT 2520.500 1703.980 2520.640 1704.180 ;
        RECT 2523.630 1704.120 2523.950 1704.180 ;
        RECT 2519.490 1703.840 2520.640 1703.980 ;
        RECT 2519.490 1703.780 2519.810 1703.840 ;
        RECT 981.710 1695.140 982.030 1695.200 ;
        RECT 1048.870 1695.140 1049.190 1695.200 ;
        RECT 981.710 1695.000 1049.190 1695.140 ;
        RECT 981.710 1694.940 982.030 1695.000 ;
        RECT 1048.870 1694.940 1049.190 1695.000 ;
        RECT 998.730 1694.800 999.050 1694.860 ;
        RECT 1069.570 1694.800 1069.890 1694.860 ;
        RECT 998.730 1694.660 1069.890 1694.800 ;
        RECT 998.730 1694.600 999.050 1694.660 ;
        RECT 1069.570 1694.600 1069.890 1694.660 ;
        RECT 999.190 1694.460 999.510 1694.520 ;
        RECT 1076.470 1694.460 1076.790 1694.520 ;
        RECT 999.190 1694.320 1076.790 1694.460 ;
        RECT 999.190 1694.260 999.510 1694.320 ;
        RECT 1076.470 1694.260 1076.790 1694.320 ;
        RECT 982.170 1694.120 982.490 1694.180 ;
        RECT 1110.970 1694.120 1111.290 1694.180 ;
        RECT 982.170 1693.980 1111.290 1694.120 ;
        RECT 982.170 1693.920 982.490 1693.980 ;
        RECT 1110.970 1693.920 1111.290 1693.980 ;
        RECT 1289.910 1694.120 1290.230 1694.180 ;
        RECT 1336.370 1694.120 1336.690 1694.180 ;
        RECT 1289.910 1693.980 1336.690 1694.120 ;
        RECT 1289.910 1693.920 1290.230 1693.980 ;
        RECT 1336.370 1693.920 1336.690 1693.980 ;
        RECT 975.270 1693.780 975.590 1693.840 ;
        RECT 1104.070 1693.780 1104.390 1693.840 ;
        RECT 975.270 1693.640 1104.390 1693.780 ;
        RECT 975.270 1693.580 975.590 1693.640 ;
        RECT 1104.070 1693.580 1104.390 1693.640 ;
        RECT 1186.410 1693.780 1186.730 1693.840 ;
        RECT 1336.830 1693.780 1337.150 1693.840 ;
        RECT 1186.410 1693.640 1337.150 1693.780 ;
        RECT 1186.410 1693.580 1186.730 1693.640 ;
        RECT 1336.830 1693.580 1337.150 1693.640 ;
        RECT 1310.610 1693.100 1310.930 1693.160 ;
        RECT 1343.730 1693.100 1344.050 1693.160 ;
        RECT 1310.610 1692.960 1344.050 1693.100 ;
        RECT 1310.610 1692.900 1310.930 1692.960 ;
        RECT 1343.730 1692.900 1344.050 1692.960 ;
        RECT 1405.370 1690.720 1405.690 1690.780 ;
        RECT 1406.290 1690.720 1406.610 1690.780 ;
        RECT 1405.370 1690.580 1406.610 1690.720 ;
        RECT 1405.370 1690.520 1405.690 1690.580 ;
        RECT 1406.290 1690.520 1406.610 1690.580 ;
        RECT 1534.170 1690.720 1534.490 1690.780 ;
        RECT 1535.090 1690.720 1535.410 1690.780 ;
        RECT 1534.170 1690.580 1535.410 1690.720 ;
        RECT 1534.170 1690.520 1534.490 1690.580 ;
        RECT 1535.090 1690.520 1535.410 1690.580 ;
        RECT 1543.830 1690.520 1544.150 1690.780 ;
        RECT 1751.290 1690.720 1751.610 1690.780 ;
        RECT 1752.670 1690.720 1752.990 1690.780 ;
        RECT 1751.290 1690.580 1752.990 1690.720 ;
        RECT 1751.290 1690.520 1751.610 1690.580 ;
        RECT 1752.670 1690.520 1752.990 1690.580 ;
        RECT 1159.270 1690.040 1159.590 1690.100 ;
        RECT 1224.130 1690.040 1224.450 1690.100 ;
        RECT 1159.270 1689.900 1224.450 1690.040 ;
        RECT 1159.270 1689.840 1159.590 1689.900 ;
        RECT 1224.130 1689.840 1224.450 1689.900 ;
        RECT 1254.950 1690.040 1255.270 1690.100 ;
        RECT 1300.950 1690.040 1301.270 1690.100 ;
        RECT 1254.950 1689.900 1301.270 1690.040 ;
        RECT 1543.920 1690.040 1544.060 1690.520 ;
        RECT 1544.290 1690.040 1544.610 1690.100 ;
        RECT 1543.920 1689.900 1544.610 1690.040 ;
        RECT 1254.950 1689.840 1255.270 1689.900 ;
        RECT 1300.950 1689.840 1301.270 1689.900 ;
        RECT 1544.290 1689.840 1544.610 1689.900 ;
        RECT 1130.750 1689.700 1131.070 1689.760 ;
        RECT 1242.530 1689.700 1242.850 1689.760 ;
        RECT 1130.750 1689.560 1242.850 1689.700 ;
        RECT 1130.750 1689.500 1131.070 1689.560 ;
        RECT 1242.530 1689.500 1242.850 1689.560 ;
        RECT 1268.750 1689.700 1269.070 1689.760 ;
        RECT 1315.670 1689.700 1315.990 1689.760 ;
        RECT 1268.750 1689.560 1315.990 1689.700 ;
        RECT 1268.750 1689.500 1269.070 1689.560 ;
        RECT 1315.670 1689.500 1315.990 1689.560 ;
        RECT 1102.230 1689.360 1102.550 1689.420 ;
        RECT 1196.990 1689.360 1197.310 1689.420 ;
        RECT 1102.230 1689.220 1197.310 1689.360 ;
        RECT 1102.230 1689.160 1102.550 1689.220 ;
        RECT 1196.990 1689.160 1197.310 1689.220 ;
        RECT 1058.990 1689.020 1059.310 1689.080 ;
        RECT 1203.890 1689.020 1204.210 1689.080 ;
        RECT 1058.990 1688.880 1204.210 1689.020 ;
        RECT 1058.990 1688.820 1059.310 1688.880 ;
        RECT 1203.890 1688.820 1204.210 1688.880 ;
        RECT 1210.790 1689.020 1211.110 1689.080 ;
        RECT 1230.110 1689.020 1230.430 1689.080 ;
        RECT 1210.790 1688.880 1230.430 1689.020 ;
        RECT 1210.790 1688.820 1211.110 1688.880 ;
        RECT 1230.110 1688.820 1230.430 1688.880 ;
        RECT 1245.290 1689.020 1245.610 1689.080 ;
        RECT 1287.150 1689.020 1287.470 1689.080 ;
        RECT 1245.290 1688.880 1287.470 1689.020 ;
        RECT 1245.290 1688.820 1245.610 1688.880 ;
        RECT 1287.150 1688.820 1287.470 1688.880 ;
        RECT 463.750 1688.680 464.070 1688.740 ;
        RECT 468.810 1688.680 469.130 1688.740 ;
        RECT 463.750 1688.540 469.130 1688.680 ;
        RECT 463.750 1688.480 464.070 1688.540 ;
        RECT 468.810 1688.480 469.130 1688.540 ;
        RECT 514.350 1688.680 514.670 1688.740 ;
        RECT 517.110 1688.680 517.430 1688.740 ;
        RECT 514.350 1688.540 517.430 1688.680 ;
        RECT 514.350 1688.480 514.670 1688.540 ;
        RECT 517.110 1688.480 517.430 1688.540 ;
        RECT 1016.670 1688.680 1016.990 1688.740 ;
        RECT 1038.290 1688.680 1038.610 1688.740 ;
        RECT 1016.670 1688.540 1038.610 1688.680 ;
        RECT 1016.670 1688.480 1016.990 1688.540 ;
        RECT 1038.290 1688.480 1038.610 1688.540 ;
        RECT 1073.710 1688.680 1074.030 1688.740 ;
        RECT 1293.590 1688.680 1293.910 1688.740 ;
        RECT 1073.710 1688.540 1293.910 1688.680 ;
        RECT 1073.710 1688.480 1074.030 1688.540 ;
        RECT 1293.590 1688.480 1293.910 1688.540 ;
        RECT 1030.470 1688.340 1030.790 1688.400 ;
        RECT 1277.950 1688.340 1278.270 1688.400 ;
        RECT 1030.470 1688.200 1278.270 1688.340 ;
        RECT 1030.470 1688.140 1030.790 1688.200 ;
        RECT 1277.950 1688.140 1278.270 1688.200 ;
        RECT 2007.510 1688.000 2007.830 1688.060 ;
        RECT 2302.830 1688.000 2303.150 1688.060 ;
        RECT 2007.510 1687.860 2303.150 1688.000 ;
        RECT 2007.510 1687.800 2007.830 1687.860 ;
        RECT 2302.830 1687.800 2303.150 1687.860 ;
        RECT 2055.810 1687.660 2056.130 1687.720 ;
        RECT 2360.790 1687.660 2361.110 1687.720 ;
        RECT 2055.810 1687.520 2361.110 1687.660 ;
        RECT 2055.810 1687.460 2056.130 1687.520 ;
        RECT 2360.790 1687.460 2361.110 1687.520 ;
        RECT 2042.010 1687.320 2042.330 1687.380 ;
        RECT 2418.750 1687.320 2419.070 1687.380 ;
        RECT 2042.010 1687.180 2419.070 1687.320 ;
        RECT 2042.010 1687.120 2042.330 1687.180 ;
        RECT 2418.750 1687.120 2419.070 1687.180 ;
        RECT 2069.610 1686.980 2069.930 1687.040 ;
        RECT 2476.710 1686.980 2477.030 1687.040 ;
        RECT 2069.610 1686.840 2477.030 1686.980 ;
        RECT 2069.610 1686.780 2069.930 1686.840 ;
        RECT 2476.710 1686.780 2477.030 1686.840 ;
        RECT 1116.030 1686.640 1116.350 1686.700 ;
        RECT 1188.250 1686.640 1188.570 1686.700 ;
        RECT 1116.030 1686.500 1188.570 1686.640 ;
        RECT 1116.030 1686.440 1116.350 1686.500 ;
        RECT 1188.250 1686.440 1188.570 1686.500 ;
        RECT 1196.990 1686.640 1197.310 1686.700 ;
        RECT 1231.490 1686.640 1231.810 1686.700 ;
        RECT 1196.990 1686.500 1231.810 1686.640 ;
        RECT 1196.990 1686.440 1197.310 1686.500 ;
        RECT 1231.490 1686.440 1231.810 1686.500 ;
        RECT 1144.550 1686.300 1144.870 1686.360 ;
        RECT 1179.970 1686.300 1180.290 1686.360 ;
        RECT 1144.550 1686.160 1180.290 1686.300 ;
        RECT 1144.550 1686.100 1144.870 1686.160 ;
        RECT 1179.970 1686.100 1180.290 1686.160 ;
        RECT 1214.010 1686.300 1214.330 1686.360 ;
        RECT 1245.290 1686.300 1245.610 1686.360 ;
        RECT 1214.010 1686.160 1245.610 1686.300 ;
        RECT 1214.010 1686.100 1214.330 1686.160 ;
        RECT 1245.290 1686.100 1245.610 1686.160 ;
        RECT 1258.630 1686.300 1258.950 1686.360 ;
        RECT 1300.490 1686.300 1300.810 1686.360 ;
        RECT 1258.630 1686.160 1300.810 1686.300 ;
        RECT 1258.630 1686.100 1258.950 1686.160 ;
        RECT 1300.490 1686.100 1300.810 1686.160 ;
        RECT 1358.910 1684.400 1359.230 1684.660 ;
        RECT 1002.870 1684.260 1003.190 1684.320 ;
        RECT 1007.010 1684.260 1007.330 1684.320 ;
        RECT 1002.870 1684.120 1007.330 1684.260 ;
        RECT 1002.870 1684.060 1003.190 1684.120 ;
        RECT 1007.010 1684.060 1007.330 1684.120 ;
        RECT 1173.070 1684.260 1173.390 1684.320 ;
        RECT 1187.330 1684.260 1187.650 1684.320 ;
        RECT 1173.070 1684.120 1187.650 1684.260 ;
        RECT 1173.070 1684.060 1173.390 1684.120 ;
        RECT 1187.330 1684.060 1187.650 1684.120 ;
        RECT 1187.790 1684.260 1188.110 1684.320 ;
        RECT 1196.990 1684.260 1197.310 1684.320 ;
        RECT 1187.790 1684.120 1197.310 1684.260 ;
        RECT 1187.790 1684.060 1188.110 1684.120 ;
        RECT 1196.990 1684.060 1197.310 1684.120 ;
        RECT 1200.210 1684.260 1200.530 1684.320 ;
        RECT 1215.390 1684.260 1215.710 1684.320 ;
        RECT 1200.210 1684.120 1215.710 1684.260 ;
        RECT 1200.210 1684.060 1200.530 1684.120 ;
        RECT 1215.390 1684.060 1215.710 1684.120 ;
        RECT 1238.390 1684.260 1238.710 1684.320 ;
        RECT 1243.910 1684.260 1244.230 1684.320 ;
        RECT 1238.390 1684.120 1244.230 1684.260 ;
        RECT 1238.390 1684.060 1238.710 1684.120 ;
        RECT 1243.910 1684.060 1244.230 1684.120 ;
        RECT 1272.430 1684.260 1272.750 1684.320 ;
        RECT 1292.210 1684.260 1292.530 1684.320 ;
        RECT 1272.430 1684.120 1292.530 1684.260 ;
        RECT 1272.430 1684.060 1272.750 1684.120 ;
        RECT 1292.210 1684.060 1292.530 1684.120 ;
        RECT 1329.470 1684.260 1329.790 1684.320 ;
        RECT 1348.330 1684.260 1348.650 1684.320 ;
        RECT 1329.470 1684.120 1348.650 1684.260 ;
        RECT 1329.470 1684.060 1329.790 1684.120 ;
        RECT 1348.330 1684.060 1348.650 1684.120 ;
        RECT 1358.450 1684.260 1358.770 1684.320 ;
        RECT 1359.000 1684.260 1359.140 1684.400 ;
        RECT 1358.450 1684.120 1359.140 1684.260 ;
        RECT 1358.450 1684.060 1358.770 1684.120 ;
        RECT 1290.830 1683.580 1291.150 1683.640 ;
        RECT 1292.210 1683.580 1292.530 1683.640 ;
        RECT 1290.830 1683.440 1292.530 1683.580 ;
        RECT 1290.830 1683.380 1291.150 1683.440 ;
        RECT 1292.210 1683.380 1292.530 1683.440 ;
        RECT 2518.110 1656.040 2518.430 1656.100 ;
        RECT 2519.950 1656.040 2520.270 1656.100 ;
        RECT 2518.110 1655.900 2520.270 1656.040 ;
        RECT 2518.110 1655.840 2518.430 1655.900 ;
        RECT 2519.950 1655.840 2520.270 1655.900 ;
        RECT 1357.070 1652.640 1357.390 1652.700 ;
        RECT 1357.990 1652.640 1358.310 1652.700 ;
        RECT 1357.070 1652.500 1358.310 1652.640 ;
        RECT 1357.070 1652.440 1357.390 1652.500 ;
        RECT 1357.990 1652.440 1358.310 1652.500 ;
        RECT 1224.130 1642.440 1224.450 1642.500 ;
        RECT 1243.450 1642.440 1243.770 1642.500 ;
        RECT 1224.130 1642.300 1243.770 1642.440 ;
        RECT 1224.130 1642.240 1224.450 1642.300 ;
        RECT 1243.450 1642.240 1243.770 1642.300 ;
        RECT 1405.830 1642.440 1406.150 1642.500 ;
        RECT 1406.290 1642.440 1406.610 1642.500 ;
        RECT 1405.830 1642.300 1406.610 1642.440 ;
        RECT 1405.830 1642.240 1406.150 1642.300 ;
        RECT 1406.290 1642.240 1406.610 1642.300 ;
        RECT 1535.090 1641.900 1535.410 1642.160 ;
        RECT 2517.650 1642.100 2517.970 1642.160 ;
        RECT 2518.570 1642.100 2518.890 1642.160 ;
        RECT 2517.650 1641.960 2518.890 1642.100 ;
        RECT 2517.650 1641.900 2517.970 1641.960 ;
        RECT 2518.570 1641.900 2518.890 1641.960 ;
        RECT 1535.180 1641.480 1535.320 1641.900 ;
        RECT 1535.090 1641.220 1535.410 1641.480 ;
        RECT 1543.830 1635.980 1544.150 1636.040 ;
        RECT 1543.830 1635.840 1544.520 1635.980 ;
        RECT 1543.830 1635.780 1544.150 1635.840 ;
        RECT 1544.380 1635.700 1544.520 1635.840 ;
        RECT 1290.830 1635.640 1291.150 1635.700 ;
        RECT 1291.750 1635.640 1292.070 1635.700 ;
        RECT 1290.830 1635.500 1292.070 1635.640 ;
        RECT 1290.830 1635.440 1291.150 1635.500 ;
        RECT 1291.750 1635.440 1292.070 1635.500 ;
        RECT 1544.290 1635.440 1544.610 1635.700 ;
        RECT 1357.070 1628.500 1357.390 1628.560 ;
        RECT 1357.530 1628.500 1357.850 1628.560 ;
        RECT 1357.070 1628.360 1357.850 1628.500 ;
        RECT 1357.070 1628.300 1357.390 1628.360 ;
        RECT 1357.530 1628.300 1357.850 1628.360 ;
        RECT 2519.950 1617.960 2520.270 1618.020 ;
        RECT 2520.870 1617.960 2521.190 1618.020 ;
        RECT 2519.950 1617.820 2521.190 1617.960 ;
        RECT 2519.950 1617.760 2520.270 1617.820 ;
        RECT 2520.870 1617.760 2521.190 1617.820 ;
        RECT 1357.530 1614.560 1357.850 1614.620 ;
        RECT 1358.450 1614.560 1358.770 1614.620 ;
        RECT 1357.530 1614.420 1358.770 1614.560 ;
        RECT 1357.530 1614.360 1357.850 1614.420 ;
        RECT 1358.450 1614.360 1358.770 1614.420 ;
        RECT 1406.290 1607.760 1406.610 1607.820 ;
        RECT 1406.750 1607.760 1407.070 1607.820 ;
        RECT 1406.290 1607.620 1407.070 1607.760 ;
        RECT 1406.290 1607.560 1406.610 1607.620 ;
        RECT 1406.750 1607.560 1407.070 1607.620 ;
        RECT 1278.870 1594.160 1279.190 1594.220 ;
        RECT 1279.330 1594.160 1279.650 1594.220 ;
        RECT 1278.870 1594.020 1279.650 1594.160 ;
        RECT 1278.870 1593.960 1279.190 1594.020 ;
        RECT 1279.330 1593.960 1279.650 1594.020 ;
        RECT 2517.650 1594.160 2517.970 1594.220 ;
        RECT 2518.570 1594.160 2518.890 1594.220 ;
        RECT 2517.650 1594.020 2518.890 1594.160 ;
        RECT 2517.650 1593.960 2517.970 1594.020 ;
        RECT 2518.570 1593.960 2518.890 1594.020 ;
        RECT 2519.950 1594.160 2520.270 1594.220 ;
        RECT 2520.870 1594.160 2521.190 1594.220 ;
        RECT 2519.950 1594.020 2521.190 1594.160 ;
        RECT 2519.950 1593.960 2520.270 1594.020 ;
        RECT 2520.870 1593.960 2521.190 1594.020 ;
        RECT 1288.530 1593.820 1288.850 1593.880 ;
        RECT 1289.910 1593.820 1290.230 1593.880 ;
        RECT 1288.530 1593.680 1290.230 1593.820 ;
        RECT 1288.530 1593.620 1288.850 1593.680 ;
        RECT 1289.910 1593.620 1290.230 1593.680 ;
        RECT 1405.370 1593.820 1405.690 1593.880 ;
        RECT 1406.750 1593.820 1407.070 1593.880 ;
        RECT 1405.370 1593.680 1407.070 1593.820 ;
        RECT 1405.370 1593.620 1405.690 1593.680 ;
        RECT 1406.750 1593.620 1407.070 1593.680 ;
        RECT 1290.830 1587.360 1291.150 1587.420 ;
        RECT 1293.130 1587.360 1293.450 1587.420 ;
        RECT 1290.830 1587.220 1293.450 1587.360 ;
        RECT 1290.830 1587.160 1291.150 1587.220 ;
        RECT 1293.130 1587.160 1293.450 1587.220 ;
        RECT 2517.190 1569.680 2517.510 1569.740 ;
        RECT 2518.570 1569.680 2518.890 1569.740 ;
        RECT 2517.190 1569.540 2518.890 1569.680 ;
        RECT 2517.190 1569.480 2517.510 1569.540 ;
        RECT 2518.570 1569.480 2518.890 1569.540 ;
        RECT 2518.110 1559.480 2518.430 1559.540 ;
        RECT 2519.950 1559.480 2520.270 1559.540 ;
        RECT 2518.110 1559.340 2520.270 1559.480 ;
        RECT 2518.110 1559.280 2518.430 1559.340 ;
        RECT 2519.950 1559.280 2520.270 1559.340 ;
        RECT 2518.110 1558.800 2518.430 1558.860 ;
        RECT 2519.950 1558.800 2520.270 1558.860 ;
        RECT 2518.110 1558.660 2520.270 1558.800 ;
        RECT 2518.110 1558.600 2518.430 1558.660 ;
        RECT 2519.950 1558.600 2520.270 1558.660 ;
        RECT 1288.530 1545.880 1288.850 1545.940 ;
        RECT 1288.990 1545.880 1289.310 1545.940 ;
        RECT 1288.530 1545.740 1289.310 1545.880 ;
        RECT 1288.530 1545.680 1288.850 1545.740 ;
        RECT 1288.990 1545.680 1289.310 1545.740 ;
        RECT 1405.370 1545.880 1405.690 1545.940 ;
        RECT 1406.290 1545.880 1406.610 1545.940 ;
        RECT 1405.370 1545.740 1406.610 1545.880 ;
        RECT 1405.370 1545.680 1405.690 1545.740 ;
        RECT 1406.290 1545.680 1406.610 1545.740 ;
        RECT 1535.090 1545.880 1535.410 1545.940 ;
        RECT 2517.190 1545.880 2517.510 1545.940 ;
        RECT 2519.030 1545.880 2519.350 1545.940 ;
        RECT 1535.090 1545.740 1535.780 1545.880 ;
        RECT 1535.090 1545.680 1535.410 1545.740 ;
        RECT 1535.640 1545.600 1535.780 1545.740 ;
        RECT 2517.190 1545.740 2519.350 1545.880 ;
        RECT 2517.190 1545.680 2517.510 1545.740 ;
        RECT 2519.030 1545.680 2519.350 1545.740 ;
        RECT 1535.550 1545.340 1535.870 1545.600 ;
        RECT 1535.550 1539.080 1535.870 1539.140 ;
        RECT 1536.010 1539.080 1536.330 1539.140 ;
        RECT 1535.550 1538.940 1536.330 1539.080 ;
        RECT 1535.550 1538.880 1535.870 1538.940 ;
        RECT 1536.010 1538.880 1536.330 1538.940 ;
        RECT 1358.910 1518.000 1359.230 1518.060 ;
        RECT 1359.830 1518.000 1360.150 1518.060 ;
        RECT 1358.910 1517.860 1360.150 1518.000 ;
        RECT 1358.910 1517.800 1359.230 1517.860 ;
        RECT 1359.830 1517.800 1360.150 1517.860 ;
        RECT 1406.290 1511.000 1406.610 1511.260 ;
        RECT 1406.380 1510.860 1406.520 1511.000 ;
        RECT 1406.750 1510.860 1407.070 1510.920 ;
        RECT 1406.380 1510.720 1407.070 1510.860 ;
        RECT 1406.750 1510.660 1407.070 1510.720 ;
        RECT 1535.090 1497.600 1535.410 1497.660 ;
        RECT 1536.010 1497.600 1536.330 1497.660 ;
        RECT 1535.090 1497.460 1536.330 1497.600 ;
        RECT 1535.090 1497.400 1535.410 1497.460 ;
        RECT 1536.010 1497.400 1536.330 1497.460 ;
        RECT 1543.370 1497.600 1543.690 1497.660 ;
        RECT 1543.830 1497.600 1544.150 1497.660 ;
        RECT 1543.370 1497.460 1544.150 1497.600 ;
        RECT 1543.370 1497.400 1543.690 1497.460 ;
        RECT 1543.830 1497.400 1544.150 1497.460 ;
        RECT 1277.490 1497.260 1277.810 1497.320 ;
        RECT 1277.950 1497.260 1278.270 1497.320 ;
        RECT 1277.490 1497.120 1278.270 1497.260 ;
        RECT 1277.490 1497.060 1277.810 1497.120 ;
        RECT 1277.950 1497.060 1278.270 1497.120 ;
        RECT 1288.530 1497.260 1288.850 1497.320 ;
        RECT 1289.450 1497.260 1289.770 1497.320 ;
        RECT 1288.530 1497.120 1289.770 1497.260 ;
        RECT 1288.530 1497.060 1288.850 1497.120 ;
        RECT 1289.450 1497.060 1289.770 1497.120 ;
        RECT 1291.290 1497.260 1291.610 1497.320 ;
        RECT 1291.750 1497.260 1292.070 1497.320 ;
        RECT 1291.290 1497.120 1292.070 1497.260 ;
        RECT 1291.290 1497.060 1291.610 1497.120 ;
        RECT 1291.750 1497.060 1292.070 1497.120 ;
        RECT 1405.370 1497.260 1405.690 1497.320 ;
        RECT 1406.750 1497.260 1407.070 1497.320 ;
        RECT 1405.370 1497.120 1407.070 1497.260 ;
        RECT 1405.370 1497.060 1405.690 1497.120 ;
        RECT 1406.750 1497.060 1407.070 1497.120 ;
        RECT 1543.370 1462.920 1543.690 1462.980 ;
        RECT 1544.290 1462.920 1544.610 1462.980 ;
        RECT 1543.370 1462.780 1544.610 1462.920 ;
        RECT 1543.370 1462.720 1543.690 1462.780 ;
        RECT 1544.290 1462.720 1544.610 1462.780 ;
        RECT 1614.210 1459.860 1614.530 1459.920 ;
        RECT 1893.430 1459.860 1893.750 1459.920 ;
        RECT 1614.210 1459.720 1893.750 1459.860 ;
        RECT 1614.210 1459.660 1614.530 1459.720 ;
        RECT 1893.430 1459.660 1893.750 1459.720 ;
        RECT 1503.810 1459.520 1504.130 1459.580 ;
        RECT 1892.970 1459.520 1893.290 1459.580 ;
        RECT 1503.810 1459.380 1893.290 1459.520 ;
        RECT 1503.810 1459.320 1504.130 1459.380 ;
        RECT 1892.970 1459.320 1893.290 1459.380 ;
        RECT 994.590 1459.180 994.910 1459.240 ;
        RECT 1159.270 1459.180 1159.590 1459.240 ;
        RECT 994.590 1459.040 1159.590 1459.180 ;
        RECT 994.590 1458.980 994.910 1459.040 ;
        RECT 1159.270 1458.980 1159.590 1459.040 ;
        RECT 1503.350 1459.180 1503.670 1459.240 ;
        RECT 1894.350 1459.180 1894.670 1459.240 ;
        RECT 1503.350 1459.040 1894.670 1459.180 ;
        RECT 1503.350 1458.980 1503.670 1459.040 ;
        RECT 1894.350 1458.980 1894.670 1459.040 ;
        RECT 1277.490 1449.660 1277.810 1449.720 ;
        RECT 1291.290 1449.660 1291.610 1449.720 ;
        RECT 1277.490 1449.520 1278.180 1449.660 ;
        RECT 1277.490 1449.460 1277.810 1449.520 ;
        RECT 1278.040 1449.380 1278.180 1449.520 ;
        RECT 1291.290 1449.520 1291.980 1449.660 ;
        RECT 1291.290 1449.460 1291.610 1449.520 ;
        RECT 1291.840 1449.380 1291.980 1449.520 ;
        RECT 1277.950 1449.120 1278.270 1449.380 ;
        RECT 1288.530 1449.320 1288.850 1449.380 ;
        RECT 1288.990 1449.320 1289.310 1449.380 ;
        RECT 1288.530 1449.180 1289.310 1449.320 ;
        RECT 1288.530 1449.120 1288.850 1449.180 ;
        RECT 1288.990 1449.120 1289.310 1449.180 ;
        RECT 1291.750 1449.120 1292.070 1449.380 ;
        RECT 1405.370 1449.320 1405.690 1449.380 ;
        RECT 1406.290 1449.320 1406.610 1449.380 ;
        RECT 1405.370 1449.180 1406.610 1449.320 ;
        RECT 1405.370 1449.120 1405.690 1449.180 ;
        RECT 1406.290 1449.120 1406.610 1449.180 ;
        RECT 1358.910 1421.440 1359.230 1421.500 ;
        RECT 1359.830 1421.440 1360.150 1421.500 ;
        RECT 1358.910 1421.300 1360.150 1421.440 ;
        RECT 1358.910 1421.240 1359.230 1421.300 ;
        RECT 1359.830 1421.240 1360.150 1421.300 ;
        RECT 1542.910 1418.040 1543.230 1418.100 ;
        RECT 1544.290 1418.040 1544.610 1418.100 ;
        RECT 1542.910 1417.900 1544.610 1418.040 ;
        RECT 1542.910 1417.840 1543.230 1417.900 ;
        RECT 1544.290 1417.840 1544.610 1417.900 ;
        RECT 2518.570 1415.320 2518.890 1415.380 ;
        RECT 2518.570 1415.180 2519.260 1415.320 ;
        RECT 2518.570 1415.120 2518.890 1415.180 ;
        RECT 2519.120 1415.040 2519.260 1415.180 ;
        RECT 2519.030 1414.780 2519.350 1415.040 ;
        RECT 1288.990 1414.640 1289.310 1414.700 ;
        RECT 1289.910 1414.640 1290.230 1414.700 ;
        RECT 1288.990 1414.500 1290.230 1414.640 ;
        RECT 1288.990 1414.440 1289.310 1414.500 ;
        RECT 1289.910 1414.440 1290.230 1414.500 ;
        RECT 1406.290 1414.440 1406.610 1414.700 ;
        RECT 1406.380 1414.300 1406.520 1414.440 ;
        RECT 1406.750 1414.300 1407.070 1414.360 ;
        RECT 1406.380 1414.160 1407.070 1414.300 ;
        RECT 1406.750 1414.100 1407.070 1414.160 ;
        RECT 1406.750 1400.700 1407.070 1400.760 ;
        RECT 1408.130 1400.700 1408.450 1400.760 ;
        RECT 1406.750 1400.560 1408.450 1400.700 ;
        RECT 1406.750 1400.500 1407.070 1400.560 ;
        RECT 1408.130 1400.500 1408.450 1400.560 ;
        RECT 1542.910 1393.900 1543.230 1393.960 ;
        RECT 1543.370 1393.900 1543.690 1393.960 ;
        RECT 1542.910 1393.760 1543.690 1393.900 ;
        RECT 1542.910 1393.700 1543.230 1393.760 ;
        RECT 1543.370 1393.700 1543.690 1393.760 ;
        RECT 1291.290 1379.960 1291.610 1380.020 ;
        RECT 1291.750 1379.960 1292.070 1380.020 ;
        RECT 1291.290 1379.820 1292.070 1379.960 ;
        RECT 1291.290 1379.760 1291.610 1379.820 ;
        RECT 1291.750 1379.760 1292.070 1379.820 ;
        RECT 2518.110 1366.700 2518.430 1366.760 ;
        RECT 2519.950 1366.700 2520.270 1366.760 ;
        RECT 2518.110 1366.560 2520.270 1366.700 ;
        RECT 2518.110 1366.500 2518.430 1366.560 ;
        RECT 2519.950 1366.500 2520.270 1366.560 ;
        RECT 2518.110 1366.020 2518.430 1366.080 ;
        RECT 2519.950 1366.020 2520.270 1366.080 ;
        RECT 2518.110 1365.880 2520.270 1366.020 ;
        RECT 2518.110 1365.820 2518.430 1365.880 ;
        RECT 2519.950 1365.820 2520.270 1365.880 ;
        RECT 1406.750 1353.100 1407.070 1353.160 ;
        RECT 1408.130 1353.100 1408.450 1353.160 ;
        RECT 1406.750 1352.960 1408.450 1353.100 ;
        RECT 1406.750 1352.900 1407.070 1352.960 ;
        RECT 1408.130 1352.900 1408.450 1352.960 ;
        RECT 1535.090 1352.760 1535.410 1352.820 ;
        RECT 1534.720 1352.620 1535.410 1352.760 ;
        RECT 1534.720 1352.480 1534.860 1352.620 ;
        RECT 1535.090 1352.560 1535.410 1352.620 ;
        RECT 1405.370 1352.420 1405.690 1352.480 ;
        RECT 1406.750 1352.420 1407.070 1352.480 ;
        RECT 1405.370 1352.280 1407.070 1352.420 ;
        RECT 1405.370 1352.220 1405.690 1352.280 ;
        RECT 1406.750 1352.220 1407.070 1352.280 ;
        RECT 1534.630 1352.220 1534.950 1352.480 ;
        RECT 1543.370 1345.620 1543.690 1345.680 ;
        RECT 1544.290 1345.620 1544.610 1345.680 ;
        RECT 1543.370 1345.480 1544.610 1345.620 ;
        RECT 1543.370 1345.420 1543.690 1345.480 ;
        RECT 1544.290 1345.420 1544.610 1345.480 ;
        RECT 1533.710 1345.280 1534.030 1345.340 ;
        RECT 1534.630 1345.280 1534.950 1345.340 ;
        RECT 1533.710 1345.140 1534.950 1345.280 ;
        RECT 1533.710 1345.080 1534.030 1345.140 ;
        RECT 1534.630 1345.080 1534.950 1345.140 ;
        RECT 1357.990 1324.540 1358.310 1324.600 ;
        RECT 1358.910 1324.540 1359.230 1324.600 ;
        RECT 1357.990 1324.400 1359.230 1324.540 ;
        RECT 1357.990 1324.340 1358.310 1324.400 ;
        RECT 1358.910 1324.340 1359.230 1324.400 ;
        RECT 2518.570 1318.420 2518.890 1318.480 ;
        RECT 2519.950 1318.420 2520.270 1318.480 ;
        RECT 2518.570 1318.280 2520.270 1318.420 ;
        RECT 2518.570 1318.220 2518.890 1318.280 ;
        RECT 2519.950 1318.220 2520.270 1318.280 ;
        RECT 2518.570 1317.740 2518.890 1317.800 ;
        RECT 2519.950 1317.740 2520.270 1317.800 ;
        RECT 2518.570 1317.600 2520.270 1317.740 ;
        RECT 2518.570 1317.540 2518.890 1317.600 ;
        RECT 2519.950 1317.540 2520.270 1317.600 ;
        RECT 1278.410 1304.280 1278.730 1304.540 ;
        RECT 1405.370 1304.480 1405.690 1304.540 ;
        RECT 1406.290 1304.480 1406.610 1304.540 ;
        RECT 1405.370 1304.340 1406.610 1304.480 ;
        RECT 1405.370 1304.280 1405.690 1304.340 ;
        RECT 1406.290 1304.280 1406.610 1304.340 ;
        RECT 1278.500 1303.860 1278.640 1304.280 ;
        RECT 1278.410 1303.600 1278.730 1303.860 ;
        RECT 1533.710 1297.340 1534.030 1297.400 ;
        RECT 1535.090 1297.340 1535.410 1297.400 ;
        RECT 1533.710 1297.200 1535.410 1297.340 ;
        RECT 1533.710 1297.140 1534.030 1297.200 ;
        RECT 1535.090 1297.140 1535.410 1297.200 ;
        RECT 1357.070 1276.260 1357.390 1276.320 ;
        RECT 1358.910 1276.260 1359.230 1276.320 ;
        RECT 1357.070 1276.120 1359.230 1276.260 ;
        RECT 1357.070 1276.060 1357.390 1276.120 ;
        RECT 1358.910 1276.060 1359.230 1276.120 ;
        RECT 2518.110 1270.140 2518.430 1270.200 ;
        RECT 2519.950 1270.140 2520.270 1270.200 ;
        RECT 2518.110 1270.000 2520.270 1270.140 ;
        RECT 2518.110 1269.940 2518.430 1270.000 ;
        RECT 2519.950 1269.940 2520.270 1270.000 ;
        RECT 2518.110 1269.460 2518.430 1269.520 ;
        RECT 2519.950 1269.460 2520.270 1269.520 ;
        RECT 2518.110 1269.320 2520.270 1269.460 ;
        RECT 2518.110 1269.260 2518.430 1269.320 ;
        RECT 2519.950 1269.260 2520.270 1269.320 ;
        RECT 1535.090 1257.360 1535.410 1257.620 ;
        RECT 1535.180 1256.940 1535.320 1257.360 ;
        RECT 1535.090 1256.680 1535.410 1256.940 ;
        RECT 1292.210 1245.460 1292.530 1245.720 ;
        RECT 1292.300 1245.040 1292.440 1245.460 ;
        RECT 1292.210 1244.780 1292.530 1245.040 ;
        RECT 1357.070 1228.320 1357.390 1228.380 ;
        RECT 1357.530 1228.320 1357.850 1228.380 ;
        RECT 1357.070 1228.180 1357.850 1228.320 ;
        RECT 1357.070 1228.120 1357.390 1228.180 ;
        RECT 1357.530 1228.120 1357.850 1228.180 ;
        RECT 1542.910 1226.960 1543.230 1227.020 ;
        RECT 1544.290 1226.960 1544.610 1227.020 ;
        RECT 1542.910 1226.820 1544.610 1226.960 ;
        RECT 1542.910 1226.760 1543.230 1226.820 ;
        RECT 1544.290 1226.760 1544.610 1226.820 ;
        RECT 2518.570 1222.200 2518.890 1222.260 ;
        RECT 2518.570 1222.060 2519.260 1222.200 ;
        RECT 2518.570 1222.000 2518.890 1222.060 ;
        RECT 2519.120 1221.920 2519.260 1222.060 ;
        RECT 2519.030 1221.660 2519.350 1221.920 ;
        RECT 1357.530 1210.980 1357.850 1211.040 ;
        RECT 1358.910 1210.980 1359.230 1211.040 ;
        RECT 1357.530 1210.840 1359.230 1210.980 ;
        RECT 1357.530 1210.780 1357.850 1210.840 ;
        RECT 1358.910 1210.780 1359.230 1210.840 ;
        RECT 1535.090 1207.920 1535.410 1207.980 ;
        RECT 1536.010 1207.920 1536.330 1207.980 ;
        RECT 1535.090 1207.780 1536.330 1207.920 ;
        RECT 1535.090 1207.720 1535.410 1207.780 ;
        RECT 1536.010 1207.720 1536.330 1207.780 ;
        RECT 1405.370 1207.580 1405.690 1207.640 ;
        RECT 1406.290 1207.580 1406.610 1207.640 ;
        RECT 1405.370 1207.440 1406.610 1207.580 ;
        RECT 1405.370 1207.380 1405.690 1207.440 ;
        RECT 1406.290 1207.380 1406.610 1207.440 ;
        RECT 1405.370 1206.900 1405.690 1206.960 ;
        RECT 1406.290 1206.900 1406.610 1206.960 ;
        RECT 1405.370 1206.760 1406.610 1206.900 ;
        RECT 1405.370 1206.700 1405.690 1206.760 ;
        RECT 1406.290 1206.700 1406.610 1206.760 ;
        RECT 1291.290 1200.780 1291.610 1200.840 ;
        RECT 1292.210 1200.780 1292.530 1200.840 ;
        RECT 1291.290 1200.640 1292.530 1200.780 ;
        RECT 1291.290 1200.580 1291.610 1200.640 ;
        RECT 1292.210 1200.580 1292.530 1200.640 ;
        RECT 1291.290 1193.640 1291.610 1193.700 ;
        RECT 1292.210 1193.640 1292.530 1193.700 ;
        RECT 1291.290 1193.500 1292.530 1193.640 ;
        RECT 1291.290 1193.440 1291.610 1193.500 ;
        RECT 1292.210 1193.440 1292.530 1193.500 ;
        RECT 1277.030 1183.440 1277.350 1183.500 ;
        RECT 1277.950 1183.440 1278.270 1183.500 ;
        RECT 1277.030 1183.300 1278.270 1183.440 ;
        RECT 1277.030 1183.240 1277.350 1183.300 ;
        RECT 1277.950 1183.240 1278.270 1183.300 ;
        RECT 1542.910 1176.640 1543.230 1176.700 ;
        RECT 1543.830 1176.640 1544.150 1176.700 ;
        RECT 1542.910 1176.500 1544.150 1176.640 ;
        RECT 1542.910 1176.440 1543.230 1176.500 ;
        RECT 1543.830 1176.440 1544.150 1176.500 ;
        RECT 2518.110 1173.580 2518.430 1173.640 ;
        RECT 2519.950 1173.580 2520.270 1173.640 ;
        RECT 2518.110 1173.440 2520.270 1173.580 ;
        RECT 2518.110 1173.380 2518.430 1173.440 ;
        RECT 2519.950 1173.380 2520.270 1173.440 ;
        RECT 2518.110 1172.900 2518.430 1172.960 ;
        RECT 2519.950 1172.900 2520.270 1172.960 ;
        RECT 2518.110 1172.760 2520.270 1172.900 ;
        RECT 2518.110 1172.700 2518.430 1172.760 ;
        RECT 2519.950 1172.700 2520.270 1172.760 ;
        RECT 1289.910 1159.300 1290.230 1159.360 ;
        RECT 1290.830 1159.300 1291.150 1159.360 ;
        RECT 1289.910 1159.160 1291.150 1159.300 ;
        RECT 1289.910 1159.100 1290.230 1159.160 ;
        RECT 1290.830 1159.100 1291.150 1159.160 ;
        RECT 1405.370 1159.300 1405.690 1159.360 ;
        RECT 1406.290 1159.300 1406.610 1159.360 ;
        RECT 1405.370 1159.160 1406.610 1159.300 ;
        RECT 1405.370 1159.100 1405.690 1159.160 ;
        RECT 1406.290 1159.100 1406.610 1159.160 ;
        RECT 1534.630 1159.100 1534.950 1159.360 ;
        RECT 1534.720 1158.960 1534.860 1159.100 ;
        RECT 1535.090 1158.960 1535.410 1159.020 ;
        RECT 1534.720 1158.820 1535.410 1158.960 ;
        RECT 1535.090 1158.760 1535.410 1158.820 ;
        RECT 1534.630 1152.500 1534.950 1152.560 ;
        RECT 1535.090 1152.500 1535.410 1152.560 ;
        RECT 1534.630 1152.360 1535.410 1152.500 ;
        RECT 1534.630 1152.300 1534.950 1152.360 ;
        RECT 1535.090 1152.300 1535.410 1152.360 ;
        RECT 1358.450 1138.560 1358.770 1138.620 ;
        RECT 1359.370 1138.560 1359.690 1138.620 ;
        RECT 1358.450 1138.420 1359.690 1138.560 ;
        RECT 1358.450 1138.360 1358.770 1138.420 ;
        RECT 1359.370 1138.360 1359.690 1138.420 ;
        RECT 2518.570 1125.640 2518.890 1125.700 ;
        RECT 2518.570 1125.500 2519.260 1125.640 ;
        RECT 2518.570 1125.440 2518.890 1125.500 ;
        RECT 2519.120 1125.360 2519.260 1125.500 ;
        RECT 2519.030 1125.100 2519.350 1125.360 ;
        RECT 1277.950 1111.020 1278.270 1111.080 ;
        RECT 1278.410 1111.020 1278.730 1111.080 ;
        RECT 1277.950 1110.880 1278.730 1111.020 ;
        RECT 1277.950 1110.820 1278.270 1110.880 ;
        RECT 1278.410 1110.820 1278.730 1110.880 ;
        RECT 1405.370 1111.020 1405.690 1111.080 ;
        RECT 1405.830 1111.020 1406.150 1111.080 ;
        RECT 1405.370 1110.880 1406.150 1111.020 ;
        RECT 1405.370 1110.820 1405.690 1110.880 ;
        RECT 1405.830 1110.820 1406.150 1110.880 ;
        RECT 1543.370 1111.020 1543.690 1111.080 ;
        RECT 1543.370 1110.880 1544.060 1111.020 ;
        RECT 1543.370 1110.820 1543.690 1110.880 ;
        RECT 1543.920 1110.740 1544.060 1110.880 ;
        RECT 1069.570 1110.680 1069.890 1110.740 ;
        RECT 1070.950 1110.680 1071.270 1110.740 ;
        RECT 1069.570 1110.540 1071.270 1110.680 ;
        RECT 1069.570 1110.480 1069.890 1110.540 ;
        RECT 1070.950 1110.480 1071.270 1110.540 ;
        RECT 1535.090 1110.680 1535.410 1110.740 ;
        RECT 1535.550 1110.680 1535.870 1110.740 ;
        RECT 1535.090 1110.540 1535.870 1110.680 ;
        RECT 1535.090 1110.480 1535.410 1110.540 ;
        RECT 1535.550 1110.480 1535.870 1110.540 ;
        RECT 1543.830 1110.480 1544.150 1110.740 ;
        RECT 1543.370 1104.220 1543.690 1104.280 ;
        RECT 1543.830 1104.220 1544.150 1104.280 ;
        RECT 1543.370 1104.080 1544.150 1104.220 ;
        RECT 1543.370 1104.020 1543.690 1104.080 ;
        RECT 1543.830 1104.020 1544.150 1104.080 ;
        RECT 1358.450 1090.280 1358.770 1090.340 ;
        RECT 1359.830 1090.280 1360.150 1090.340 ;
        RECT 1358.450 1090.140 1360.150 1090.280 ;
        RECT 1358.450 1090.080 1358.770 1090.140 ;
        RECT 1359.830 1090.080 1360.150 1090.140 ;
        RECT 1541.530 1080.080 1541.850 1080.140 ;
        RECT 1543.370 1080.080 1543.690 1080.140 ;
        RECT 1541.530 1079.940 1543.690 1080.080 ;
        RECT 1541.530 1079.880 1541.850 1079.940 ;
        RECT 1543.370 1079.880 1543.690 1079.940 ;
        RECT 1292.670 1077.020 1292.990 1077.080 ;
        RECT 1292.300 1076.880 1292.990 1077.020 ;
        RECT 1292.300 1076.400 1292.440 1076.880 ;
        RECT 1292.670 1076.820 1292.990 1076.880 ;
        RECT 2518.110 1077.020 2518.430 1077.080 ;
        RECT 2519.950 1077.020 2520.270 1077.080 ;
        RECT 2518.110 1076.880 2520.270 1077.020 ;
        RECT 2518.110 1076.820 2518.430 1076.880 ;
        RECT 2519.950 1076.820 2520.270 1076.880 ;
        RECT 1405.830 1076.480 1406.150 1076.740 ;
        RECT 1292.210 1076.140 1292.530 1076.400 ;
        RECT 1405.920 1076.000 1406.060 1076.480 ;
        RECT 1486.330 1076.340 1486.650 1076.400 ;
        RECT 1490.010 1076.340 1490.330 1076.400 ;
        RECT 1486.330 1076.200 1490.330 1076.340 ;
        RECT 1486.330 1076.140 1486.650 1076.200 ;
        RECT 1490.010 1076.140 1490.330 1076.200 ;
        RECT 2518.110 1076.340 2518.430 1076.400 ;
        RECT 2519.950 1076.340 2520.270 1076.400 ;
        RECT 2518.110 1076.200 2520.270 1076.340 ;
        RECT 2518.110 1076.140 2518.430 1076.200 ;
        RECT 2519.950 1076.140 2520.270 1076.200 ;
        RECT 1406.290 1076.000 1406.610 1076.060 ;
        RECT 1405.920 1075.860 1406.610 1076.000 ;
        RECT 1406.290 1075.800 1406.610 1075.860 ;
        RECT 1070.950 1062.740 1071.270 1062.800 ;
        RECT 1071.870 1062.740 1072.190 1062.800 ;
        RECT 1070.950 1062.600 1072.190 1062.740 ;
        RECT 1070.950 1062.540 1071.270 1062.600 ;
        RECT 1071.870 1062.540 1072.190 1062.600 ;
        RECT 1277.950 1062.740 1278.270 1062.800 ;
        RECT 1278.410 1062.740 1278.730 1062.800 ;
        RECT 1277.950 1062.600 1278.730 1062.740 ;
        RECT 1277.950 1062.540 1278.270 1062.600 ;
        RECT 1278.410 1062.540 1278.730 1062.600 ;
        RECT 1288.990 1062.740 1289.310 1062.800 ;
        RECT 1289.910 1062.740 1290.230 1062.800 ;
        RECT 1288.990 1062.600 1290.230 1062.740 ;
        RECT 1288.990 1062.540 1289.310 1062.600 ;
        RECT 1289.910 1062.540 1290.230 1062.600 ;
        RECT 1357.530 1062.740 1357.850 1062.800 ;
        RECT 1359.830 1062.740 1360.150 1062.800 ;
        RECT 1357.530 1062.600 1360.150 1062.740 ;
        RECT 1357.530 1062.540 1357.850 1062.600 ;
        RECT 1359.830 1062.540 1360.150 1062.600 ;
        RECT 1378.230 1062.740 1378.550 1062.800 ;
        RECT 1379.610 1062.740 1379.930 1062.800 ;
        RECT 1378.230 1062.600 1379.930 1062.740 ;
        RECT 1378.230 1062.540 1378.550 1062.600 ;
        RECT 1379.610 1062.540 1379.930 1062.600 ;
        RECT 1535.090 1062.740 1535.410 1062.800 ;
        RECT 1536.010 1062.740 1536.330 1062.800 ;
        RECT 1535.090 1062.600 1536.330 1062.740 ;
        RECT 1535.090 1062.540 1535.410 1062.600 ;
        RECT 1536.010 1062.540 1536.330 1062.600 ;
        RECT 1277.950 1057.640 1278.270 1057.700 ;
        RECT 1280.710 1057.640 1281.030 1057.700 ;
        RECT 1277.950 1057.500 1281.030 1057.640 ;
        RECT 1277.950 1057.440 1278.270 1057.500 ;
        RECT 1280.710 1057.440 1281.030 1057.500 ;
        RECT 1489.090 1055.600 1489.410 1055.660 ;
        RECT 1519.450 1055.600 1519.770 1055.660 ;
        RECT 1489.090 1055.460 1519.770 1055.600 ;
        RECT 1489.090 1055.400 1489.410 1055.460 ;
        RECT 1519.450 1055.400 1519.770 1055.460 ;
        RECT 1342.350 1052.200 1342.670 1052.260 ;
        RECT 1344.190 1052.200 1344.510 1052.260 ;
        RECT 1342.350 1052.060 1344.510 1052.200 ;
        RECT 1342.350 1052.000 1342.670 1052.060 ;
        RECT 1344.190 1052.000 1344.510 1052.060 ;
        RECT 1454.590 1052.200 1454.910 1052.260 ;
        RECT 1455.510 1052.200 1455.830 1052.260 ;
        RECT 1454.590 1052.060 1455.830 1052.200 ;
        RECT 1454.590 1052.000 1454.910 1052.060 ;
        RECT 1455.510 1052.000 1455.830 1052.060 ;
        RECT 1488.630 1052.200 1488.950 1052.260 ;
        RECT 1559.930 1052.200 1560.250 1052.260 ;
        RECT 1488.630 1052.060 1560.250 1052.200 ;
        RECT 1488.630 1052.000 1488.950 1052.060 ;
        RECT 1559.930 1052.000 1560.250 1052.060 ;
        RECT 2518.570 1029.080 2518.890 1029.140 ;
        RECT 2518.570 1028.940 2519.260 1029.080 ;
        RECT 2518.570 1028.880 2518.890 1028.940 ;
        RECT 2519.120 1028.800 2519.260 1028.940 ;
        RECT 2519.030 1028.540 2519.350 1028.800 ;
        RECT 1486.330 1028.400 1486.650 1028.460 ;
        RECT 1489.090 1028.400 1489.410 1028.460 ;
        RECT 1486.330 1028.260 1489.410 1028.400 ;
        RECT 1486.330 1028.200 1486.650 1028.260 ;
        RECT 1489.090 1028.200 1489.410 1028.260 ;
        RECT 2518.570 1028.400 2518.890 1028.460 ;
        RECT 2519.950 1028.400 2520.270 1028.460 ;
        RECT 2518.570 1028.260 2520.270 1028.400 ;
        RECT 2518.570 1028.200 2518.890 1028.260 ;
        RECT 2519.950 1028.200 2520.270 1028.260 ;
        RECT 1541.990 1028.060 1542.310 1028.120 ;
        RECT 1542.910 1028.060 1543.230 1028.120 ;
        RECT 1541.990 1027.920 1543.230 1028.060 ;
        RECT 1541.990 1027.860 1542.310 1027.920 ;
        RECT 1542.910 1027.860 1543.230 1027.920 ;
        RECT 983.090 1025.680 983.410 1025.740 ;
        RECT 1152.830 1025.680 1153.150 1025.740 ;
        RECT 983.090 1025.540 1153.150 1025.680 ;
        RECT 983.090 1025.480 983.410 1025.540 ;
        RECT 1152.830 1025.480 1153.150 1025.540 ;
        RECT 975.730 1025.340 976.050 1025.400 ;
        RECT 1147.770 1025.340 1148.090 1025.400 ;
        RECT 975.730 1025.200 1148.090 1025.340 ;
        RECT 975.730 1025.140 976.050 1025.200 ;
        RECT 1147.770 1025.140 1148.090 1025.200 ;
        RECT 976.190 1025.000 976.510 1025.060 ;
        RECT 1156.050 1025.000 1156.370 1025.060 ;
        RECT 976.190 1024.860 1156.370 1025.000 ;
        RECT 976.190 1024.800 976.510 1024.860 ;
        RECT 1156.050 1024.800 1156.370 1024.860 ;
        RECT 1474.370 1025.000 1474.690 1025.060 ;
        RECT 1891.590 1025.000 1891.910 1025.060 ;
        RECT 1474.370 1024.860 1891.910 1025.000 ;
        RECT 1474.370 1024.800 1474.690 1024.860 ;
        RECT 1891.590 1024.800 1891.910 1024.860 ;
        RECT 982.630 1024.660 982.950 1024.720 ;
        RECT 1166.170 1024.660 1166.490 1024.720 ;
        RECT 982.630 1024.520 1166.490 1024.660 ;
        RECT 982.630 1024.460 982.950 1024.520 ;
        RECT 1166.170 1024.460 1166.490 1024.520 ;
        RECT 1187.330 1024.660 1187.650 1024.720 ;
        RECT 1188.710 1024.660 1189.030 1024.720 ;
        RECT 1187.330 1024.520 1189.030 1024.660 ;
        RECT 1187.330 1024.460 1187.650 1024.520 ;
        RECT 1188.710 1024.460 1189.030 1024.520 ;
        RECT 1431.130 1024.660 1431.450 1024.720 ;
        RECT 1891.130 1024.660 1891.450 1024.720 ;
        RECT 1431.130 1024.520 1891.450 1024.660 ;
        RECT 1431.130 1024.460 1431.450 1024.520 ;
        RECT 1891.130 1024.460 1891.450 1024.520 ;
        RECT 997.350 1021.260 997.670 1021.320 ;
        RECT 1223.670 1021.260 1223.990 1021.320 ;
        RECT 997.350 1021.120 1223.990 1021.260 ;
        RECT 997.350 1021.060 997.670 1021.120 ;
        RECT 1223.670 1021.060 1223.990 1021.120 ;
        RECT 1278.870 1021.260 1279.190 1021.320 ;
        RECT 1334.530 1021.260 1334.850 1021.320 ;
        RECT 1278.870 1021.120 1334.850 1021.260 ;
        RECT 1278.870 1021.060 1279.190 1021.120 ;
        RECT 1334.530 1021.060 1334.850 1021.120 ;
        RECT 1595.810 1021.260 1596.130 1021.320 ;
        RECT 1900.330 1021.260 1900.650 1021.320 ;
        RECT 1595.810 1021.120 1900.650 1021.260 ;
        RECT 1595.810 1021.060 1596.130 1021.120 ;
        RECT 1900.330 1021.060 1900.650 1021.120 ;
        RECT 988.150 1020.920 988.470 1020.980 ;
        RECT 1228.270 1020.920 1228.590 1020.980 ;
        RECT 988.150 1020.780 1228.590 1020.920 ;
        RECT 988.150 1020.720 988.470 1020.780 ;
        RECT 1228.270 1020.720 1228.590 1020.780 ;
        RECT 1252.650 1020.920 1252.970 1020.980 ;
        RECT 1339.130 1020.920 1339.450 1020.980 ;
        RECT 1252.650 1020.780 1339.450 1020.920 ;
        RECT 1252.650 1020.720 1252.970 1020.780 ;
        RECT 1339.130 1020.720 1339.450 1020.780 ;
        RECT 1567.750 1020.920 1568.070 1020.980 ;
        RECT 1890.670 1020.920 1890.990 1020.980 ;
        RECT 1567.750 1020.780 1890.990 1020.920 ;
        RECT 1567.750 1020.720 1568.070 1020.780 ;
        RECT 1890.670 1020.720 1890.990 1020.780 ;
        RECT 987.230 1020.580 987.550 1020.640 ;
        RECT 1259.550 1020.580 1259.870 1020.640 ;
        RECT 987.230 1020.440 1259.870 1020.580 ;
        RECT 987.230 1020.380 987.550 1020.440 ;
        RECT 1259.550 1020.380 1259.870 1020.440 ;
        RECT 1267.830 1020.580 1268.150 1020.640 ;
        RECT 1343.270 1020.580 1343.590 1020.640 ;
        RECT 1267.830 1020.440 1343.590 1020.580 ;
        RECT 1267.830 1020.380 1268.150 1020.440 ;
        RECT 1343.270 1020.380 1343.590 1020.440 ;
        RECT 1574.650 1020.580 1574.970 1020.640 ;
        RECT 1900.790 1020.580 1901.110 1020.640 ;
        RECT 1574.650 1020.440 1901.110 1020.580 ;
        RECT 1574.650 1020.380 1574.970 1020.440 ;
        RECT 1900.790 1020.380 1901.110 1020.440 ;
        RECT 996.890 1020.240 997.210 1020.300 ;
        RECT 1270.130 1020.240 1270.450 1020.300 ;
        RECT 996.890 1020.100 1270.450 1020.240 ;
        RECT 996.890 1020.040 997.210 1020.100 ;
        RECT 1270.130 1020.040 1270.450 1020.100 ;
        RECT 1279.790 1020.240 1280.110 1020.300 ;
        RECT 1341.890 1020.240 1342.210 1020.300 ;
        RECT 1279.790 1020.100 1342.210 1020.240 ;
        RECT 1279.790 1020.040 1280.110 1020.100 ;
        RECT 1341.890 1020.040 1342.210 1020.100 ;
        RECT 1541.990 1020.240 1542.310 1020.300 ;
        RECT 1886.070 1020.240 1886.390 1020.300 ;
        RECT 1541.990 1020.100 1886.390 1020.240 ;
        RECT 1541.990 1020.040 1542.310 1020.100 ;
        RECT 1886.070 1020.040 1886.390 1020.100 ;
        RECT 995.970 1019.900 996.290 1019.960 ;
        RECT 1292.210 1019.900 1292.530 1019.960 ;
        RECT 995.970 1019.760 1292.530 1019.900 ;
        RECT 995.970 1019.700 996.290 1019.760 ;
        RECT 1292.210 1019.700 1292.530 1019.760 ;
        RECT 1533.250 1019.900 1533.570 1019.960 ;
        RECT 1903.550 1019.900 1903.870 1019.960 ;
        RECT 1533.250 1019.760 1903.870 1019.900 ;
        RECT 1533.250 1019.700 1533.570 1019.760 ;
        RECT 1903.550 1019.700 1903.870 1019.760 ;
        RECT 988.610 1019.560 988.930 1019.620 ;
        RECT 1285.770 1019.560 1286.090 1019.620 ;
        RECT 988.610 1019.420 1286.090 1019.560 ;
        RECT 988.610 1019.360 988.930 1019.420 ;
        RECT 1285.770 1019.360 1286.090 1019.420 ;
        RECT 1299.110 1019.560 1299.430 1019.620 ;
        RECT 1335.910 1019.560 1336.230 1019.620 ;
        RECT 1299.110 1019.420 1336.230 1019.560 ;
        RECT 1299.110 1019.360 1299.430 1019.420 ;
        RECT 1335.910 1019.360 1336.230 1019.420 ;
        RECT 1507.030 1019.560 1507.350 1019.620 ;
        RECT 1897.570 1019.560 1897.890 1019.620 ;
        RECT 1507.030 1019.420 1897.890 1019.560 ;
        RECT 1507.030 1019.360 1507.350 1019.420 ;
        RECT 1897.570 1019.360 1897.890 1019.420 ;
        RECT 989.530 1019.220 989.850 1019.280 ;
        RECT 1301.870 1019.220 1302.190 1019.280 ;
        RECT 989.530 1019.080 1302.190 1019.220 ;
        RECT 989.530 1019.020 989.850 1019.080 ;
        RECT 1301.870 1019.020 1302.190 1019.080 ;
        RECT 1496.910 1019.220 1497.230 1019.280 ;
        RECT 1901.250 1019.220 1901.570 1019.280 ;
        RECT 1496.910 1019.080 1901.570 1019.220 ;
        RECT 1496.910 1019.020 1497.230 1019.080 ;
        RECT 1901.250 1019.020 1901.570 1019.080 ;
        RECT 990.910 1018.880 991.230 1018.940 ;
        RECT 1313.830 1018.880 1314.150 1018.940 ;
        RECT 990.910 1018.740 1314.150 1018.880 ;
        RECT 990.910 1018.680 991.230 1018.740 ;
        RECT 1313.830 1018.680 1314.150 1018.740 ;
        RECT 1462.410 1018.880 1462.730 1018.940 ;
        RECT 1898.950 1018.880 1899.270 1018.940 ;
        RECT 1462.410 1018.740 1899.270 1018.880 ;
        RECT 1462.410 1018.680 1462.730 1018.740 ;
        RECT 1898.950 1018.680 1899.270 1018.740 ;
        RECT 987.690 1018.540 988.010 1018.600 ;
        RECT 1314.750 1018.540 1315.070 1018.600 ;
        RECT 987.690 1018.400 1315.070 1018.540 ;
        RECT 987.690 1018.340 988.010 1018.400 ;
        RECT 1314.750 1018.340 1315.070 1018.400 ;
        RECT 1437.570 1018.540 1437.890 1018.600 ;
        RECT 1898.030 1018.540 1898.350 1018.600 ;
        RECT 1437.570 1018.400 1898.350 1018.540 ;
        RECT 1437.570 1018.340 1437.890 1018.400 ;
        RECT 1898.030 1018.340 1898.350 1018.400 ;
        RECT 989.070 1018.200 989.390 1018.260 ;
        RECT 1327.170 1018.200 1327.490 1018.260 ;
        RECT 989.070 1018.060 1327.490 1018.200 ;
        RECT 989.070 1018.000 989.390 1018.060 ;
        RECT 1327.170 1018.000 1327.490 1018.060 ;
        RECT 1358.910 1018.200 1359.230 1018.260 ;
        RECT 1849.270 1018.200 1849.590 1018.260 ;
        RECT 1358.910 1018.060 1849.590 1018.200 ;
        RECT 1358.910 1018.000 1359.230 1018.060 ;
        RECT 1849.270 1018.000 1849.590 1018.060 ;
        RECT 989.990 1017.860 990.310 1017.920 ;
        RECT 1335.910 1017.860 1336.230 1017.920 ;
        RECT 989.990 1017.720 1336.230 1017.860 ;
        RECT 989.990 1017.660 990.310 1017.720 ;
        RECT 1335.910 1017.660 1336.230 1017.720 ;
        RECT 1402.610 1017.860 1402.930 1017.920 ;
        RECT 1899.410 1017.860 1899.730 1017.920 ;
        RECT 1402.610 1017.720 1899.730 1017.860 ;
        RECT 1402.610 1017.660 1402.930 1017.720 ;
        RECT 1899.410 1017.660 1899.730 1017.720 ;
        RECT 990.450 1017.520 990.770 1017.580 ;
        RECT 1193.770 1017.520 1194.090 1017.580 ;
        RECT 990.450 1017.380 1194.090 1017.520 ;
        RECT 990.450 1017.320 990.770 1017.380 ;
        RECT 1193.770 1017.320 1194.090 1017.380 ;
        RECT 1204.810 1017.520 1205.130 1017.580 ;
        RECT 1342.810 1017.520 1343.130 1017.580 ;
        RECT 1204.810 1017.380 1343.130 1017.520 ;
        RECT 1204.810 1017.320 1205.130 1017.380 ;
        RECT 1342.810 1017.320 1343.130 1017.380 ;
        RECT 1480.810 1017.520 1481.130 1017.580 ;
        RECT 1766.470 1017.520 1766.790 1017.580 ;
        RECT 1480.810 1017.380 1766.790 1017.520 ;
        RECT 1480.810 1017.320 1481.130 1017.380 ;
        RECT 1766.470 1017.320 1766.790 1017.380 ;
        RECT 1048.410 1017.180 1048.730 1017.240 ;
        RECT 1215.850 1017.180 1216.170 1017.240 ;
        RECT 1048.410 1017.040 1216.170 1017.180 ;
        RECT 1048.410 1016.980 1048.730 1017.040 ;
        RECT 1215.850 1016.980 1216.170 1017.040 ;
        RECT 1472.070 1017.180 1472.390 1017.240 ;
        RECT 1704.370 1017.180 1704.690 1017.240 ;
        RECT 1472.070 1017.040 1704.690 1017.180 ;
        RECT 1472.070 1016.980 1472.390 1017.040 ;
        RECT 1704.370 1016.980 1704.690 1017.040 ;
        RECT 991.830 1016.840 992.150 1016.900 ;
        RECT 1125.690 1016.840 1126.010 1016.900 ;
        RECT 991.830 1016.700 1126.010 1016.840 ;
        RECT 991.830 1016.640 992.150 1016.700 ;
        RECT 1125.690 1016.640 1126.010 1016.700 ;
        RECT 1514.390 1016.840 1514.710 1016.900 ;
        RECT 1656.070 1016.840 1656.390 1016.900 ;
        RECT 1514.390 1016.700 1656.390 1016.840 ;
        RECT 1514.390 1016.640 1514.710 1016.700 ;
        RECT 1656.070 1016.640 1656.390 1016.700 ;
        RECT 1489.550 1016.500 1489.870 1016.560 ;
        RECT 1625.710 1016.500 1626.030 1016.560 ;
        RECT 1489.550 1016.360 1626.030 1016.500 ;
        RECT 1489.550 1016.300 1489.870 1016.360 ;
        RECT 1625.710 1016.300 1626.030 1016.360 ;
        RECT 1576.030 1016.160 1576.350 1016.220 ;
        RECT 1679.990 1016.160 1680.310 1016.220 ;
        RECT 1576.030 1016.020 1680.310 1016.160 ;
        RECT 1576.030 1015.960 1576.350 1016.020 ;
        RECT 1679.990 1015.960 1680.310 1016.020 ;
        RECT 1544.750 1015.820 1545.070 1015.880 ;
        RECT 1608.690 1015.820 1609.010 1015.880 ;
        RECT 1544.750 1015.680 1609.010 1015.820 ;
        RECT 1544.750 1015.620 1545.070 1015.680 ;
        RECT 1608.690 1015.620 1609.010 1015.680 ;
        RECT 1294.050 1014.460 1294.370 1014.520 ;
        RECT 1292.760 1014.320 1294.370 1014.460 ;
        RECT 983.550 1014.120 983.870 1014.180 ;
        RECT 1104.070 1014.120 1104.390 1014.180 ;
        RECT 1106.370 1014.120 1106.690 1014.180 ;
        RECT 983.550 1013.980 1103.840 1014.120 ;
        RECT 983.550 1013.920 983.870 1013.980 ;
        RECT 976.650 1013.780 976.970 1013.840 ;
        RECT 1103.150 1013.780 1103.470 1013.840 ;
        RECT 976.650 1013.640 1103.470 1013.780 ;
        RECT 1103.700 1013.780 1103.840 1013.980 ;
        RECT 1104.070 1013.980 1106.690 1014.120 ;
        RECT 1104.070 1013.920 1104.390 1013.980 ;
        RECT 1106.370 1013.920 1106.690 1013.980 ;
        RECT 1198.370 1014.120 1198.690 1014.180 ;
        RECT 1200.670 1014.120 1200.990 1014.180 ;
        RECT 1198.370 1013.980 1200.990 1014.120 ;
        RECT 1198.370 1013.920 1198.690 1013.980 ;
        RECT 1200.670 1013.920 1200.990 1013.980 ;
        RECT 1202.510 1014.120 1202.830 1014.180 ;
        RECT 1210.790 1014.120 1211.110 1014.180 ;
        RECT 1202.510 1013.980 1211.110 1014.120 ;
        RECT 1202.510 1013.920 1202.830 1013.980 ;
        RECT 1210.790 1013.920 1211.110 1013.980 ;
        RECT 1211.250 1014.120 1211.570 1014.180 ;
        RECT 1214.010 1014.120 1214.330 1014.180 ;
        RECT 1211.250 1013.980 1214.330 1014.120 ;
        RECT 1211.250 1013.920 1211.570 1013.980 ;
        RECT 1214.010 1013.920 1214.330 1013.980 ;
        RECT 1257.250 1014.120 1257.570 1014.180 ;
        RECT 1292.760 1014.120 1292.900 1014.320 ;
        RECT 1294.050 1014.260 1294.370 1014.320 ;
        RECT 1294.970 1014.120 1295.290 1014.180 ;
        RECT 1257.250 1013.980 1292.900 1014.120 ;
        RECT 1293.220 1013.980 1295.290 1014.120 ;
        RECT 1257.250 1013.920 1257.570 1013.980 ;
        RECT 1134.430 1013.780 1134.750 1013.840 ;
        RECT 1103.700 1013.640 1134.750 1013.780 ;
        RECT 976.650 1013.580 976.970 1013.640 ;
        RECT 1103.150 1013.580 1103.470 1013.640 ;
        RECT 1134.430 1013.580 1134.750 1013.640 ;
        RECT 1181.810 1013.780 1182.130 1013.840 ;
        RECT 1293.220 1013.780 1293.360 1013.980 ;
        RECT 1294.970 1013.920 1295.290 1013.980 ;
        RECT 1300.490 1014.120 1300.810 1014.180 ;
        RECT 1317.970 1014.120 1318.290 1014.180 ;
        RECT 1300.490 1013.980 1318.290 1014.120 ;
        RECT 1300.490 1013.920 1300.810 1013.980 ;
        RECT 1317.970 1013.920 1318.290 1013.980 ;
        RECT 1331.310 1014.120 1331.630 1014.180 ;
        RECT 1346.950 1014.120 1347.270 1014.180 ;
        RECT 1331.310 1013.980 1347.270 1014.120 ;
        RECT 1331.310 1013.920 1331.630 1013.980 ;
        RECT 1346.950 1013.920 1347.270 1013.980 ;
        RECT 1446.310 1014.120 1446.630 1014.180 ;
        RECT 1448.610 1014.120 1448.930 1014.180 ;
        RECT 1446.310 1013.980 1448.930 1014.120 ;
        RECT 1446.310 1013.920 1446.630 1013.980 ;
        RECT 1448.610 1013.920 1448.930 1013.980 ;
        RECT 1452.750 1014.120 1453.070 1014.180 ;
        RECT 1455.050 1014.120 1455.370 1014.180 ;
        RECT 1452.750 1013.980 1455.370 1014.120 ;
        RECT 1452.750 1013.920 1453.070 1013.980 ;
        RECT 1455.050 1013.920 1455.370 1013.980 ;
        RECT 1456.890 1014.120 1457.210 1014.180 ;
        RECT 1461.950 1014.120 1462.270 1014.180 ;
        RECT 1456.890 1013.980 1462.270 1014.120 ;
        RECT 1456.890 1013.920 1457.210 1013.980 ;
        RECT 1461.950 1013.920 1462.270 1013.980 ;
        RECT 1465.630 1014.120 1465.950 1014.180 ;
        RECT 1469.310 1014.120 1469.630 1014.180 ;
        RECT 1465.630 1013.980 1469.630 1014.120 ;
        RECT 1465.630 1013.920 1465.950 1013.980 ;
        RECT 1469.310 1013.920 1469.630 1013.980 ;
        RECT 1478.970 1014.120 1479.290 1014.180 ;
        RECT 1482.190 1014.120 1482.510 1014.180 ;
        RECT 1478.970 1013.980 1482.510 1014.120 ;
        RECT 1478.970 1013.920 1479.290 1013.980 ;
        RECT 1482.190 1013.920 1482.510 1013.980 ;
        RECT 1500.590 1014.120 1500.910 1014.180 ;
        RECT 1503.350 1014.120 1503.670 1014.180 ;
        RECT 1535.550 1014.120 1535.870 1014.180 ;
        RECT 1500.590 1013.980 1503.670 1014.120 ;
        RECT 1500.590 1013.920 1500.910 1013.980 ;
        RECT 1503.350 1013.920 1503.670 1013.980 ;
        RECT 1504.820 1013.980 1535.870 1014.120 ;
        RECT 1181.810 1013.640 1293.360 1013.780 ;
        RECT 1293.590 1013.780 1293.910 1013.840 ;
        RECT 1319.350 1013.780 1319.670 1013.840 ;
        RECT 1293.590 1013.640 1319.670 1013.780 ;
        RECT 1181.810 1013.580 1182.130 1013.640 ;
        RECT 1293.590 1013.580 1293.910 1013.640 ;
        RECT 1319.350 1013.580 1319.670 1013.640 ;
        RECT 1324.410 1013.780 1324.730 1013.840 ;
        RECT 1347.410 1013.780 1347.730 1013.840 ;
        RECT 1324.410 1013.640 1347.730 1013.780 ;
        RECT 1324.410 1013.580 1324.730 1013.640 ;
        RECT 1347.410 1013.580 1347.730 1013.640 ;
        RECT 1497.370 1013.780 1497.690 1013.840 ;
        RECT 1504.820 1013.780 1504.960 1013.980 ;
        RECT 1535.550 1013.920 1535.870 1013.980 ;
        RECT 1559.470 1014.120 1559.790 1014.180 ;
        RECT 1562.690 1014.120 1563.010 1014.180 ;
        RECT 1559.470 1013.980 1563.010 1014.120 ;
        RECT 1559.470 1013.920 1559.790 1013.980 ;
        RECT 1562.690 1013.920 1563.010 1013.980 ;
        RECT 1563.150 1014.120 1563.470 1014.180 ;
        RECT 1595.810 1014.120 1596.130 1014.180 ;
        RECT 1563.150 1013.980 1596.130 1014.120 ;
        RECT 1563.150 1013.920 1563.470 1013.980 ;
        RECT 1595.810 1013.920 1596.130 1013.980 ;
        RECT 1596.270 1014.120 1596.590 1014.180 ;
        RECT 1600.410 1014.120 1600.730 1014.180 ;
        RECT 1596.270 1013.980 1600.730 1014.120 ;
        RECT 1596.270 1013.920 1596.590 1013.980 ;
        RECT 1600.410 1013.920 1600.730 1013.980 ;
        RECT 1754.970 1014.120 1755.290 1014.180 ;
        RECT 1759.110 1014.120 1759.430 1014.180 ;
        RECT 1754.970 1013.980 1759.430 1014.120 ;
        RECT 1754.970 1013.920 1755.290 1013.980 ;
        RECT 1759.110 1013.920 1759.430 1013.980 ;
        RECT 1763.710 1014.120 1764.030 1014.180 ;
        RECT 1766.010 1014.120 1766.330 1014.180 ;
        RECT 1763.710 1013.980 1766.330 1014.120 ;
        RECT 1763.710 1013.920 1764.030 1013.980 ;
        RECT 1766.010 1013.920 1766.330 1013.980 ;
        RECT 1766.470 1014.120 1766.790 1014.180 ;
        RECT 2065.010 1014.120 2065.330 1014.180 ;
        RECT 1766.470 1013.980 2065.330 1014.120 ;
        RECT 1766.470 1013.920 1766.790 1013.980 ;
        RECT 2065.010 1013.920 2065.330 1013.980 ;
        RECT 2065.470 1014.120 2065.790 1014.180 ;
        RECT 2073.290 1014.120 2073.610 1014.180 ;
        RECT 2065.470 1013.980 2073.610 1014.120 ;
        RECT 2065.470 1013.920 2065.790 1013.980 ;
        RECT 2073.290 1013.920 2073.610 1013.980 ;
        RECT 2075.130 1014.120 2075.450 1014.180 ;
        RECT 2087.090 1014.120 2087.410 1014.180 ;
        RECT 2075.130 1013.980 2087.410 1014.120 ;
        RECT 2075.130 1013.920 2075.450 1013.980 ;
        RECT 2087.090 1013.920 2087.410 1013.980 ;
        RECT 2087.550 1014.120 2087.870 1014.180 ;
        RECT 2090.310 1014.120 2090.630 1014.180 ;
        RECT 2087.550 1013.980 2090.630 1014.120 ;
        RECT 2087.550 1013.920 2087.870 1013.980 ;
        RECT 2090.310 1013.920 2090.630 1013.980 ;
        RECT 1497.370 1013.640 1504.960 1013.780 ;
        RECT 1505.190 1013.780 1505.510 1013.840 ;
        RECT 1536.010 1013.780 1536.330 1013.840 ;
        RECT 1505.190 1013.640 1536.330 1013.780 ;
        RECT 1497.370 1013.580 1497.690 1013.640 ;
        RECT 1505.190 1013.580 1505.510 1013.640 ;
        RECT 1536.010 1013.580 1536.330 1013.640 ;
        RECT 1552.110 1013.780 1552.430 1013.840 ;
        RECT 1878.250 1013.780 1878.570 1013.840 ;
        RECT 1552.110 1013.640 1878.570 1013.780 ;
        RECT 1552.110 1013.580 1552.430 1013.640 ;
        RECT 1878.250 1013.580 1878.570 1013.640 ;
        RECT 1878.710 1013.780 1879.030 1013.840 ;
        RECT 1893.890 1013.780 1894.210 1013.840 ;
        RECT 1878.710 1013.640 1894.210 1013.780 ;
        RECT 1878.710 1013.580 1879.030 1013.640 ;
        RECT 1893.890 1013.580 1894.210 1013.640 ;
        RECT 2002.910 1013.780 2003.230 1013.840 ;
        RECT 2007.510 1013.780 2007.830 1013.840 ;
        RECT 2002.910 1013.640 2007.830 1013.780 ;
        RECT 2002.910 1013.580 2003.230 1013.640 ;
        RECT 2007.510 1013.580 2007.830 1013.640 ;
        RECT 2007.970 1013.780 2008.290 1013.840 ;
        RECT 2294.090 1013.780 2294.410 1013.840 ;
        RECT 2007.970 1013.640 2294.410 1013.780 ;
        RECT 2007.970 1013.580 2008.290 1013.640 ;
        RECT 2294.090 1013.580 2294.410 1013.640 ;
        RECT 1000.110 1013.440 1000.430 1013.500 ;
        RECT 1191.010 1013.440 1191.330 1013.500 ;
        RECT 1000.110 1013.300 1191.330 1013.440 ;
        RECT 1000.110 1013.240 1000.430 1013.300 ;
        RECT 1191.010 1013.240 1191.330 1013.300 ;
        RECT 1203.890 1013.440 1204.210 1013.500 ;
        RECT 1211.710 1013.440 1212.030 1013.500 ;
        RECT 1203.890 1013.300 1212.030 1013.440 ;
        RECT 1203.890 1013.240 1204.210 1013.300 ;
        RECT 1211.710 1013.240 1212.030 1013.300 ;
        RECT 1254.490 1013.440 1254.810 1013.500 ;
        RECT 1346.030 1013.440 1346.350 1013.500 ;
        RECT 1254.490 1013.300 1346.350 1013.440 ;
        RECT 1254.490 1013.240 1254.810 1013.300 ;
        RECT 1346.030 1013.240 1346.350 1013.300 ;
        RECT 1495.530 1013.440 1495.850 1013.500 ;
        RECT 1524.970 1013.440 1525.290 1013.500 ;
        RECT 1495.530 1013.300 1525.290 1013.440 ;
        RECT 1495.530 1013.240 1495.850 1013.300 ;
        RECT 1524.970 1013.240 1525.290 1013.300 ;
        RECT 1534.630 1013.440 1534.950 1013.500 ;
        RECT 1603.170 1013.440 1603.490 1013.500 ;
        RECT 1534.630 1013.300 1603.490 1013.440 ;
        RECT 1534.630 1013.240 1534.950 1013.300 ;
        RECT 1603.170 1013.240 1603.490 1013.300 ;
        RECT 1720.010 1013.440 1720.330 1013.500 ;
        RECT 1749.910 1013.440 1750.230 1013.500 ;
        RECT 1752.210 1013.440 1752.530 1013.500 ;
        RECT 1720.010 1013.300 1739.100 1013.440 ;
        RECT 1720.010 1013.240 1720.330 1013.300 ;
        RECT 782.990 1013.100 783.310 1013.160 ;
        RECT 845.550 1013.100 845.870 1013.160 ;
        RECT 782.990 1012.960 845.870 1013.100 ;
        RECT 782.990 1012.900 783.310 1012.960 ;
        RECT 845.550 1012.900 845.870 1012.960 ;
        RECT 991.370 1013.100 991.690 1013.160 ;
        RECT 1014.370 1013.100 1014.690 1013.160 ;
        RECT 991.370 1012.960 1014.690 1013.100 ;
        RECT 991.370 1012.900 991.690 1012.960 ;
        RECT 1014.370 1012.900 1014.690 1012.960 ;
        RECT 1038.290 1013.100 1038.610 1013.160 ;
        RECT 1196.530 1013.100 1196.850 1013.160 ;
        RECT 1038.290 1012.960 1196.850 1013.100 ;
        RECT 1038.290 1012.900 1038.610 1012.960 ;
        RECT 1196.530 1012.900 1196.850 1012.960 ;
        RECT 1196.990 1013.100 1197.310 1013.160 ;
        RECT 1219.070 1013.100 1219.390 1013.160 ;
        RECT 1196.990 1012.960 1219.390 1013.100 ;
        RECT 1196.990 1012.900 1197.310 1012.960 ;
        RECT 1219.070 1012.900 1219.390 1012.960 ;
        RECT 1244.830 1013.100 1245.150 1013.160 ;
        RECT 1340.510 1013.100 1340.830 1013.160 ;
        RECT 1244.830 1012.960 1340.830 1013.100 ;
        RECT 1244.830 1012.900 1245.150 1012.960 ;
        RECT 1340.510 1012.900 1340.830 1012.960 ;
        RECT 1419.630 1013.100 1419.950 1013.160 ;
        RECT 1421.010 1013.100 1421.330 1013.160 ;
        RECT 1419.630 1012.960 1421.330 1013.100 ;
        RECT 1419.630 1012.900 1419.950 1012.960 ;
        RECT 1421.010 1012.900 1421.330 1012.960 ;
        RECT 1495.070 1013.100 1495.390 1013.160 ;
        RECT 1528.190 1013.100 1528.510 1013.160 ;
        RECT 1495.070 1012.960 1528.510 1013.100 ;
        RECT 1495.070 1012.900 1495.390 1012.960 ;
        RECT 1528.190 1012.900 1528.510 1012.960 ;
        RECT 1536.010 1013.100 1536.330 1013.160 ;
        RECT 1547.510 1013.100 1547.830 1013.160 ;
        RECT 1536.010 1012.960 1547.830 1013.100 ;
        RECT 1536.010 1012.900 1536.330 1012.960 ;
        RECT 1547.510 1012.900 1547.830 1012.960 ;
        RECT 1555.790 1013.100 1556.110 1013.160 ;
        RECT 1659.290 1013.100 1659.610 1013.160 ;
        RECT 1555.790 1012.960 1659.610 1013.100 ;
        RECT 1555.790 1012.900 1556.110 1012.960 ;
        RECT 1659.290 1012.900 1659.610 1012.960 ;
        RECT 1710.350 1013.100 1710.670 1013.160 ;
        RECT 1710.350 1012.960 1738.640 1013.100 ;
        RECT 1710.350 1012.900 1710.670 1012.960 ;
        RECT 769.190 1012.760 769.510 1012.820 ;
        RECT 890.170 1012.760 890.490 1012.820 ;
        RECT 769.190 1012.620 890.490 1012.760 ;
        RECT 769.190 1012.560 769.510 1012.620 ;
        RECT 890.170 1012.560 890.490 1012.620 ;
        RECT 984.930 1012.760 985.250 1012.820 ;
        RECT 1207.570 1012.760 1207.890 1012.820 ;
        RECT 984.930 1012.620 1207.890 1012.760 ;
        RECT 984.930 1012.560 985.250 1012.620 ;
        RECT 1207.570 1012.560 1207.890 1012.620 ;
        RECT 1237.470 1012.760 1237.790 1012.820 ;
        RECT 1269.210 1012.760 1269.530 1012.820 ;
        RECT 1339.590 1012.760 1339.910 1012.820 ;
        RECT 1237.470 1012.620 1268.980 1012.760 ;
        RECT 1237.470 1012.560 1237.790 1012.620 ;
        RECT 650.510 1012.420 650.830 1012.480 ;
        RECT 672.130 1012.420 672.450 1012.480 ;
        RECT 650.510 1012.280 672.450 1012.420 ;
        RECT 650.510 1012.220 650.830 1012.280 ;
        RECT 672.130 1012.220 672.450 1012.280 ;
        RECT 762.290 1012.420 762.610 1012.480 ;
        RECT 884.650 1012.420 884.970 1012.480 ;
        RECT 762.290 1012.280 884.970 1012.420 ;
        RECT 762.290 1012.220 762.610 1012.280 ;
        RECT 884.650 1012.220 884.970 1012.280 ;
        RECT 977.570 1012.420 977.890 1012.480 ;
        RECT 1205.270 1012.420 1205.590 1012.480 ;
        RECT 977.570 1012.280 1205.590 1012.420 ;
        RECT 977.570 1012.220 977.890 1012.280 ;
        RECT 1205.270 1012.220 1205.590 1012.280 ;
        RECT 1218.610 1012.420 1218.930 1012.480 ;
        RECT 1263.230 1012.420 1263.550 1012.480 ;
        RECT 1218.610 1012.280 1263.550 1012.420 ;
        RECT 1268.840 1012.420 1268.980 1012.620 ;
        RECT 1269.210 1012.620 1339.910 1012.760 ;
        RECT 1269.210 1012.560 1269.530 1012.620 ;
        RECT 1339.590 1012.560 1339.910 1012.620 ;
        RECT 1496.450 1012.760 1496.770 1012.820 ;
        RECT 1511.170 1012.760 1511.490 1012.820 ;
        RECT 1496.450 1012.620 1511.490 1012.760 ;
        RECT 1496.450 1012.560 1496.770 1012.620 ;
        RECT 1511.170 1012.560 1511.490 1012.620 ;
        RECT 1511.630 1012.760 1511.950 1012.820 ;
        RECT 1514.850 1012.760 1515.170 1012.820 ;
        RECT 1511.630 1012.620 1515.170 1012.760 ;
        RECT 1511.630 1012.560 1511.950 1012.620 ;
        RECT 1514.850 1012.560 1515.170 1012.620 ;
        RECT 1536.470 1012.760 1536.790 1012.820 ;
        RECT 1628.470 1012.760 1628.790 1012.820 ;
        RECT 1536.470 1012.620 1628.790 1012.760 ;
        RECT 1536.470 1012.560 1536.790 1012.620 ;
        RECT 1628.470 1012.560 1628.790 1012.620 ;
        RECT 1270.590 1012.420 1270.910 1012.480 ;
        RECT 1331.310 1012.420 1331.630 1012.480 ;
        RECT 1268.840 1012.280 1269.440 1012.420 ;
        RECT 1218.610 1012.220 1218.930 1012.280 ;
        RECT 1263.230 1012.220 1263.550 1012.280 ;
        RECT 755.390 1012.080 755.710 1012.140 ;
        RECT 910.870 1012.080 911.190 1012.140 ;
        RECT 755.390 1011.940 911.190 1012.080 ;
        RECT 755.390 1011.880 755.710 1011.940 ;
        RECT 910.870 1011.880 911.190 1011.940 ;
        RECT 999.650 1012.080 999.970 1012.140 ;
        RECT 1232.410 1012.080 1232.730 1012.140 ;
        RECT 999.650 1011.940 1232.730 1012.080 ;
        RECT 999.650 1011.880 999.970 1011.940 ;
        RECT 1232.410 1011.880 1232.730 1011.940 ;
        RECT 686.390 1011.740 686.710 1011.800 ;
        RECT 841.870 1011.740 842.190 1011.800 ;
        RECT 686.390 1011.600 842.190 1011.740 ;
        RECT 686.390 1011.540 686.710 1011.600 ;
        RECT 841.870 1011.540 842.190 1011.600 ;
        RECT 978.030 1011.740 978.350 1011.800 ;
        RECT 1225.970 1011.740 1226.290 1011.800 ;
        RECT 978.030 1011.600 1226.290 1011.740 ;
        RECT 978.030 1011.540 978.350 1011.600 ;
        RECT 1225.970 1011.540 1226.290 1011.600 ;
        RECT 1237.930 1011.740 1238.250 1011.800 ;
        RECT 1267.370 1011.740 1267.690 1011.800 ;
        RECT 1237.930 1011.600 1267.690 1011.740 ;
        RECT 1269.300 1011.740 1269.440 1012.280 ;
        RECT 1270.590 1012.280 1331.630 1012.420 ;
        RECT 1270.590 1012.220 1270.910 1012.280 ;
        RECT 1331.310 1012.220 1331.630 1012.280 ;
        RECT 1338.210 1012.420 1338.530 1012.480 ;
        RECT 1346.490 1012.420 1346.810 1012.480 ;
        RECT 1338.210 1012.280 1346.810 1012.420 ;
        RECT 1338.210 1012.220 1338.530 1012.280 ;
        RECT 1346.490 1012.220 1346.810 1012.280 ;
        RECT 1369.950 1012.420 1370.270 1012.480 ;
        RECT 1372.710 1012.420 1373.030 1012.480 ;
        RECT 1369.950 1012.280 1373.030 1012.420 ;
        RECT 1369.950 1012.220 1370.270 1012.280 ;
        RECT 1372.710 1012.220 1373.030 1012.280 ;
        RECT 1404.910 1012.420 1405.230 1012.480 ;
        RECT 1406.290 1012.420 1406.610 1012.480 ;
        RECT 1404.910 1012.280 1406.610 1012.420 ;
        RECT 1404.910 1012.220 1405.230 1012.280 ;
        RECT 1406.290 1012.220 1406.610 1012.280 ;
        RECT 1411.350 1012.420 1411.670 1012.480 ;
        RECT 1413.650 1012.420 1413.970 1012.480 ;
        RECT 1411.350 1012.280 1413.970 1012.420 ;
        RECT 1411.350 1012.220 1411.670 1012.280 ;
        RECT 1413.650 1012.220 1413.970 1012.280 ;
        RECT 1444.010 1012.420 1444.330 1012.480 ;
        RECT 1576.490 1012.420 1576.810 1012.480 ;
        RECT 1444.010 1012.280 1576.810 1012.420 ;
        RECT 1444.010 1012.220 1444.330 1012.280 ;
        RECT 1576.490 1012.220 1576.810 1012.280 ;
        RECT 1665.730 1012.420 1666.050 1012.480 ;
        RECT 1669.410 1012.420 1669.730 1012.480 ;
        RECT 1665.730 1012.280 1669.730 1012.420 ;
        RECT 1665.730 1012.220 1666.050 1012.280 ;
        RECT 1669.410 1012.220 1669.730 1012.280 ;
        RECT 1707.130 1012.420 1707.450 1012.480 ;
        RECT 1710.810 1012.420 1711.130 1012.480 ;
        RECT 1707.130 1012.280 1711.130 1012.420 ;
        RECT 1707.130 1012.220 1707.450 1012.280 ;
        RECT 1710.810 1012.220 1711.130 1012.280 ;
        RECT 1715.870 1012.420 1716.190 1012.480 ;
        RECT 1717.710 1012.420 1718.030 1012.480 ;
        RECT 1715.870 1012.280 1718.030 1012.420 ;
        RECT 1715.870 1012.220 1716.190 1012.280 ;
        RECT 1717.710 1012.220 1718.030 1012.280 ;
        RECT 1733.350 1012.420 1733.670 1012.480 ;
        RECT 1737.950 1012.420 1738.270 1012.480 ;
        RECT 1733.350 1012.280 1738.270 1012.420 ;
        RECT 1738.500 1012.420 1738.640 1012.960 ;
        RECT 1738.960 1012.760 1739.100 1013.300 ;
        RECT 1749.910 1013.300 1752.530 1013.440 ;
        RECT 1749.910 1013.240 1750.230 1013.300 ;
        RECT 1752.210 1013.240 1752.530 1013.300 ;
        RECT 1758.650 1013.440 1758.970 1013.500 ;
        RECT 1766.470 1013.440 1766.790 1013.500 ;
        RECT 2064.550 1013.440 2064.870 1013.500 ;
        RECT 1758.650 1013.300 1766.790 1013.440 ;
        RECT 1758.650 1013.240 1758.970 1013.300 ;
        RECT 1766.470 1013.240 1766.790 1013.300 ;
        RECT 1767.020 1013.300 2064.870 1013.440 ;
        RECT 1741.630 1013.100 1741.950 1013.160 ;
        RECT 1767.020 1013.100 1767.160 1013.300 ;
        RECT 2064.550 1013.240 2064.870 1013.300 ;
        RECT 2065.010 1013.440 2065.330 1013.500 ;
        RECT 2086.630 1013.440 2086.950 1013.500 ;
        RECT 2065.010 1013.300 2086.950 1013.440 ;
        RECT 2065.010 1013.240 2065.330 1013.300 ;
        RECT 2086.630 1013.240 2086.950 1013.300 ;
        RECT 1741.630 1012.960 1767.160 1013.100 ;
        RECT 1767.390 1013.100 1767.710 1013.160 ;
        RECT 2085.710 1013.100 2086.030 1013.160 ;
        RECT 1767.390 1012.960 2086.030 1013.100 ;
        RECT 1741.630 1012.900 1741.950 1012.960 ;
        RECT 1767.390 1012.900 1767.710 1012.960 ;
        RECT 2085.710 1012.900 2086.030 1012.960 ;
        RECT 2084.330 1012.760 2084.650 1012.820 ;
        RECT 1738.960 1012.620 2084.650 1012.760 ;
        RECT 2084.330 1012.560 2084.650 1012.620 ;
        RECT 2064.090 1012.420 2064.410 1012.480 ;
        RECT 1738.500 1012.280 2064.410 1012.420 ;
        RECT 1733.350 1012.220 1733.670 1012.280 ;
        RECT 1737.950 1012.220 1738.270 1012.280 ;
        RECT 2064.090 1012.220 2064.410 1012.280 ;
        RECT 2064.550 1012.420 2064.870 1012.480 ;
        RECT 2086.170 1012.420 2086.490 1012.480 ;
        RECT 2064.550 1012.280 2086.490 1012.420 ;
        RECT 2064.550 1012.220 2064.870 1012.280 ;
        RECT 2086.170 1012.220 2086.490 1012.280 ;
        RECT 1269.670 1012.080 1269.990 1012.140 ;
        RECT 1340.050 1012.080 1340.370 1012.140 ;
        RECT 1269.670 1011.940 1340.370 1012.080 ;
        RECT 1269.670 1011.880 1269.990 1011.940 ;
        RECT 1340.050 1011.880 1340.370 1011.940 ;
        RECT 1495.990 1012.080 1496.310 1012.140 ;
        RECT 1534.630 1012.080 1534.950 1012.140 ;
        RECT 1495.990 1011.940 1534.950 1012.080 ;
        RECT 1495.990 1011.880 1496.310 1011.940 ;
        RECT 1534.630 1011.880 1534.950 1011.940 ;
        RECT 1535.090 1012.080 1535.410 1012.140 ;
        RECT 1537.850 1012.080 1538.170 1012.140 ;
        RECT 1535.090 1011.940 1538.170 1012.080 ;
        RECT 1535.090 1011.880 1535.410 1011.940 ;
        RECT 1537.850 1011.880 1538.170 1011.940 ;
        RECT 1552.570 1012.080 1552.890 1012.140 ;
        RECT 1556.250 1012.080 1556.570 1012.140 ;
        RECT 1552.570 1011.940 1556.570 1012.080 ;
        RECT 1552.570 1011.880 1552.890 1011.940 ;
        RECT 1556.250 1011.880 1556.570 1011.940 ;
        RECT 1556.710 1012.080 1557.030 1012.140 ;
        RECT 1628.470 1012.080 1628.790 1012.140 ;
        RECT 1556.710 1011.940 1628.790 1012.080 ;
        RECT 1556.710 1011.880 1557.030 1011.940 ;
        RECT 1628.470 1011.880 1628.790 1011.940 ;
        RECT 1662.510 1012.080 1662.830 1012.140 ;
        RECT 2075.130 1012.080 2075.450 1012.140 ;
        RECT 1662.510 1011.940 2075.450 1012.080 ;
        RECT 1662.510 1011.880 1662.830 1011.940 ;
        RECT 2075.130 1011.880 2075.450 1011.940 ;
        RECT 2078.810 1012.080 2079.130 1012.140 ;
        RECT 2083.410 1012.080 2083.730 1012.140 ;
        RECT 2078.810 1011.940 2083.730 1012.080 ;
        RECT 2078.810 1011.880 2079.130 1011.940 ;
        RECT 2083.410 1011.880 2083.730 1011.940 ;
        RECT 1330.390 1011.740 1330.710 1011.800 ;
        RECT 1269.300 1011.600 1330.710 1011.740 ;
        RECT 1237.930 1011.540 1238.250 1011.600 ;
        RECT 1267.370 1011.540 1267.690 1011.600 ;
        RECT 1330.390 1011.540 1330.710 1011.600 ;
        RECT 1330.850 1011.740 1331.170 1011.800 ;
        RECT 1347.870 1011.740 1348.190 1011.800 ;
        RECT 1330.850 1011.600 1348.190 1011.740 ;
        RECT 1330.850 1011.540 1331.170 1011.600 ;
        RECT 1347.870 1011.540 1348.190 1011.600 ;
        RECT 1487.710 1011.740 1488.030 1011.800 ;
        RECT 1511.170 1011.740 1511.490 1011.800 ;
        RECT 1487.710 1011.600 1511.490 1011.740 ;
        RECT 1487.710 1011.540 1488.030 1011.600 ;
        RECT 1511.170 1011.540 1511.490 1011.600 ;
        RECT 1527.730 1011.740 1528.050 1011.800 ;
        RECT 1878.250 1011.740 1878.570 1011.800 ;
        RECT 1886.530 1011.740 1886.850 1011.800 ;
        RECT 1527.730 1011.600 1878.020 1011.740 ;
        RECT 1527.730 1011.540 1528.050 1011.600 ;
        RECT 700.190 1011.400 700.510 1011.460 ;
        RECT 893.390 1011.400 893.710 1011.460 ;
        RECT 700.190 1011.260 893.710 1011.400 ;
        RECT 700.190 1011.200 700.510 1011.260 ;
        RECT 893.390 1011.200 893.710 1011.260 ;
        RECT 1007.010 1011.400 1007.330 1011.460 ;
        RECT 1292.670 1011.400 1292.990 1011.460 ;
        RECT 1348.790 1011.400 1349.110 1011.460 ;
        RECT 1007.010 1011.260 1292.990 1011.400 ;
        RECT 1007.010 1011.200 1007.330 1011.260 ;
        RECT 1292.670 1011.200 1292.990 1011.260 ;
        RECT 1294.140 1011.260 1349.110 1011.400 ;
        RECT 517.110 1011.060 517.430 1011.120 ;
        RECT 712.610 1011.060 712.930 1011.120 ;
        RECT 517.110 1010.920 712.930 1011.060 ;
        RECT 517.110 1010.860 517.430 1010.920 ;
        RECT 712.610 1010.860 712.930 1010.920 ;
        RECT 720.890 1011.060 721.210 1011.120 ;
        RECT 906.270 1011.060 906.590 1011.120 ;
        RECT 720.890 1010.920 906.590 1011.060 ;
        RECT 720.890 1010.860 721.210 1010.920 ;
        RECT 906.270 1010.860 906.590 1010.920 ;
        RECT 995.510 1011.060 995.830 1011.120 ;
        RECT 1282.550 1011.060 1282.870 1011.120 ;
        RECT 995.510 1010.920 1282.870 1011.060 ;
        RECT 995.510 1010.860 995.830 1010.920 ;
        RECT 1282.550 1010.860 1282.870 1010.920 ;
        RECT 468.810 1010.720 469.130 1010.780 ;
        RECT 673.510 1010.720 673.830 1010.780 ;
        RECT 468.810 1010.580 673.830 1010.720 ;
        RECT 468.810 1010.520 469.130 1010.580 ;
        RECT 673.510 1010.520 673.830 1010.580 ;
        RECT 707.090 1010.720 707.410 1010.780 ;
        RECT 901.670 1010.720 901.990 1010.780 ;
        RECT 707.090 1010.580 901.990 1010.720 ;
        RECT 707.090 1010.520 707.410 1010.580 ;
        RECT 901.670 1010.520 901.990 1010.580 ;
        RECT 996.430 1010.720 996.750 1010.780 ;
        RECT 1294.140 1010.720 1294.280 1011.260 ;
        RECT 1348.790 1011.200 1349.110 1011.260 ;
        RECT 1461.490 1011.400 1461.810 1011.460 ;
        RECT 1877.880 1011.400 1878.020 1011.600 ;
        RECT 1878.250 1011.600 1886.850 1011.740 ;
        RECT 1878.250 1011.540 1878.570 1011.600 ;
        RECT 1886.530 1011.540 1886.850 1011.600 ;
        RECT 2050.750 1011.740 2051.070 1011.800 ;
        RECT 2055.810 1011.740 2056.130 1011.800 ;
        RECT 2050.750 1011.600 2056.130 1011.740 ;
        RECT 2050.750 1011.540 2051.070 1011.600 ;
        RECT 2055.810 1011.540 2056.130 1011.600 ;
        RECT 2085.710 1011.740 2086.030 1011.800 ;
        RECT 2519.490 1011.740 2519.810 1011.800 ;
        RECT 2085.710 1011.600 2519.810 1011.740 ;
        RECT 2085.710 1011.540 2086.030 1011.600 ;
        RECT 2519.490 1011.540 2519.810 1011.600 ;
        RECT 1892.510 1011.400 1892.830 1011.460 ;
        RECT 1461.490 1011.260 1877.560 1011.400 ;
        RECT 1877.880 1011.260 1892.830 1011.400 ;
        RECT 1461.490 1011.200 1461.810 1011.260 ;
        RECT 1294.970 1011.060 1295.290 1011.120 ;
        RECT 1333.610 1011.060 1333.930 1011.120 ;
        RECT 1294.970 1010.920 1333.930 1011.060 ;
        RECT 1294.970 1010.860 1295.290 1010.920 ;
        RECT 1333.610 1010.860 1333.930 1010.920 ;
        RECT 1354.770 1011.060 1355.090 1011.120 ;
        RECT 1871.810 1011.060 1872.130 1011.120 ;
        RECT 1354.770 1010.920 1872.130 1011.060 ;
        RECT 1354.770 1010.860 1355.090 1010.920 ;
        RECT 1871.810 1010.860 1872.130 1010.920 ;
        RECT 1872.270 1011.060 1872.590 1011.120 ;
        RECT 1876.410 1011.060 1876.730 1011.120 ;
        RECT 1872.270 1010.920 1876.730 1011.060 ;
        RECT 1877.420 1011.060 1877.560 1011.260 ;
        RECT 1892.510 1011.200 1892.830 1011.260 ;
        RECT 2055.350 1011.400 2055.670 1011.460 ;
        RECT 2519.030 1011.400 2519.350 1011.460 ;
        RECT 2055.350 1011.260 2519.350 1011.400 ;
        RECT 2055.350 1011.200 2055.670 1011.260 ;
        RECT 2519.030 1011.200 2519.350 1011.260 ;
        RECT 1898.490 1011.060 1898.810 1011.120 ;
        RECT 1877.420 1010.920 1898.810 1011.060 ;
        RECT 1872.270 1010.860 1872.590 1010.920 ;
        RECT 1876.410 1010.860 1876.730 1010.920 ;
        RECT 1898.490 1010.860 1898.810 1010.920 ;
        RECT 2046.150 1011.060 2046.470 1011.120 ;
        RECT 2518.570 1011.060 2518.890 1011.120 ;
        RECT 2046.150 1010.920 2518.890 1011.060 ;
        RECT 2046.150 1010.860 2046.470 1010.920 ;
        RECT 2518.570 1010.860 2518.890 1010.920 ;
        RECT 996.430 1010.580 1294.280 1010.720 ;
        RECT 1294.510 1010.720 1294.830 1010.780 ;
        RECT 1341.430 1010.720 1341.750 1010.780 ;
        RECT 1294.510 1010.580 1341.750 1010.720 ;
        RECT 996.430 1010.520 996.750 1010.580 ;
        RECT 1294.510 1010.520 1294.830 1010.580 ;
        RECT 1341.430 1010.520 1341.750 1010.580 ;
        RECT 1417.790 1010.720 1418.110 1010.780 ;
        RECT 1728.750 1010.720 1729.070 1010.780 ;
        RECT 1767.390 1010.720 1767.710 1010.780 ;
        RECT 1417.790 1010.580 1631.920 1010.720 ;
        RECT 1417.790 1010.520 1418.110 1010.580 ;
        RECT 984.470 1010.380 984.790 1010.440 ;
        RECT 1084.290 1010.380 1084.610 1010.440 ;
        RECT 984.470 1010.240 1084.610 1010.380 ;
        RECT 984.470 1010.180 984.790 1010.240 ;
        RECT 1084.290 1010.180 1084.610 1010.240 ;
        RECT 1089.810 1010.380 1090.130 1010.440 ;
        RECT 1196.070 1010.380 1196.390 1010.440 ;
        RECT 1200.210 1010.380 1200.530 1010.440 ;
        RECT 1089.810 1010.240 1195.840 1010.380 ;
        RECT 1089.810 1010.180 1090.130 1010.240 ;
        RECT 977.110 1010.040 977.430 1010.100 ;
        RECT 1115.110 1010.040 1115.430 1010.100 ;
        RECT 977.110 1009.900 1115.430 1010.040 ;
        RECT 977.110 1009.840 977.430 1009.900 ;
        RECT 1115.110 1009.840 1115.430 1009.900 ;
        RECT 979.410 1009.700 979.730 1009.760 ;
        RECT 1090.270 1009.700 1090.590 1009.760 ;
        RECT 979.410 1009.560 1090.590 1009.700 ;
        RECT 979.410 1009.500 979.730 1009.560 ;
        RECT 1090.270 1009.500 1090.590 1009.560 ;
        RECT 1103.150 1009.700 1103.470 1009.760 ;
        RECT 1139.030 1009.700 1139.350 1009.760 ;
        RECT 1103.150 1009.560 1139.350 1009.700 ;
        RECT 1103.150 1009.500 1103.470 1009.560 ;
        RECT 1139.030 1009.500 1139.350 1009.560 ;
        RECT 998.270 1009.360 998.590 1009.420 ;
        RECT 1097.630 1009.360 1097.950 1009.420 ;
        RECT 998.270 1009.220 1097.950 1009.360 ;
        RECT 998.270 1009.160 998.590 1009.220 ;
        RECT 1097.630 1009.160 1097.950 1009.220 ;
        RECT 984.010 1009.020 984.330 1009.080 ;
        RECT 1093.030 1009.020 1093.350 1009.080 ;
        RECT 984.010 1008.880 1093.350 1009.020 ;
        RECT 1195.700 1009.020 1195.840 1010.240 ;
        RECT 1196.070 1010.240 1200.530 1010.380 ;
        RECT 1196.070 1010.180 1196.390 1010.240 ;
        RECT 1200.210 1010.180 1200.530 1010.240 ;
        RECT 1259.090 1010.380 1259.410 1010.440 ;
        RECT 1338.670 1010.380 1338.990 1010.440 ;
        RECT 1259.090 1010.240 1338.990 1010.380 ;
        RECT 1259.090 1010.180 1259.410 1010.240 ;
        RECT 1338.670 1010.180 1338.990 1010.240 ;
        RECT 1487.250 1010.380 1487.570 1010.440 ;
        RECT 1519.450 1010.380 1519.770 1010.440 ;
        RECT 1487.250 1010.240 1519.770 1010.380 ;
        RECT 1487.250 1010.180 1487.570 1010.240 ;
        RECT 1519.450 1010.180 1519.770 1010.240 ;
        RECT 1534.630 1010.380 1534.950 1010.440 ;
        RECT 1576.490 1010.380 1576.810 1010.440 ;
        RECT 1534.630 1010.240 1576.810 1010.380 ;
        RECT 1534.630 1010.180 1534.950 1010.240 ;
        RECT 1576.490 1010.180 1576.810 1010.240 ;
        RECT 1231.490 1010.040 1231.810 1010.100 ;
        RECT 1265.530 1010.040 1265.850 1010.100 ;
        RECT 1268.290 1010.040 1268.610 1010.100 ;
        RECT 1231.490 1009.900 1240.000 1010.040 ;
        RECT 1231.490 1009.840 1231.810 1009.900 ;
        RECT 1215.390 1009.700 1215.710 1009.760 ;
        RECT 1238.390 1009.700 1238.710 1009.760 ;
        RECT 1215.390 1009.560 1238.710 1009.700 ;
        RECT 1239.860 1009.700 1240.000 1009.900 ;
        RECT 1265.530 1009.900 1268.610 1010.040 ;
        RECT 1265.530 1009.840 1265.850 1009.900 ;
        RECT 1268.290 1009.840 1268.610 1009.900 ;
        RECT 1268.750 1010.040 1269.070 1010.100 ;
        RECT 1293.590 1010.040 1293.910 1010.100 ;
        RECT 1268.750 1009.900 1293.910 1010.040 ;
        RECT 1268.750 1009.840 1269.070 1009.900 ;
        RECT 1293.590 1009.840 1293.910 1009.900 ;
        RECT 1294.050 1010.040 1294.370 1010.100 ;
        RECT 1332.230 1010.040 1332.550 1010.100 ;
        RECT 1294.050 1009.900 1332.550 1010.040 ;
        RECT 1294.050 1009.840 1294.370 1009.900 ;
        RECT 1332.230 1009.840 1332.550 1009.900 ;
        RECT 1502.430 1010.040 1502.750 1010.100 ;
        RECT 1585.690 1010.040 1586.010 1010.100 ;
        RECT 1502.430 1009.900 1586.010 1010.040 ;
        RECT 1502.430 1009.840 1502.750 1009.900 ;
        RECT 1585.690 1009.840 1586.010 1009.900 ;
        RECT 1602.710 1010.040 1603.030 1010.100 ;
        RECT 1607.310 1010.040 1607.630 1010.100 ;
        RECT 1602.710 1009.900 1607.630 1010.040 ;
        RECT 1602.710 1009.840 1603.030 1009.900 ;
        RECT 1607.310 1009.840 1607.630 1009.900 ;
        RECT 1620.190 1010.040 1620.510 1010.100 ;
        RECT 1624.790 1010.040 1625.110 1010.100 ;
        RECT 1620.190 1009.900 1625.110 1010.040 ;
        RECT 1631.780 1010.040 1631.920 1010.580 ;
        RECT 1728.750 1010.580 1767.710 1010.720 ;
        RECT 1728.750 1010.520 1729.070 1010.580 ;
        RECT 1767.390 1010.520 1767.710 1010.580 ;
        RECT 1767.850 1010.720 1768.170 1010.780 ;
        RECT 1772.910 1010.720 1773.230 1010.780 ;
        RECT 1767.850 1010.580 1773.230 1010.720 ;
        RECT 1767.850 1010.520 1768.170 1010.580 ;
        RECT 1772.910 1010.520 1773.230 1010.580 ;
        RECT 1824.430 1010.720 1824.750 1010.780 ;
        RECT 1827.650 1010.720 1827.970 1010.780 ;
        RECT 1824.430 1010.580 1827.970 1010.720 ;
        RECT 1824.430 1010.520 1824.750 1010.580 ;
        RECT 1827.650 1010.520 1827.970 1010.580 ;
        RECT 1830.870 1010.720 1831.190 1010.780 ;
        RECT 1835.010 1010.720 1835.330 1010.780 ;
        RECT 1830.870 1010.580 1835.330 1010.720 ;
        RECT 1830.870 1010.520 1831.190 1010.580 ;
        RECT 1835.010 1010.520 1835.330 1010.580 ;
        RECT 1882.390 1010.720 1882.710 1010.780 ;
        RECT 2528.690 1010.720 2529.010 1010.780 ;
        RECT 1882.390 1010.580 2529.010 1010.720 ;
        RECT 1882.390 1010.520 1882.710 1010.580 ;
        RECT 2528.690 1010.520 2529.010 1010.580 ;
        RECT 1789.470 1010.380 1789.790 1010.440 ;
        RECT 2074.670 1010.380 2074.990 1010.440 ;
        RECT 2085.710 1010.380 2086.030 1010.440 ;
        RECT 1789.470 1010.240 2073.980 1010.380 ;
        RECT 1789.470 1010.180 1789.790 1010.240 ;
        RECT 1673.090 1010.040 1673.410 1010.100 ;
        RECT 1631.780 1009.900 1673.410 1010.040 ;
        RECT 1620.190 1009.840 1620.510 1009.900 ;
        RECT 1624.790 1009.840 1625.110 1009.900 ;
        RECT 1673.090 1009.840 1673.410 1009.900 ;
        RECT 1834.550 1010.040 1834.870 1010.100 ;
        RECT 2073.290 1010.040 2073.610 1010.100 ;
        RECT 1834.550 1009.900 2073.610 1010.040 ;
        RECT 2073.840 1010.040 2073.980 1010.240 ;
        RECT 2074.670 1010.240 2086.030 1010.380 ;
        RECT 2074.670 1010.180 2074.990 1010.240 ;
        RECT 2085.710 1010.180 2086.030 1010.240 ;
        RECT 2084.790 1010.040 2085.110 1010.100 ;
        RECT 2073.840 1009.900 2085.110 1010.040 ;
        RECT 1834.550 1009.840 1834.870 1009.900 ;
        RECT 2073.290 1009.840 2073.610 1009.900 ;
        RECT 2084.790 1009.840 2085.110 1009.900 ;
        RECT 1304.170 1009.700 1304.490 1009.760 ;
        RECT 1239.860 1009.560 1304.490 1009.700 ;
        RECT 1215.390 1009.500 1215.710 1009.560 ;
        RECT 1238.390 1009.500 1238.710 1009.560 ;
        RECT 1304.170 1009.500 1304.490 1009.560 ;
        RECT 1326.710 1009.700 1327.030 1009.760 ;
        RECT 1334.070 1009.700 1334.390 1009.760 ;
        RECT 1326.710 1009.560 1334.390 1009.700 ;
        RECT 1326.710 1009.500 1327.030 1009.560 ;
        RECT 1334.070 1009.500 1334.390 1009.560 ;
        RECT 1334.990 1009.700 1335.310 1009.760 ;
        RECT 1340.970 1009.700 1341.290 1009.760 ;
        RECT 1334.990 1009.560 1341.290 1009.700 ;
        RECT 1334.990 1009.500 1335.310 1009.560 ;
        RECT 1340.970 1009.500 1341.290 1009.560 ;
        RECT 1495.990 1009.700 1496.310 1009.760 ;
        RECT 1521.290 1009.700 1521.610 1009.760 ;
        RECT 1577.870 1009.700 1578.190 1009.760 ;
        RECT 1495.990 1009.560 1521.610 1009.700 ;
        RECT 1495.990 1009.500 1496.310 1009.560 ;
        RECT 1521.290 1009.500 1521.610 1009.560 ;
        RECT 1529.660 1009.560 1578.190 1009.700 ;
        RECT 1196.530 1009.360 1196.850 1009.420 ;
        RECT 1238.850 1009.360 1239.170 1009.420 ;
        RECT 1196.530 1009.220 1239.170 1009.360 ;
        RECT 1196.530 1009.160 1196.850 1009.220 ;
        RECT 1238.850 1009.160 1239.170 1009.220 ;
        RECT 1285.310 1009.360 1285.630 1009.420 ;
        RECT 1329.930 1009.360 1330.250 1009.420 ;
        RECT 1285.310 1009.220 1330.250 1009.360 ;
        RECT 1285.310 1009.160 1285.630 1009.220 ;
        RECT 1329.930 1009.160 1330.250 1009.220 ;
        RECT 1330.390 1009.360 1330.710 1009.420 ;
        RECT 1353.390 1009.360 1353.710 1009.420 ;
        RECT 1330.390 1009.220 1353.710 1009.360 ;
        RECT 1330.390 1009.160 1330.710 1009.220 ;
        RECT 1353.390 1009.160 1353.710 1009.220 ;
        RECT 1486.330 1009.360 1486.650 1009.420 ;
        RECT 1527.730 1009.360 1528.050 1009.420 ;
        RECT 1486.330 1009.220 1528.050 1009.360 ;
        RECT 1486.330 1009.160 1486.650 1009.220 ;
        RECT 1527.730 1009.160 1528.050 1009.220 ;
        RECT 1230.110 1009.020 1230.430 1009.080 ;
        RECT 1195.700 1008.880 1230.430 1009.020 ;
        RECT 984.010 1008.820 984.330 1008.880 ;
        RECT 1093.030 1008.820 1093.350 1008.880 ;
        RECT 1230.110 1008.820 1230.430 1008.880 ;
        RECT 1282.550 1009.020 1282.870 1009.080 ;
        RECT 1299.570 1009.020 1299.890 1009.080 ;
        RECT 1332.230 1009.020 1332.550 1009.080 ;
        RECT 1354.310 1009.020 1354.630 1009.080 ;
        RECT 1282.550 1008.880 1299.890 1009.020 ;
        RECT 1282.550 1008.820 1282.870 1008.880 ;
        RECT 1299.570 1008.820 1299.890 1008.880 ;
        RECT 1300.120 1008.880 1332.550 1009.020 ;
        RECT 993.670 1008.680 993.990 1008.740 ;
        RECT 1080.150 1008.680 1080.470 1008.740 ;
        RECT 993.670 1008.540 1080.470 1008.680 ;
        RECT 993.670 1008.480 993.990 1008.540 ;
        RECT 1080.150 1008.480 1080.470 1008.540 ;
        RECT 1250.350 1008.680 1250.670 1008.740 ;
        RECT 1254.950 1008.680 1255.270 1008.740 ;
        RECT 1250.350 1008.540 1255.270 1008.680 ;
        RECT 1250.350 1008.480 1250.670 1008.540 ;
        RECT 1254.950 1008.480 1255.270 1008.540 ;
        RECT 1274.270 1008.680 1274.590 1008.740 ;
        RECT 1300.120 1008.680 1300.260 1008.880 ;
        RECT 1332.230 1008.820 1332.550 1008.880 ;
        RECT 1333.930 1008.880 1354.630 1009.020 ;
        RECT 1274.270 1008.540 1300.260 1008.680 ;
        RECT 1313.370 1008.680 1313.690 1008.740 ;
        RECT 1329.470 1008.680 1329.790 1008.740 ;
        RECT 1313.370 1008.540 1329.790 1008.680 ;
        RECT 1274.270 1008.480 1274.590 1008.540 ;
        RECT 1313.370 1008.480 1313.690 1008.540 ;
        RECT 1329.470 1008.480 1329.790 1008.540 ;
        RECT 1329.930 1008.680 1330.250 1008.740 ;
        RECT 1333.930 1008.680 1334.070 1008.880 ;
        RECT 1354.310 1008.820 1354.630 1008.880 ;
        RECT 1501.970 1009.020 1502.290 1009.080 ;
        RECT 1529.660 1009.020 1529.800 1009.560 ;
        RECT 1577.870 1009.500 1578.190 1009.560 ;
        RECT 1871.810 1009.700 1872.130 1009.760 ;
        RECT 1899.870 1009.700 1900.190 1009.760 ;
        RECT 1871.810 1009.560 1900.190 1009.700 ;
        RECT 1871.810 1009.500 1872.130 1009.560 ;
        RECT 1899.870 1009.500 1900.190 1009.560 ;
        RECT 2061.330 1009.700 2061.650 1009.760 ;
        RECT 2287.190 1009.700 2287.510 1009.760 ;
        RECT 2061.330 1009.560 2287.510 1009.700 ;
        RECT 2061.330 1009.500 2061.650 1009.560 ;
        RECT 2287.190 1009.500 2287.510 1009.560 ;
        RECT 2064.090 1009.360 2064.410 1009.420 ;
        RECT 2085.250 1009.360 2085.570 1009.420 ;
        RECT 2064.090 1009.220 2085.570 1009.360 ;
        RECT 2064.090 1009.160 2064.410 1009.220 ;
        RECT 2085.250 1009.160 2085.570 1009.220 ;
        RECT 1501.970 1008.880 1529.800 1009.020 ;
        RECT 1535.550 1009.020 1535.870 1009.080 ;
        RECT 1568.210 1009.020 1568.530 1009.080 ;
        RECT 1535.550 1008.880 1568.530 1009.020 ;
        RECT 1501.970 1008.820 1502.290 1008.880 ;
        RECT 1535.550 1008.820 1535.870 1008.880 ;
        RECT 1568.210 1008.820 1568.530 1008.880 ;
        RECT 2073.290 1009.020 2073.610 1009.080 ;
        RECT 2093.990 1009.020 2094.310 1009.080 ;
        RECT 2073.290 1008.880 2094.310 1009.020 ;
        RECT 2073.290 1008.820 2073.610 1008.880 ;
        RECT 2093.990 1008.820 2094.310 1008.880 ;
        RECT 1329.930 1008.540 1334.070 1008.680 ;
        RECT 1340.510 1008.680 1340.830 1008.740 ;
        RECT 1352.930 1008.680 1353.250 1008.740 ;
        RECT 1340.510 1008.540 1353.250 1008.680 ;
        RECT 1329.930 1008.480 1330.250 1008.540 ;
        RECT 1340.510 1008.480 1340.830 1008.540 ;
        RECT 1352.930 1008.480 1353.250 1008.540 ;
        RECT 1361.210 1008.680 1361.530 1008.740 ;
        RECT 1365.810 1008.680 1366.130 1008.740 ;
        RECT 1361.210 1008.540 1366.130 1008.680 ;
        RECT 1361.210 1008.480 1361.530 1008.540 ;
        RECT 1365.810 1008.480 1366.130 1008.540 ;
        RECT 1368.110 1008.680 1368.430 1008.740 ;
        RECT 1372.250 1008.680 1372.570 1008.740 ;
        RECT 1368.110 1008.540 1372.570 1008.680 ;
        RECT 1368.110 1008.480 1368.430 1008.540 ;
        RECT 1372.250 1008.480 1372.570 1008.540 ;
        RECT 1376.390 1008.680 1376.710 1008.740 ;
        RECT 1379.150 1008.680 1379.470 1008.740 ;
        RECT 1376.390 1008.540 1379.470 1008.680 ;
        RECT 1376.390 1008.480 1376.710 1008.540 ;
        RECT 1379.150 1008.480 1379.470 1008.540 ;
        RECT 1396.170 1008.680 1396.490 1008.740 ;
        RECT 1400.310 1008.680 1400.630 1008.740 ;
        RECT 1396.170 1008.540 1400.630 1008.680 ;
        RECT 1396.170 1008.480 1396.490 1008.540 ;
        RECT 1400.310 1008.480 1400.630 1008.540 ;
        RECT 1491.850 1008.680 1492.170 1008.740 ;
        RECT 1505.190 1008.680 1505.510 1008.740 ;
        RECT 1556.710 1008.680 1557.030 1008.740 ;
        RECT 1491.850 1008.540 1505.510 1008.680 ;
        RECT 1491.850 1008.480 1492.170 1008.540 ;
        RECT 1505.190 1008.480 1505.510 1008.540 ;
        RECT 1505.740 1008.540 1557.030 1008.680 ;
        RECT 992.750 1008.340 993.070 1008.400 ;
        RECT 1062.670 1008.340 1062.990 1008.400 ;
        RECT 992.750 1008.200 1062.990 1008.340 ;
        RECT 992.750 1008.140 993.070 1008.200 ;
        RECT 1062.670 1008.140 1062.990 1008.200 ;
        RECT 1223.210 1008.340 1223.530 1008.400 ;
        RECT 1269.210 1008.340 1269.530 1008.400 ;
        RECT 1223.210 1008.200 1269.530 1008.340 ;
        RECT 1223.210 1008.140 1223.530 1008.200 ;
        RECT 1269.210 1008.140 1269.530 1008.200 ;
        RECT 1291.750 1008.340 1292.070 1008.400 ;
        RECT 1333.610 1008.340 1333.930 1008.400 ;
        RECT 1353.850 1008.340 1354.170 1008.400 ;
        RECT 1291.750 1008.200 1333.930 1008.340 ;
        RECT 1291.750 1008.140 1292.070 1008.200 ;
        RECT 1333.610 1008.140 1333.930 1008.200 ;
        RECT 1334.160 1008.200 1354.170 1008.340 ;
        RECT 638.090 1008.000 638.410 1008.060 ;
        RECT 670.750 1008.000 671.070 1008.060 ;
        RECT 638.090 1007.860 671.070 1008.000 ;
        RECT 638.090 1007.800 638.410 1007.860 ;
        RECT 670.750 1007.800 671.070 1007.860 ;
        RECT 992.290 1008.000 992.610 1008.060 ;
        RECT 1055.770 1008.000 1056.090 1008.060 ;
        RECT 992.290 1007.860 1056.090 1008.000 ;
        RECT 992.290 1007.800 992.610 1007.860 ;
        RECT 1055.770 1007.800 1056.090 1007.860 ;
        RECT 1293.590 1008.000 1293.910 1008.060 ;
        RECT 1331.770 1008.000 1332.090 1008.060 ;
        RECT 1334.160 1008.000 1334.300 1008.200 ;
        RECT 1353.850 1008.140 1354.170 1008.200 ;
        RECT 1486.790 1008.340 1487.110 1008.400 ;
        RECT 1505.740 1008.340 1505.880 1008.540 ;
        RECT 1556.710 1008.480 1557.030 1008.540 ;
        RECT 1486.790 1008.200 1505.880 1008.340 ;
        RECT 1509.330 1008.340 1509.650 1008.400 ;
        RECT 1563.150 1008.340 1563.470 1008.400 ;
        RECT 1509.330 1008.200 1563.470 1008.340 ;
        RECT 1486.790 1008.140 1487.110 1008.200 ;
        RECT 1509.330 1008.140 1509.650 1008.200 ;
        RECT 1563.150 1008.140 1563.470 1008.200 ;
        RECT 1293.590 1007.860 1332.090 1008.000 ;
        RECT 1293.590 1007.800 1293.910 1007.860 ;
        RECT 1331.770 1007.800 1332.090 1007.860 ;
        RECT 1332.780 1007.860 1334.300 1008.000 ;
        RECT 1335.450 1008.000 1335.770 1008.060 ;
        RECT 1352.470 1008.000 1352.790 1008.060 ;
        RECT 1335.450 1007.860 1352.790 1008.000 ;
        RECT 994.130 1007.660 994.450 1007.720 ;
        RECT 1058.530 1007.660 1058.850 1007.720 ;
        RECT 1332.230 1007.660 1332.550 1007.720 ;
        RECT 994.130 1007.520 1058.850 1007.660 ;
        RECT 994.130 1007.460 994.450 1007.520 ;
        RECT 1058.530 1007.460 1058.850 1007.520 ;
        RECT 1294.600 1007.520 1332.550 1007.660 ;
        RECT 1263.690 1007.320 1264.010 1007.380 ;
        RECT 1294.600 1007.320 1294.740 1007.520 ;
        RECT 1332.230 1007.460 1332.550 1007.520 ;
        RECT 1263.690 1007.180 1294.740 1007.320 ;
        RECT 1329.470 1007.320 1329.790 1007.380 ;
        RECT 1332.780 1007.320 1332.920 1007.860 ;
        RECT 1335.450 1007.800 1335.770 1007.860 ;
        RECT 1352.470 1007.800 1352.790 1007.860 ;
        RECT 1493.690 1008.000 1494.010 1008.060 ;
        RECT 1536.470 1008.000 1536.790 1008.060 ;
        RECT 1493.690 1007.860 1536.790 1008.000 ;
        RECT 1493.690 1007.800 1494.010 1007.860 ;
        RECT 1536.470 1007.800 1536.790 1007.860 ;
        RECT 1333.150 1007.660 1333.470 1007.720 ;
        RECT 1340.050 1007.660 1340.370 1007.720 ;
        RECT 1333.150 1007.520 1340.370 1007.660 ;
        RECT 1333.150 1007.460 1333.470 1007.520 ;
        RECT 1340.050 1007.460 1340.370 1007.520 ;
        RECT 1488.170 1007.660 1488.490 1007.720 ;
        RECT 1534.630 1007.660 1534.950 1007.720 ;
        RECT 1488.170 1007.520 1534.950 1007.660 ;
        RECT 1488.170 1007.460 1488.490 1007.520 ;
        RECT 1534.630 1007.460 1534.950 1007.520 ;
        RECT 1776.590 1007.660 1776.910 1007.720 ;
        RECT 1779.810 1007.660 1780.130 1007.720 ;
        RECT 1776.590 1007.520 1780.130 1007.660 ;
        RECT 1776.590 1007.460 1776.910 1007.520 ;
        RECT 1779.810 1007.460 1780.130 1007.520 ;
        RECT 1798.210 1007.660 1798.530 1007.720 ;
        RECT 1800.510 1007.660 1800.830 1007.720 ;
        RECT 1798.210 1007.520 1800.830 1007.660 ;
        RECT 1798.210 1007.460 1798.530 1007.520 ;
        RECT 1800.510 1007.460 1800.830 1007.520 ;
        RECT 1802.810 1007.660 1803.130 1007.720 ;
        RECT 1806.950 1007.660 1807.270 1007.720 ;
        RECT 1802.810 1007.520 1807.270 1007.660 ;
        RECT 1802.810 1007.460 1803.130 1007.520 ;
        RECT 1806.950 1007.460 1807.270 1007.520 ;
        RECT 1811.550 1007.660 1811.870 1007.720 ;
        RECT 1813.850 1007.660 1814.170 1007.720 ;
        RECT 1811.550 1007.520 1814.170 1007.660 ;
        RECT 1811.550 1007.460 1811.870 1007.520 ;
        RECT 1813.850 1007.460 1814.170 1007.520 ;
        RECT 2004.750 1007.660 2005.070 1007.720 ;
        RECT 2007.510 1007.660 2007.830 1007.720 ;
        RECT 2004.750 1007.520 2007.830 1007.660 ;
        RECT 2004.750 1007.460 2005.070 1007.520 ;
        RECT 2007.510 1007.460 2007.830 1007.520 ;
        RECT 1329.470 1007.180 1332.920 1007.320 ;
        RECT 1263.690 1007.120 1264.010 1007.180 ;
        RECT 1329.470 1007.120 1329.790 1007.180 ;
        RECT 1243.450 1001.200 1243.770 1001.260 ;
        RECT 1246.900 1001.200 1247.220 1001.260 ;
        RECT 1243.450 1001.060 1247.220 1001.200 ;
        RECT 1243.450 1001.000 1243.770 1001.060 ;
        RECT 1246.900 1001.000 1247.220 1001.060 ;
        RECT 1274.960 1001.200 1275.280 1001.260 ;
        RECT 1294.510 1001.200 1294.830 1001.260 ;
        RECT 1274.960 1001.060 1294.830 1001.200 ;
        RECT 1274.960 1001.000 1275.280 1001.060 ;
        RECT 1294.510 1001.000 1294.830 1001.060 ;
        RECT 1542.680 1001.200 1543.000 1001.260 ;
        RECT 1543.830 1001.200 1544.150 1001.260 ;
        RECT 1542.680 1001.060 1544.150 1001.200 ;
        RECT 1542.680 1001.000 1543.000 1001.060 ;
        RECT 1543.830 1001.000 1544.150 1001.060 ;
        RECT 1193.770 999.500 1194.090 999.560 ;
        RECT 1197.450 999.500 1197.770 999.560 ;
        RECT 1193.770 999.360 1197.770 999.500 ;
        RECT 1193.770 999.300 1194.090 999.360 ;
        RECT 1197.450 999.300 1197.770 999.360 ;
      LAYER met1 ;
        RECT 670.990 604.460 2169.070 998.780 ;
      LAYER via ;
        RECT 1352.040 2917.920 1352.300 2918.180 ;
        RECT 1535.120 2917.920 1535.380 2918.180 ;
        RECT 1414.140 2917.580 1414.400 2917.840 ;
        RECT 1567.320 2917.580 1567.580 2917.840 ;
        RECT 1448.640 2915.880 1448.900 2916.140 ;
        RECT 1641.840 2915.880 1642.100 2916.140 ;
        RECT 1379.640 2915.540 1379.900 2915.800 ;
        RECT 1598.600 2915.540 1598.860 2915.800 ;
        RECT 1405.860 2915.200 1406.120 2915.460 ;
        RECT 1630.800 2915.200 1631.060 2915.460 ;
        RECT 1469.340 2914.860 1469.600 2915.120 ;
        RECT 1694.280 2914.860 1694.540 2915.120 ;
        RECT 1502.000 2914.520 1502.260 2914.780 ;
        RECT 1768.800 2914.520 1769.060 2914.780 ;
        RECT 1502.460 2914.180 1502.720 2914.440 ;
        RECT 1779.840 2914.180 1780.100 2914.440 ;
        RECT 1455.540 2913.840 1455.800 2914.100 ;
        RECT 1758.680 2913.840 1758.940 2914.100 ;
        RECT 1372.740 2913.500 1373.000 2913.760 ;
        RECT 1843.320 2913.500 1843.580 2913.760 ;
        RECT 1494.640 2913.160 1494.900 2913.420 ;
        RECT 1705.320 2913.160 1705.580 2913.420 ;
        RECT 1789.960 2913.160 1790.220 2913.420 ;
        RECT 1895.300 2913.160 1895.560 2913.420 ;
        RECT 1501.540 2912.820 1501.800 2913.080 ;
        RECT 1812.040 2912.820 1812.300 2913.080 ;
        RECT 1833.200 2912.820 1833.460 2913.080 ;
        RECT 1887.940 2912.820 1888.200 2913.080 ;
        RECT 1496.480 2912.480 1496.740 2912.740 ;
        RECT 1663.000 2912.480 1663.260 2912.740 ;
        RECT 1854.360 2912.480 1854.620 2912.740 ;
        RECT 1886.560 2912.480 1886.820 2912.740 ;
        RECT 1493.720 2912.140 1493.980 2912.400 ;
        RECT 1609.640 2912.140 1609.900 2912.400 ;
        RECT 1864.480 2912.140 1864.740 2912.400 ;
        RECT 1887.480 2912.140 1887.740 2912.400 ;
        RECT 1494.180 2911.800 1494.440 2912.060 ;
        RECT 1546.160 2911.800 1546.420 2912.060 ;
        RECT 1496.020 2898.200 1496.280 2898.460 ;
        RECT 1524.080 2898.200 1524.340 2898.460 ;
        RECT 1652.880 2897.180 1653.140 2897.440 ;
        RECT 1693.360 2897.180 1693.620 2897.440 ;
        RECT 1497.400 2896.500 1497.660 2896.760 ;
        RECT 1503.380 2896.500 1503.640 2896.760 ;
        RECT 1490.040 2894.120 1490.300 2894.380 ;
        RECT 1652.880 2896.500 1653.140 2896.760 ;
        RECT 1693.360 2896.500 1693.620 2896.760 ;
        RECT 1801.920 2896.500 1802.180 2896.760 ;
        RECT 1876.900 2896.500 1877.160 2896.760 ;
        RECT 1894.840 2896.500 1895.100 2896.760 ;
        RECT 1406.320 2863.520 1406.580 2863.780 ;
        RECT 1406.320 2862.840 1406.580 2863.100 ;
        RECT 1358.940 2849.580 1359.200 2849.840 ;
        RECT 1483.600 2849.580 1483.860 2849.840 ;
        RECT 1405.400 2848.900 1405.660 2849.160 ;
        RECT 1406.320 2848.900 1406.580 2849.160 ;
        RECT 1000.600 2810.480 1000.860 2810.740 ;
        RECT 1048.440 2810.480 1048.700 2810.740 ;
        RECT 978.980 2810.140 979.240 2810.400 ;
        RECT 1073.740 2810.140 1074.000 2810.400 ;
        RECT 978.520 2809.800 978.780 2810.060 ;
        RECT 1027.740 2809.800 1028.000 2810.060 ;
        RECT 986.340 2809.460 986.600 2809.720 ;
        RECT 1043.380 2809.460 1043.640 2809.720 ;
        RECT 979.440 2809.120 979.700 2809.380 ;
        RECT 1058.100 2809.120 1058.360 2809.380 ;
        RECT 985.880 2808.780 986.140 2809.040 ;
        RECT 1000.600 2808.780 1000.860 2809.040 ;
        RECT 1048.440 2808.440 1048.700 2808.700 ;
        RECT 1089.380 2808.440 1089.640 2808.700 ;
        RECT 1405.400 2801.300 1405.660 2801.560 ;
        RECT 1406.320 2801.300 1406.580 2801.560 ;
        RECT 985.420 2800.960 985.680 2801.220 ;
        RECT 1010.260 2800.960 1010.520 2801.220 ;
        RECT 445.840 2769.340 446.100 2769.600 ;
        RECT 783.020 2769.340 783.280 2769.600 ;
        RECT 532.320 2767.980 532.580 2768.240 ;
        RECT 686.420 2767.980 686.680 2768.240 ;
        RECT 518.520 2767.640 518.780 2767.900 ;
        RECT 707.120 2767.640 707.380 2767.900 ;
        RECT 489.080 2767.300 489.340 2767.560 ;
        RECT 755.420 2767.300 755.680 2767.560 ;
        RECT 588.900 2684.000 589.160 2684.260 ;
        RECT 700.220 2684.000 700.480 2684.260 ;
        RECT 588.900 2663.600 589.160 2663.860 ;
        RECT 769.220 2663.600 769.480 2663.860 ;
        RECT 1365.840 2780.900 1366.100 2781.160 ;
        RECT 1489.120 2780.900 1489.380 2781.160 ;
        RECT 1406.320 2766.960 1406.580 2767.220 ;
        RECT 1406.780 2766.620 1407.040 2766.880 ;
        RECT 1357.560 2753.020 1357.820 2753.280 ;
        RECT 1358.940 2753.020 1359.200 2753.280 ;
        RECT 1406.320 2753.020 1406.580 2753.280 ;
        RECT 1406.780 2753.020 1407.040 2753.280 ;
        RECT 1405.400 2752.340 1405.660 2752.600 ;
        RECT 1406.320 2752.340 1406.580 2752.600 ;
        RECT 1357.560 2728.880 1357.820 2729.140 ;
        RECT 1358.940 2728.880 1359.200 2729.140 ;
        RECT 1357.560 2704.740 1357.820 2705.000 ;
        RECT 1358.020 2704.740 1358.280 2705.000 ;
        RECT 1405.400 2704.740 1405.660 2705.000 ;
        RECT 1406.320 2704.740 1406.580 2705.000 ;
        RECT 1434.840 2691.140 1435.100 2691.400 ;
        RECT 1488.200 2691.140 1488.460 2691.400 ;
        RECT 1406.320 2670.400 1406.580 2670.660 ;
        RECT 1406.780 2670.060 1407.040 2670.320 ;
        RECT 1358.940 2656.460 1359.200 2656.720 ;
        RECT 1359.860 2656.460 1360.120 2656.720 ;
        RECT 1406.320 2656.460 1406.580 2656.720 ;
        RECT 1406.780 2656.460 1407.040 2656.720 ;
        RECT 1358.940 2622.460 1359.200 2622.720 ;
        RECT 1406.320 2622.460 1406.580 2622.720 ;
        RECT 1358.940 2621.780 1359.200 2622.040 ;
        RECT 1406.320 2621.780 1406.580 2622.040 ;
        RECT 1400.340 2608.180 1400.600 2608.440 ;
        RECT 1487.740 2608.180 1488.000 2608.440 ;
        RECT 998.760 2605.460 999.020 2605.720 ;
        RECT 1111.920 2605.460 1112.180 2605.720 ;
        RECT 999.220 2605.120 999.480 2605.380 ;
        RECT 1112.840 2605.120 1113.100 2605.380 ;
        RECT 982.200 2604.780 982.460 2605.040 ;
        RECT 1112.380 2604.780 1112.640 2605.040 ;
        RECT 975.300 2604.440 975.560 2604.700 ;
        RECT 1113.300 2604.440 1113.560 2604.700 ;
        RECT 1393.440 2594.580 1393.700 2594.840 ;
        RECT 1487.280 2594.580 1487.540 2594.840 ;
        RECT 533.240 2591.520 533.500 2591.780 ;
        RECT 720.920 2591.520 721.180 2591.780 ;
        RECT 504.720 2591.180 504.980 2591.440 ;
        RECT 762.320 2591.180 762.580 2591.440 ;
        RECT 981.740 2591.180 982.000 2591.440 ;
        RECT 1094.900 2591.180 1095.160 2591.440 ;
        RECT 1028.200 2587.440 1028.460 2587.700 ;
        RECT 1033.260 2587.440 1033.520 2587.700 ;
        RECT 1413.680 2580.640 1413.940 2580.900 ;
        RECT 1487.280 2580.640 1487.540 2580.900 ;
        RECT 1358.940 2573.840 1359.200 2574.100 ;
        RECT 1406.320 2573.840 1406.580 2574.100 ;
        RECT 1358.480 2573.500 1358.740 2573.760 ;
        RECT 1406.780 2573.500 1407.040 2573.760 ;
        RECT 1358.480 2559.900 1358.740 2560.160 ;
        RECT 1358.940 2559.900 1359.200 2560.160 ;
        RECT 1406.320 2559.900 1406.580 2560.160 ;
        RECT 1406.780 2559.900 1407.040 2560.160 ;
        RECT 1405.400 2559.220 1405.660 2559.480 ;
        RECT 1406.320 2559.220 1406.580 2559.480 ;
        RECT 1468.880 2546.300 1469.140 2546.560 ;
        RECT 1483.600 2546.300 1483.860 2546.560 ;
        RECT 1357.560 2535.760 1357.820 2536.020 ;
        RECT 1358.940 2535.760 1359.200 2536.020 ;
        RECT 1485.900 2525.220 1486.160 2525.480 ;
        RECT 1490.040 2525.220 1490.300 2525.480 ;
        RECT 1357.560 2511.620 1357.820 2511.880 ;
        RECT 1358.020 2511.620 1358.280 2511.880 ;
        RECT 1405.400 2511.620 1405.660 2511.880 ;
        RECT 1406.320 2511.620 1406.580 2511.880 ;
        RECT 2094.020 2781.240 2094.280 2781.500 ;
        RECT 2556.320 2781.240 2556.580 2781.500 ;
        RECT 1893.920 2780.900 1894.180 2781.160 ;
        RECT 2422.000 2780.900 2422.260 2781.160 ;
        RECT 2528.720 2587.440 2528.980 2587.700 ;
        RECT 2534.240 2587.440 2534.500 2587.700 ;
        RECT 1494.180 2497.000 1494.440 2497.260 ;
        RECT 1512.120 2497.000 1512.380 2497.260 ;
        RECT 1621.140 2495.300 1621.400 2495.560 ;
        RECT 1895.300 2495.300 1895.560 2495.560 ;
        RECT 1494.640 2494.960 1494.900 2495.220 ;
        RECT 1552.600 2494.960 1552.860 2495.220 ;
        RECT 1607.340 2494.960 1607.600 2495.220 ;
        RECT 1894.840 2494.960 1895.100 2495.220 ;
        RECT 1501.540 2494.620 1501.800 2494.880 ;
        RECT 1559.500 2494.620 1559.760 2494.880 ;
        RECT 1586.640 2494.620 1586.900 2494.880 ;
        RECT 1887.940 2494.620 1888.200 2494.880 ;
        RECT 1545.240 2494.280 1545.500 2494.540 ;
        RECT 1887.480 2494.280 1887.740 2494.540 ;
        RECT 1876.440 2493.940 1876.700 2494.200 ;
        RECT 2394.400 2493.940 2394.660 2494.200 ;
        RECT 1680.020 2489.520 1680.280 2489.780 ;
        RECT 1746.720 2489.520 1746.980 2489.780 ;
        RECT 1593.540 2489.180 1593.800 2489.440 ;
        RECT 1778.920 2489.180 1779.180 2489.440 ;
        RECT 1600.440 2488.840 1600.700 2489.100 ;
        RECT 1789.960 2488.840 1790.220 2489.100 ;
        RECT 1421.040 2488.500 1421.300 2488.760 ;
        RECT 1842.400 2488.500 1842.660 2488.760 ;
        RECT 1455.080 2488.160 1455.340 2488.420 ;
        RECT 1885.640 2488.160 1885.900 2488.420 ;
        RECT 1405.400 2487.820 1405.660 2488.080 ;
        RECT 1406.320 2487.820 1406.580 2488.080 ;
        RECT 1420.580 2487.820 1420.840 2488.080 ;
        RECT 1874.600 2487.820 1874.860 2488.080 ;
        RECT 1448.180 2486.800 1448.440 2487.060 ;
        RECT 1832.280 2486.800 1832.540 2487.060 ;
        RECT 1427.940 2486.460 1428.200 2486.720 ;
        RECT 1725.560 2486.460 1725.820 2486.720 ;
        RECT 1461.980 2486.120 1462.240 2486.380 ;
        RECT 1757.760 2486.120 1758.020 2486.380 ;
        RECT 1379.180 2485.780 1379.440 2486.040 ;
        RECT 1534.200 2485.780 1534.460 2486.040 ;
        RECT 1535.120 2485.780 1535.380 2486.040 ;
        RECT 1811.120 2485.780 1811.380 2486.040 ;
        RECT 1386.540 2485.440 1386.800 2485.700 ;
        RECT 1587.560 2485.440 1587.820 2485.700 ;
        RECT 1673.120 2485.440 1673.380 2485.700 ;
        RECT 1715.440 2485.440 1715.700 2485.700 ;
        RECT 1441.280 2485.100 1441.540 2485.360 ;
        RECT 1608.720 2485.100 1608.980 2485.360 ;
        RECT 1537.880 2484.760 1538.140 2485.020 ;
        RECT 1575.140 2484.760 1575.400 2485.020 ;
        RECT 1576.520 2484.760 1576.780 2485.020 ;
        RECT 1619.760 2484.760 1620.020 2485.020 ;
        RECT 1524.080 2484.420 1524.340 2484.680 ;
        RECT 1546.620 2484.420 1546.880 2484.680 ;
        RECT 1624.820 2484.420 1625.080 2484.680 ;
        RECT 1640.920 2484.420 1641.180 2484.680 ;
        RECT 1659.320 2484.420 1659.580 2484.680 ;
        RECT 1683.240 2484.420 1683.500 2484.680 ;
        RECT 1485.900 2477.280 1486.160 2477.540 ;
        RECT 1490.040 2477.280 1490.300 2477.540 ;
        RECT 1544.320 2463.680 1544.580 2463.940 ;
        RECT 1545.240 2463.680 1545.500 2463.940 ;
        RECT 1357.560 2438.860 1357.820 2439.120 ;
        RECT 1358.940 2438.860 1359.200 2439.120 ;
        RECT 1406.320 2429.340 1406.580 2429.600 ;
        RECT 1406.320 2428.660 1406.580 2428.920 ;
        RECT 1357.560 2415.400 1357.820 2415.660 ;
        RECT 1358.480 2415.400 1358.740 2415.660 ;
        RECT 1358.480 2414.720 1358.740 2414.980 ;
        RECT 1358.940 2414.720 1359.200 2414.980 ;
        RECT 1543.860 2407.920 1544.120 2408.180 ;
        RECT 1544.320 2407.920 1544.580 2408.180 ;
        RECT 1358.940 2380.380 1359.200 2380.640 ;
        RECT 1406.320 2380.380 1406.580 2380.640 ;
        RECT 1406.780 2380.380 1407.040 2380.640 ;
        RECT 1358.480 2380.040 1358.740 2380.300 ;
        RECT 1406.320 2366.780 1406.580 2367.040 ;
        RECT 1406.780 2366.780 1407.040 2367.040 ;
        RECT 1544.320 2366.780 1544.580 2367.040 ;
        RECT 1543.860 2366.440 1544.120 2366.700 ;
        RECT 1357.560 2342.300 1357.820 2342.560 ;
        RECT 1358.940 2342.300 1359.200 2342.560 ;
        RECT 1406.320 2332.440 1406.580 2332.700 ;
        RECT 1406.320 2331.760 1406.580 2332.020 ;
        RECT 1357.560 2318.840 1357.820 2319.100 ;
        RECT 1358.480 2318.840 1358.740 2319.100 ;
        RECT 1358.480 2318.160 1358.740 2318.420 ;
        RECT 1358.940 2318.160 1359.200 2318.420 ;
        RECT 1534.200 2318.160 1534.460 2318.420 ;
        RECT 1535.120 2318.160 1535.380 2318.420 ;
        RECT 1405.400 2294.020 1405.660 2294.280 ;
        RECT 1406.320 2294.020 1406.580 2294.280 ;
        RECT 1358.940 2283.820 1359.200 2284.080 ;
        RECT 1358.480 2283.480 1358.740 2283.740 ;
        RECT 1357.560 2245.740 1357.820 2246.000 ;
        RECT 1358.940 2245.740 1359.200 2246.000 ;
        RECT 1406.320 2235.880 1406.580 2236.140 ;
        RECT 1406.320 2235.200 1406.580 2235.460 ;
        RECT 1357.560 2222.280 1357.820 2222.540 ;
        RECT 1358.480 2222.280 1358.740 2222.540 ;
        RECT 1358.480 2221.600 1358.740 2221.860 ;
        RECT 1358.940 2221.600 1359.200 2221.860 ;
        RECT 1534.200 2221.600 1534.460 2221.860 ;
        RECT 1535.120 2221.600 1535.380 2221.860 ;
        RECT 1543.860 2214.800 1544.120 2215.060 ;
        RECT 1544.320 2214.800 1544.580 2215.060 ;
        RECT 1405.400 2197.460 1405.660 2197.720 ;
        RECT 1406.320 2197.460 1406.580 2197.720 ;
        RECT 1358.940 2187.260 1359.200 2187.520 ;
        RECT 1358.480 2186.920 1358.740 2187.180 ;
        RECT 1534.200 2173.660 1534.460 2173.920 ;
        RECT 1535.120 2173.660 1535.380 2173.920 ;
        RECT 1357.560 2149.180 1357.820 2149.440 ;
        RECT 1358.940 2149.180 1359.200 2149.440 ;
        RECT 1406.320 2139.320 1406.580 2139.580 ;
        RECT 1406.320 2138.640 1406.580 2138.900 ;
        RECT 1357.560 2125.720 1357.820 2125.980 ;
        RECT 1358.480 2125.720 1358.740 2125.980 ;
        RECT 1358.480 2125.040 1358.740 2125.300 ;
        RECT 1358.940 2125.040 1359.200 2125.300 ;
        RECT 1543.860 2118.240 1544.120 2118.500 ;
        RECT 1544.320 2118.240 1544.580 2118.500 ;
        RECT 1406.320 2117.900 1406.580 2118.160 ;
        RECT 1407.700 2117.900 1407.960 2118.160 ;
        RECT 1408.160 2069.620 1408.420 2069.880 ;
        RECT 1409.080 2069.620 1409.340 2069.880 ;
        RECT 1272.920 2055.340 1273.180 2055.600 ;
        RECT 1347.900 2055.340 1348.160 2055.600 ;
        RECT 1273.380 2055.000 1273.640 2055.260 ;
        RECT 1331.800 2055.000 1332.060 2055.260 ;
        RECT 1293.620 2054.660 1293.880 2054.920 ;
        RECT 1335.020 2054.660 1335.280 2054.920 ;
        RECT 1130.780 2054.320 1131.040 2054.580 ;
        RECT 1353.880 2054.320 1354.140 2054.580 ;
        RECT 1116.980 2053.980 1117.240 2054.240 ;
        RECT 1332.720 2053.980 1332.980 2054.240 ;
        RECT 1230.140 2053.640 1230.400 2053.900 ;
        RECT 1353.420 2053.640 1353.680 2053.900 ;
        RECT 1059.940 2053.300 1060.200 2053.560 ;
        RECT 1293.620 2053.300 1293.880 2053.560 ;
        RECT 1294.080 2053.300 1294.340 2053.560 ;
        RECT 1333.640 2053.300 1333.900 2053.560 ;
        RECT 1031.420 2052.960 1031.680 2053.220 ;
        RECT 1352.500 2052.960 1352.760 2053.220 ;
        RECT 1016.700 2052.620 1016.960 2052.880 ;
        RECT 1272.920 2052.620 1273.180 2052.880 ;
        RECT 1286.260 2052.620 1286.520 2052.880 ;
        RECT 1346.060 2052.620 1346.320 2052.880 ;
        RECT 1201.620 2052.280 1201.880 2052.540 ;
        RECT 1332.260 2052.280 1332.520 2052.540 ;
        RECT 1187.820 2051.940 1188.080 2052.200 ;
        RECT 1294.080 2051.940 1294.340 2052.200 ;
        RECT 1301.900 2051.940 1302.160 2052.200 ;
        RECT 1336.400 2051.940 1336.660 2052.200 ;
        RECT 1173.100 2051.600 1173.360 2051.860 ;
        RECT 1286.260 2051.600 1286.520 2051.860 ;
        RECT 1286.720 2051.600 1286.980 2051.860 ;
        RECT 1346.520 2051.600 1346.780 2051.860 ;
        RECT 1159.300 2051.260 1159.560 2051.520 ;
        RECT 1354.340 2051.260 1354.600 2051.520 ;
        RECT 1144.580 2050.920 1144.840 2051.180 ;
        RECT 1352.960 2050.920 1353.220 2051.180 ;
        RECT 1000.140 2050.580 1000.400 2050.840 ;
        RECT 1088.460 2050.580 1088.720 2050.840 ;
        RECT 1258.660 2050.580 1258.920 2050.840 ;
        RECT 1286.720 2050.580 1286.980 2050.840 ;
        RECT 1287.180 2050.580 1287.440 2050.840 ;
        RECT 1346.980 2050.580 1347.240 2050.840 ;
        RECT 977.600 2050.240 977.860 2050.500 ;
        RECT 1102.260 2050.240 1102.520 2050.500 ;
        RECT 978.060 2049.900 978.320 2050.160 ;
        RECT 1073.740 2049.900 1074.000 2050.160 ;
        RECT 1244.860 2049.900 1245.120 2050.160 ;
        RECT 1347.440 2050.240 1347.700 2050.500 ;
        RECT 999.680 2049.560 999.940 2049.820 ;
        RECT 1045.220 2049.560 1045.480 2049.820 ;
        RECT 1216.340 2049.560 1216.600 2049.820 ;
        RECT 1333.180 2049.900 1333.440 2050.160 ;
        RECT 1315.700 2049.560 1315.960 2049.820 ;
        RECT 1336.860 2049.560 1337.120 2049.820 ;
        RECT 984.960 2049.220 985.220 2049.480 ;
        RECT 1002.900 2049.220 1003.160 2049.480 ;
        RECT 1329.500 2049.220 1329.760 2049.480 ;
        RECT 1343.760 2049.220 1344.020 2049.480 ;
        RECT 984.040 2048.200 984.300 2048.460 ;
        RECT 1014.400 2048.200 1014.660 2048.460 ;
        RECT 984.500 2047.860 984.760 2048.120 ;
        RECT 1028.200 2047.860 1028.460 2048.120 ;
        RECT 977.140 2047.520 977.400 2047.780 ;
        RECT 1048.900 2047.520 1049.160 2047.780 ;
        RECT 975.760 2047.180 976.020 2047.440 ;
        RECT 1062.700 2047.180 1062.960 2047.440 ;
        RECT 983.120 2046.840 983.380 2047.100 ;
        RECT 1076.500 2046.840 1076.760 2047.100 ;
        RECT 983.580 2046.500 983.840 2046.760 ;
        RECT 1097.200 2046.500 1097.460 2046.760 ;
        RECT 976.680 2046.160 976.940 2046.420 ;
        RECT 1097.660 2046.160 1097.920 2046.420 ;
        RECT 982.660 2045.820 982.920 2046.080 ;
        RECT 1111.000 2045.820 1111.260 2046.080 ;
        RECT 976.220 2045.480 976.480 2045.740 ;
        RECT 1111.460 2045.480 1111.720 2045.740 ;
        RECT 1358.020 2042.420 1358.280 2042.680 ;
        RECT 1359.860 2042.420 1360.120 2042.680 ;
        RECT 530.020 1988.360 530.280 1988.620 ;
        RECT 650.540 1988.360 650.800 1988.620 ;
        RECT 579.240 1987.340 579.500 1987.600 ;
        RECT 638.120 1987.340 638.380 1987.600 ;
        RECT 420.540 1978.500 420.800 1978.760 ;
        RECT 420.080 1978.160 420.340 1978.420 ;
        RECT 843.280 1977.820 843.540 1978.080 ;
        RECT 897.560 1977.480 897.820 1977.740 ;
        RECT 998.300 1713.640 998.560 1713.900 ;
        RECT 1001.060 1713.640 1001.320 1713.900 ;
        RECT 1543.860 2021.680 1544.120 2021.940 ;
        RECT 1544.320 2021.680 1544.580 2021.940 ;
        RECT 1358.020 1993.800 1358.280 1994.060 ;
        RECT 1358.940 1993.800 1359.200 1994.060 ;
        RECT 1542.940 1972.720 1543.200 1972.980 ;
        RECT 1544.320 1972.720 1544.580 1972.980 ;
        RECT 2294.120 1946.880 2294.380 1947.140 ;
        RECT 2379.220 1946.880 2379.480 1947.140 ;
        RECT 2083.440 1946.540 2083.700 1946.800 ;
        RECT 2321.260 1946.540 2321.520 1946.800 ;
        RECT 2090.340 1946.200 2090.600 1946.460 ;
        RECT 2437.180 1946.200 2437.440 1946.460 ;
        RECT 2082.980 1945.860 2083.240 1946.120 ;
        RECT 2495.140 1945.860 2495.400 1946.120 ;
        RECT 1357.560 1945.520 1357.820 1945.780 ;
        RECT 1358.020 1945.520 1358.280 1945.780 ;
        RECT 1485.900 1945.520 1486.160 1945.780 ;
        RECT 1490.040 1945.520 1490.300 1945.780 ;
        RECT 1406.780 1931.580 1407.040 1931.840 ;
        RECT 1407.700 1931.580 1407.960 1931.840 ;
        RECT 1534.200 1931.580 1534.460 1931.840 ;
        RECT 1535.120 1931.580 1535.380 1931.840 ;
        RECT 1724.640 1928.520 1724.900 1928.780 ;
        RECT 2044.340 1928.520 2044.600 1928.780 ;
        RECT 1828.140 1927.840 1828.400 1928.100 ;
        RECT 1964.300 1927.840 1964.560 1928.100 ;
        RECT 1745.340 1927.500 1745.600 1927.760 ;
        RECT 1929.340 1927.500 1929.600 1927.760 ;
        RECT 1779.380 1927.160 1779.640 1927.420 ;
        RECT 1998.340 1927.160 1998.600 1927.420 ;
        RECT 1766.040 1926.820 1766.300 1927.080 ;
        RECT 2010.300 1926.820 2010.560 1927.080 ;
        RECT 1786.740 1926.480 1787.000 1926.740 ;
        RECT 2033.300 1926.480 2033.560 1926.740 ;
        RECT 1738.440 1926.140 1738.700 1926.400 ;
        RECT 1987.300 1926.140 1987.560 1926.400 ;
        RECT 1717.740 1925.800 1718.000 1926.060 ;
        RECT 1975.340 1925.800 1975.600 1926.060 ;
        RECT 1779.840 1925.460 1780.100 1925.720 ;
        RECT 2067.340 1925.460 2067.600 1925.720 ;
        RECT 1835.040 1925.120 1835.300 1925.380 ;
        RECT 1952.340 1925.120 1952.600 1925.380 ;
        RECT 1357.560 1921.040 1357.820 1921.300 ;
        RECT 1358.480 1921.040 1358.740 1921.300 ;
        RECT 1485.900 1897.580 1486.160 1897.840 ;
        RECT 1490.040 1897.580 1490.300 1897.840 ;
        RECT 1358.480 1897.240 1358.740 1897.500 ;
        RECT 1358.940 1897.240 1359.200 1897.500 ;
        RECT 1405.860 1883.980 1406.120 1884.240 ;
        RECT 1407.700 1883.980 1407.960 1884.240 ;
        RECT 1534.200 1883.640 1534.460 1883.900 ;
        RECT 1535.120 1883.640 1535.380 1883.900 ;
        RECT 1542.940 1883.640 1543.200 1883.900 ;
        RECT 1543.400 1883.640 1543.660 1883.900 ;
        RECT 1759.140 1883.640 1759.400 1883.900 ;
        RECT 1904.500 1883.640 1904.760 1883.900 ;
        RECT 1405.400 1883.300 1405.660 1883.560 ;
        RECT 1405.860 1883.300 1406.120 1883.560 ;
        RECT 1821.240 1870.040 1821.500 1870.300 ;
        RECT 1904.500 1870.040 1904.760 1870.300 ;
        RECT 1737.980 1849.300 1738.240 1849.560 ;
        RECT 1904.500 1849.300 1904.760 1849.560 ;
        RECT 1405.400 1835.700 1405.660 1835.960 ;
        RECT 1406.780 1835.700 1407.040 1835.960 ;
        RECT 1405.400 1835.020 1405.660 1835.280 ;
        RECT 1406.780 1835.020 1407.040 1835.280 ;
        RECT 1534.200 1835.020 1534.460 1835.280 ;
        RECT 1535.120 1835.020 1535.380 1835.280 ;
        RECT 1543.400 1828.900 1543.660 1829.160 ;
        RECT 1544.320 1828.900 1544.580 1829.160 ;
        RECT 1543.400 1828.220 1543.660 1828.480 ;
        RECT 1544.320 1828.220 1544.580 1828.480 ;
        RECT 1669.440 1814.620 1669.700 1814.880 ;
        RECT 1904.500 1814.620 1904.760 1814.880 ;
        RECT 1358.480 1801.020 1358.740 1801.280 ;
        RECT 1358.940 1801.020 1359.200 1801.280 ;
        RECT 1405.400 1787.420 1405.660 1787.680 ;
        RECT 1405.860 1787.420 1406.120 1787.680 ;
        RECT 1534.200 1787.080 1534.460 1787.340 ;
        RECT 1535.120 1787.080 1535.380 1787.340 ;
        RECT 1543.400 1787.080 1543.660 1787.340 ;
        RECT 1405.400 1786.740 1405.660 1787.000 ;
        RECT 1405.860 1786.740 1406.120 1787.000 ;
        RECT 1544.320 1786.740 1544.580 1787.000 ;
        RECT 1772.940 1766.340 1773.200 1766.600 ;
        RECT 1904.500 1766.340 1904.760 1766.600 ;
        RECT 2073.320 1870.040 2073.580 1870.300 ;
        RECT 2284.000 1870.040 2284.260 1870.300 ;
        RECT 1405.400 1739.140 1405.660 1739.400 ;
        RECT 1406.780 1739.140 1407.040 1739.400 ;
        RECT 1405.400 1738.460 1405.660 1738.720 ;
        RECT 1406.780 1738.460 1407.040 1738.720 ;
        RECT 1534.200 1738.460 1534.460 1738.720 ;
        RECT 1534.660 1738.460 1534.920 1738.720 ;
        RECT 1827.680 1738.460 1827.940 1738.720 ;
        RECT 1933.940 1738.460 1934.200 1738.720 ;
        RECT 1800.540 1738.120 1800.800 1738.380 ;
        RECT 1956.940 1738.120 1957.200 1738.380 ;
        RECT 1793.640 1737.780 1793.900 1738.040 ;
        RECT 1967.980 1737.780 1968.240 1738.040 ;
        RECT 1814.340 1737.440 1814.600 1737.700 ;
        RECT 1990.980 1737.440 1991.240 1737.700 ;
        RECT 1813.880 1737.100 1814.140 1737.360 ;
        RECT 2013.980 1737.100 2014.240 1737.360 ;
        RECT 1752.700 1736.760 1752.960 1737.020 ;
        RECT 1979.940 1736.760 1980.200 1737.020 ;
        RECT 1710.840 1736.420 1711.100 1736.680 ;
        RECT 1944.980 1736.420 1945.240 1736.680 ;
        RECT 1807.440 1736.080 1807.700 1736.340 ;
        RECT 2036.980 1736.080 2037.240 1736.340 ;
        RECT 1772.480 1735.740 1772.740 1736.000 ;
        RECT 2002.940 1735.740 2003.200 1736.000 ;
        RECT 1806.980 1735.400 1807.240 1735.660 ;
        RECT 2071.940 1735.400 2072.200 1735.660 ;
        RECT 1372.280 1735.060 1372.540 1735.320 ;
        RECT 1553.060 1735.060 1553.320 1735.320 ;
        RECT 1668.980 1735.060 1669.240 1735.320 ;
        RECT 2059.980 1735.060 2060.240 1735.320 ;
        RECT 1543.400 1732.000 1543.660 1732.260 ;
        RECT 1543.860 1732.000 1544.120 1732.260 ;
        RECT 2519.060 1709.900 2519.320 1710.160 ;
        RECT 2520.900 1709.900 2521.160 1710.160 ;
        RECT 2519.520 1703.780 2519.780 1704.040 ;
        RECT 2523.660 1704.120 2523.920 1704.380 ;
        RECT 981.740 1694.940 982.000 1695.200 ;
        RECT 1048.900 1694.940 1049.160 1695.200 ;
        RECT 998.760 1694.600 999.020 1694.860 ;
        RECT 1069.600 1694.600 1069.860 1694.860 ;
        RECT 999.220 1694.260 999.480 1694.520 ;
        RECT 1076.500 1694.260 1076.760 1694.520 ;
        RECT 982.200 1693.920 982.460 1694.180 ;
        RECT 1111.000 1693.920 1111.260 1694.180 ;
        RECT 1289.940 1693.920 1290.200 1694.180 ;
        RECT 1336.400 1693.920 1336.660 1694.180 ;
        RECT 975.300 1693.580 975.560 1693.840 ;
        RECT 1104.100 1693.580 1104.360 1693.840 ;
        RECT 1186.440 1693.580 1186.700 1693.840 ;
        RECT 1336.860 1693.580 1337.120 1693.840 ;
        RECT 1310.640 1692.900 1310.900 1693.160 ;
        RECT 1343.760 1692.900 1344.020 1693.160 ;
        RECT 1405.400 1690.520 1405.660 1690.780 ;
        RECT 1406.320 1690.520 1406.580 1690.780 ;
        RECT 1534.200 1690.520 1534.460 1690.780 ;
        RECT 1535.120 1690.520 1535.380 1690.780 ;
        RECT 1543.860 1690.520 1544.120 1690.780 ;
        RECT 1751.320 1690.520 1751.580 1690.780 ;
        RECT 1752.700 1690.520 1752.960 1690.780 ;
        RECT 1159.300 1689.840 1159.560 1690.100 ;
        RECT 1224.160 1689.840 1224.420 1690.100 ;
        RECT 1254.980 1689.840 1255.240 1690.100 ;
        RECT 1300.980 1689.840 1301.240 1690.100 ;
        RECT 1544.320 1689.840 1544.580 1690.100 ;
        RECT 1130.780 1689.500 1131.040 1689.760 ;
        RECT 1242.560 1689.500 1242.820 1689.760 ;
        RECT 1268.780 1689.500 1269.040 1689.760 ;
        RECT 1315.700 1689.500 1315.960 1689.760 ;
        RECT 1102.260 1689.160 1102.520 1689.420 ;
        RECT 1197.020 1689.160 1197.280 1689.420 ;
        RECT 1059.020 1688.820 1059.280 1689.080 ;
        RECT 1203.920 1688.820 1204.180 1689.080 ;
        RECT 1210.820 1688.820 1211.080 1689.080 ;
        RECT 1230.140 1688.820 1230.400 1689.080 ;
        RECT 1245.320 1688.820 1245.580 1689.080 ;
        RECT 1287.180 1688.820 1287.440 1689.080 ;
        RECT 463.780 1688.480 464.040 1688.740 ;
        RECT 468.840 1688.480 469.100 1688.740 ;
        RECT 514.380 1688.480 514.640 1688.740 ;
        RECT 517.140 1688.480 517.400 1688.740 ;
        RECT 1016.700 1688.480 1016.960 1688.740 ;
        RECT 1038.320 1688.480 1038.580 1688.740 ;
        RECT 1073.740 1688.480 1074.000 1688.740 ;
        RECT 1293.620 1688.480 1293.880 1688.740 ;
        RECT 1030.500 1688.140 1030.760 1688.400 ;
        RECT 1277.980 1688.140 1278.240 1688.400 ;
        RECT 2007.540 1687.800 2007.800 1688.060 ;
        RECT 2302.860 1687.800 2303.120 1688.060 ;
        RECT 2055.840 1687.460 2056.100 1687.720 ;
        RECT 2360.820 1687.460 2361.080 1687.720 ;
        RECT 2042.040 1687.120 2042.300 1687.380 ;
        RECT 2418.780 1687.120 2419.040 1687.380 ;
        RECT 2069.640 1686.780 2069.900 1687.040 ;
        RECT 2476.740 1686.780 2477.000 1687.040 ;
        RECT 1116.060 1686.440 1116.320 1686.700 ;
        RECT 1188.280 1686.440 1188.540 1686.700 ;
        RECT 1197.020 1686.440 1197.280 1686.700 ;
        RECT 1231.520 1686.440 1231.780 1686.700 ;
        RECT 1144.580 1686.100 1144.840 1686.360 ;
        RECT 1180.000 1686.100 1180.260 1686.360 ;
        RECT 1214.040 1686.100 1214.300 1686.360 ;
        RECT 1245.320 1686.100 1245.580 1686.360 ;
        RECT 1258.660 1686.100 1258.920 1686.360 ;
        RECT 1300.520 1686.100 1300.780 1686.360 ;
        RECT 1358.940 1684.400 1359.200 1684.660 ;
        RECT 1002.900 1684.060 1003.160 1684.320 ;
        RECT 1007.040 1684.060 1007.300 1684.320 ;
        RECT 1173.100 1684.060 1173.360 1684.320 ;
        RECT 1187.360 1684.060 1187.620 1684.320 ;
        RECT 1187.820 1684.060 1188.080 1684.320 ;
        RECT 1197.020 1684.060 1197.280 1684.320 ;
        RECT 1200.240 1684.060 1200.500 1684.320 ;
        RECT 1215.420 1684.060 1215.680 1684.320 ;
        RECT 1238.420 1684.060 1238.680 1684.320 ;
        RECT 1243.940 1684.060 1244.200 1684.320 ;
        RECT 1272.460 1684.060 1272.720 1684.320 ;
        RECT 1292.240 1684.060 1292.500 1684.320 ;
        RECT 1329.500 1684.060 1329.760 1684.320 ;
        RECT 1348.360 1684.060 1348.620 1684.320 ;
        RECT 1358.480 1684.060 1358.740 1684.320 ;
        RECT 1290.860 1683.380 1291.120 1683.640 ;
        RECT 1292.240 1683.380 1292.500 1683.640 ;
        RECT 2518.140 1655.840 2518.400 1656.100 ;
        RECT 2519.980 1655.840 2520.240 1656.100 ;
        RECT 1357.100 1652.440 1357.360 1652.700 ;
        RECT 1358.020 1652.440 1358.280 1652.700 ;
        RECT 1224.160 1642.240 1224.420 1642.500 ;
        RECT 1243.480 1642.240 1243.740 1642.500 ;
        RECT 1405.860 1642.240 1406.120 1642.500 ;
        RECT 1406.320 1642.240 1406.580 1642.500 ;
        RECT 1535.120 1641.900 1535.380 1642.160 ;
        RECT 2517.680 1641.900 2517.940 1642.160 ;
        RECT 2518.600 1641.900 2518.860 1642.160 ;
        RECT 1535.120 1641.220 1535.380 1641.480 ;
        RECT 1543.860 1635.780 1544.120 1636.040 ;
        RECT 1290.860 1635.440 1291.120 1635.700 ;
        RECT 1291.780 1635.440 1292.040 1635.700 ;
        RECT 1544.320 1635.440 1544.580 1635.700 ;
        RECT 1357.100 1628.300 1357.360 1628.560 ;
        RECT 1357.560 1628.300 1357.820 1628.560 ;
        RECT 2519.980 1617.760 2520.240 1618.020 ;
        RECT 2520.900 1617.760 2521.160 1618.020 ;
        RECT 1357.560 1614.360 1357.820 1614.620 ;
        RECT 1358.480 1614.360 1358.740 1614.620 ;
        RECT 1406.320 1607.560 1406.580 1607.820 ;
        RECT 1406.780 1607.560 1407.040 1607.820 ;
        RECT 1278.900 1593.960 1279.160 1594.220 ;
        RECT 1279.360 1593.960 1279.620 1594.220 ;
        RECT 2517.680 1593.960 2517.940 1594.220 ;
        RECT 2518.600 1593.960 2518.860 1594.220 ;
        RECT 2519.980 1593.960 2520.240 1594.220 ;
        RECT 2520.900 1593.960 2521.160 1594.220 ;
        RECT 1288.560 1593.620 1288.820 1593.880 ;
        RECT 1289.940 1593.620 1290.200 1593.880 ;
        RECT 1405.400 1593.620 1405.660 1593.880 ;
        RECT 1406.780 1593.620 1407.040 1593.880 ;
        RECT 1290.860 1587.160 1291.120 1587.420 ;
        RECT 1293.160 1587.160 1293.420 1587.420 ;
        RECT 2517.220 1569.480 2517.480 1569.740 ;
        RECT 2518.600 1569.480 2518.860 1569.740 ;
        RECT 2518.140 1559.280 2518.400 1559.540 ;
        RECT 2519.980 1559.280 2520.240 1559.540 ;
        RECT 2518.140 1558.600 2518.400 1558.860 ;
        RECT 2519.980 1558.600 2520.240 1558.860 ;
        RECT 1288.560 1545.680 1288.820 1545.940 ;
        RECT 1289.020 1545.680 1289.280 1545.940 ;
        RECT 1405.400 1545.680 1405.660 1545.940 ;
        RECT 1406.320 1545.680 1406.580 1545.940 ;
        RECT 1535.120 1545.680 1535.380 1545.940 ;
        RECT 2517.220 1545.680 2517.480 1545.940 ;
        RECT 2519.060 1545.680 2519.320 1545.940 ;
        RECT 1535.580 1545.340 1535.840 1545.600 ;
        RECT 1535.580 1538.880 1535.840 1539.140 ;
        RECT 1536.040 1538.880 1536.300 1539.140 ;
        RECT 1358.940 1517.800 1359.200 1518.060 ;
        RECT 1359.860 1517.800 1360.120 1518.060 ;
        RECT 1406.320 1511.000 1406.580 1511.260 ;
        RECT 1406.780 1510.660 1407.040 1510.920 ;
        RECT 1535.120 1497.400 1535.380 1497.660 ;
        RECT 1536.040 1497.400 1536.300 1497.660 ;
        RECT 1543.400 1497.400 1543.660 1497.660 ;
        RECT 1543.860 1497.400 1544.120 1497.660 ;
        RECT 1277.520 1497.060 1277.780 1497.320 ;
        RECT 1277.980 1497.060 1278.240 1497.320 ;
        RECT 1288.560 1497.060 1288.820 1497.320 ;
        RECT 1289.480 1497.060 1289.740 1497.320 ;
        RECT 1291.320 1497.060 1291.580 1497.320 ;
        RECT 1291.780 1497.060 1292.040 1497.320 ;
        RECT 1405.400 1497.060 1405.660 1497.320 ;
        RECT 1406.780 1497.060 1407.040 1497.320 ;
        RECT 1543.400 1462.720 1543.660 1462.980 ;
        RECT 1544.320 1462.720 1544.580 1462.980 ;
        RECT 1614.240 1459.660 1614.500 1459.920 ;
        RECT 1893.460 1459.660 1893.720 1459.920 ;
        RECT 1503.840 1459.320 1504.100 1459.580 ;
        RECT 1893.000 1459.320 1893.260 1459.580 ;
        RECT 994.620 1458.980 994.880 1459.240 ;
        RECT 1159.300 1458.980 1159.560 1459.240 ;
        RECT 1503.380 1458.980 1503.640 1459.240 ;
        RECT 1894.380 1458.980 1894.640 1459.240 ;
        RECT 1277.520 1449.460 1277.780 1449.720 ;
        RECT 1291.320 1449.460 1291.580 1449.720 ;
        RECT 1277.980 1449.120 1278.240 1449.380 ;
        RECT 1288.560 1449.120 1288.820 1449.380 ;
        RECT 1289.020 1449.120 1289.280 1449.380 ;
        RECT 1291.780 1449.120 1292.040 1449.380 ;
        RECT 1405.400 1449.120 1405.660 1449.380 ;
        RECT 1406.320 1449.120 1406.580 1449.380 ;
        RECT 1358.940 1421.240 1359.200 1421.500 ;
        RECT 1359.860 1421.240 1360.120 1421.500 ;
        RECT 1542.940 1417.840 1543.200 1418.100 ;
        RECT 1544.320 1417.840 1544.580 1418.100 ;
        RECT 2518.600 1415.120 2518.860 1415.380 ;
        RECT 2519.060 1414.780 2519.320 1415.040 ;
        RECT 1289.020 1414.440 1289.280 1414.700 ;
        RECT 1289.940 1414.440 1290.200 1414.700 ;
        RECT 1406.320 1414.440 1406.580 1414.700 ;
        RECT 1406.780 1414.100 1407.040 1414.360 ;
        RECT 1406.780 1400.500 1407.040 1400.760 ;
        RECT 1408.160 1400.500 1408.420 1400.760 ;
        RECT 1542.940 1393.700 1543.200 1393.960 ;
        RECT 1543.400 1393.700 1543.660 1393.960 ;
        RECT 1291.320 1379.760 1291.580 1380.020 ;
        RECT 1291.780 1379.760 1292.040 1380.020 ;
        RECT 2518.140 1366.500 2518.400 1366.760 ;
        RECT 2519.980 1366.500 2520.240 1366.760 ;
        RECT 2518.140 1365.820 2518.400 1366.080 ;
        RECT 2519.980 1365.820 2520.240 1366.080 ;
        RECT 1406.780 1352.900 1407.040 1353.160 ;
        RECT 1408.160 1352.900 1408.420 1353.160 ;
        RECT 1535.120 1352.560 1535.380 1352.820 ;
        RECT 1405.400 1352.220 1405.660 1352.480 ;
        RECT 1406.780 1352.220 1407.040 1352.480 ;
        RECT 1534.660 1352.220 1534.920 1352.480 ;
        RECT 1543.400 1345.420 1543.660 1345.680 ;
        RECT 1544.320 1345.420 1544.580 1345.680 ;
        RECT 1533.740 1345.080 1534.000 1345.340 ;
        RECT 1534.660 1345.080 1534.920 1345.340 ;
        RECT 1358.020 1324.340 1358.280 1324.600 ;
        RECT 1358.940 1324.340 1359.200 1324.600 ;
        RECT 2518.600 1318.220 2518.860 1318.480 ;
        RECT 2519.980 1318.220 2520.240 1318.480 ;
        RECT 2518.600 1317.540 2518.860 1317.800 ;
        RECT 2519.980 1317.540 2520.240 1317.800 ;
        RECT 1278.440 1304.280 1278.700 1304.540 ;
        RECT 1405.400 1304.280 1405.660 1304.540 ;
        RECT 1406.320 1304.280 1406.580 1304.540 ;
        RECT 1278.440 1303.600 1278.700 1303.860 ;
        RECT 1533.740 1297.140 1534.000 1297.400 ;
        RECT 1535.120 1297.140 1535.380 1297.400 ;
        RECT 1357.100 1276.060 1357.360 1276.320 ;
        RECT 1358.940 1276.060 1359.200 1276.320 ;
        RECT 2518.140 1269.940 2518.400 1270.200 ;
        RECT 2519.980 1269.940 2520.240 1270.200 ;
        RECT 2518.140 1269.260 2518.400 1269.520 ;
        RECT 2519.980 1269.260 2520.240 1269.520 ;
        RECT 1535.120 1257.360 1535.380 1257.620 ;
        RECT 1535.120 1256.680 1535.380 1256.940 ;
        RECT 1292.240 1245.460 1292.500 1245.720 ;
        RECT 1292.240 1244.780 1292.500 1245.040 ;
        RECT 1357.100 1228.120 1357.360 1228.380 ;
        RECT 1357.560 1228.120 1357.820 1228.380 ;
        RECT 1542.940 1226.760 1543.200 1227.020 ;
        RECT 1544.320 1226.760 1544.580 1227.020 ;
        RECT 2518.600 1222.000 2518.860 1222.260 ;
        RECT 2519.060 1221.660 2519.320 1221.920 ;
        RECT 1357.560 1210.780 1357.820 1211.040 ;
        RECT 1358.940 1210.780 1359.200 1211.040 ;
        RECT 1535.120 1207.720 1535.380 1207.980 ;
        RECT 1536.040 1207.720 1536.300 1207.980 ;
        RECT 1405.400 1207.380 1405.660 1207.640 ;
        RECT 1406.320 1207.380 1406.580 1207.640 ;
        RECT 1405.400 1206.700 1405.660 1206.960 ;
        RECT 1406.320 1206.700 1406.580 1206.960 ;
        RECT 1291.320 1200.580 1291.580 1200.840 ;
        RECT 1292.240 1200.580 1292.500 1200.840 ;
        RECT 1291.320 1193.440 1291.580 1193.700 ;
        RECT 1292.240 1193.440 1292.500 1193.700 ;
        RECT 1277.060 1183.240 1277.320 1183.500 ;
        RECT 1277.980 1183.240 1278.240 1183.500 ;
        RECT 1542.940 1176.440 1543.200 1176.700 ;
        RECT 1543.860 1176.440 1544.120 1176.700 ;
        RECT 2518.140 1173.380 2518.400 1173.640 ;
        RECT 2519.980 1173.380 2520.240 1173.640 ;
        RECT 2518.140 1172.700 2518.400 1172.960 ;
        RECT 2519.980 1172.700 2520.240 1172.960 ;
        RECT 1289.940 1159.100 1290.200 1159.360 ;
        RECT 1290.860 1159.100 1291.120 1159.360 ;
        RECT 1405.400 1159.100 1405.660 1159.360 ;
        RECT 1406.320 1159.100 1406.580 1159.360 ;
        RECT 1534.660 1159.100 1534.920 1159.360 ;
        RECT 1535.120 1158.760 1535.380 1159.020 ;
        RECT 1534.660 1152.300 1534.920 1152.560 ;
        RECT 1535.120 1152.300 1535.380 1152.560 ;
        RECT 1358.480 1138.360 1358.740 1138.620 ;
        RECT 1359.400 1138.360 1359.660 1138.620 ;
        RECT 2518.600 1125.440 2518.860 1125.700 ;
        RECT 2519.060 1125.100 2519.320 1125.360 ;
        RECT 1277.980 1110.820 1278.240 1111.080 ;
        RECT 1278.440 1110.820 1278.700 1111.080 ;
        RECT 1405.400 1110.820 1405.660 1111.080 ;
        RECT 1405.860 1110.820 1406.120 1111.080 ;
        RECT 1543.400 1110.820 1543.660 1111.080 ;
        RECT 1069.600 1110.480 1069.860 1110.740 ;
        RECT 1070.980 1110.480 1071.240 1110.740 ;
        RECT 1535.120 1110.480 1535.380 1110.740 ;
        RECT 1535.580 1110.480 1535.840 1110.740 ;
        RECT 1543.860 1110.480 1544.120 1110.740 ;
        RECT 1543.400 1104.020 1543.660 1104.280 ;
        RECT 1543.860 1104.020 1544.120 1104.280 ;
        RECT 1358.480 1090.080 1358.740 1090.340 ;
        RECT 1359.860 1090.080 1360.120 1090.340 ;
        RECT 1541.560 1079.880 1541.820 1080.140 ;
        RECT 1543.400 1079.880 1543.660 1080.140 ;
        RECT 1292.700 1076.820 1292.960 1077.080 ;
        RECT 2518.140 1076.820 2518.400 1077.080 ;
        RECT 2519.980 1076.820 2520.240 1077.080 ;
        RECT 1405.860 1076.480 1406.120 1076.740 ;
        RECT 1292.240 1076.140 1292.500 1076.400 ;
        RECT 1486.360 1076.140 1486.620 1076.400 ;
        RECT 1490.040 1076.140 1490.300 1076.400 ;
        RECT 2518.140 1076.140 2518.400 1076.400 ;
        RECT 2519.980 1076.140 2520.240 1076.400 ;
        RECT 1406.320 1075.800 1406.580 1076.060 ;
        RECT 1070.980 1062.540 1071.240 1062.800 ;
        RECT 1071.900 1062.540 1072.160 1062.800 ;
        RECT 1277.980 1062.540 1278.240 1062.800 ;
        RECT 1278.440 1062.540 1278.700 1062.800 ;
        RECT 1289.020 1062.540 1289.280 1062.800 ;
        RECT 1289.940 1062.540 1290.200 1062.800 ;
        RECT 1357.560 1062.540 1357.820 1062.800 ;
        RECT 1359.860 1062.540 1360.120 1062.800 ;
        RECT 1378.260 1062.540 1378.520 1062.800 ;
        RECT 1379.640 1062.540 1379.900 1062.800 ;
        RECT 1535.120 1062.540 1535.380 1062.800 ;
        RECT 1536.040 1062.540 1536.300 1062.800 ;
        RECT 1277.980 1057.440 1278.240 1057.700 ;
        RECT 1280.740 1057.440 1281.000 1057.700 ;
        RECT 1489.120 1055.400 1489.380 1055.660 ;
        RECT 1519.480 1055.400 1519.740 1055.660 ;
        RECT 1342.380 1052.000 1342.640 1052.260 ;
        RECT 1344.220 1052.000 1344.480 1052.260 ;
        RECT 1454.620 1052.000 1454.880 1052.260 ;
        RECT 1455.540 1052.000 1455.800 1052.260 ;
        RECT 1488.660 1052.000 1488.920 1052.260 ;
        RECT 1559.960 1052.000 1560.220 1052.260 ;
        RECT 2518.600 1028.880 2518.860 1029.140 ;
        RECT 2519.060 1028.540 2519.320 1028.800 ;
        RECT 1486.360 1028.200 1486.620 1028.460 ;
        RECT 1489.120 1028.200 1489.380 1028.460 ;
        RECT 2518.600 1028.200 2518.860 1028.460 ;
        RECT 2519.980 1028.200 2520.240 1028.460 ;
        RECT 1542.020 1027.860 1542.280 1028.120 ;
        RECT 1542.940 1027.860 1543.200 1028.120 ;
        RECT 983.120 1025.480 983.380 1025.740 ;
        RECT 1152.860 1025.480 1153.120 1025.740 ;
        RECT 975.760 1025.140 976.020 1025.400 ;
        RECT 1147.800 1025.140 1148.060 1025.400 ;
        RECT 976.220 1024.800 976.480 1025.060 ;
        RECT 1156.080 1024.800 1156.340 1025.060 ;
        RECT 1474.400 1024.800 1474.660 1025.060 ;
        RECT 1891.620 1024.800 1891.880 1025.060 ;
        RECT 982.660 1024.460 982.920 1024.720 ;
        RECT 1166.200 1024.460 1166.460 1024.720 ;
        RECT 1187.360 1024.460 1187.620 1024.720 ;
        RECT 1188.740 1024.460 1189.000 1024.720 ;
        RECT 1431.160 1024.460 1431.420 1024.720 ;
        RECT 1891.160 1024.460 1891.420 1024.720 ;
        RECT 997.380 1021.060 997.640 1021.320 ;
        RECT 1223.700 1021.060 1223.960 1021.320 ;
        RECT 1278.900 1021.060 1279.160 1021.320 ;
        RECT 1334.560 1021.060 1334.820 1021.320 ;
        RECT 1595.840 1021.060 1596.100 1021.320 ;
        RECT 1900.360 1021.060 1900.620 1021.320 ;
        RECT 988.180 1020.720 988.440 1020.980 ;
        RECT 1228.300 1020.720 1228.560 1020.980 ;
        RECT 1252.680 1020.720 1252.940 1020.980 ;
        RECT 1339.160 1020.720 1339.420 1020.980 ;
        RECT 1567.780 1020.720 1568.040 1020.980 ;
        RECT 1890.700 1020.720 1890.960 1020.980 ;
        RECT 987.260 1020.380 987.520 1020.640 ;
        RECT 1259.580 1020.380 1259.840 1020.640 ;
        RECT 1267.860 1020.380 1268.120 1020.640 ;
        RECT 1343.300 1020.380 1343.560 1020.640 ;
        RECT 1574.680 1020.380 1574.940 1020.640 ;
        RECT 1900.820 1020.380 1901.080 1020.640 ;
        RECT 996.920 1020.040 997.180 1020.300 ;
        RECT 1270.160 1020.040 1270.420 1020.300 ;
        RECT 1279.820 1020.040 1280.080 1020.300 ;
        RECT 1341.920 1020.040 1342.180 1020.300 ;
        RECT 1542.020 1020.040 1542.280 1020.300 ;
        RECT 1886.100 1020.040 1886.360 1020.300 ;
        RECT 996.000 1019.700 996.260 1019.960 ;
        RECT 1292.240 1019.700 1292.500 1019.960 ;
        RECT 1533.280 1019.700 1533.540 1019.960 ;
        RECT 1903.580 1019.700 1903.840 1019.960 ;
        RECT 988.640 1019.360 988.900 1019.620 ;
        RECT 1285.800 1019.360 1286.060 1019.620 ;
        RECT 1299.140 1019.360 1299.400 1019.620 ;
        RECT 1335.940 1019.360 1336.200 1019.620 ;
        RECT 1507.060 1019.360 1507.320 1019.620 ;
        RECT 1897.600 1019.360 1897.860 1019.620 ;
        RECT 989.560 1019.020 989.820 1019.280 ;
        RECT 1301.900 1019.020 1302.160 1019.280 ;
        RECT 1496.940 1019.020 1497.200 1019.280 ;
        RECT 1901.280 1019.020 1901.540 1019.280 ;
        RECT 990.940 1018.680 991.200 1018.940 ;
        RECT 1313.860 1018.680 1314.120 1018.940 ;
        RECT 1462.440 1018.680 1462.700 1018.940 ;
        RECT 1898.980 1018.680 1899.240 1018.940 ;
        RECT 987.720 1018.340 987.980 1018.600 ;
        RECT 1314.780 1018.340 1315.040 1018.600 ;
        RECT 1437.600 1018.340 1437.860 1018.600 ;
        RECT 1898.060 1018.340 1898.320 1018.600 ;
        RECT 989.100 1018.000 989.360 1018.260 ;
        RECT 1327.200 1018.000 1327.460 1018.260 ;
        RECT 1358.940 1018.000 1359.200 1018.260 ;
        RECT 1849.300 1018.000 1849.560 1018.260 ;
        RECT 990.020 1017.660 990.280 1017.920 ;
        RECT 1335.940 1017.660 1336.200 1017.920 ;
        RECT 1402.640 1017.660 1402.900 1017.920 ;
        RECT 1899.440 1017.660 1899.700 1017.920 ;
        RECT 990.480 1017.320 990.740 1017.580 ;
        RECT 1193.800 1017.320 1194.060 1017.580 ;
        RECT 1204.840 1017.320 1205.100 1017.580 ;
        RECT 1342.840 1017.320 1343.100 1017.580 ;
        RECT 1480.840 1017.320 1481.100 1017.580 ;
        RECT 1766.500 1017.320 1766.760 1017.580 ;
        RECT 1048.440 1016.980 1048.700 1017.240 ;
        RECT 1215.880 1016.980 1216.140 1017.240 ;
        RECT 1472.100 1016.980 1472.360 1017.240 ;
        RECT 1704.400 1016.980 1704.660 1017.240 ;
        RECT 991.860 1016.640 992.120 1016.900 ;
        RECT 1125.720 1016.640 1125.980 1016.900 ;
        RECT 1514.420 1016.640 1514.680 1016.900 ;
        RECT 1656.100 1016.640 1656.360 1016.900 ;
        RECT 1489.580 1016.300 1489.840 1016.560 ;
        RECT 1625.740 1016.300 1626.000 1016.560 ;
        RECT 1576.060 1015.960 1576.320 1016.220 ;
        RECT 1680.020 1015.960 1680.280 1016.220 ;
        RECT 1544.780 1015.620 1545.040 1015.880 ;
        RECT 1608.720 1015.620 1608.980 1015.880 ;
        RECT 983.580 1013.920 983.840 1014.180 ;
        RECT 976.680 1013.580 976.940 1013.840 ;
        RECT 1103.180 1013.580 1103.440 1013.840 ;
        RECT 1104.100 1013.920 1104.360 1014.180 ;
        RECT 1106.400 1013.920 1106.660 1014.180 ;
        RECT 1198.400 1013.920 1198.660 1014.180 ;
        RECT 1200.700 1013.920 1200.960 1014.180 ;
        RECT 1202.540 1013.920 1202.800 1014.180 ;
        RECT 1210.820 1013.920 1211.080 1014.180 ;
        RECT 1211.280 1013.920 1211.540 1014.180 ;
        RECT 1214.040 1013.920 1214.300 1014.180 ;
        RECT 1257.280 1013.920 1257.540 1014.180 ;
        RECT 1294.080 1014.260 1294.340 1014.520 ;
        RECT 1134.460 1013.580 1134.720 1013.840 ;
        RECT 1181.840 1013.580 1182.100 1013.840 ;
        RECT 1295.000 1013.920 1295.260 1014.180 ;
        RECT 1300.520 1013.920 1300.780 1014.180 ;
        RECT 1318.000 1013.920 1318.260 1014.180 ;
        RECT 1331.340 1013.920 1331.600 1014.180 ;
        RECT 1346.980 1013.920 1347.240 1014.180 ;
        RECT 1446.340 1013.920 1446.600 1014.180 ;
        RECT 1448.640 1013.920 1448.900 1014.180 ;
        RECT 1452.780 1013.920 1453.040 1014.180 ;
        RECT 1455.080 1013.920 1455.340 1014.180 ;
        RECT 1456.920 1013.920 1457.180 1014.180 ;
        RECT 1461.980 1013.920 1462.240 1014.180 ;
        RECT 1465.660 1013.920 1465.920 1014.180 ;
        RECT 1469.340 1013.920 1469.600 1014.180 ;
        RECT 1479.000 1013.920 1479.260 1014.180 ;
        RECT 1482.220 1013.920 1482.480 1014.180 ;
        RECT 1500.620 1013.920 1500.880 1014.180 ;
        RECT 1503.380 1013.920 1503.640 1014.180 ;
        RECT 1293.620 1013.580 1293.880 1013.840 ;
        RECT 1319.380 1013.580 1319.640 1013.840 ;
        RECT 1324.440 1013.580 1324.700 1013.840 ;
        RECT 1347.440 1013.580 1347.700 1013.840 ;
        RECT 1497.400 1013.580 1497.660 1013.840 ;
        RECT 1535.580 1013.920 1535.840 1014.180 ;
        RECT 1559.500 1013.920 1559.760 1014.180 ;
        RECT 1562.720 1013.920 1562.980 1014.180 ;
        RECT 1563.180 1013.920 1563.440 1014.180 ;
        RECT 1595.840 1013.920 1596.100 1014.180 ;
        RECT 1596.300 1013.920 1596.560 1014.180 ;
        RECT 1600.440 1013.920 1600.700 1014.180 ;
        RECT 1755.000 1013.920 1755.260 1014.180 ;
        RECT 1759.140 1013.920 1759.400 1014.180 ;
        RECT 1763.740 1013.920 1764.000 1014.180 ;
        RECT 1766.040 1013.920 1766.300 1014.180 ;
        RECT 1766.500 1013.920 1766.760 1014.180 ;
        RECT 2065.040 1013.920 2065.300 1014.180 ;
        RECT 2065.500 1013.920 2065.760 1014.180 ;
        RECT 2073.320 1013.920 2073.580 1014.180 ;
        RECT 2075.160 1013.920 2075.420 1014.180 ;
        RECT 2087.120 1013.920 2087.380 1014.180 ;
        RECT 2087.580 1013.920 2087.840 1014.180 ;
        RECT 2090.340 1013.920 2090.600 1014.180 ;
        RECT 1505.220 1013.580 1505.480 1013.840 ;
        RECT 1536.040 1013.580 1536.300 1013.840 ;
        RECT 1552.140 1013.580 1552.400 1013.840 ;
        RECT 1878.280 1013.580 1878.540 1013.840 ;
        RECT 1878.740 1013.580 1879.000 1013.840 ;
        RECT 1893.920 1013.580 1894.180 1013.840 ;
        RECT 2002.940 1013.580 2003.200 1013.840 ;
        RECT 2007.540 1013.580 2007.800 1013.840 ;
        RECT 2008.000 1013.580 2008.260 1013.840 ;
        RECT 2294.120 1013.580 2294.380 1013.840 ;
        RECT 1000.140 1013.240 1000.400 1013.500 ;
        RECT 1191.040 1013.240 1191.300 1013.500 ;
        RECT 1203.920 1013.240 1204.180 1013.500 ;
        RECT 1211.740 1013.240 1212.000 1013.500 ;
        RECT 1254.520 1013.240 1254.780 1013.500 ;
        RECT 1346.060 1013.240 1346.320 1013.500 ;
        RECT 1495.560 1013.240 1495.820 1013.500 ;
        RECT 1525.000 1013.240 1525.260 1013.500 ;
        RECT 1534.660 1013.240 1534.920 1013.500 ;
        RECT 1603.200 1013.240 1603.460 1013.500 ;
        RECT 1720.040 1013.240 1720.300 1013.500 ;
        RECT 783.020 1012.900 783.280 1013.160 ;
        RECT 845.580 1012.900 845.840 1013.160 ;
        RECT 991.400 1012.900 991.660 1013.160 ;
        RECT 1014.400 1012.900 1014.660 1013.160 ;
        RECT 1038.320 1012.900 1038.580 1013.160 ;
        RECT 1196.560 1012.900 1196.820 1013.160 ;
        RECT 1197.020 1012.900 1197.280 1013.160 ;
        RECT 1219.100 1012.900 1219.360 1013.160 ;
        RECT 1244.860 1012.900 1245.120 1013.160 ;
        RECT 1340.540 1012.900 1340.800 1013.160 ;
        RECT 1419.660 1012.900 1419.920 1013.160 ;
        RECT 1421.040 1012.900 1421.300 1013.160 ;
        RECT 1495.100 1012.900 1495.360 1013.160 ;
        RECT 1528.220 1012.900 1528.480 1013.160 ;
        RECT 1536.040 1012.900 1536.300 1013.160 ;
        RECT 1547.540 1012.900 1547.800 1013.160 ;
        RECT 1555.820 1012.900 1556.080 1013.160 ;
        RECT 1659.320 1012.900 1659.580 1013.160 ;
        RECT 1710.380 1012.900 1710.640 1013.160 ;
        RECT 769.220 1012.560 769.480 1012.820 ;
        RECT 890.200 1012.560 890.460 1012.820 ;
        RECT 984.960 1012.560 985.220 1012.820 ;
        RECT 1207.600 1012.560 1207.860 1012.820 ;
        RECT 1237.500 1012.560 1237.760 1012.820 ;
        RECT 650.540 1012.220 650.800 1012.480 ;
        RECT 672.160 1012.220 672.420 1012.480 ;
        RECT 762.320 1012.220 762.580 1012.480 ;
        RECT 884.680 1012.220 884.940 1012.480 ;
        RECT 977.600 1012.220 977.860 1012.480 ;
        RECT 1205.300 1012.220 1205.560 1012.480 ;
        RECT 1218.640 1012.220 1218.900 1012.480 ;
        RECT 1263.260 1012.220 1263.520 1012.480 ;
        RECT 1269.240 1012.560 1269.500 1012.820 ;
        RECT 1339.620 1012.560 1339.880 1012.820 ;
        RECT 1496.480 1012.560 1496.740 1012.820 ;
        RECT 1511.200 1012.560 1511.460 1012.820 ;
        RECT 1511.660 1012.560 1511.920 1012.820 ;
        RECT 1514.880 1012.560 1515.140 1012.820 ;
        RECT 1536.500 1012.560 1536.760 1012.820 ;
        RECT 1628.500 1012.560 1628.760 1012.820 ;
        RECT 755.420 1011.880 755.680 1012.140 ;
        RECT 910.900 1011.880 911.160 1012.140 ;
        RECT 999.680 1011.880 999.940 1012.140 ;
        RECT 1232.440 1011.880 1232.700 1012.140 ;
        RECT 686.420 1011.540 686.680 1011.800 ;
        RECT 841.900 1011.540 842.160 1011.800 ;
        RECT 978.060 1011.540 978.320 1011.800 ;
        RECT 1226.000 1011.540 1226.260 1011.800 ;
        RECT 1237.960 1011.540 1238.220 1011.800 ;
        RECT 1267.400 1011.540 1267.660 1011.800 ;
        RECT 1270.620 1012.220 1270.880 1012.480 ;
        RECT 1331.340 1012.220 1331.600 1012.480 ;
        RECT 1338.240 1012.220 1338.500 1012.480 ;
        RECT 1346.520 1012.220 1346.780 1012.480 ;
        RECT 1369.980 1012.220 1370.240 1012.480 ;
        RECT 1372.740 1012.220 1373.000 1012.480 ;
        RECT 1404.940 1012.220 1405.200 1012.480 ;
        RECT 1406.320 1012.220 1406.580 1012.480 ;
        RECT 1411.380 1012.220 1411.640 1012.480 ;
        RECT 1413.680 1012.220 1413.940 1012.480 ;
        RECT 1444.040 1012.220 1444.300 1012.480 ;
        RECT 1576.520 1012.220 1576.780 1012.480 ;
        RECT 1665.760 1012.220 1666.020 1012.480 ;
        RECT 1669.440 1012.220 1669.700 1012.480 ;
        RECT 1707.160 1012.220 1707.420 1012.480 ;
        RECT 1710.840 1012.220 1711.100 1012.480 ;
        RECT 1715.900 1012.220 1716.160 1012.480 ;
        RECT 1717.740 1012.220 1718.000 1012.480 ;
        RECT 1733.380 1012.220 1733.640 1012.480 ;
        RECT 1737.980 1012.220 1738.240 1012.480 ;
        RECT 1749.940 1013.240 1750.200 1013.500 ;
        RECT 1752.240 1013.240 1752.500 1013.500 ;
        RECT 1758.680 1013.240 1758.940 1013.500 ;
        RECT 1766.500 1013.240 1766.760 1013.500 ;
        RECT 1741.660 1012.900 1741.920 1013.160 ;
        RECT 2064.580 1013.240 2064.840 1013.500 ;
        RECT 2065.040 1013.240 2065.300 1013.500 ;
        RECT 2086.660 1013.240 2086.920 1013.500 ;
        RECT 1767.420 1012.900 1767.680 1013.160 ;
        RECT 2085.740 1012.900 2086.000 1013.160 ;
        RECT 2084.360 1012.560 2084.620 1012.820 ;
        RECT 2064.120 1012.220 2064.380 1012.480 ;
        RECT 2064.580 1012.220 2064.840 1012.480 ;
        RECT 2086.200 1012.220 2086.460 1012.480 ;
        RECT 1269.700 1011.880 1269.960 1012.140 ;
        RECT 1340.080 1011.880 1340.340 1012.140 ;
        RECT 1496.020 1011.880 1496.280 1012.140 ;
        RECT 1534.660 1011.880 1534.920 1012.140 ;
        RECT 1535.120 1011.880 1535.380 1012.140 ;
        RECT 1537.880 1011.880 1538.140 1012.140 ;
        RECT 1552.600 1011.880 1552.860 1012.140 ;
        RECT 1556.280 1011.880 1556.540 1012.140 ;
        RECT 1556.740 1011.880 1557.000 1012.140 ;
        RECT 1628.500 1011.880 1628.760 1012.140 ;
        RECT 1662.540 1011.880 1662.800 1012.140 ;
        RECT 2075.160 1011.880 2075.420 1012.140 ;
        RECT 2078.840 1011.880 2079.100 1012.140 ;
        RECT 2083.440 1011.880 2083.700 1012.140 ;
        RECT 1330.420 1011.540 1330.680 1011.800 ;
        RECT 1330.880 1011.540 1331.140 1011.800 ;
        RECT 1347.900 1011.540 1348.160 1011.800 ;
        RECT 1487.740 1011.540 1488.000 1011.800 ;
        RECT 1511.200 1011.540 1511.460 1011.800 ;
        RECT 1527.760 1011.540 1528.020 1011.800 ;
        RECT 700.220 1011.200 700.480 1011.460 ;
        RECT 893.420 1011.200 893.680 1011.460 ;
        RECT 1007.040 1011.200 1007.300 1011.460 ;
        RECT 1292.700 1011.200 1292.960 1011.460 ;
        RECT 517.140 1010.860 517.400 1011.120 ;
        RECT 712.640 1010.860 712.900 1011.120 ;
        RECT 720.920 1010.860 721.180 1011.120 ;
        RECT 906.300 1010.860 906.560 1011.120 ;
        RECT 995.540 1010.860 995.800 1011.120 ;
        RECT 1282.580 1010.860 1282.840 1011.120 ;
        RECT 468.840 1010.520 469.100 1010.780 ;
        RECT 673.540 1010.520 673.800 1010.780 ;
        RECT 707.120 1010.520 707.380 1010.780 ;
        RECT 901.700 1010.520 901.960 1010.780 ;
        RECT 996.460 1010.520 996.720 1010.780 ;
        RECT 1348.820 1011.200 1349.080 1011.460 ;
        RECT 1461.520 1011.200 1461.780 1011.460 ;
        RECT 1878.280 1011.540 1878.540 1011.800 ;
        RECT 1886.560 1011.540 1886.820 1011.800 ;
        RECT 2050.780 1011.540 2051.040 1011.800 ;
        RECT 2055.840 1011.540 2056.100 1011.800 ;
        RECT 2085.740 1011.540 2086.000 1011.800 ;
        RECT 2519.520 1011.540 2519.780 1011.800 ;
        RECT 1295.000 1010.860 1295.260 1011.120 ;
        RECT 1333.640 1010.860 1333.900 1011.120 ;
        RECT 1354.800 1010.860 1355.060 1011.120 ;
        RECT 1871.840 1010.860 1872.100 1011.120 ;
        RECT 1872.300 1010.860 1872.560 1011.120 ;
        RECT 1876.440 1010.860 1876.700 1011.120 ;
        RECT 1892.540 1011.200 1892.800 1011.460 ;
        RECT 2055.380 1011.200 2055.640 1011.460 ;
        RECT 2519.060 1011.200 2519.320 1011.460 ;
        RECT 1898.520 1010.860 1898.780 1011.120 ;
        RECT 2046.180 1010.860 2046.440 1011.120 ;
        RECT 2518.600 1010.860 2518.860 1011.120 ;
        RECT 1294.540 1010.520 1294.800 1010.780 ;
        RECT 1341.460 1010.520 1341.720 1010.780 ;
        RECT 1417.820 1010.520 1418.080 1010.780 ;
        RECT 984.500 1010.180 984.760 1010.440 ;
        RECT 1084.320 1010.180 1084.580 1010.440 ;
        RECT 1089.840 1010.180 1090.100 1010.440 ;
        RECT 977.140 1009.840 977.400 1010.100 ;
        RECT 1115.140 1009.840 1115.400 1010.100 ;
        RECT 979.440 1009.500 979.700 1009.760 ;
        RECT 1090.300 1009.500 1090.560 1009.760 ;
        RECT 1103.180 1009.500 1103.440 1009.760 ;
        RECT 1139.060 1009.500 1139.320 1009.760 ;
        RECT 998.300 1009.160 998.560 1009.420 ;
        RECT 1097.660 1009.160 1097.920 1009.420 ;
        RECT 984.040 1008.820 984.300 1009.080 ;
        RECT 1093.060 1008.820 1093.320 1009.080 ;
        RECT 1196.100 1010.180 1196.360 1010.440 ;
        RECT 1200.240 1010.180 1200.500 1010.440 ;
        RECT 1259.120 1010.180 1259.380 1010.440 ;
        RECT 1338.700 1010.180 1338.960 1010.440 ;
        RECT 1487.280 1010.180 1487.540 1010.440 ;
        RECT 1519.480 1010.180 1519.740 1010.440 ;
        RECT 1534.660 1010.180 1534.920 1010.440 ;
        RECT 1576.520 1010.180 1576.780 1010.440 ;
        RECT 1231.520 1009.840 1231.780 1010.100 ;
        RECT 1215.420 1009.500 1215.680 1009.760 ;
        RECT 1238.420 1009.500 1238.680 1009.760 ;
        RECT 1265.560 1009.840 1265.820 1010.100 ;
        RECT 1268.320 1009.840 1268.580 1010.100 ;
        RECT 1268.780 1009.840 1269.040 1010.100 ;
        RECT 1293.620 1009.840 1293.880 1010.100 ;
        RECT 1294.080 1009.840 1294.340 1010.100 ;
        RECT 1332.260 1009.840 1332.520 1010.100 ;
        RECT 1502.460 1009.840 1502.720 1010.100 ;
        RECT 1585.720 1009.840 1585.980 1010.100 ;
        RECT 1602.740 1009.840 1603.000 1010.100 ;
        RECT 1607.340 1009.840 1607.600 1010.100 ;
        RECT 1620.220 1009.840 1620.480 1010.100 ;
        RECT 1624.820 1009.840 1625.080 1010.100 ;
        RECT 1728.780 1010.520 1729.040 1010.780 ;
        RECT 1767.420 1010.520 1767.680 1010.780 ;
        RECT 1767.880 1010.520 1768.140 1010.780 ;
        RECT 1772.940 1010.520 1773.200 1010.780 ;
        RECT 1824.460 1010.520 1824.720 1010.780 ;
        RECT 1827.680 1010.520 1827.940 1010.780 ;
        RECT 1830.900 1010.520 1831.160 1010.780 ;
        RECT 1835.040 1010.520 1835.300 1010.780 ;
        RECT 1882.420 1010.520 1882.680 1010.780 ;
        RECT 2528.720 1010.520 2528.980 1010.780 ;
        RECT 1789.500 1010.180 1789.760 1010.440 ;
        RECT 1673.120 1009.840 1673.380 1010.100 ;
        RECT 1834.580 1009.840 1834.840 1010.100 ;
        RECT 2073.320 1009.840 2073.580 1010.100 ;
        RECT 2074.700 1010.180 2074.960 1010.440 ;
        RECT 2085.740 1010.180 2086.000 1010.440 ;
        RECT 2084.820 1009.840 2085.080 1010.100 ;
        RECT 1304.200 1009.500 1304.460 1009.760 ;
        RECT 1326.740 1009.500 1327.000 1009.760 ;
        RECT 1334.100 1009.500 1334.360 1009.760 ;
        RECT 1335.020 1009.500 1335.280 1009.760 ;
        RECT 1341.000 1009.500 1341.260 1009.760 ;
        RECT 1496.020 1009.500 1496.280 1009.760 ;
        RECT 1521.320 1009.500 1521.580 1009.760 ;
        RECT 1196.560 1009.160 1196.820 1009.420 ;
        RECT 1238.880 1009.160 1239.140 1009.420 ;
        RECT 1285.340 1009.160 1285.600 1009.420 ;
        RECT 1329.960 1009.160 1330.220 1009.420 ;
        RECT 1330.420 1009.160 1330.680 1009.420 ;
        RECT 1353.420 1009.160 1353.680 1009.420 ;
        RECT 1486.360 1009.160 1486.620 1009.420 ;
        RECT 1527.760 1009.160 1528.020 1009.420 ;
        RECT 1230.140 1008.820 1230.400 1009.080 ;
        RECT 1282.580 1008.820 1282.840 1009.080 ;
        RECT 1299.600 1008.820 1299.860 1009.080 ;
        RECT 993.700 1008.480 993.960 1008.740 ;
        RECT 1080.180 1008.480 1080.440 1008.740 ;
        RECT 1250.380 1008.480 1250.640 1008.740 ;
        RECT 1254.980 1008.480 1255.240 1008.740 ;
        RECT 1274.300 1008.480 1274.560 1008.740 ;
        RECT 1332.260 1008.820 1332.520 1009.080 ;
        RECT 1313.400 1008.480 1313.660 1008.740 ;
        RECT 1329.500 1008.480 1329.760 1008.740 ;
        RECT 1329.960 1008.480 1330.220 1008.740 ;
        RECT 1354.340 1008.820 1354.600 1009.080 ;
        RECT 1502.000 1008.820 1502.260 1009.080 ;
        RECT 1577.900 1009.500 1578.160 1009.760 ;
        RECT 1871.840 1009.500 1872.100 1009.760 ;
        RECT 1899.900 1009.500 1900.160 1009.760 ;
        RECT 2061.360 1009.500 2061.620 1009.760 ;
        RECT 2287.220 1009.500 2287.480 1009.760 ;
        RECT 2064.120 1009.160 2064.380 1009.420 ;
        RECT 2085.280 1009.160 2085.540 1009.420 ;
        RECT 1535.580 1008.820 1535.840 1009.080 ;
        RECT 1568.240 1008.820 1568.500 1009.080 ;
        RECT 2073.320 1008.820 2073.580 1009.080 ;
        RECT 2094.020 1008.820 2094.280 1009.080 ;
        RECT 1340.540 1008.480 1340.800 1008.740 ;
        RECT 1352.960 1008.480 1353.220 1008.740 ;
        RECT 1361.240 1008.480 1361.500 1008.740 ;
        RECT 1365.840 1008.480 1366.100 1008.740 ;
        RECT 1368.140 1008.480 1368.400 1008.740 ;
        RECT 1372.280 1008.480 1372.540 1008.740 ;
        RECT 1376.420 1008.480 1376.680 1008.740 ;
        RECT 1379.180 1008.480 1379.440 1008.740 ;
        RECT 1396.200 1008.480 1396.460 1008.740 ;
        RECT 1400.340 1008.480 1400.600 1008.740 ;
        RECT 1491.880 1008.480 1492.140 1008.740 ;
        RECT 1505.220 1008.480 1505.480 1008.740 ;
        RECT 992.780 1008.140 993.040 1008.400 ;
        RECT 1062.700 1008.140 1062.960 1008.400 ;
        RECT 1223.240 1008.140 1223.500 1008.400 ;
        RECT 1269.240 1008.140 1269.500 1008.400 ;
        RECT 1291.780 1008.140 1292.040 1008.400 ;
        RECT 1333.640 1008.140 1333.900 1008.400 ;
        RECT 638.120 1007.800 638.380 1008.060 ;
        RECT 670.780 1007.800 671.040 1008.060 ;
        RECT 992.320 1007.800 992.580 1008.060 ;
        RECT 1055.800 1007.800 1056.060 1008.060 ;
        RECT 1293.620 1007.800 1293.880 1008.060 ;
        RECT 1331.800 1007.800 1332.060 1008.060 ;
        RECT 1353.880 1008.140 1354.140 1008.400 ;
        RECT 1486.820 1008.140 1487.080 1008.400 ;
        RECT 1556.740 1008.480 1557.000 1008.740 ;
        RECT 1509.360 1008.140 1509.620 1008.400 ;
        RECT 1563.180 1008.140 1563.440 1008.400 ;
        RECT 994.160 1007.460 994.420 1007.720 ;
        RECT 1058.560 1007.460 1058.820 1007.720 ;
        RECT 1263.720 1007.120 1263.980 1007.380 ;
        RECT 1332.260 1007.460 1332.520 1007.720 ;
        RECT 1329.500 1007.120 1329.760 1007.380 ;
        RECT 1335.480 1007.800 1335.740 1008.060 ;
        RECT 1352.500 1007.800 1352.760 1008.060 ;
        RECT 1493.720 1007.800 1493.980 1008.060 ;
        RECT 1536.500 1007.800 1536.760 1008.060 ;
        RECT 1333.180 1007.460 1333.440 1007.720 ;
        RECT 1340.080 1007.460 1340.340 1007.720 ;
        RECT 1488.200 1007.460 1488.460 1007.720 ;
        RECT 1534.660 1007.460 1534.920 1007.720 ;
        RECT 1776.620 1007.460 1776.880 1007.720 ;
        RECT 1779.840 1007.460 1780.100 1007.720 ;
        RECT 1798.240 1007.460 1798.500 1007.720 ;
        RECT 1800.540 1007.460 1800.800 1007.720 ;
        RECT 1802.840 1007.460 1803.100 1007.720 ;
        RECT 1806.980 1007.460 1807.240 1007.720 ;
        RECT 1811.580 1007.460 1811.840 1007.720 ;
        RECT 1813.880 1007.460 1814.140 1007.720 ;
        RECT 2004.780 1007.460 2005.040 1007.720 ;
        RECT 2007.540 1007.460 2007.800 1007.720 ;
        RECT 1243.480 1001.000 1243.740 1001.260 ;
        RECT 1246.930 1001.000 1247.190 1001.260 ;
        RECT 1274.990 1001.000 1275.250 1001.260 ;
        RECT 1294.540 1001.000 1294.800 1001.260 ;
        RECT 1542.710 1001.000 1542.970 1001.260 ;
        RECT 1543.860 1001.000 1544.120 1001.260 ;
        RECT 1193.800 999.300 1194.060 999.560 ;
        RECT 1197.480 999.300 1197.740 999.560 ;
      LAYER met2 ;
        RECT 1352.040 2917.890 1352.300 2918.210 ;
        RECT 1535.120 2917.890 1535.380 2918.210 ;
        RECT 1000.600 2810.450 1000.860 2810.770 ;
        RECT 1048.440 2810.450 1048.700 2810.770 ;
        RECT 978.980 2810.110 979.240 2810.430 ;
        RECT 978.520 2809.770 978.780 2810.090 ;
        RECT 445.840 2769.310 446.100 2769.630 ;
        RECT 783.020 2769.310 783.280 2769.630 ;
        RECT 445.900 2759.520 446.040 2769.310 ;
        RECT 532.320 2767.950 532.580 2768.270 ;
        RECT 686.420 2767.950 686.680 2768.270 ;
        RECT 518.520 2767.610 518.780 2767.930 ;
        RECT 489.080 2767.270 489.340 2767.590 ;
        RECT 489.140 2759.520 489.280 2767.270 ;
        RECT 518.580 2759.520 518.720 2767.610 ;
        RECT 532.380 2759.520 532.520 2767.950 ;
        RECT 445.730 2759.100 446.040 2759.520 ;
        RECT 488.970 2759.100 489.280 2759.520 ;
        RECT 518.410 2759.100 518.720 2759.520 ;
        RECT 532.210 2759.100 532.520 2759.520 ;
        RECT 445.730 2755.520 446.010 2759.100 ;
        RECT 488.970 2755.520 489.250 2759.100 ;
        RECT 518.410 2755.520 518.690 2759.100 ;
        RECT 532.210 2755.520 532.490 2759.100 ;
      LAYER met2 ;
        RECT 432.860 2755.240 445.450 2755.520 ;
        RECT 446.290 2755.240 460.170 2755.520 ;
        RECT 461.010 2755.240 474.890 2755.520 ;
        RECT 475.730 2755.240 488.690 2755.520 ;
        RECT 489.530 2755.240 503.410 2755.520 ;
        RECT 504.250 2755.240 518.130 2755.520 ;
        RECT 518.970 2755.240 531.930 2755.520 ;
        RECT 532.770 2755.240 546.650 2755.520 ;
        RECT 547.490 2755.240 561.370 2755.520 ;
        RECT 562.210 2755.240 575.170 2755.520 ;
      LAYER met2 ;
        RECT 420.530 2728.995 420.810 2729.365 ;
        RECT 420.070 2707.235 420.350 2707.605 ;
        RECT 420.140 1978.450 420.280 2707.235 ;
        RECT 420.600 1978.790 420.740 2728.995 ;
      LAYER met2 ;
        RECT 432.860 2604.280 575.720 2755.240 ;
      LAYER met2 ;
        RECT 588.890 2686.835 589.170 2687.205 ;
        RECT 588.960 2684.290 589.100 2686.835 ;
        RECT 588.900 2683.970 589.160 2684.290 ;
        RECT 588.890 2666.435 589.170 2666.805 ;
        RECT 588.960 2663.890 589.100 2666.435 ;
        RECT 588.900 2663.570 589.160 2663.890 ;
      LAYER met2 ;
        RECT 433.410 2604.000 446.370 2604.280 ;
        RECT 447.210 2604.000 461.090 2604.280 ;
        RECT 461.930 2604.000 475.810 2604.280 ;
        RECT 476.650 2604.000 489.610 2604.280 ;
        RECT 490.450 2604.000 504.330 2604.280 ;
        RECT 505.170 2604.000 519.050 2604.280 ;
        RECT 519.890 2604.000 532.850 2604.280 ;
        RECT 533.690 2604.000 547.570 2604.280 ;
        RECT 548.410 2604.000 562.290 2604.280 ;
        RECT 563.130 2604.000 575.720 2604.280 ;
      LAYER met2 ;
        RECT 504.610 2600.660 504.890 2604.000 ;
        RECT 533.130 2600.660 533.410 2604.000 ;
        RECT 504.610 2600.000 504.920 2600.660 ;
        RECT 533.130 2600.000 533.440 2600.660 ;
        RECT 504.780 2591.470 504.920 2600.000 ;
        RECT 533.300 2591.810 533.440 2600.000 ;
        RECT 533.240 2591.490 533.500 2591.810 ;
        RECT 504.720 2591.150 504.980 2591.470 ;
        RECT 530.020 1988.330 530.280 1988.650 ;
        RECT 650.540 1988.330 650.800 1988.650 ;
        RECT 528.450 1981.250 528.730 1981.750 ;
        RECT 530.080 1981.250 530.220 1988.330 ;
        RECT 579.240 1987.310 579.500 1987.630 ;
        RECT 638.120 1987.310 638.380 1987.630 ;
        RECT 528.450 1981.110 530.220 1981.250 ;
        RECT 578.130 1981.250 578.410 1981.750 ;
        RECT 579.300 1981.250 579.440 1987.310 ;
        RECT 578.130 1981.110 579.440 1981.250 ;
        RECT 420.540 1978.470 420.800 1978.790 ;
        RECT 420.080 1978.130 420.340 1978.450 ;
        RECT 528.450 1977.750 528.730 1981.110 ;
        RECT 578.130 1977.750 578.410 1981.110 ;
      LAYER met2 ;
        RECT 362.860 1977.470 377.290 1977.750 ;
        RECT 378.130 1977.470 402.130 1977.750 ;
        RECT 402.970 1977.470 427.890 1977.750 ;
        RECT 428.730 1977.470 452.730 1977.750 ;
        RECT 453.570 1977.470 477.570 1977.750 ;
        RECT 478.410 1977.470 502.410 1977.750 ;
        RECT 503.250 1977.470 528.170 1977.750 ;
        RECT 529.010 1977.470 553.010 1977.750 ;
        RECT 553.850 1977.470 577.850 1977.750 ;
        RECT 578.690 1977.470 602.690 1977.750 ;
        RECT 603.530 1977.470 627.530 1977.750 ;
        RECT 362.860 1704.280 628.080 1977.470 ;
        RECT 363.410 1704.000 387.410 1704.280 ;
        RECT 388.250 1704.000 412.250 1704.280 ;
        RECT 413.090 1704.000 437.090 1704.280 ;
        RECT 437.930 1704.000 461.930 1704.280 ;
        RECT 462.770 1704.000 487.690 1704.280 ;
        RECT 488.530 1704.000 512.530 1704.280 ;
        RECT 513.370 1704.000 537.370 1704.280 ;
        RECT 538.210 1704.000 562.210 1704.280 ;
        RECT 563.050 1704.000 587.970 1704.280 ;
        RECT 588.810 1704.000 612.810 1704.280 ;
        RECT 613.650 1704.000 628.080 1704.280 ;
      LAYER met2 ;
        RECT 462.210 1700.410 462.490 1704.000 ;
        RECT 512.810 1700.410 513.090 1704.000 ;
        RECT 462.210 1700.270 463.980 1700.410 ;
        RECT 462.210 1700.000 462.490 1700.270 ;
        RECT 463.840 1688.770 463.980 1700.270 ;
        RECT 512.810 1700.270 514.580 1700.410 ;
        RECT 512.810 1700.000 513.090 1700.270 ;
        RECT 514.440 1688.770 514.580 1700.270 ;
        RECT 463.780 1688.450 464.040 1688.770 ;
        RECT 468.840 1688.450 469.100 1688.770 ;
        RECT 514.380 1688.450 514.640 1688.770 ;
        RECT 517.140 1688.450 517.400 1688.770 ;
        RECT 468.900 1010.810 469.040 1688.450 ;
        RECT 517.200 1011.150 517.340 1688.450 ;
        RECT 517.140 1010.830 517.400 1011.150 ;
        RECT 468.840 1010.490 469.100 1010.810 ;
        RECT 638.180 1008.090 638.320 1987.310 ;
        RECT 650.600 1012.510 650.740 1988.330 ;
        RECT 650.540 1012.190 650.800 1012.510 ;
        RECT 672.160 1012.190 672.420 1012.510 ;
        RECT 638.120 1007.770 638.380 1008.090 ;
        RECT 670.780 1007.770 671.040 1008.090 ;
        RECT 670.840 1000.010 670.980 1007.770 ;
        RECT 672.220 1000.010 672.360 1012.190 ;
        RECT 686.480 1011.830 686.620 2767.950 ;
        RECT 707.120 2767.610 707.380 2767.930 ;
        RECT 700.220 2683.970 700.480 2684.290 ;
        RECT 686.420 1011.510 686.680 1011.830 ;
        RECT 700.280 1011.490 700.420 2683.970 ;
        RECT 700.220 1011.170 700.480 1011.490 ;
        RECT 707.180 1010.810 707.320 2767.610 ;
        RECT 755.420 2767.270 755.680 2767.590 ;
        RECT 720.920 2591.490 721.180 2591.810 ;
        RECT 720.980 1011.150 721.120 2591.490 ;
        RECT 755.480 1012.170 755.620 2767.270 ;
        RECT 769.220 2663.570 769.480 2663.890 ;
        RECT 762.320 2591.150 762.580 2591.470 ;
        RECT 762.380 1012.510 762.520 2591.150 ;
        RECT 769.280 1012.850 769.420 2663.570 ;
        RECT 783.080 1013.190 783.220 2769.310 ;
        RECT 975.300 2604.410 975.560 2604.730 ;
        RECT 843.280 1977.790 843.540 1978.110 ;
        RECT 783.020 1012.870 783.280 1013.190 ;
        RECT 769.220 1012.530 769.480 1012.850 ;
        RECT 762.320 1012.190 762.580 1012.510 ;
        RECT 755.420 1011.850 755.680 1012.170 ;
        RECT 841.900 1011.510 842.160 1011.830 ;
        RECT 712.640 1010.830 712.900 1011.150 ;
        RECT 720.920 1010.830 721.180 1011.150 ;
        RECT 673.540 1010.490 673.800 1010.810 ;
        RECT 707.120 1010.490 707.380 1010.810 ;
        RECT 673.600 1000.010 673.740 1010.490 ;
        RECT 712.700 1000.010 712.840 1010.830 ;
        RECT 841.960 1000.010 842.100 1011.510 ;
        RECT 843.340 1000.010 843.480 1977.790 ;
        RECT 897.560 1977.450 897.820 1977.770 ;
        RECT 845.580 1012.870 845.840 1013.190 ;
        RECT 845.640 1000.010 845.780 1012.870 ;
        RECT 890.200 1012.530 890.460 1012.850 ;
        RECT 884.680 1012.190 884.940 1012.510 ;
        RECT 884.740 1000.010 884.880 1012.190 ;
        RECT 890.260 1000.010 890.400 1012.530 ;
        RECT 893.420 1011.170 893.680 1011.490 ;
        RECT 893.480 1000.010 893.620 1011.170 ;
        RECT 897.620 1000.010 897.760 1977.450 ;
        RECT 975.360 1693.870 975.500 2604.410 ;
        RECT 977.600 2050.210 977.860 2050.530 ;
        RECT 977.140 2047.490 977.400 2047.810 ;
        RECT 975.760 2047.150 976.020 2047.470 ;
        RECT 975.300 1693.550 975.560 1693.870 ;
        RECT 975.820 1025.430 975.960 2047.150 ;
        RECT 976.680 2046.130 976.940 2046.450 ;
        RECT 976.220 2045.450 976.480 2045.770 ;
        RECT 975.760 1025.110 976.020 1025.430 ;
        RECT 976.280 1025.090 976.420 2045.450 ;
        RECT 976.220 1024.770 976.480 1025.090 ;
        RECT 976.740 1013.870 976.880 2046.130 ;
        RECT 976.680 1013.550 976.940 1013.870 ;
        RECT 910.900 1011.850 911.160 1012.170 ;
        RECT 906.300 1010.830 906.560 1011.150 ;
        RECT 901.700 1010.490 901.960 1010.810 ;
        RECT 901.760 1000.010 901.900 1010.490 ;
        RECT 906.360 1000.010 906.500 1010.830 ;
        RECT 910.960 1000.010 911.100 1011.850 ;
        RECT 977.200 1010.130 977.340 2047.490 ;
        RECT 977.660 1012.510 977.800 2050.210 ;
        RECT 978.060 2049.870 978.320 2050.190 ;
        RECT 977.600 1012.190 977.860 1012.510 ;
        RECT 978.120 1011.830 978.260 2049.870 ;
        RECT 978.580 1013.725 978.720 2809.770 ;
        RECT 978.510 1013.355 978.790 1013.725 ;
        RECT 979.040 1013.045 979.180 2810.110 ;
        RECT 986.340 2809.430 986.600 2809.750 ;
        RECT 979.440 2809.090 979.700 2809.410 ;
        RECT 978.970 1012.675 979.250 1013.045 ;
        RECT 978.060 1011.510 978.320 1011.830 ;
        RECT 977.140 1009.810 977.400 1010.130 ;
        RECT 979.500 1009.790 979.640 2809.090 ;
        RECT 985.880 2808.750 986.140 2809.070 ;
        RECT 985.420 2800.930 985.680 2801.250 ;
        RECT 982.200 2604.750 982.460 2605.070 ;
        RECT 981.740 2591.150 982.000 2591.470 ;
        RECT 981.800 1695.230 981.940 2591.150 ;
        RECT 981.740 1694.910 982.000 1695.230 ;
        RECT 982.260 1694.210 982.400 2604.750 ;
        RECT 984.960 2049.190 985.220 2049.510 ;
        RECT 984.040 2048.170 984.300 2048.490 ;
        RECT 983.120 2046.810 983.380 2047.130 ;
        RECT 982.660 2045.790 982.920 2046.110 ;
        RECT 982.200 1693.890 982.460 1694.210 ;
        RECT 982.720 1024.750 982.860 2045.790 ;
        RECT 983.180 1025.770 983.320 2046.810 ;
        RECT 983.580 2046.470 983.840 2046.790 ;
        RECT 983.120 1025.450 983.380 1025.770 ;
        RECT 982.660 1024.430 982.920 1024.750 ;
        RECT 983.640 1014.210 983.780 2046.470 ;
        RECT 983.580 1013.890 983.840 1014.210 ;
        RECT 979.440 1009.470 979.700 1009.790 ;
        RECT 984.100 1009.110 984.240 2048.170 ;
        RECT 984.500 2047.830 984.760 2048.150 ;
        RECT 984.560 1010.470 984.700 2047.830 ;
        RECT 985.020 1012.850 985.160 2049.190 ;
        RECT 984.960 1012.530 985.220 1012.850 ;
        RECT 985.480 1011.685 985.620 2800.930 ;
        RECT 985.940 1012.365 986.080 2808.750 ;
        RECT 986.400 1014.405 986.540 2809.430 ;
        RECT 1000.660 2809.070 1000.800 2810.450 ;
        RECT 1027.740 2809.770 1028.000 2810.090 ;
        RECT 1000.600 2808.750 1000.860 2809.070 ;
        RECT 1010.260 2800.930 1010.520 2801.250 ;
        RECT 1010.320 2799.970 1010.460 2800.930 ;
        RECT 1027.800 2800.000 1027.940 2809.770 ;
        RECT 1043.380 2809.430 1043.640 2809.750 ;
        RECT 1043.440 2800.000 1043.580 2809.430 ;
        RECT 1048.500 2808.730 1048.640 2810.450 ;
        RECT 1073.740 2810.110 1074.000 2810.430 ;
        RECT 1058.100 2809.090 1058.360 2809.410 ;
        RECT 1048.440 2808.410 1048.700 2808.730 ;
        RECT 1058.160 2800.000 1058.300 2809.090 ;
        RECT 1073.800 2800.000 1073.940 2810.110 ;
        RECT 1089.380 2808.410 1089.640 2808.730 ;
        RECT 1089.440 2800.000 1089.580 2808.410 ;
        RECT 1012.050 2799.970 1012.330 2800.000 ;
        RECT 1010.320 2799.830 1012.330 2799.970 ;
        RECT 1012.050 2796.000 1012.330 2799.830 ;
        RECT 1027.690 2796.000 1027.970 2800.000 ;
        RECT 1043.330 2796.000 1043.610 2800.000 ;
        RECT 1058.050 2796.000 1058.330 2800.000 ;
        RECT 1073.690 2796.000 1073.970 2800.000 ;
        RECT 1089.330 2796.000 1089.610 2800.000 ;
      LAYER met2 ;
        RECT 1002.860 2795.720 1011.770 2796.000 ;
        RECT 1012.610 2795.720 1027.410 2796.000 ;
        RECT 1028.250 2795.720 1043.050 2796.000 ;
        RECT 1043.890 2795.720 1057.770 2796.000 ;
        RECT 1058.610 2795.720 1073.410 2796.000 ;
        RECT 1074.250 2795.720 1089.050 2796.000 ;
        RECT 1089.890 2795.720 1095.120 2796.000 ;
      LAYER met2 ;
        RECT 993.230 2783.395 993.510 2783.765 ;
        RECT 992.770 2760.275 993.050 2760.645 ;
        RECT 992.310 2718.795 992.590 2719.165 ;
        RECT 991.850 2692.275 992.130 2692.645 ;
        RECT 991.390 2622.915 991.670 2623.285 ;
        RECT 990.930 1997.995 991.210 1998.365 ;
        RECT 990.470 1955.835 990.750 1956.205 ;
        RECT 990.010 1935.435 990.290 1935.805 ;
        RECT 989.550 1893.275 989.830 1893.645 ;
        RECT 989.090 1851.115 989.370 1851.485 ;
        RECT 988.630 1808.955 988.910 1809.325 ;
        RECT 988.170 1787.195 988.450 1787.565 ;
        RECT 987.710 1766.795 987.990 1767.165 ;
        RECT 987.250 1745.035 987.530 1745.405 ;
        RECT 987.320 1020.670 987.460 1745.035 ;
        RECT 987.260 1020.350 987.520 1020.670 ;
        RECT 987.780 1018.630 987.920 1766.795 ;
        RECT 988.240 1021.010 988.380 1787.195 ;
        RECT 988.180 1020.690 988.440 1021.010 ;
        RECT 988.700 1019.650 988.840 1808.955 ;
        RECT 988.640 1019.330 988.900 1019.650 ;
        RECT 987.720 1018.310 987.980 1018.630 ;
        RECT 989.160 1018.290 989.300 1851.115 ;
        RECT 989.620 1019.310 989.760 1893.275 ;
        RECT 989.560 1018.990 989.820 1019.310 ;
        RECT 989.100 1017.970 989.360 1018.290 ;
        RECT 990.080 1017.950 990.220 1935.435 ;
        RECT 990.020 1017.630 990.280 1017.950 ;
        RECT 990.540 1017.610 990.680 1955.835 ;
        RECT 991.000 1018.970 991.140 1997.995 ;
        RECT 990.940 1018.650 991.200 1018.970 ;
        RECT 990.480 1017.290 990.740 1017.610 ;
        RECT 986.330 1014.035 986.610 1014.405 ;
        RECT 991.460 1013.190 991.600 2622.915 ;
        RECT 991.920 1016.930 992.060 2692.275 ;
        RECT 991.860 1016.610 992.120 1016.930 ;
        RECT 991.400 1012.870 991.660 1013.190 ;
        RECT 985.870 1011.995 986.150 1012.365 ;
        RECT 985.410 1011.315 985.690 1011.685 ;
        RECT 984.500 1010.150 984.760 1010.470 ;
        RECT 984.040 1008.790 984.300 1009.110 ;
        RECT 992.380 1008.090 992.520 2718.795 ;
        RECT 992.840 1008.430 992.980 2760.275 ;
        RECT 993.300 1010.325 993.440 2783.395 ;
        RECT 994.610 2739.195 994.890 2739.565 ;
        RECT 993.690 2670.515 993.970 2670.885 ;
        RECT 993.230 1009.955 993.510 1010.325 ;
        RECT 993.760 1008.770 993.900 2670.515 ;
        RECT 994.150 2646.035 994.430 2646.405 ;
        RECT 993.700 1008.450 993.960 1008.770 ;
        RECT 992.780 1008.110 993.040 1008.430 ;
        RECT 992.320 1007.770 992.580 1008.090 ;
        RECT 994.220 1007.750 994.360 2646.035 ;
        RECT 994.680 1459.270 994.820 2739.195 ;
        RECT 998.760 2605.430 999.020 2605.750 ;
        RECT 995.070 2018.395 995.350 2018.765 ;
        RECT 994.620 1458.950 994.880 1459.270 ;
        RECT 995.140 1011.005 995.280 2018.395 ;
        RECT 995.530 1976.235 995.810 1976.605 ;
        RECT 995.600 1011.150 995.740 1976.235 ;
        RECT 995.990 1913.675 996.270 1914.045 ;
        RECT 996.060 1019.990 996.200 1913.675 ;
        RECT 996.450 1871.515 996.730 1871.885 ;
        RECT 996.000 1019.670 996.260 1019.990 ;
        RECT 995.070 1010.635 995.350 1011.005 ;
        RECT 995.540 1010.830 995.800 1011.150 ;
        RECT 996.520 1010.810 996.660 1871.515 ;
        RECT 996.910 1829.355 997.190 1829.725 ;
        RECT 996.980 1020.330 997.120 1829.355 ;
        RECT 997.370 1724.635 997.650 1725.005 ;
        RECT 997.440 1021.350 997.580 1724.635 ;
        RECT 998.300 1713.610 998.560 1713.930 ;
        RECT 997.380 1021.030 997.640 1021.350 ;
        RECT 996.920 1020.010 997.180 1020.330 ;
        RECT 996.460 1010.490 996.720 1010.810 ;
        RECT 998.360 1009.450 998.500 1713.610 ;
        RECT 998.820 1694.890 998.960 2605.430 ;
        RECT 999.220 2605.090 999.480 2605.410 ;
        RECT 998.760 1694.570 999.020 1694.890 ;
        RECT 999.280 1694.550 999.420 2605.090 ;
      LAYER met2 ;
        RECT 1002.860 2604.280 1095.120 2795.720 ;
      LAYER met2 ;
        RECT 1110.990 2780.675 1111.270 2781.045 ;
        RECT 1097.190 2644.675 1097.470 2645.045 ;
      LAYER met2 ;
        RECT 1003.410 2604.000 1017.290 2604.280 ;
        RECT 1018.130 2604.000 1032.930 2604.280 ;
        RECT 1033.770 2604.000 1048.570 2604.280 ;
        RECT 1049.410 2604.000 1064.210 2604.280 ;
        RECT 1065.050 2604.000 1079.850 2604.280 ;
        RECT 1080.690 2604.000 1094.570 2604.280 ;
      LAYER met2 ;
        RECT 1002.850 2600.730 1003.130 2604.000 ;
        RECT 1017.570 2600.730 1017.850 2604.000 ;
        RECT 1001.120 2600.590 1003.130 2600.730 ;
        RECT 1000.140 2050.550 1000.400 2050.870 ;
        RECT 999.680 2049.530 999.940 2049.850 ;
        RECT 999.220 1694.230 999.480 1694.550 ;
        RECT 999.740 1012.170 999.880 2049.530 ;
        RECT 1000.200 1013.530 1000.340 2050.550 ;
        RECT 1001.120 1713.930 1001.260 2600.590 ;
        RECT 1002.850 2600.000 1003.130 2600.590 ;
        RECT 1014.460 2600.590 1017.850 2600.730 ;
        RECT 1002.900 2049.190 1003.160 2049.510 ;
        RECT 1002.960 2044.110 1003.100 2049.190 ;
        RECT 1014.460 2048.490 1014.600 2600.590 ;
        RECT 1017.570 2600.000 1017.850 2600.590 ;
        RECT 1033.210 2600.000 1033.490 2604.000 ;
        RECT 1048.850 2600.000 1049.130 2604.000 ;
        RECT 1064.490 2600.730 1064.770 2604.000 ;
        RECT 1080.130 2600.730 1080.410 2604.000 ;
        RECT 1062.760 2600.590 1064.770 2600.730 ;
        RECT 1033.320 2587.730 1033.460 2600.000 ;
        RECT 1028.200 2587.410 1028.460 2587.730 ;
        RECT 1033.260 2587.410 1033.520 2587.730 ;
        RECT 1016.700 2052.590 1016.960 2052.910 ;
        RECT 1014.400 2048.170 1014.660 2048.490 ;
        RECT 1016.760 2044.110 1016.900 2052.590 ;
        RECT 1028.260 2048.150 1028.400 2587.410 ;
        RECT 1031.420 2052.930 1031.680 2053.250 ;
        RECT 1028.200 2047.830 1028.460 2048.150 ;
        RECT 1031.480 2044.110 1031.620 2052.930 ;
        RECT 1045.220 2049.530 1045.480 2049.850 ;
        RECT 1045.280 2044.110 1045.420 2049.530 ;
        RECT 1048.960 2047.810 1049.100 2600.000 ;
        RECT 1059.940 2053.270 1060.200 2053.590 ;
        RECT 1048.900 2047.490 1049.160 2047.810 ;
        RECT 1060.000 2044.110 1060.140 2053.270 ;
        RECT 1062.760 2047.470 1062.900 2600.590 ;
        RECT 1064.490 2600.000 1064.770 2600.590 ;
        RECT 1076.560 2600.590 1080.410 2600.730 ;
        RECT 1073.740 2049.870 1074.000 2050.190 ;
        RECT 1062.700 2047.150 1062.960 2047.470 ;
        RECT 1073.800 2044.110 1073.940 2049.870 ;
        RECT 1076.560 2047.130 1076.700 2600.590 ;
        RECT 1080.130 2600.000 1080.410 2600.590 ;
        RECT 1094.850 2600.000 1095.130 2604.000 ;
        RECT 1094.960 2591.470 1095.100 2600.000 ;
        RECT 1094.900 2591.150 1095.160 2591.470 ;
        RECT 1088.460 2050.550 1088.720 2050.870 ;
        RECT 1076.500 2046.810 1076.760 2047.130 ;
        RECT 1088.520 2044.110 1088.660 2050.550 ;
        RECT 1097.260 2046.790 1097.400 2644.675 ;
        RECT 1097.650 2622.235 1097.930 2622.605 ;
        RECT 1097.200 2046.470 1097.460 2046.790 ;
        RECT 1097.720 2046.450 1097.860 2622.235 ;
        RECT 1102.260 2050.210 1102.520 2050.530 ;
        RECT 1097.660 2046.130 1097.920 2046.450 ;
        RECT 1102.320 2044.110 1102.460 2050.210 ;
        RECT 1111.060 2046.110 1111.200 2780.675 ;
        RECT 1111.450 2760.275 1111.730 2760.645 ;
        RECT 1111.000 2045.790 1111.260 2046.110 ;
        RECT 1111.520 2045.770 1111.660 2760.275 ;
        RECT 1111.910 2734.435 1112.190 2734.805 ;
        RECT 1111.980 2605.750 1112.120 2734.435 ;
        RECT 1112.370 2712.675 1112.650 2713.045 ;
        RECT 1111.920 2605.430 1112.180 2605.750 ;
        RECT 1112.440 2605.070 1112.580 2712.675 ;
        RECT 1112.830 2691.595 1113.110 2691.965 ;
        RECT 1112.900 2605.410 1113.040 2691.595 ;
        RECT 1113.290 2666.435 1113.570 2666.805 ;
        RECT 1112.840 2605.090 1113.100 2605.410 ;
        RECT 1112.380 2604.750 1112.640 2605.070 ;
        RECT 1113.360 2604.730 1113.500 2666.435 ;
        RECT 1113.300 2604.410 1113.560 2604.730 ;
        RECT 1272.920 2055.310 1273.180 2055.630 ;
        RECT 1347.900 2055.310 1348.160 2055.630 ;
        RECT 1130.780 2054.290 1131.040 2054.610 ;
        RECT 1116.980 2053.950 1117.240 2054.270 ;
        RECT 1111.460 2045.450 1111.720 2045.770 ;
        RECT 1117.040 2044.110 1117.180 2053.950 ;
        RECT 1130.840 2044.110 1130.980 2054.290 ;
        RECT 1230.140 2053.610 1230.400 2053.930 ;
        RECT 1201.620 2052.250 1201.880 2052.570 ;
        RECT 1187.820 2051.910 1188.080 2052.230 ;
        RECT 1173.100 2051.570 1173.360 2051.890 ;
        RECT 1159.300 2051.230 1159.560 2051.550 ;
        RECT 1144.580 2050.890 1144.840 2051.210 ;
        RECT 1144.640 2044.110 1144.780 2050.890 ;
        RECT 1159.360 2044.110 1159.500 2051.230 ;
        RECT 1173.160 2044.110 1173.300 2051.570 ;
        RECT 1187.880 2044.110 1188.020 2051.910 ;
        RECT 1201.680 2044.110 1201.820 2052.250 ;
        RECT 1216.340 2049.530 1216.600 2049.850 ;
        RECT 1216.400 2044.110 1216.540 2049.530 ;
        RECT 1230.200 2044.110 1230.340 2053.610 ;
        RECT 1272.980 2052.910 1273.120 2055.310 ;
        RECT 1273.380 2054.970 1273.640 2055.290 ;
        RECT 1331.800 2054.970 1332.060 2055.290 ;
        RECT 1272.920 2052.590 1273.180 2052.910 ;
        RECT 1258.660 2050.550 1258.920 2050.870 ;
        RECT 1244.860 2049.870 1245.120 2050.190 ;
        RECT 1244.920 2044.110 1245.060 2049.870 ;
        RECT 1258.720 2044.110 1258.860 2050.550 ;
        RECT 1273.440 2044.110 1273.580 2054.970 ;
        RECT 1293.620 2054.630 1293.880 2054.950 ;
        RECT 1293.680 2053.590 1293.820 2054.630 ;
        RECT 1293.620 2053.270 1293.880 2053.590 ;
        RECT 1294.080 2053.270 1294.340 2053.590 ;
        RECT 1286.260 2052.590 1286.520 2052.910 ;
        RECT 1286.320 2051.890 1286.460 2052.590 ;
        RECT 1294.140 2052.230 1294.280 2053.270 ;
        RECT 1294.080 2051.910 1294.340 2052.230 ;
        RECT 1301.900 2051.910 1302.160 2052.230 ;
        RECT 1286.260 2051.570 1286.520 2051.890 ;
        RECT 1286.720 2051.570 1286.980 2051.890 ;
        RECT 1286.780 2050.870 1286.920 2051.570 ;
        RECT 1286.720 2050.550 1286.980 2050.870 ;
        RECT 1287.180 2050.550 1287.440 2050.870 ;
        RECT 1287.240 2044.110 1287.380 2050.550 ;
        RECT 1301.960 2044.110 1302.100 2051.910 ;
        RECT 1315.700 2049.530 1315.960 2049.850 ;
        RECT 1315.760 2044.110 1315.900 2049.530 ;
        RECT 1329.500 2049.190 1329.760 2049.510 ;
        RECT 1329.560 2044.110 1329.700 2049.190 ;
        RECT 1002.850 2040.110 1003.130 2044.110 ;
        RECT 1016.650 2040.110 1016.930 2044.110 ;
        RECT 1031.370 2040.110 1031.650 2044.110 ;
        RECT 1045.170 2040.110 1045.450 2044.110 ;
        RECT 1059.890 2040.110 1060.170 2044.110 ;
        RECT 1073.690 2040.110 1073.970 2044.110 ;
        RECT 1088.410 2040.110 1088.690 2044.110 ;
        RECT 1102.210 2040.110 1102.490 2044.110 ;
        RECT 1116.930 2040.110 1117.210 2044.110 ;
        RECT 1130.730 2040.110 1131.010 2044.110 ;
        RECT 1144.530 2040.110 1144.810 2044.110 ;
        RECT 1159.250 2040.110 1159.530 2044.110 ;
        RECT 1173.050 2040.110 1173.330 2044.110 ;
        RECT 1187.770 2040.110 1188.050 2044.110 ;
        RECT 1201.570 2040.110 1201.850 2044.110 ;
        RECT 1216.290 2040.110 1216.570 2044.110 ;
        RECT 1230.090 2040.110 1230.370 2044.110 ;
        RECT 1244.810 2040.110 1245.090 2044.110 ;
        RECT 1258.610 2040.110 1258.890 2044.110 ;
        RECT 1273.330 2040.110 1273.610 2044.110 ;
        RECT 1287.130 2040.110 1287.410 2044.110 ;
        RECT 1301.850 2040.110 1302.130 2044.110 ;
        RECT 1315.650 2040.110 1315.930 2044.110 ;
        RECT 1329.450 2040.110 1329.730 2044.110 ;
      LAYER met2 ;
        RECT 1003.410 2039.830 1016.370 2040.110 ;
        RECT 1017.210 2039.830 1031.090 2040.110 ;
        RECT 1031.930 2039.830 1044.890 2040.110 ;
        RECT 1045.730 2039.830 1059.610 2040.110 ;
        RECT 1060.450 2039.830 1073.410 2040.110 ;
        RECT 1074.250 2039.830 1088.130 2040.110 ;
        RECT 1088.970 2039.830 1101.930 2040.110 ;
        RECT 1102.770 2039.830 1116.650 2040.110 ;
        RECT 1117.490 2039.830 1130.450 2040.110 ;
        RECT 1131.290 2039.830 1144.250 2040.110 ;
        RECT 1145.090 2039.830 1158.970 2040.110 ;
        RECT 1159.810 2039.830 1172.770 2040.110 ;
        RECT 1173.610 2039.830 1187.490 2040.110 ;
        RECT 1188.330 2039.830 1201.290 2040.110 ;
        RECT 1202.130 2039.830 1216.010 2040.110 ;
        RECT 1216.850 2039.830 1229.810 2040.110 ;
        RECT 1230.650 2039.830 1244.530 2040.110 ;
        RECT 1245.370 2039.830 1258.330 2040.110 ;
        RECT 1259.170 2039.830 1273.050 2040.110 ;
        RECT 1273.890 2039.830 1286.850 2040.110 ;
        RECT 1287.690 2039.830 1301.570 2040.110 ;
        RECT 1302.410 2039.830 1315.370 2040.110 ;
        RECT 1316.210 2039.830 1329.170 2040.110 ;
      LAYER met2 ;
        RECT 1001.060 1713.610 1001.320 1713.930 ;
      LAYER met2 ;
        RECT 1002.860 1704.280 1329.720 2039.830 ;
        RECT 1003.410 1704.000 1016.370 1704.280 ;
        RECT 1017.210 1704.000 1030.170 1704.280 ;
        RECT 1031.010 1704.000 1044.890 1704.280 ;
        RECT 1045.730 1704.000 1058.690 1704.280 ;
        RECT 1059.530 1704.000 1073.410 1704.280 ;
        RECT 1074.250 1704.000 1087.210 1704.280 ;
        RECT 1088.050 1704.000 1101.930 1704.280 ;
        RECT 1102.770 1704.000 1115.730 1704.280 ;
        RECT 1116.570 1704.000 1130.450 1704.280 ;
        RECT 1131.290 1704.000 1144.250 1704.280 ;
        RECT 1145.090 1704.000 1158.970 1704.280 ;
        RECT 1159.810 1704.000 1172.770 1704.280 ;
        RECT 1173.610 1704.000 1187.490 1704.280 ;
        RECT 1188.330 1704.000 1201.290 1704.280 ;
        RECT 1202.130 1704.000 1215.090 1704.280 ;
        RECT 1215.930 1704.000 1229.810 1704.280 ;
        RECT 1230.650 1704.000 1243.610 1704.280 ;
        RECT 1244.450 1704.000 1258.330 1704.280 ;
        RECT 1259.170 1704.000 1272.130 1704.280 ;
        RECT 1272.970 1704.000 1286.850 1704.280 ;
        RECT 1287.690 1704.000 1300.650 1704.280 ;
        RECT 1301.490 1704.000 1315.370 1704.280 ;
        RECT 1316.210 1704.000 1329.170 1704.280 ;
      LAYER met2 ;
        RECT 1002.850 1700.000 1003.130 1704.000 ;
        RECT 1016.650 1700.000 1016.930 1704.000 ;
        RECT 1030.450 1700.000 1030.730 1704.000 ;
        RECT 1045.170 1700.410 1045.450 1704.000 ;
        RECT 1045.170 1700.270 1048.640 1700.410 ;
        RECT 1045.170 1700.000 1045.450 1700.270 ;
        RECT 1002.960 1684.350 1003.100 1700.000 ;
        RECT 1016.760 1688.770 1016.900 1700.000 ;
        RECT 1016.700 1688.450 1016.960 1688.770 ;
        RECT 1030.560 1688.430 1030.700 1700.000 ;
        RECT 1038.320 1688.450 1038.580 1688.770 ;
        RECT 1030.500 1688.110 1030.760 1688.430 ;
        RECT 1002.900 1684.030 1003.160 1684.350 ;
        RECT 1007.040 1684.030 1007.300 1684.350 ;
        RECT 1000.140 1013.210 1000.400 1013.530 ;
        RECT 999.680 1011.850 999.940 1012.170 ;
        RECT 1007.100 1011.490 1007.240 1684.030 ;
        RECT 1038.380 1013.190 1038.520 1688.450 ;
        RECT 1048.500 1017.270 1048.640 1700.270 ;
        RECT 1058.970 1700.000 1059.250 1704.000 ;
        RECT 1073.690 1700.000 1073.970 1704.000 ;
        RECT 1087.490 1700.410 1087.770 1704.000 ;
        RECT 1087.490 1700.270 1090.040 1700.410 ;
        RECT 1087.490 1700.000 1087.770 1700.270 ;
        RECT 1048.900 1694.910 1049.160 1695.230 ;
        RECT 1048.960 1076.170 1049.100 1694.910 ;
        RECT 1059.080 1689.110 1059.220 1700.000 ;
        RECT 1069.600 1694.570 1069.860 1694.890 ;
        RECT 1059.020 1688.790 1059.280 1689.110 ;
        RECT 1069.660 1110.770 1069.800 1694.570 ;
        RECT 1073.800 1688.770 1073.940 1700.000 ;
        RECT 1076.500 1694.230 1076.760 1694.550 ;
        RECT 1073.740 1688.450 1074.000 1688.770 ;
        RECT 1069.600 1110.450 1069.860 1110.770 ;
        RECT 1070.980 1110.450 1071.240 1110.770 ;
        RECT 1048.960 1076.030 1049.560 1076.170 ;
        RECT 1049.420 1028.570 1049.560 1076.030 ;
        RECT 1071.040 1062.830 1071.180 1110.450 ;
        RECT 1070.980 1062.510 1071.240 1062.830 ;
        RECT 1071.900 1062.510 1072.160 1062.830 ;
        RECT 1049.420 1028.430 1050.020 1028.570 ;
        RECT 1048.440 1016.950 1048.700 1017.270 ;
        RECT 1014.400 1012.870 1014.660 1013.190 ;
        RECT 1038.320 1012.870 1038.580 1013.190 ;
        RECT 1007.040 1011.170 1007.300 1011.490 ;
        RECT 998.300 1009.130 998.560 1009.450 ;
        RECT 994.160 1007.430 994.420 1007.750 ;
        RECT 1014.460 1000.010 1014.600 1012.870 ;
        RECT 670.840 1000.000 671.140 1000.010 ;
        RECT 672.220 1000.000 672.980 1000.010 ;
        RECT 673.600 1000.000 675.280 1000.010 ;
        RECT 712.700 1000.000 714.380 1000.010 ;
        RECT 841.960 1000.000 842.720 1000.010 ;
        RECT 843.340 1000.000 845.020 1000.010 ;
        RECT 845.640 1000.000 846.860 1000.010 ;
        RECT 884.740 1000.000 885.960 1000.010 ;
        RECT 890.260 1000.000 890.560 1000.010 ;
        RECT 893.480 1000.000 894.700 1000.010 ;
        RECT 897.620 1000.000 899.300 1000.010 ;
        RECT 901.760 1000.000 903.440 1000.010 ;
        RECT 906.360 1000.000 908.040 1000.010 ;
        RECT 910.960 1000.000 912.180 1000.010 ;
        RECT 1014.300 1000.000 1014.600 1000.010 ;
        RECT 1049.880 1000.010 1050.020 1028.430 ;
        RECT 1067.290 1009.955 1067.570 1010.325 ;
        RECT 1062.700 1008.110 1062.960 1008.430 ;
        RECT 1055.800 1007.770 1056.060 1008.090 ;
        RECT 1055.860 1000.010 1056.000 1007.770 ;
        RECT 1058.560 1007.430 1058.820 1007.750 ;
        RECT 1049.880 1000.000 1051.560 1000.010 ;
        RECT 1055.700 1000.000 1056.000 1000.010 ;
        RECT 1058.620 1000.010 1058.760 1007.430 ;
        RECT 1062.760 1000.010 1062.900 1008.110 ;
        RECT 1067.360 1000.010 1067.500 1009.955 ;
        RECT 1071.960 1000.010 1072.100 1062.510 ;
        RECT 1076.560 1000.010 1076.700 1694.230 ;
        RECT 1089.900 1010.470 1090.040 1700.270 ;
        RECT 1102.210 1700.000 1102.490 1704.000 ;
        RECT 1116.010 1700.000 1116.290 1704.000 ;
        RECT 1130.730 1700.000 1131.010 1704.000 ;
        RECT 1144.530 1700.000 1144.810 1704.000 ;
        RECT 1159.250 1700.000 1159.530 1704.000 ;
        RECT 1173.050 1700.000 1173.330 1704.000 ;
        RECT 1187.770 1700.000 1188.050 1704.000 ;
        RECT 1201.570 1700.410 1201.850 1704.000 ;
        RECT 1200.760 1700.270 1201.850 1700.410 ;
        RECT 1102.320 1689.450 1102.460 1700.000 ;
        RECT 1111.000 1693.890 1111.260 1694.210 ;
        RECT 1104.100 1693.550 1104.360 1693.870 ;
        RECT 1102.260 1689.130 1102.520 1689.450 ;
        RECT 1101.790 1014.035 1102.070 1014.405 ;
        RECT 1104.160 1014.210 1104.300 1693.550 ;
        RECT 1084.320 1010.150 1084.580 1010.470 ;
        RECT 1089.840 1010.150 1090.100 1010.470 ;
        RECT 1080.180 1008.450 1080.440 1008.770 ;
        RECT 1080.240 1000.010 1080.380 1008.450 ;
        RECT 1084.380 1000.010 1084.520 1010.150 ;
        RECT 1090.300 1009.470 1090.560 1009.790 ;
        RECT 1090.360 1000.010 1090.500 1009.470 ;
        RECT 1097.660 1009.130 1097.920 1009.450 ;
        RECT 1093.060 1008.790 1093.320 1009.110 ;
        RECT 1093.120 1000.010 1093.260 1008.790 ;
        RECT 1097.720 1000.010 1097.860 1009.130 ;
        RECT 1101.860 1000.010 1102.000 1014.035 ;
        RECT 1104.100 1013.890 1104.360 1014.210 ;
        RECT 1106.400 1013.890 1106.660 1014.210 ;
        RECT 1103.180 1013.550 1103.440 1013.870 ;
        RECT 1103.240 1009.790 1103.380 1013.550 ;
        RECT 1103.180 1009.470 1103.440 1009.790 ;
        RECT 1106.460 1000.010 1106.600 1013.890 ;
        RECT 1111.060 1000.010 1111.200 1693.890 ;
        RECT 1116.120 1686.730 1116.260 1700.000 ;
        RECT 1130.840 1689.790 1130.980 1700.000 ;
        RECT 1130.780 1689.470 1131.040 1689.790 ;
        RECT 1116.060 1686.410 1116.320 1686.730 ;
        RECT 1144.640 1686.390 1144.780 1700.000 ;
        RECT 1159.360 1690.130 1159.500 1700.000 ;
        RECT 1159.300 1689.810 1159.560 1690.130 ;
        RECT 1144.580 1686.070 1144.840 1686.390 ;
        RECT 1173.160 1684.350 1173.300 1700.000 ;
        RECT 1186.440 1693.550 1186.700 1693.870 ;
        RECT 1180.000 1686.070 1180.260 1686.390 ;
        RECT 1173.100 1684.030 1173.360 1684.350 ;
        RECT 1159.300 1458.950 1159.560 1459.270 ;
        RECT 1159.360 1076.170 1159.500 1458.950 ;
        RECT 1159.360 1076.030 1159.960 1076.170 ;
        RECT 1159.820 1028.570 1159.960 1076.030 ;
        RECT 1159.820 1028.430 1160.880 1028.570 ;
        RECT 1152.860 1025.450 1153.120 1025.770 ;
        RECT 1147.800 1025.110 1148.060 1025.430 ;
        RECT 1125.720 1016.610 1125.980 1016.930 ;
        RECT 1119.270 1013.355 1119.550 1013.725 ;
        RECT 1115.140 1009.810 1115.400 1010.130 ;
        RECT 1115.200 1000.010 1115.340 1009.810 ;
        RECT 1119.340 1000.010 1119.480 1013.355 ;
        RECT 1125.780 1000.010 1125.920 1016.610 ;
        RECT 1134.460 1013.550 1134.720 1013.870 ;
        RECT 1131.690 1012.675 1131.970 1013.045 ;
        RECT 1131.760 1000.010 1131.900 1012.675 ;
        RECT 1058.620 1000.000 1059.840 1000.010 ;
        RECT 1062.760 1000.000 1064.440 1000.010 ;
        RECT 1067.360 1000.000 1068.580 1000.010 ;
        RECT 1071.960 1000.000 1073.180 1000.010 ;
        RECT 1076.560 1000.000 1077.320 1000.010 ;
        RECT 1080.240 1000.000 1081.920 1000.010 ;
        RECT 1084.380 1000.000 1086.060 1000.010 ;
        RECT 1090.360 1000.000 1090.660 1000.010 ;
        RECT 1093.120 1000.000 1094.800 1000.010 ;
        RECT 1097.720 1000.000 1099.400 1000.010 ;
        RECT 1101.860 1000.000 1103.540 1000.010 ;
        RECT 1106.460 1000.000 1107.680 1000.010 ;
        RECT 1111.060 1000.000 1112.280 1000.010 ;
        RECT 1115.200 1000.000 1116.420 1000.010 ;
        RECT 1119.340 1000.000 1121.020 1000.010 ;
        RECT 1125.780 1000.000 1127.460 1000.010 ;
        RECT 1131.600 1000.000 1131.900 1000.010 ;
        RECT 1134.520 1000.010 1134.660 1013.550 ;
        RECT 1143.190 1011.995 1143.470 1012.365 ;
        RECT 1139.060 1009.470 1139.320 1009.790 ;
        RECT 1139.120 1000.010 1139.260 1009.470 ;
        RECT 1143.260 1000.010 1143.400 1011.995 ;
        RECT 1147.860 1000.010 1148.000 1025.110 ;
        RECT 1152.920 1000.010 1153.060 1025.450 ;
        RECT 1156.080 1024.770 1156.340 1025.090 ;
        RECT 1156.140 1000.010 1156.280 1024.770 ;
        RECT 1160.740 1000.010 1160.880 1028.430 ;
        RECT 1166.200 1024.430 1166.460 1024.750 ;
        RECT 1180.060 1024.490 1180.200 1686.070 ;
        RECT 1166.260 1000.010 1166.400 1024.430 ;
        RECT 1180.060 1024.350 1182.500 1024.490 ;
        RECT 1181.840 1013.550 1182.100 1013.870 ;
        RECT 1167.110 1011.315 1167.390 1011.685 ;
        RECT 1167.180 1000.010 1167.320 1011.315 ;
        RECT 1181.900 1000.010 1182.040 1013.550 ;
        RECT 1134.520 1000.000 1136.200 1000.010 ;
        RECT 1139.120 1000.000 1140.340 1000.010 ;
        RECT 1143.260 1000.000 1144.940 1000.010 ;
        RECT 1147.860 1000.000 1149.080 1000.010 ;
        RECT 1152.920 1000.000 1153.680 1000.010 ;
        RECT 1156.140 1000.000 1157.820 1000.010 ;
        RECT 1160.740 1000.000 1162.420 1000.010 ;
        RECT 1166.260 1000.000 1166.560 1000.010 ;
        RECT 1167.180 1000.000 1168.860 1000.010 ;
        RECT 1181.740 1000.000 1182.040 1000.010 ;
        RECT 670.840 999.870 671.290 1000.000 ;
        RECT 672.220 999.870 673.130 1000.000 ;
        RECT 673.600 999.870 675.430 1000.000 ;
        RECT 671.010 996.000 671.290 999.870 ;
      LAYER met2 ;
        RECT 671.570 995.720 672.570 998.810 ;
      LAYER met2 ;
        RECT 672.850 996.000 673.130 999.870 ;
      LAYER met2 ;
        RECT 673.410 995.720 674.870 998.810 ;
      LAYER met2 ;
        RECT 675.150 996.000 675.430 999.870 ;
      LAYER met2 ;
        RECT 675.710 995.720 677.170 998.810 ;
      LAYER met2 ;
        RECT 677.450 996.000 677.730 1000.000 ;
      LAYER met2 ;
        RECT 678.010 995.720 679.010 998.810 ;
      LAYER met2 ;
        RECT 679.290 996.000 679.570 1000.000 ;
      LAYER met2 ;
        RECT 679.850 995.720 681.310 998.810 ;
      LAYER met2 ;
        RECT 681.590 996.000 681.870 1000.000 ;
      LAYER met2 ;
        RECT 682.150 995.720 683.610 998.810 ;
      LAYER met2 ;
        RECT 683.890 996.000 684.170 1000.000 ;
      LAYER met2 ;
        RECT 684.450 995.720 685.910 998.810 ;
      LAYER met2 ;
        RECT 686.190 996.000 686.470 1000.000 ;
      LAYER met2 ;
        RECT 686.750 995.720 687.750 998.810 ;
      LAYER met2 ;
        RECT 688.030 996.000 688.310 1000.000 ;
      LAYER met2 ;
        RECT 688.590 995.720 690.050 998.810 ;
      LAYER met2 ;
        RECT 690.330 996.000 690.610 1000.000 ;
      LAYER met2 ;
        RECT 690.890 995.720 692.350 998.810 ;
      LAYER met2 ;
        RECT 692.630 996.000 692.910 1000.000 ;
      LAYER met2 ;
        RECT 693.190 995.720 694.190 998.810 ;
      LAYER met2 ;
        RECT 694.470 996.000 694.750 1000.000 ;
      LAYER met2 ;
        RECT 695.030 995.720 696.490 998.810 ;
      LAYER met2 ;
        RECT 696.770 996.000 697.050 1000.000 ;
      LAYER met2 ;
        RECT 697.330 995.720 698.790 998.810 ;
      LAYER met2 ;
        RECT 699.070 996.000 699.350 1000.000 ;
      LAYER met2 ;
        RECT 699.630 995.720 701.090 998.810 ;
      LAYER met2 ;
        RECT 701.370 996.000 701.650 1000.000 ;
      LAYER met2 ;
        RECT 701.930 995.720 702.930 998.810 ;
      LAYER met2 ;
        RECT 703.210 996.000 703.490 1000.000 ;
      LAYER met2 ;
        RECT 703.770 995.720 705.230 998.810 ;
      LAYER met2 ;
        RECT 705.510 996.000 705.790 1000.000 ;
      LAYER met2 ;
        RECT 706.070 995.720 707.530 998.810 ;
      LAYER met2 ;
        RECT 707.810 996.000 708.090 1000.000 ;
      LAYER met2 ;
        RECT 708.370 995.720 709.830 998.810 ;
      LAYER met2 ;
        RECT 710.110 996.000 710.390 1000.000 ;
      LAYER met2 ;
        RECT 710.670 995.720 711.670 998.810 ;
      LAYER met2 ;
        RECT 711.950 996.000 712.230 1000.000 ;
        RECT 712.700 999.870 714.530 1000.000 ;
      LAYER met2 ;
        RECT 712.510 995.720 713.970 998.810 ;
      LAYER met2 ;
        RECT 714.250 996.000 714.530 999.870 ;
      LAYER met2 ;
        RECT 714.810 995.720 716.270 998.810 ;
      LAYER met2 ;
        RECT 716.550 996.000 716.830 1000.000 ;
      LAYER met2 ;
        RECT 717.110 995.720 718.110 998.810 ;
      LAYER met2 ;
        RECT 718.390 996.000 718.670 1000.000 ;
      LAYER met2 ;
        RECT 718.950 995.720 720.410 998.810 ;
      LAYER met2 ;
        RECT 720.690 996.000 720.970 1000.000 ;
      LAYER met2 ;
        RECT 721.250 995.720 722.710 998.810 ;
      LAYER met2 ;
        RECT 722.990 996.000 723.270 1000.000 ;
      LAYER met2 ;
        RECT 723.550 995.720 725.010 998.810 ;
      LAYER met2 ;
        RECT 725.290 996.000 725.570 1000.000 ;
      LAYER met2 ;
        RECT 725.850 995.720 726.850 998.810 ;
      LAYER met2 ;
        RECT 727.130 996.000 727.410 1000.000 ;
      LAYER met2 ;
        RECT 727.690 995.720 729.150 998.810 ;
      LAYER met2 ;
        RECT 729.430 996.000 729.710 1000.000 ;
      LAYER met2 ;
        RECT 729.990 995.720 731.450 998.810 ;
      LAYER met2 ;
        RECT 731.730 996.000 732.010 1000.000 ;
      LAYER met2 ;
        RECT 732.290 995.720 733.750 998.810 ;
      LAYER met2 ;
        RECT 734.030 996.000 734.310 1000.000 ;
      LAYER met2 ;
        RECT 734.590 995.720 735.590 998.810 ;
      LAYER met2 ;
        RECT 735.870 996.000 736.150 1000.000 ;
      LAYER met2 ;
        RECT 736.430 995.720 737.890 998.810 ;
      LAYER met2 ;
        RECT 738.170 996.000 738.450 1000.000 ;
      LAYER met2 ;
        RECT 738.730 995.720 740.190 998.810 ;
      LAYER met2 ;
        RECT 740.470 996.000 740.750 1000.000 ;
      LAYER met2 ;
        RECT 741.030 995.720 742.030 998.810 ;
      LAYER met2 ;
        RECT 742.310 996.000 742.590 1000.000 ;
      LAYER met2 ;
        RECT 742.870 995.720 744.330 998.810 ;
      LAYER met2 ;
        RECT 744.610 996.000 744.890 1000.000 ;
      LAYER met2 ;
        RECT 745.170 995.720 746.630 998.810 ;
      LAYER met2 ;
        RECT 746.910 996.000 747.190 1000.000 ;
      LAYER met2 ;
        RECT 747.470 995.720 748.930 998.810 ;
      LAYER met2 ;
        RECT 749.210 996.000 749.490 1000.000 ;
      LAYER met2 ;
        RECT 749.770 995.720 750.770 998.810 ;
      LAYER met2 ;
        RECT 751.050 996.000 751.330 1000.000 ;
      LAYER met2 ;
        RECT 751.610 995.720 753.070 998.810 ;
      LAYER met2 ;
        RECT 753.350 996.000 753.630 1000.000 ;
      LAYER met2 ;
        RECT 753.910 995.720 755.370 998.810 ;
      LAYER met2 ;
        RECT 755.650 996.000 755.930 1000.000 ;
      LAYER met2 ;
        RECT 756.210 995.720 757.670 998.810 ;
      LAYER met2 ;
        RECT 757.950 996.000 758.230 1000.000 ;
      LAYER met2 ;
        RECT 758.510 995.720 759.510 998.810 ;
      LAYER met2 ;
        RECT 759.790 996.000 760.070 1000.000 ;
      LAYER met2 ;
        RECT 760.350 995.720 761.810 998.810 ;
      LAYER met2 ;
        RECT 762.090 996.000 762.370 1000.000 ;
      LAYER met2 ;
        RECT 762.650 995.720 764.110 998.810 ;
      LAYER met2 ;
        RECT 764.390 996.000 764.670 1000.000 ;
      LAYER met2 ;
        RECT 764.950 995.720 765.950 998.810 ;
      LAYER met2 ;
        RECT 766.230 996.000 766.510 1000.000 ;
      LAYER met2 ;
        RECT 766.790 995.720 768.250 998.810 ;
      LAYER met2 ;
        RECT 768.530 996.000 768.810 1000.000 ;
      LAYER met2 ;
        RECT 769.090 995.720 770.550 998.810 ;
      LAYER met2 ;
        RECT 770.830 996.000 771.110 1000.000 ;
      LAYER met2 ;
        RECT 771.390 995.720 772.850 998.810 ;
      LAYER met2 ;
        RECT 773.130 996.000 773.410 1000.000 ;
      LAYER met2 ;
        RECT 773.690 995.720 774.690 998.810 ;
      LAYER met2 ;
        RECT 774.970 996.000 775.250 1000.000 ;
      LAYER met2 ;
        RECT 775.530 995.720 776.990 998.810 ;
      LAYER met2 ;
        RECT 777.270 996.000 777.550 1000.000 ;
      LAYER met2 ;
        RECT 777.830 995.720 779.290 998.810 ;
      LAYER met2 ;
        RECT 779.570 996.000 779.850 1000.000 ;
      LAYER met2 ;
        RECT 780.130 995.720 781.590 998.810 ;
      LAYER met2 ;
        RECT 781.870 996.000 782.150 1000.000 ;
      LAYER met2 ;
        RECT 782.430 995.720 783.430 998.810 ;
      LAYER met2 ;
        RECT 783.710 996.000 783.990 1000.000 ;
      LAYER met2 ;
        RECT 784.270 995.720 785.730 998.810 ;
      LAYER met2 ;
        RECT 786.010 996.000 786.290 1000.000 ;
      LAYER met2 ;
        RECT 786.570 995.720 788.030 998.810 ;
      LAYER met2 ;
        RECT 788.310 996.000 788.590 1000.000 ;
      LAYER met2 ;
        RECT 788.870 995.720 789.870 998.810 ;
      LAYER met2 ;
        RECT 790.150 996.000 790.430 1000.000 ;
      LAYER met2 ;
        RECT 790.710 995.720 792.170 998.810 ;
      LAYER met2 ;
        RECT 792.450 996.000 792.730 1000.000 ;
      LAYER met2 ;
        RECT 793.010 995.720 794.470 998.810 ;
      LAYER met2 ;
        RECT 794.750 996.000 795.030 1000.000 ;
      LAYER met2 ;
        RECT 795.310 995.720 796.770 998.810 ;
      LAYER met2 ;
        RECT 797.050 996.000 797.330 1000.000 ;
      LAYER met2 ;
        RECT 797.610 995.720 798.610 998.810 ;
      LAYER met2 ;
        RECT 798.890 996.000 799.170 1000.000 ;
      LAYER met2 ;
        RECT 799.450 995.720 800.910 998.810 ;
      LAYER met2 ;
        RECT 801.190 996.000 801.470 1000.000 ;
      LAYER met2 ;
        RECT 801.750 995.720 803.210 998.810 ;
      LAYER met2 ;
        RECT 803.490 996.000 803.770 1000.000 ;
      LAYER met2 ;
        RECT 804.050 995.720 805.510 998.810 ;
      LAYER met2 ;
        RECT 805.790 996.000 806.070 1000.000 ;
      LAYER met2 ;
        RECT 806.350 995.720 807.350 998.810 ;
      LAYER met2 ;
        RECT 807.630 996.000 807.910 1000.000 ;
      LAYER met2 ;
        RECT 808.190 995.720 809.650 998.810 ;
      LAYER met2 ;
        RECT 809.930 996.000 810.210 1000.000 ;
      LAYER met2 ;
        RECT 810.490 995.720 811.950 998.810 ;
      LAYER met2 ;
        RECT 812.230 996.000 812.510 1000.000 ;
      LAYER met2 ;
        RECT 812.790 995.720 813.790 998.810 ;
      LAYER met2 ;
        RECT 814.070 996.000 814.350 1000.000 ;
      LAYER met2 ;
        RECT 814.630 995.720 816.090 998.810 ;
      LAYER met2 ;
        RECT 816.370 996.000 816.650 1000.000 ;
      LAYER met2 ;
        RECT 816.930 995.720 818.390 998.810 ;
      LAYER met2 ;
        RECT 818.670 996.000 818.950 1000.000 ;
      LAYER met2 ;
        RECT 819.230 995.720 820.690 998.810 ;
      LAYER met2 ;
        RECT 820.970 996.000 821.250 1000.000 ;
      LAYER met2 ;
        RECT 821.530 995.720 822.530 998.810 ;
      LAYER met2 ;
        RECT 822.810 996.000 823.090 1000.000 ;
      LAYER met2 ;
        RECT 823.370 995.720 824.830 998.810 ;
      LAYER met2 ;
        RECT 825.110 996.000 825.390 1000.000 ;
      LAYER met2 ;
        RECT 825.670 995.720 827.130 998.810 ;
      LAYER met2 ;
        RECT 827.410 996.000 827.690 1000.000 ;
      LAYER met2 ;
        RECT 827.970 995.720 829.430 998.810 ;
      LAYER met2 ;
        RECT 829.710 996.000 829.990 1000.000 ;
      LAYER met2 ;
        RECT 830.270 995.720 831.270 998.810 ;
      LAYER met2 ;
        RECT 831.550 996.000 831.830 1000.000 ;
      LAYER met2 ;
        RECT 832.110 995.720 833.570 998.810 ;
      LAYER met2 ;
        RECT 833.850 996.000 834.130 1000.000 ;
      LAYER met2 ;
        RECT 834.410 995.720 835.870 998.810 ;
      LAYER met2 ;
        RECT 836.150 996.000 836.430 1000.000 ;
      LAYER met2 ;
        RECT 836.710 995.720 837.710 998.810 ;
      LAYER met2 ;
        RECT 837.990 996.000 838.270 1000.000 ;
      LAYER met2 ;
        RECT 838.550 995.720 840.010 998.810 ;
      LAYER met2 ;
        RECT 840.290 996.000 840.570 1000.000 ;
        RECT 841.960 999.870 842.870 1000.000 ;
        RECT 843.340 999.870 845.170 1000.000 ;
        RECT 845.640 999.870 847.010 1000.000 ;
      LAYER met2 ;
        RECT 840.850 995.720 842.310 998.810 ;
      LAYER met2 ;
        RECT 842.590 996.000 842.870 999.870 ;
      LAYER met2 ;
        RECT 843.150 995.720 844.610 998.810 ;
      LAYER met2 ;
        RECT 844.890 996.000 845.170 999.870 ;
      LAYER met2 ;
        RECT 845.450 995.720 846.450 998.810 ;
      LAYER met2 ;
        RECT 846.730 996.000 847.010 999.870 ;
      LAYER met2 ;
        RECT 847.290 995.720 848.750 998.810 ;
      LAYER met2 ;
        RECT 849.030 996.000 849.310 1000.000 ;
      LAYER met2 ;
        RECT 849.590 995.720 851.050 998.810 ;
      LAYER met2 ;
        RECT 851.330 996.000 851.610 1000.000 ;
      LAYER met2 ;
        RECT 851.890 995.720 852.890 998.810 ;
      LAYER met2 ;
        RECT 853.170 996.000 853.450 1000.000 ;
      LAYER met2 ;
        RECT 853.730 995.720 855.190 998.810 ;
      LAYER met2 ;
        RECT 855.470 996.000 855.750 1000.000 ;
      LAYER met2 ;
        RECT 856.030 995.720 857.490 998.810 ;
      LAYER met2 ;
        RECT 857.770 996.000 858.050 1000.000 ;
      LAYER met2 ;
        RECT 858.330 995.720 859.790 998.810 ;
      LAYER met2 ;
        RECT 860.070 996.000 860.350 1000.000 ;
      LAYER met2 ;
        RECT 860.630 995.720 861.630 998.810 ;
      LAYER met2 ;
        RECT 861.910 996.000 862.190 1000.000 ;
      LAYER met2 ;
        RECT 862.470 995.720 863.930 998.810 ;
      LAYER met2 ;
        RECT 864.210 996.000 864.490 1000.000 ;
      LAYER met2 ;
        RECT 864.770 995.720 866.230 998.810 ;
      LAYER met2 ;
        RECT 866.510 996.000 866.790 1000.000 ;
      LAYER met2 ;
        RECT 867.070 995.720 868.530 998.810 ;
      LAYER met2 ;
        RECT 868.810 996.000 869.090 1000.000 ;
      LAYER met2 ;
        RECT 869.370 995.720 870.370 998.810 ;
      LAYER met2 ;
        RECT 870.650 996.000 870.930 1000.000 ;
      LAYER met2 ;
        RECT 871.210 995.720 872.670 998.810 ;
      LAYER met2 ;
        RECT 872.950 996.000 873.230 1000.000 ;
      LAYER met2 ;
        RECT 873.510 995.720 874.970 998.810 ;
      LAYER met2 ;
        RECT 875.250 996.000 875.530 1000.000 ;
      LAYER met2 ;
        RECT 875.810 995.720 876.810 998.810 ;
      LAYER met2 ;
        RECT 877.090 996.000 877.370 1000.000 ;
      LAYER met2 ;
        RECT 877.650 995.720 879.110 998.810 ;
      LAYER met2 ;
        RECT 879.390 996.000 879.670 1000.000 ;
      LAYER met2 ;
        RECT 879.950 995.720 881.410 998.810 ;
      LAYER met2 ;
        RECT 881.690 996.000 881.970 1000.000 ;
      LAYER met2 ;
        RECT 882.250 995.720 883.710 998.810 ;
      LAYER met2 ;
        RECT 883.990 996.000 884.270 1000.000 ;
        RECT 884.740 999.870 886.110 1000.000 ;
      LAYER met2 ;
        RECT 884.550 995.720 885.550 998.810 ;
      LAYER met2 ;
        RECT 885.830 996.000 886.110 999.870 ;
      LAYER met2 ;
        RECT 886.390 995.720 887.850 998.810 ;
      LAYER met2 ;
        RECT 888.130 996.000 888.410 1000.000 ;
        RECT 890.260 999.870 890.710 1000.000 ;
      LAYER met2 ;
        RECT 888.690 995.720 890.150 998.810 ;
      LAYER met2 ;
        RECT 890.430 996.000 890.710 999.870 ;
      LAYER met2 ;
        RECT 890.990 995.720 892.450 998.810 ;
      LAYER met2 ;
        RECT 892.730 996.000 893.010 1000.000 ;
        RECT 893.480 999.870 894.850 1000.000 ;
      LAYER met2 ;
        RECT 893.290 995.720 894.290 998.810 ;
      LAYER met2 ;
        RECT 894.570 996.000 894.850 999.870 ;
      LAYER met2 ;
        RECT 895.130 995.720 896.590 998.810 ;
      LAYER met2 ;
        RECT 896.870 996.000 897.150 1000.000 ;
        RECT 897.620 999.870 899.450 1000.000 ;
      LAYER met2 ;
        RECT 897.430 995.720 898.890 998.810 ;
      LAYER met2 ;
        RECT 899.170 996.000 899.450 999.870 ;
      LAYER met2 ;
        RECT 899.730 995.720 900.730 998.810 ;
      LAYER met2 ;
        RECT 901.010 996.000 901.290 1000.000 ;
        RECT 901.760 999.870 903.590 1000.000 ;
      LAYER met2 ;
        RECT 901.570 995.720 903.030 998.810 ;
      LAYER met2 ;
        RECT 903.310 996.000 903.590 999.870 ;
      LAYER met2 ;
        RECT 903.870 995.720 905.330 998.810 ;
      LAYER met2 ;
        RECT 905.610 996.000 905.890 1000.000 ;
        RECT 906.360 999.870 908.190 1000.000 ;
      LAYER met2 ;
        RECT 906.170 995.720 907.630 998.810 ;
      LAYER met2 ;
        RECT 907.910 996.000 908.190 999.870 ;
      LAYER met2 ;
        RECT 908.470 995.720 909.470 998.810 ;
      LAYER met2 ;
        RECT 909.750 996.000 910.030 1000.000 ;
        RECT 910.960 999.870 912.330 1000.000 ;
      LAYER met2 ;
        RECT 910.310 995.720 911.770 998.810 ;
      LAYER met2 ;
        RECT 912.050 996.000 912.330 999.870 ;
      LAYER met2 ;
        RECT 912.610 995.720 914.070 998.810 ;
      LAYER met2 ;
        RECT 914.350 996.000 914.630 1000.000 ;
      LAYER met2 ;
        RECT 914.910 995.720 916.370 998.810 ;
      LAYER met2 ;
        RECT 916.650 996.000 916.930 1000.000 ;
      LAYER met2 ;
        RECT 917.210 995.720 918.210 998.810 ;
      LAYER met2 ;
        RECT 918.490 996.000 918.770 1000.000 ;
      LAYER met2 ;
        RECT 919.050 995.720 920.510 998.810 ;
      LAYER met2 ;
        RECT 920.790 996.000 921.070 1000.000 ;
      LAYER met2 ;
        RECT 921.350 995.720 922.810 998.810 ;
      LAYER met2 ;
        RECT 923.090 996.000 923.370 1000.000 ;
      LAYER met2 ;
        RECT 923.650 995.720 924.650 998.810 ;
      LAYER met2 ;
        RECT 924.930 996.000 925.210 1000.000 ;
      LAYER met2 ;
        RECT 925.490 995.720 926.950 998.810 ;
      LAYER met2 ;
        RECT 927.230 996.000 927.510 1000.000 ;
      LAYER met2 ;
        RECT 927.790 995.720 929.250 998.810 ;
      LAYER met2 ;
        RECT 929.530 996.000 929.810 1000.000 ;
      LAYER met2 ;
        RECT 930.090 995.720 931.550 998.810 ;
      LAYER met2 ;
        RECT 931.830 996.000 932.110 1000.000 ;
      LAYER met2 ;
        RECT 932.390 995.720 933.390 998.810 ;
      LAYER met2 ;
        RECT 933.670 996.000 933.950 1000.000 ;
      LAYER met2 ;
        RECT 934.230 995.720 935.690 998.810 ;
      LAYER met2 ;
        RECT 935.970 996.000 936.250 1000.000 ;
      LAYER met2 ;
        RECT 936.530 995.720 937.990 998.810 ;
      LAYER met2 ;
        RECT 938.270 996.000 938.550 1000.000 ;
      LAYER met2 ;
        RECT 938.830 995.720 940.290 998.810 ;
      LAYER met2 ;
        RECT 940.570 996.000 940.850 1000.000 ;
      LAYER met2 ;
        RECT 941.130 995.720 942.130 998.810 ;
      LAYER met2 ;
        RECT 942.410 996.000 942.690 1000.000 ;
      LAYER met2 ;
        RECT 942.970 995.720 944.430 998.810 ;
      LAYER met2 ;
        RECT 944.710 996.000 944.990 1000.000 ;
      LAYER met2 ;
        RECT 945.270 995.720 946.730 998.810 ;
      LAYER met2 ;
        RECT 947.010 996.000 947.290 1000.000 ;
      LAYER met2 ;
        RECT 947.570 995.720 948.570 998.810 ;
      LAYER met2 ;
        RECT 948.850 996.000 949.130 1000.000 ;
      LAYER met2 ;
        RECT 949.410 995.720 950.870 998.810 ;
      LAYER met2 ;
        RECT 951.150 996.000 951.430 1000.000 ;
      LAYER met2 ;
        RECT 951.710 995.720 953.170 998.810 ;
      LAYER met2 ;
        RECT 953.450 996.000 953.730 1000.000 ;
      LAYER met2 ;
        RECT 954.010 995.720 955.470 998.810 ;
      LAYER met2 ;
        RECT 955.750 996.000 956.030 1000.000 ;
      LAYER met2 ;
        RECT 956.310 995.720 957.310 998.810 ;
      LAYER met2 ;
        RECT 957.590 996.000 957.870 1000.000 ;
      LAYER met2 ;
        RECT 958.150 995.720 959.610 998.810 ;
      LAYER met2 ;
        RECT 959.890 996.000 960.170 1000.000 ;
      LAYER met2 ;
        RECT 960.450 995.720 961.910 998.810 ;
      LAYER met2 ;
        RECT 962.190 996.000 962.470 1000.000 ;
      LAYER met2 ;
        RECT 962.750 995.720 964.210 998.810 ;
      LAYER met2 ;
        RECT 964.490 996.000 964.770 1000.000 ;
      LAYER met2 ;
        RECT 965.050 995.720 966.050 998.810 ;
      LAYER met2 ;
        RECT 966.330 996.000 966.610 1000.000 ;
      LAYER met2 ;
        RECT 966.890 995.720 968.350 998.810 ;
      LAYER met2 ;
        RECT 968.630 996.000 968.910 1000.000 ;
      LAYER met2 ;
        RECT 969.190 995.720 970.650 998.810 ;
      LAYER met2 ;
        RECT 970.930 996.000 971.210 1000.000 ;
      LAYER met2 ;
        RECT 971.490 995.720 972.490 998.810 ;
      LAYER met2 ;
        RECT 972.770 996.000 973.050 1000.000 ;
      LAYER met2 ;
        RECT 973.330 995.720 974.790 998.810 ;
      LAYER met2 ;
        RECT 975.070 996.000 975.350 1000.000 ;
      LAYER met2 ;
        RECT 975.630 995.720 977.090 998.810 ;
      LAYER met2 ;
        RECT 977.370 996.000 977.650 1000.000 ;
      LAYER met2 ;
        RECT 977.930 995.720 979.390 998.810 ;
      LAYER met2 ;
        RECT 979.670 996.000 979.950 1000.000 ;
      LAYER met2 ;
        RECT 980.230 995.720 981.230 998.810 ;
      LAYER met2 ;
        RECT 981.510 996.000 981.790 1000.000 ;
      LAYER met2 ;
        RECT 982.070 995.720 983.530 998.810 ;
      LAYER met2 ;
        RECT 983.810 996.000 984.090 1000.000 ;
      LAYER met2 ;
        RECT 984.370 995.720 985.830 998.810 ;
      LAYER met2 ;
        RECT 986.110 996.000 986.390 1000.000 ;
      LAYER met2 ;
        RECT 986.670 995.720 988.130 998.810 ;
      LAYER met2 ;
        RECT 988.410 996.000 988.690 1000.000 ;
      LAYER met2 ;
        RECT 988.970 995.720 989.970 998.810 ;
      LAYER met2 ;
        RECT 990.250 996.000 990.530 1000.000 ;
      LAYER met2 ;
        RECT 990.810 995.720 992.270 998.810 ;
      LAYER met2 ;
        RECT 992.550 996.000 992.830 1000.000 ;
      LAYER met2 ;
        RECT 993.110 995.720 994.570 998.810 ;
      LAYER met2 ;
        RECT 994.850 996.000 995.130 1000.000 ;
      LAYER met2 ;
        RECT 995.410 995.720 996.410 998.810 ;
      LAYER met2 ;
        RECT 996.690 996.000 996.970 1000.000 ;
      LAYER met2 ;
        RECT 997.250 995.720 998.710 998.810 ;
      LAYER met2 ;
        RECT 998.990 996.000 999.270 1000.000 ;
      LAYER met2 ;
        RECT 999.550 995.720 1001.010 998.810 ;
      LAYER met2 ;
        RECT 1001.290 996.000 1001.570 1000.000 ;
      LAYER met2 ;
        RECT 1001.850 995.720 1003.310 998.810 ;
      LAYER met2 ;
        RECT 1003.590 996.000 1003.870 1000.000 ;
      LAYER met2 ;
        RECT 1004.150 995.720 1005.150 998.810 ;
      LAYER met2 ;
        RECT 1005.430 996.000 1005.710 1000.000 ;
      LAYER met2 ;
        RECT 1005.990 995.720 1007.450 998.810 ;
      LAYER met2 ;
        RECT 1007.730 996.000 1008.010 1000.000 ;
      LAYER met2 ;
        RECT 1008.290 995.720 1009.750 998.810 ;
      LAYER met2 ;
        RECT 1010.030 996.000 1010.310 1000.000 ;
      LAYER met2 ;
        RECT 1010.590 995.720 1011.590 998.810 ;
      LAYER met2 ;
        RECT 1011.870 996.000 1012.150 1000.000 ;
        RECT 1014.170 999.870 1014.600 1000.000 ;
      LAYER met2 ;
        RECT 1012.430 995.720 1013.890 998.810 ;
      LAYER met2 ;
        RECT 1014.170 996.000 1014.450 999.870 ;
      LAYER met2 ;
        RECT 1014.730 995.720 1016.190 998.810 ;
      LAYER met2 ;
        RECT 1016.470 996.000 1016.750 1000.000 ;
      LAYER met2 ;
        RECT 1017.030 995.720 1018.490 998.810 ;
      LAYER met2 ;
        RECT 1018.770 996.000 1019.050 1000.000 ;
      LAYER met2 ;
        RECT 1019.330 995.720 1020.330 998.810 ;
      LAYER met2 ;
        RECT 1020.610 996.000 1020.890 1000.000 ;
      LAYER met2 ;
        RECT 1021.170 995.720 1022.630 998.810 ;
      LAYER met2 ;
        RECT 1022.910 996.000 1023.190 1000.000 ;
      LAYER met2 ;
        RECT 1023.470 995.720 1024.930 998.810 ;
      LAYER met2 ;
        RECT 1025.210 996.000 1025.490 1000.000 ;
      LAYER met2 ;
        RECT 1025.770 995.720 1027.230 998.810 ;
      LAYER met2 ;
        RECT 1027.510 996.000 1027.790 1000.000 ;
      LAYER met2 ;
        RECT 1028.070 995.720 1029.070 998.810 ;
      LAYER met2 ;
        RECT 1029.350 996.000 1029.630 1000.000 ;
      LAYER met2 ;
        RECT 1029.910 995.720 1031.370 998.810 ;
      LAYER met2 ;
        RECT 1031.650 996.000 1031.930 1000.000 ;
      LAYER met2 ;
        RECT 1032.210 995.720 1033.670 998.810 ;
      LAYER met2 ;
        RECT 1033.950 996.000 1034.230 1000.000 ;
      LAYER met2 ;
        RECT 1034.510 995.720 1035.510 998.810 ;
      LAYER met2 ;
        RECT 1035.790 996.000 1036.070 1000.000 ;
      LAYER met2 ;
        RECT 1036.350 995.720 1037.810 998.810 ;
      LAYER met2 ;
        RECT 1038.090 996.000 1038.370 1000.000 ;
      LAYER met2 ;
        RECT 1038.650 995.720 1040.110 998.810 ;
      LAYER met2 ;
        RECT 1040.390 996.000 1040.670 1000.000 ;
      LAYER met2 ;
        RECT 1040.950 995.720 1042.410 998.810 ;
      LAYER met2 ;
        RECT 1042.690 996.000 1042.970 1000.000 ;
      LAYER met2 ;
        RECT 1043.250 995.720 1044.250 998.810 ;
      LAYER met2 ;
        RECT 1044.530 996.000 1044.810 1000.000 ;
      LAYER met2 ;
        RECT 1045.090 995.720 1046.550 998.810 ;
      LAYER met2 ;
        RECT 1046.830 996.000 1047.110 1000.000 ;
      LAYER met2 ;
        RECT 1047.390 995.720 1048.850 998.810 ;
      LAYER met2 ;
        RECT 1049.130 996.000 1049.410 1000.000 ;
        RECT 1049.880 999.870 1051.710 1000.000 ;
      LAYER met2 ;
        RECT 1049.690 995.720 1051.150 998.810 ;
      LAYER met2 ;
        RECT 1051.430 996.000 1051.710 999.870 ;
      LAYER met2 ;
        RECT 1051.990 995.720 1052.990 998.810 ;
      LAYER met2 ;
        RECT 1053.270 996.000 1053.550 1000.000 ;
        RECT 1055.570 999.870 1056.000 1000.000 ;
      LAYER met2 ;
        RECT 1053.830 995.720 1055.290 998.810 ;
      LAYER met2 ;
        RECT 1055.570 996.000 1055.850 999.870 ;
      LAYER met2 ;
        RECT 1056.130 995.720 1057.590 998.810 ;
      LAYER met2 ;
        RECT 1057.870 996.000 1058.150 1000.000 ;
        RECT 1058.620 999.870 1059.990 1000.000 ;
      LAYER met2 ;
        RECT 1058.430 995.720 1059.430 998.810 ;
      LAYER met2 ;
        RECT 1059.710 996.000 1059.990 999.870 ;
      LAYER met2 ;
        RECT 1060.270 995.720 1061.730 998.810 ;
      LAYER met2 ;
        RECT 1062.010 996.000 1062.290 1000.000 ;
        RECT 1062.760 999.870 1064.590 1000.000 ;
      LAYER met2 ;
        RECT 1062.570 995.720 1064.030 998.810 ;
      LAYER met2 ;
        RECT 1064.310 996.000 1064.590 999.870 ;
      LAYER met2 ;
        RECT 1064.870 995.720 1066.330 998.810 ;
      LAYER met2 ;
        RECT 1066.610 996.000 1066.890 1000.000 ;
        RECT 1067.360 999.870 1068.730 1000.000 ;
      LAYER met2 ;
        RECT 1067.170 995.720 1068.170 998.810 ;
      LAYER met2 ;
        RECT 1068.450 996.000 1068.730 999.870 ;
      LAYER met2 ;
        RECT 1069.010 995.720 1070.470 998.810 ;
      LAYER met2 ;
        RECT 1070.750 996.000 1071.030 1000.000 ;
        RECT 1071.960 999.870 1073.330 1000.000 ;
      LAYER met2 ;
        RECT 1071.310 995.720 1072.770 998.810 ;
      LAYER met2 ;
        RECT 1073.050 996.000 1073.330 999.870 ;
      LAYER met2 ;
        RECT 1073.610 995.720 1075.070 998.810 ;
      LAYER met2 ;
        RECT 1075.350 996.000 1075.630 1000.000 ;
        RECT 1076.560 999.870 1077.470 1000.000 ;
      LAYER met2 ;
        RECT 1075.910 995.720 1076.910 998.810 ;
      LAYER met2 ;
        RECT 1077.190 996.000 1077.470 999.870 ;
      LAYER met2 ;
        RECT 1077.750 995.720 1079.210 998.810 ;
      LAYER met2 ;
        RECT 1079.490 996.000 1079.770 1000.000 ;
        RECT 1080.240 999.870 1082.070 1000.000 ;
      LAYER met2 ;
        RECT 1080.050 995.720 1081.510 998.810 ;
      LAYER met2 ;
        RECT 1081.790 996.000 1082.070 999.870 ;
      LAYER met2 ;
        RECT 1082.350 995.720 1083.350 998.810 ;
      LAYER met2 ;
        RECT 1083.630 996.000 1083.910 1000.000 ;
        RECT 1084.380 999.870 1086.210 1000.000 ;
      LAYER met2 ;
        RECT 1084.190 995.720 1085.650 998.810 ;
      LAYER met2 ;
        RECT 1085.930 996.000 1086.210 999.870 ;
      LAYER met2 ;
        RECT 1086.490 995.720 1087.950 998.810 ;
      LAYER met2 ;
        RECT 1088.230 996.000 1088.510 1000.000 ;
        RECT 1090.360 999.870 1090.810 1000.000 ;
      LAYER met2 ;
        RECT 1088.790 995.720 1090.250 998.810 ;
      LAYER met2 ;
        RECT 1090.530 996.000 1090.810 999.870 ;
      LAYER met2 ;
        RECT 1091.090 995.720 1092.090 998.810 ;
      LAYER met2 ;
        RECT 1092.370 996.000 1092.650 1000.000 ;
        RECT 1093.120 999.870 1094.950 1000.000 ;
      LAYER met2 ;
        RECT 1092.930 995.720 1094.390 998.810 ;
      LAYER met2 ;
        RECT 1094.670 996.000 1094.950 999.870 ;
      LAYER met2 ;
        RECT 1095.230 995.720 1096.690 998.810 ;
      LAYER met2 ;
        RECT 1096.970 996.000 1097.250 1000.000 ;
        RECT 1097.720 999.870 1099.550 1000.000 ;
      LAYER met2 ;
        RECT 1097.530 995.720 1098.990 998.810 ;
      LAYER met2 ;
        RECT 1099.270 996.000 1099.550 999.870 ;
      LAYER met2 ;
        RECT 1099.830 995.720 1100.830 998.810 ;
      LAYER met2 ;
        RECT 1101.110 996.000 1101.390 1000.000 ;
        RECT 1101.860 999.870 1103.690 1000.000 ;
      LAYER met2 ;
        RECT 1101.670 995.720 1103.130 998.810 ;
      LAYER met2 ;
        RECT 1103.410 996.000 1103.690 999.870 ;
      LAYER met2 ;
        RECT 1103.970 995.720 1105.430 998.810 ;
      LAYER met2 ;
        RECT 1105.710 996.000 1105.990 1000.000 ;
        RECT 1106.460 999.870 1107.830 1000.000 ;
      LAYER met2 ;
        RECT 1106.270 995.720 1107.270 998.810 ;
      LAYER met2 ;
        RECT 1107.550 996.000 1107.830 999.870 ;
      LAYER met2 ;
        RECT 1108.110 995.720 1109.570 998.810 ;
      LAYER met2 ;
        RECT 1109.850 996.000 1110.130 1000.000 ;
        RECT 1111.060 999.870 1112.430 1000.000 ;
      LAYER met2 ;
        RECT 1110.410 995.720 1111.870 998.810 ;
      LAYER met2 ;
        RECT 1112.150 996.000 1112.430 999.870 ;
      LAYER met2 ;
        RECT 1112.710 995.720 1114.170 998.810 ;
      LAYER met2 ;
        RECT 1114.450 996.000 1114.730 1000.000 ;
        RECT 1115.200 999.870 1116.570 1000.000 ;
      LAYER met2 ;
        RECT 1115.010 995.720 1116.010 998.810 ;
      LAYER met2 ;
        RECT 1116.290 996.000 1116.570 999.870 ;
      LAYER met2 ;
        RECT 1116.850 995.720 1118.310 998.810 ;
      LAYER met2 ;
        RECT 1118.590 996.000 1118.870 1000.000 ;
        RECT 1119.340 999.870 1121.170 1000.000 ;
      LAYER met2 ;
        RECT 1119.150 995.720 1120.610 998.810 ;
      LAYER met2 ;
        RECT 1120.890 996.000 1121.170 999.870 ;
      LAYER met2 ;
        RECT 1121.450 995.720 1122.910 998.810 ;
      LAYER met2 ;
        RECT 1123.190 996.000 1123.470 1000.000 ;
      LAYER met2 ;
        RECT 1123.750 995.720 1124.750 998.810 ;
      LAYER met2 ;
        RECT 1125.030 996.000 1125.310 1000.000 ;
        RECT 1125.780 999.870 1127.610 1000.000 ;
      LAYER met2 ;
        RECT 1125.590 995.720 1127.050 998.810 ;
      LAYER met2 ;
        RECT 1127.330 996.000 1127.610 999.870 ;
      LAYER met2 ;
        RECT 1127.890 995.720 1129.350 998.810 ;
      LAYER met2 ;
        RECT 1129.630 996.000 1129.910 1000.000 ;
        RECT 1131.470 999.870 1131.900 1000.000 ;
      LAYER met2 ;
        RECT 1130.190 995.720 1131.190 998.810 ;
      LAYER met2 ;
        RECT 1131.470 996.000 1131.750 999.870 ;
      LAYER met2 ;
        RECT 1132.030 995.720 1133.490 998.810 ;
      LAYER met2 ;
        RECT 1133.770 996.000 1134.050 1000.000 ;
        RECT 1134.520 999.870 1136.350 1000.000 ;
      LAYER met2 ;
        RECT 1134.330 995.720 1135.790 998.810 ;
      LAYER met2 ;
        RECT 1136.070 996.000 1136.350 999.870 ;
      LAYER met2 ;
        RECT 1136.630 995.720 1138.090 998.810 ;
      LAYER met2 ;
        RECT 1138.370 996.000 1138.650 1000.000 ;
        RECT 1139.120 999.870 1140.490 1000.000 ;
      LAYER met2 ;
        RECT 1138.930 995.720 1139.930 998.810 ;
      LAYER met2 ;
        RECT 1140.210 996.000 1140.490 999.870 ;
      LAYER met2 ;
        RECT 1140.770 995.720 1142.230 998.810 ;
      LAYER met2 ;
        RECT 1142.510 996.000 1142.790 1000.000 ;
        RECT 1143.260 999.870 1145.090 1000.000 ;
      LAYER met2 ;
        RECT 1143.070 995.720 1144.530 998.810 ;
      LAYER met2 ;
        RECT 1144.810 996.000 1145.090 999.870 ;
      LAYER met2 ;
        RECT 1145.370 995.720 1146.830 998.810 ;
      LAYER met2 ;
        RECT 1147.110 996.000 1147.390 1000.000 ;
        RECT 1147.860 999.870 1149.230 1000.000 ;
      LAYER met2 ;
        RECT 1147.670 995.720 1148.670 998.810 ;
      LAYER met2 ;
        RECT 1148.950 996.000 1149.230 999.870 ;
      LAYER met2 ;
        RECT 1149.510 995.720 1150.970 998.810 ;
      LAYER met2 ;
        RECT 1151.250 996.000 1151.530 1000.000 ;
        RECT 1152.920 999.870 1153.830 1000.000 ;
      LAYER met2 ;
        RECT 1151.810 995.720 1153.270 998.810 ;
      LAYER met2 ;
        RECT 1153.550 996.000 1153.830 999.870 ;
      LAYER met2 ;
        RECT 1154.110 995.720 1155.110 998.810 ;
      LAYER met2 ;
        RECT 1155.390 996.000 1155.670 1000.000 ;
        RECT 1156.140 999.870 1157.970 1000.000 ;
      LAYER met2 ;
        RECT 1155.950 995.720 1157.410 998.810 ;
      LAYER met2 ;
        RECT 1157.690 996.000 1157.970 999.870 ;
      LAYER met2 ;
        RECT 1158.250 995.720 1159.710 998.810 ;
      LAYER met2 ;
        RECT 1159.990 996.000 1160.270 1000.000 ;
        RECT 1160.740 999.870 1162.570 1000.000 ;
      LAYER met2 ;
        RECT 1160.550 995.720 1162.010 998.810 ;
      LAYER met2 ;
        RECT 1162.290 996.000 1162.570 999.870 ;
      LAYER met2 ;
        RECT 1162.850 995.720 1163.850 998.810 ;
      LAYER met2 ;
        RECT 1164.130 996.000 1164.410 1000.000 ;
        RECT 1166.260 999.870 1166.710 1000.000 ;
        RECT 1167.180 999.870 1169.010 1000.000 ;
      LAYER met2 ;
        RECT 1164.690 995.720 1166.150 998.810 ;
      LAYER met2 ;
        RECT 1166.430 996.000 1166.710 999.870 ;
      LAYER met2 ;
        RECT 1166.990 995.720 1168.450 998.810 ;
      LAYER met2 ;
        RECT 1168.730 996.000 1169.010 999.870 ;
      LAYER met2 ;
        RECT 1169.290 995.720 1170.750 998.810 ;
      LAYER met2 ;
        RECT 1171.030 996.000 1171.310 1000.000 ;
      LAYER met2 ;
        RECT 1171.590 995.720 1172.590 998.810 ;
      LAYER met2 ;
        RECT 1172.870 996.000 1173.150 1000.000 ;
      LAYER met2 ;
        RECT 1173.430 995.720 1174.890 998.810 ;
      LAYER met2 ;
        RECT 1175.170 996.000 1175.450 1000.000 ;
      LAYER met2 ;
        RECT 1175.730 995.720 1177.190 998.810 ;
      LAYER met2 ;
        RECT 1177.470 996.000 1177.750 1000.000 ;
      LAYER met2 ;
        RECT 1178.030 995.720 1179.030 998.810 ;
      LAYER met2 ;
        RECT 1179.310 996.000 1179.590 1000.000 ;
        RECT 1181.610 999.870 1182.040 1000.000 ;
        RECT 1182.360 1000.010 1182.500 1024.350 ;
        RECT 1186.500 1000.010 1186.640 1693.550 ;
        RECT 1187.880 1684.350 1188.020 1700.000 ;
        RECT 1197.020 1689.130 1197.280 1689.450 ;
        RECT 1197.080 1686.730 1197.220 1689.130 ;
        RECT 1188.280 1686.410 1188.540 1686.730 ;
        RECT 1197.020 1686.410 1197.280 1686.730 ;
        RECT 1187.360 1684.030 1187.620 1684.350 ;
        RECT 1187.820 1684.030 1188.080 1684.350 ;
        RECT 1187.420 1024.750 1187.560 1684.030 ;
        RECT 1187.360 1024.430 1187.620 1024.750 ;
        RECT 1188.340 1000.010 1188.480 1686.410 ;
        RECT 1197.020 1684.030 1197.280 1684.350 ;
        RECT 1200.240 1684.030 1200.500 1684.350 ;
        RECT 1188.740 1024.430 1189.000 1024.750 ;
        RECT 1182.360 1000.000 1184.040 1000.010 ;
        RECT 1186.340 1000.000 1186.640 1000.010 ;
        RECT 1188.180 1000.000 1188.480 1000.010 ;
        RECT 1182.360 999.870 1184.190 1000.000 ;
      LAYER met2 ;
        RECT 1179.870 995.720 1181.330 998.810 ;
      LAYER met2 ;
        RECT 1181.610 996.000 1181.890 999.870 ;
      LAYER met2 ;
        RECT 1182.170 995.720 1183.630 998.810 ;
      LAYER met2 ;
        RECT 1183.910 996.000 1184.190 999.870 ;
        RECT 1186.210 999.870 1186.640 1000.000 ;
        RECT 1188.050 999.870 1188.480 1000.000 ;
        RECT 1188.800 1000.010 1188.940 1024.430 ;
        RECT 1193.800 1017.290 1194.060 1017.610 ;
        RECT 1191.040 1013.210 1191.300 1013.530 ;
        RECT 1191.100 1000.010 1191.240 1013.210 ;
        RECT 1188.800 1000.000 1190.480 1000.010 ;
        RECT 1191.100 1000.000 1192.780 1000.010 ;
        RECT 1188.800 999.870 1190.630 1000.000 ;
        RECT 1191.100 999.870 1192.930 1000.000 ;
      LAYER met2 ;
        RECT 1184.470 995.720 1185.930 998.810 ;
      LAYER met2 ;
        RECT 1186.210 996.000 1186.490 999.870 ;
      LAYER met2 ;
        RECT 1186.770 995.720 1187.770 998.810 ;
      LAYER met2 ;
        RECT 1188.050 996.000 1188.330 999.870 ;
      LAYER met2 ;
        RECT 1188.610 995.720 1190.070 998.810 ;
      LAYER met2 ;
        RECT 1190.350 996.000 1190.630 999.870 ;
      LAYER met2 ;
        RECT 1190.910 995.720 1192.370 998.810 ;
      LAYER met2 ;
        RECT 1192.650 996.000 1192.930 999.870 ;
        RECT 1193.860 999.590 1194.000 1017.290 ;
        RECT 1197.080 1013.190 1197.220 1684.030 ;
        RECT 1198.400 1013.890 1198.660 1014.210 ;
        RECT 1196.560 1012.870 1196.820 1013.190 ;
        RECT 1197.020 1012.870 1197.280 1013.190 ;
        RECT 1196.100 1010.150 1196.360 1010.470 ;
        RECT 1196.160 1000.010 1196.300 1010.150 ;
        RECT 1196.620 1009.450 1196.760 1012.870 ;
        RECT 1196.560 1009.130 1196.820 1009.450 ;
        RECT 1198.460 1000.010 1198.600 1013.890 ;
        RECT 1200.300 1010.470 1200.440 1684.030 ;
        RECT 1200.760 1014.210 1200.900 1700.270 ;
        RECT 1201.570 1700.000 1201.850 1700.270 ;
        RECT 1215.370 1700.000 1215.650 1704.000 ;
        RECT 1230.090 1700.000 1230.370 1704.000 ;
        RECT 1243.890 1700.000 1244.170 1704.000 ;
        RECT 1258.610 1700.000 1258.890 1704.000 ;
        RECT 1272.410 1700.000 1272.690 1704.000 ;
        RECT 1287.130 1700.000 1287.410 1704.000 ;
        RECT 1300.930 1700.000 1301.210 1704.000 ;
        RECT 1315.650 1700.000 1315.930 1704.000 ;
        RECT 1329.450 1700.000 1329.730 1704.000 ;
        RECT 1203.920 1688.790 1204.180 1689.110 ;
        RECT 1210.820 1688.790 1211.080 1689.110 ;
        RECT 1200.700 1013.890 1200.960 1014.210 ;
        RECT 1202.540 1013.890 1202.800 1014.210 ;
        RECT 1200.240 1010.150 1200.500 1010.470 ;
        RECT 1202.600 1000.010 1202.740 1013.890 ;
        RECT 1203.980 1013.530 1204.120 1688.790 ;
        RECT 1204.840 1017.290 1205.100 1017.610 ;
        RECT 1203.920 1013.210 1204.180 1013.530 ;
        RECT 1204.900 1000.010 1205.040 1017.290 ;
        RECT 1210.880 1014.210 1211.020 1688.790 ;
        RECT 1214.040 1686.070 1214.300 1686.390 ;
        RECT 1214.100 1014.210 1214.240 1686.070 ;
        RECT 1215.480 1684.350 1215.620 1700.000 ;
        RECT 1224.160 1689.810 1224.420 1690.130 ;
        RECT 1215.420 1684.030 1215.680 1684.350 ;
        RECT 1224.220 1642.530 1224.360 1689.810 ;
        RECT 1230.200 1689.110 1230.340 1700.000 ;
        RECT 1242.560 1689.470 1242.820 1689.790 ;
        RECT 1230.140 1688.790 1230.400 1689.110 ;
        RECT 1231.520 1686.410 1231.780 1686.730 ;
        RECT 1224.160 1642.210 1224.420 1642.530 ;
        RECT 1223.700 1021.030 1223.960 1021.350 ;
        RECT 1215.880 1016.950 1216.140 1017.270 ;
        RECT 1210.820 1013.890 1211.080 1014.210 ;
        RECT 1211.280 1013.890 1211.540 1014.210 ;
        RECT 1214.040 1013.890 1214.300 1014.210 ;
        RECT 1207.600 1012.530 1207.860 1012.850 ;
        RECT 1205.300 1012.190 1205.560 1012.510 ;
        RECT 1194.620 1000.000 1196.300 1000.010 ;
        RECT 1196.920 1000.000 1198.600 1000.010 ;
        RECT 1201.520 1000.000 1202.740 1000.010 ;
        RECT 1203.360 1000.000 1205.040 1000.010 ;
        RECT 1194.490 999.870 1196.300 1000.000 ;
        RECT 1196.790 999.870 1198.600 1000.000 ;
        RECT 1193.800 999.270 1194.060 999.590 ;
      LAYER met2 ;
        RECT 1193.210 995.720 1194.210 998.810 ;
      LAYER met2 ;
        RECT 1194.490 996.000 1194.770 999.870 ;
      LAYER met2 ;
        RECT 1195.050 995.720 1196.510 998.810 ;
      LAYER met2 ;
        RECT 1196.790 996.000 1197.070 999.870 ;
        RECT 1197.480 999.330 1197.740 999.590 ;
        RECT 1199.090 999.330 1199.370 1000.000 ;
        RECT 1197.480 999.270 1199.370 999.330 ;
        RECT 1197.540 999.190 1199.370 999.270 ;
      LAYER met2 ;
        RECT 1197.350 995.720 1198.810 998.810 ;
      LAYER met2 ;
        RECT 1199.090 996.000 1199.370 999.190 ;
        RECT 1201.390 999.870 1202.740 1000.000 ;
        RECT 1203.230 999.870 1205.040 1000.000 ;
        RECT 1205.360 1000.010 1205.500 1012.190 ;
        RECT 1207.660 1000.010 1207.800 1012.530 ;
        RECT 1211.340 1000.010 1211.480 1013.890 ;
        RECT 1211.740 1013.210 1212.000 1013.530 ;
        RECT 1205.360 1000.000 1205.660 1000.010 ;
        RECT 1207.660 1000.000 1207.960 1000.010 ;
        RECT 1210.260 1000.000 1211.480 1000.010 ;
        RECT 1205.360 999.870 1205.810 1000.000 ;
        RECT 1207.660 999.870 1208.110 1000.000 ;
      LAYER met2 ;
        RECT 1199.650 995.720 1201.110 998.810 ;
      LAYER met2 ;
        RECT 1201.390 996.000 1201.670 999.870 ;
      LAYER met2 ;
        RECT 1201.950 995.720 1202.950 998.810 ;
      LAYER met2 ;
        RECT 1203.230 996.000 1203.510 999.870 ;
      LAYER met2 ;
        RECT 1203.790 995.720 1205.250 998.810 ;
      LAYER met2 ;
        RECT 1205.530 996.000 1205.810 999.870 ;
      LAYER met2 ;
        RECT 1206.090 995.720 1207.550 998.810 ;
      LAYER met2 ;
        RECT 1207.830 996.000 1208.110 999.870 ;
        RECT 1210.130 999.870 1211.480 1000.000 ;
        RECT 1211.800 1000.010 1211.940 1013.210 ;
        RECT 1215.420 1009.470 1215.680 1009.790 ;
        RECT 1215.480 1000.010 1215.620 1009.470 ;
        RECT 1211.800 1000.000 1212.100 1000.010 ;
        RECT 1214.400 1000.000 1215.620 1000.010 ;
        RECT 1211.800 999.870 1212.250 1000.000 ;
      LAYER met2 ;
        RECT 1208.390 995.720 1209.850 998.810 ;
      LAYER met2 ;
        RECT 1210.130 996.000 1210.410 999.870 ;
      LAYER met2 ;
        RECT 1210.690 995.720 1211.690 998.810 ;
      LAYER met2 ;
        RECT 1211.970 996.000 1212.250 999.870 ;
        RECT 1214.270 999.870 1215.620 1000.000 ;
        RECT 1215.940 1000.010 1216.080 1016.950 ;
        RECT 1219.100 1012.870 1219.360 1013.190 ;
        RECT 1218.640 1012.190 1218.900 1012.510 ;
        RECT 1218.700 1000.010 1218.840 1012.190 ;
        RECT 1215.940 1000.000 1216.700 1000.010 ;
        RECT 1218.540 1000.000 1218.840 1000.010 ;
        RECT 1215.940 999.870 1216.850 1000.000 ;
      LAYER met2 ;
        RECT 1212.530 995.720 1213.990 998.810 ;
      LAYER met2 ;
        RECT 1214.270 996.000 1214.550 999.870 ;
      LAYER met2 ;
        RECT 1214.830 995.720 1216.290 998.810 ;
      LAYER met2 ;
        RECT 1216.570 996.000 1216.850 999.870 ;
        RECT 1218.410 999.870 1218.840 1000.000 ;
        RECT 1219.160 1000.010 1219.300 1012.870 ;
        RECT 1223.240 1008.110 1223.500 1008.430 ;
        RECT 1223.300 1000.010 1223.440 1008.110 ;
        RECT 1219.160 1000.000 1220.840 1000.010 ;
        RECT 1223.140 1000.000 1223.440 1000.010 ;
        RECT 1219.160 999.870 1220.990 1000.000 ;
      LAYER met2 ;
        RECT 1217.130 995.720 1218.130 998.810 ;
      LAYER met2 ;
        RECT 1218.410 996.000 1218.690 999.870 ;
      LAYER met2 ;
        RECT 1218.970 995.720 1220.430 998.810 ;
      LAYER met2 ;
        RECT 1220.710 996.000 1220.990 999.870 ;
        RECT 1223.010 999.870 1223.440 1000.000 ;
        RECT 1223.760 1000.010 1223.900 1021.030 ;
        RECT 1228.300 1020.690 1228.560 1021.010 ;
        RECT 1226.000 1011.510 1226.260 1011.830 ;
        RECT 1226.060 1000.010 1226.200 1011.510 ;
        RECT 1228.360 1000.010 1228.500 1020.690 ;
        RECT 1231.580 1010.130 1231.720 1686.410 ;
        RECT 1238.420 1684.030 1238.680 1684.350 ;
        RECT 1237.500 1012.530 1237.760 1012.850 ;
        RECT 1232.440 1011.850 1232.700 1012.170 ;
        RECT 1231.520 1009.810 1231.780 1010.130 ;
        RECT 1230.140 1008.790 1230.400 1009.110 ;
        RECT 1230.200 1000.010 1230.340 1008.790 ;
        RECT 1232.500 1000.010 1232.640 1011.850 ;
        RECT 1237.560 1000.010 1237.700 1012.530 ;
        RECT 1237.960 1011.510 1238.220 1011.830 ;
        RECT 1223.760 1000.000 1225.440 1000.010 ;
        RECT 1226.060 1000.000 1227.280 1000.010 ;
        RECT 1228.360 1000.000 1229.580 1000.010 ;
        RECT 1230.200 1000.000 1231.880 1000.010 ;
        RECT 1232.500 1000.000 1234.180 1000.010 ;
        RECT 1236.020 1000.000 1237.700 1000.010 ;
        RECT 1223.760 999.870 1225.590 1000.000 ;
        RECT 1226.060 999.870 1227.430 1000.000 ;
        RECT 1228.360 999.870 1229.730 1000.000 ;
        RECT 1230.200 999.870 1232.030 1000.000 ;
        RECT 1232.500 999.870 1234.330 1000.000 ;
      LAYER met2 ;
        RECT 1221.270 995.720 1222.730 998.810 ;
      LAYER met2 ;
        RECT 1223.010 996.000 1223.290 999.870 ;
      LAYER met2 ;
        RECT 1223.570 995.720 1225.030 998.810 ;
      LAYER met2 ;
        RECT 1225.310 996.000 1225.590 999.870 ;
      LAYER met2 ;
        RECT 1225.870 995.720 1226.870 998.810 ;
      LAYER met2 ;
        RECT 1227.150 996.000 1227.430 999.870 ;
      LAYER met2 ;
        RECT 1227.710 995.720 1229.170 998.810 ;
      LAYER met2 ;
        RECT 1229.450 996.000 1229.730 999.870 ;
      LAYER met2 ;
        RECT 1230.010 995.720 1231.470 998.810 ;
      LAYER met2 ;
        RECT 1231.750 996.000 1232.030 999.870 ;
      LAYER met2 ;
        RECT 1232.310 995.720 1233.770 998.810 ;
      LAYER met2 ;
        RECT 1234.050 996.000 1234.330 999.870 ;
        RECT 1235.890 999.870 1237.700 1000.000 ;
        RECT 1238.020 1000.010 1238.160 1011.510 ;
        RECT 1238.480 1009.790 1238.620 1684.030 ;
        RECT 1238.420 1009.470 1238.680 1009.790 ;
        RECT 1238.880 1009.130 1239.140 1009.450 ;
        RECT 1238.940 1000.010 1239.080 1009.130 ;
        RECT 1242.620 1000.010 1242.760 1689.470 ;
        RECT 1244.000 1684.350 1244.140 1700.000 ;
        RECT 1254.980 1689.810 1255.240 1690.130 ;
        RECT 1245.320 1688.790 1245.580 1689.110 ;
        RECT 1245.380 1686.390 1245.520 1688.790 ;
        RECT 1245.320 1686.070 1245.580 1686.390 ;
        RECT 1243.940 1684.030 1244.200 1684.350 ;
        RECT 1243.480 1642.210 1243.740 1642.530 ;
        RECT 1243.540 1001.290 1243.680 1642.210 ;
        RECT 1252.680 1020.690 1252.940 1021.010 ;
        RECT 1244.860 1012.870 1245.120 1013.190 ;
        RECT 1243.480 1000.970 1243.740 1001.290 ;
        RECT 1244.920 1000.010 1245.060 1012.870 ;
        RECT 1250.380 1008.450 1250.640 1008.770 ;
        RECT 1246.930 1000.970 1247.190 1001.290 ;
        RECT 1238.020 1000.000 1238.320 1000.010 ;
        RECT 1238.940 1000.000 1240.620 1000.010 ;
        RECT 1242.460 1000.000 1242.760 1000.010 ;
        RECT 1244.760 1000.000 1245.060 1000.010 ;
        RECT 1246.990 1000.000 1247.130 1000.970 ;
        RECT 1250.440 1000.010 1250.580 1008.450 ;
        RECT 1252.740 1000.010 1252.880 1020.690 ;
        RECT 1254.520 1013.210 1254.780 1013.530 ;
        RECT 1254.580 1000.010 1254.720 1013.210 ;
        RECT 1255.040 1008.770 1255.180 1689.810 ;
        RECT 1258.720 1686.390 1258.860 1700.000 ;
        RECT 1268.780 1689.470 1269.040 1689.790 ;
        RECT 1258.660 1686.070 1258.920 1686.390 ;
        RECT 1259.580 1020.350 1259.840 1020.670 ;
        RECT 1267.860 1020.350 1268.120 1020.670 ;
        RECT 1257.280 1013.890 1257.540 1014.210 ;
        RECT 1254.980 1008.450 1255.240 1008.770 ;
        RECT 1257.340 1000.010 1257.480 1013.890 ;
        RECT 1259.120 1010.150 1259.380 1010.470 ;
        RECT 1259.180 1000.010 1259.320 1010.150 ;
        RECT 1249.360 1000.000 1250.580 1000.010 ;
        RECT 1251.200 1000.000 1252.880 1000.010 ;
        RECT 1253.500 1000.000 1254.720 1000.010 ;
        RECT 1255.800 1000.000 1257.480 1000.010 ;
        RECT 1258.100 1000.000 1259.320 1000.010 ;
        RECT 1238.020 999.870 1238.470 1000.000 ;
        RECT 1238.940 999.870 1240.770 1000.000 ;
      LAYER met2 ;
        RECT 1234.610 995.720 1235.610 998.810 ;
      LAYER met2 ;
        RECT 1235.890 996.000 1236.170 999.870 ;
      LAYER met2 ;
        RECT 1236.450 995.720 1237.910 998.810 ;
      LAYER met2 ;
        RECT 1238.190 996.000 1238.470 999.870 ;
      LAYER met2 ;
        RECT 1238.750 995.720 1240.210 998.810 ;
      LAYER met2 ;
        RECT 1240.490 996.000 1240.770 999.870 ;
        RECT 1242.330 999.870 1242.760 1000.000 ;
        RECT 1244.630 999.870 1245.060 1000.000 ;
      LAYER met2 ;
        RECT 1241.050 995.720 1242.050 998.810 ;
      LAYER met2 ;
        RECT 1242.330 996.000 1242.610 999.870 ;
      LAYER met2 ;
        RECT 1242.890 995.720 1244.350 998.810 ;
      LAYER met2 ;
        RECT 1244.630 996.000 1244.910 999.870 ;
      LAYER met2 ;
        RECT 1245.190 995.720 1246.650 998.810 ;
      LAYER met2 ;
        RECT 1246.930 996.000 1247.210 1000.000 ;
        RECT 1249.230 999.870 1250.580 1000.000 ;
        RECT 1251.070 999.870 1252.880 1000.000 ;
        RECT 1253.370 999.870 1254.720 1000.000 ;
        RECT 1255.670 999.870 1257.480 1000.000 ;
        RECT 1257.970 999.870 1259.320 1000.000 ;
        RECT 1259.640 1000.010 1259.780 1020.350 ;
        RECT 1263.260 1012.365 1263.520 1012.510 ;
        RECT 1263.250 1011.995 1263.530 1012.365 ;
        RECT 1267.400 1011.685 1267.660 1011.830 ;
        RECT 1267.390 1011.315 1267.670 1011.685 ;
        RECT 1265.560 1009.810 1265.820 1010.130 ;
        RECT 1263.720 1007.090 1263.980 1007.410 ;
        RECT 1263.780 1000.010 1263.920 1007.090 ;
        RECT 1265.620 1000.010 1265.760 1009.810 ;
        RECT 1267.920 1000.010 1268.060 1020.350 ;
        RECT 1268.840 1010.890 1268.980 1689.470 ;
        RECT 1272.520 1684.350 1272.660 1700.000 ;
        RECT 1287.240 1689.110 1287.380 1700.000 ;
        RECT 1289.940 1693.890 1290.200 1694.210 ;
        RECT 1287.180 1688.790 1287.440 1689.110 ;
        RECT 1277.980 1688.110 1278.240 1688.430 ;
        RECT 1272.460 1684.030 1272.720 1684.350 ;
        RECT 1278.040 1618.130 1278.180 1688.110 ;
        RECT 1278.040 1617.990 1279.100 1618.130 ;
        RECT 1278.960 1594.250 1279.100 1617.990 ;
        RECT 1278.900 1593.930 1279.160 1594.250 ;
        RECT 1279.360 1593.930 1279.620 1594.250 ;
        RECT 1279.420 1546.165 1279.560 1593.930 ;
        RECT 1290.000 1593.910 1290.140 1693.890 ;
        RECT 1301.040 1690.130 1301.180 1700.000 ;
        RECT 1310.640 1692.870 1310.900 1693.190 ;
        RECT 1300.980 1689.810 1301.240 1690.130 ;
        RECT 1293.620 1688.450 1293.880 1688.770 ;
        RECT 1292.240 1684.030 1292.500 1684.350 ;
        RECT 1292.300 1683.670 1292.440 1684.030 ;
        RECT 1290.860 1683.350 1291.120 1683.670 ;
        RECT 1292.240 1683.350 1292.500 1683.670 ;
        RECT 1290.920 1635.730 1291.060 1683.350 ;
        RECT 1290.860 1635.410 1291.120 1635.730 ;
        RECT 1291.780 1635.410 1292.040 1635.730 ;
        RECT 1291.840 1635.245 1291.980 1635.410 ;
        RECT 1290.850 1634.875 1291.130 1635.245 ;
        RECT 1291.770 1634.875 1292.050 1635.245 ;
        RECT 1288.560 1593.590 1288.820 1593.910 ;
        RECT 1289.940 1593.590 1290.200 1593.910 ;
        RECT 1277.970 1545.795 1278.250 1546.165 ;
        RECT 1279.350 1545.795 1279.630 1546.165 ;
        RECT 1288.620 1545.970 1288.760 1593.590 ;
        RECT 1290.920 1587.450 1291.060 1634.875 ;
        RECT 1290.860 1587.130 1291.120 1587.450 ;
        RECT 1293.160 1587.130 1293.420 1587.450 ;
        RECT 1293.220 1546.165 1293.360 1587.130 ;
        RECT 1278.040 1497.350 1278.180 1545.795 ;
        RECT 1288.560 1545.650 1288.820 1545.970 ;
        RECT 1289.020 1545.650 1289.280 1545.970 ;
        RECT 1291.770 1545.795 1292.050 1546.165 ;
        RECT 1293.150 1545.795 1293.430 1546.165 ;
        RECT 1289.080 1510.690 1289.220 1545.650 ;
        RECT 1289.080 1510.550 1289.680 1510.690 ;
        RECT 1289.540 1497.350 1289.680 1510.550 ;
        RECT 1291.840 1497.350 1291.980 1545.795 ;
        RECT 1277.520 1497.030 1277.780 1497.350 ;
        RECT 1277.980 1497.030 1278.240 1497.350 ;
        RECT 1288.560 1497.030 1288.820 1497.350 ;
        RECT 1289.480 1497.030 1289.740 1497.350 ;
        RECT 1291.320 1497.030 1291.580 1497.350 ;
        RECT 1291.780 1497.030 1292.040 1497.350 ;
        RECT 1277.580 1449.750 1277.720 1497.030 ;
        RECT 1277.520 1449.430 1277.780 1449.750 ;
        RECT 1288.620 1449.410 1288.760 1497.030 ;
        RECT 1291.380 1449.750 1291.520 1497.030 ;
        RECT 1291.320 1449.430 1291.580 1449.750 ;
        RECT 1277.980 1449.090 1278.240 1449.410 ;
        RECT 1288.560 1449.090 1288.820 1449.410 ;
        RECT 1289.020 1449.090 1289.280 1449.410 ;
        RECT 1291.780 1449.090 1292.040 1449.410 ;
        RECT 1278.040 1345.450 1278.180 1449.090 ;
        RECT 1289.080 1414.730 1289.220 1449.090 ;
        RECT 1289.020 1414.410 1289.280 1414.730 ;
        RECT 1289.940 1414.410 1290.200 1414.730 ;
        RECT 1278.040 1345.310 1278.640 1345.450 ;
        RECT 1278.500 1304.570 1278.640 1345.310 ;
        RECT 1278.440 1304.250 1278.700 1304.570 ;
        RECT 1278.440 1303.570 1278.700 1303.890 ;
        RECT 1278.500 1255.010 1278.640 1303.570 ;
        RECT 1277.120 1254.870 1278.640 1255.010 ;
        RECT 1277.120 1183.530 1277.260 1254.870 ;
        RECT 1290.000 1207.525 1290.140 1414.410 ;
        RECT 1291.840 1386.930 1291.980 1449.090 ;
        RECT 1291.380 1386.790 1291.980 1386.930 ;
        RECT 1291.380 1380.050 1291.520 1386.790 ;
        RECT 1291.320 1379.730 1291.580 1380.050 ;
        RECT 1291.780 1379.730 1292.040 1380.050 ;
        RECT 1291.840 1290.370 1291.980 1379.730 ;
        RECT 1291.840 1290.230 1292.440 1290.370 ;
        RECT 1292.300 1245.750 1292.440 1290.230 ;
        RECT 1292.240 1245.430 1292.500 1245.750 ;
        RECT 1292.240 1244.750 1292.500 1245.070 ;
        RECT 1289.930 1207.155 1290.210 1207.525 ;
        RECT 1290.850 1207.155 1291.130 1207.525 ;
        RECT 1277.060 1183.210 1277.320 1183.530 ;
        RECT 1277.980 1183.210 1278.240 1183.530 ;
        RECT 1278.040 1111.110 1278.180 1183.210 ;
        RECT 1290.920 1159.390 1291.060 1207.155 ;
        RECT 1292.300 1200.870 1292.440 1244.750 ;
        RECT 1291.320 1200.550 1291.580 1200.870 ;
        RECT 1292.240 1200.550 1292.500 1200.870 ;
        RECT 1291.380 1193.730 1291.520 1200.550 ;
        RECT 1291.320 1193.410 1291.580 1193.730 ;
        RECT 1292.240 1193.410 1292.500 1193.730 ;
        RECT 1289.940 1159.070 1290.200 1159.390 ;
        RECT 1290.860 1159.070 1291.120 1159.390 ;
        RECT 1290.000 1124.450 1290.140 1159.070 ;
        RECT 1292.300 1145.530 1292.440 1193.410 ;
        RECT 1292.300 1145.390 1292.900 1145.530 ;
        RECT 1289.540 1124.310 1290.140 1124.450 ;
        RECT 1277.980 1110.790 1278.240 1111.110 ;
        RECT 1278.440 1110.790 1278.700 1111.110 ;
        RECT 1289.540 1110.850 1289.680 1124.310 ;
        RECT 1278.500 1062.830 1278.640 1110.790 ;
        RECT 1289.540 1110.710 1290.140 1110.850 ;
        RECT 1290.000 1062.830 1290.140 1110.710 ;
        RECT 1292.760 1077.110 1292.900 1145.390 ;
        RECT 1292.700 1076.790 1292.960 1077.110 ;
        RECT 1292.240 1076.110 1292.500 1076.430 ;
        RECT 1277.980 1062.510 1278.240 1062.830 ;
        RECT 1278.440 1062.510 1278.700 1062.830 ;
        RECT 1289.020 1062.510 1289.280 1062.830 ;
        RECT 1289.940 1062.510 1290.200 1062.830 ;
        RECT 1278.040 1057.730 1278.180 1062.510 ;
        RECT 1277.980 1057.410 1278.240 1057.730 ;
        RECT 1280.740 1057.410 1281.000 1057.730 ;
        RECT 1278.900 1021.030 1279.160 1021.350 ;
        RECT 1270.160 1020.010 1270.420 1020.330 ;
        RECT 1269.240 1012.530 1269.500 1012.850 ;
        RECT 1268.380 1010.750 1268.980 1010.890 ;
        RECT 1268.380 1010.130 1268.520 1010.750 ;
        RECT 1268.320 1009.810 1268.580 1010.130 ;
        RECT 1268.780 1009.810 1269.040 1010.130 ;
        RECT 1268.840 1000.010 1268.980 1009.810 ;
        RECT 1269.300 1008.430 1269.440 1012.530 ;
        RECT 1269.700 1011.850 1269.960 1012.170 ;
        RECT 1269.760 1011.685 1269.900 1011.850 ;
        RECT 1269.690 1011.315 1269.970 1011.685 ;
        RECT 1269.240 1008.110 1269.500 1008.430 ;
        RECT 1259.640 1000.000 1259.940 1000.010 ;
        RECT 1262.240 1000.000 1263.920 1000.010 ;
        RECT 1264.540 1000.000 1265.760 1000.010 ;
        RECT 1266.380 1000.000 1268.060 1000.010 ;
        RECT 1268.680 1000.000 1268.980 1000.010 ;
        RECT 1259.640 999.870 1260.090 1000.000 ;
      LAYER met2 ;
        RECT 1247.490 995.720 1248.950 998.810 ;
      LAYER met2 ;
        RECT 1249.230 996.000 1249.510 999.870 ;
      LAYER met2 ;
        RECT 1249.790 995.720 1250.790 998.810 ;
      LAYER met2 ;
        RECT 1251.070 996.000 1251.350 999.870 ;
      LAYER met2 ;
        RECT 1251.630 995.720 1253.090 998.810 ;
      LAYER met2 ;
        RECT 1253.370 996.000 1253.650 999.870 ;
      LAYER met2 ;
        RECT 1253.930 995.720 1255.390 998.810 ;
      LAYER met2 ;
        RECT 1255.670 996.000 1255.950 999.870 ;
      LAYER met2 ;
        RECT 1256.230 995.720 1257.690 998.810 ;
      LAYER met2 ;
        RECT 1257.970 996.000 1258.250 999.870 ;
      LAYER met2 ;
        RECT 1258.530 995.720 1259.530 998.810 ;
      LAYER met2 ;
        RECT 1259.810 996.000 1260.090 999.870 ;
        RECT 1262.110 999.870 1263.920 1000.000 ;
        RECT 1264.410 999.870 1265.760 1000.000 ;
        RECT 1266.250 999.870 1268.060 1000.000 ;
        RECT 1268.550 999.870 1268.980 1000.000 ;
        RECT 1270.220 1000.010 1270.360 1020.010 ;
        RECT 1270.620 1012.365 1270.880 1012.510 ;
        RECT 1270.610 1011.995 1270.890 1012.365 ;
        RECT 1274.300 1008.450 1274.560 1008.770 ;
        RECT 1274.360 1000.010 1274.500 1008.450 ;
        RECT 1274.990 1000.970 1275.250 1001.290 ;
        RECT 1270.220 1000.000 1270.980 1000.010 ;
        RECT 1273.280 1000.000 1274.500 1000.010 ;
        RECT 1275.050 1000.000 1275.190 1000.970 ;
        RECT 1278.960 1000.010 1279.100 1021.030 ;
        RECT 1279.820 1020.010 1280.080 1020.330 ;
        RECT 1279.880 1000.010 1280.020 1020.010 ;
        RECT 1277.420 1000.000 1279.100 1000.010 ;
        RECT 1279.720 1000.000 1280.020 1000.010 ;
        RECT 1270.220 999.870 1271.130 1000.000 ;
      LAYER met2 ;
        RECT 1260.370 995.720 1261.830 998.810 ;
      LAYER met2 ;
        RECT 1262.110 996.000 1262.390 999.870 ;
      LAYER met2 ;
        RECT 1262.670 995.720 1264.130 998.810 ;
      LAYER met2 ;
        RECT 1264.410 996.000 1264.690 999.870 ;
      LAYER met2 ;
        RECT 1264.970 995.720 1265.970 998.810 ;
      LAYER met2 ;
        RECT 1266.250 996.000 1266.530 999.870 ;
      LAYER met2 ;
        RECT 1266.810 995.720 1268.270 998.810 ;
      LAYER met2 ;
        RECT 1268.550 996.000 1268.830 999.870 ;
      LAYER met2 ;
        RECT 1269.110 995.720 1270.570 998.810 ;
      LAYER met2 ;
        RECT 1270.850 996.000 1271.130 999.870 ;
        RECT 1273.150 999.870 1274.500 1000.000 ;
      LAYER met2 ;
        RECT 1271.410 995.720 1272.870 998.810 ;
      LAYER met2 ;
        RECT 1273.150 996.000 1273.430 999.870 ;
      LAYER met2 ;
        RECT 1273.710 995.720 1274.710 998.810 ;
      LAYER met2 ;
        RECT 1274.990 996.000 1275.270 1000.000 ;
        RECT 1277.290 999.870 1279.100 1000.000 ;
        RECT 1279.590 999.870 1280.020 1000.000 ;
        RECT 1280.800 1000.010 1280.940 1057.410 ;
        RECT 1289.080 1028.570 1289.220 1062.510 ;
        RECT 1289.080 1028.430 1289.680 1028.570 ;
        RECT 1289.540 1027.890 1289.680 1028.430 ;
        RECT 1288.620 1027.750 1289.680 1027.890 ;
        RECT 1285.800 1019.330 1286.060 1019.650 ;
        RECT 1282.580 1010.830 1282.840 1011.150 ;
        RECT 1282.640 1009.110 1282.780 1010.830 ;
        RECT 1285.340 1009.130 1285.600 1009.450 ;
        RECT 1282.580 1008.790 1282.840 1009.110 ;
        RECT 1285.400 1000.010 1285.540 1009.130 ;
        RECT 1280.800 1000.000 1282.020 1000.010 ;
        RECT 1283.860 1000.000 1285.540 1000.010 ;
        RECT 1280.800 999.870 1282.170 1000.000 ;
      LAYER met2 ;
        RECT 1275.550 995.720 1277.010 998.810 ;
      LAYER met2 ;
        RECT 1277.290 996.000 1277.570 999.870 ;
      LAYER met2 ;
        RECT 1277.850 995.720 1279.310 998.810 ;
      LAYER met2 ;
        RECT 1279.590 996.000 1279.870 999.870 ;
      LAYER met2 ;
        RECT 1280.150 995.720 1281.610 998.810 ;
      LAYER met2 ;
        RECT 1281.890 996.000 1282.170 999.870 ;
        RECT 1283.730 999.870 1285.540 1000.000 ;
        RECT 1285.860 1000.010 1286.000 1019.330 ;
        RECT 1288.620 1014.120 1288.760 1027.750 ;
        RECT 1292.300 1020.410 1292.440 1076.110 ;
        RECT 1292.300 1020.270 1293.360 1020.410 ;
        RECT 1292.240 1019.670 1292.500 1019.990 ;
        RECT 1288.160 1013.980 1288.760 1014.120 ;
        RECT 1288.160 1000.690 1288.300 1013.980 ;
        RECT 1291.780 1008.110 1292.040 1008.430 ;
        RECT 1288.160 1000.550 1288.530 1000.690 ;
        RECT 1285.860 1000.000 1286.160 1000.010 ;
        RECT 1288.390 1000.000 1288.530 1000.550 ;
        RECT 1291.840 1000.010 1291.980 1008.110 ;
        RECT 1290.300 1000.000 1291.980 1000.010 ;
        RECT 1285.860 999.870 1286.310 1000.000 ;
      LAYER met2 ;
        RECT 1282.450 995.720 1283.450 998.810 ;
      LAYER met2 ;
        RECT 1283.730 996.000 1284.010 999.870 ;
      LAYER met2 ;
        RECT 1284.290 995.720 1285.750 998.810 ;
      LAYER met2 ;
        RECT 1286.030 996.000 1286.310 999.870 ;
      LAYER met2 ;
        RECT 1286.590 995.720 1288.050 998.810 ;
      LAYER met2 ;
        RECT 1288.330 996.000 1288.610 1000.000 ;
        RECT 1290.170 999.870 1291.980 1000.000 ;
        RECT 1292.300 1000.010 1292.440 1019.670 ;
        RECT 1292.690 1011.315 1292.970 1011.685 ;
        RECT 1292.700 1011.170 1292.960 1011.315 ;
        RECT 1293.220 1000.690 1293.360 1020.270 ;
        RECT 1293.680 1013.870 1293.820 1688.450 ;
        RECT 1300.520 1686.070 1300.780 1686.390 ;
        RECT 1299.140 1019.330 1299.400 1019.650 ;
        RECT 1294.080 1014.230 1294.340 1014.550 ;
        RECT 1293.620 1013.550 1293.880 1013.870 ;
        RECT 1294.140 1010.130 1294.280 1014.230 ;
        RECT 1295.000 1013.890 1295.260 1014.210 ;
        RECT 1295.060 1011.150 1295.200 1013.890 ;
        RECT 1297.290 1011.315 1297.570 1011.685 ;
        RECT 1295.000 1010.830 1295.260 1011.150 ;
        RECT 1294.540 1010.490 1294.800 1010.810 ;
        RECT 1293.620 1009.810 1293.880 1010.130 ;
        RECT 1294.080 1009.810 1294.340 1010.130 ;
        RECT 1293.680 1008.090 1293.820 1009.810 ;
        RECT 1293.620 1007.770 1293.880 1008.090 ;
        RECT 1294.600 1001.290 1294.740 1010.490 ;
        RECT 1294.540 1000.970 1294.800 1001.290 ;
        RECT 1293.220 1000.550 1293.820 1000.690 ;
        RECT 1293.680 1000.010 1293.820 1000.550 ;
        RECT 1297.360 1000.010 1297.500 1011.315 ;
        RECT 1299.200 1000.010 1299.340 1019.330 ;
        RECT 1300.580 1014.210 1300.720 1686.070 ;
        RECT 1301.900 1018.990 1302.160 1019.310 ;
        RECT 1300.520 1013.890 1300.780 1014.210 ;
        RECT 1299.600 1008.790 1299.860 1009.110 ;
        RECT 1292.300 1000.000 1292.600 1000.010 ;
        RECT 1293.680 1000.000 1294.900 1000.010 ;
        RECT 1297.200 1000.000 1297.500 1000.010 ;
        RECT 1299.040 1000.000 1299.340 1000.010 ;
        RECT 1292.300 999.870 1292.750 1000.000 ;
        RECT 1293.680 999.870 1295.050 1000.000 ;
      LAYER met2 ;
        RECT 1288.890 995.720 1289.890 998.810 ;
      LAYER met2 ;
        RECT 1290.170 996.000 1290.450 999.870 ;
      LAYER met2 ;
        RECT 1290.730 995.720 1292.190 998.810 ;
      LAYER met2 ;
        RECT 1292.470 996.000 1292.750 999.870 ;
      LAYER met2 ;
        RECT 1293.030 995.720 1294.490 998.810 ;
      LAYER met2 ;
        RECT 1294.770 996.000 1295.050 999.870 ;
        RECT 1297.070 999.870 1297.500 1000.000 ;
        RECT 1298.910 999.870 1299.340 1000.000 ;
        RECT 1299.660 1000.010 1299.800 1008.790 ;
        RECT 1301.960 1000.010 1302.100 1018.990 ;
        RECT 1310.700 1011.570 1310.840 1692.870 ;
        RECT 1315.760 1689.790 1315.900 1700.000 ;
        RECT 1315.700 1689.470 1315.960 1689.790 ;
        RECT 1329.560 1684.350 1329.700 1700.000 ;
        RECT 1329.500 1684.030 1329.760 1684.350 ;
        RECT 1313.860 1018.650 1314.120 1018.970 ;
        RECT 1308.860 1011.430 1310.840 1011.570 ;
        RECT 1304.200 1009.470 1304.460 1009.790 ;
        RECT 1304.260 1000.010 1304.400 1009.470 ;
        RECT 1308.860 1000.010 1309.000 1011.430 ;
        RECT 1309.710 1010.635 1309.990 1011.005 ;
        RECT 1299.660 1000.000 1301.340 1000.010 ;
        RECT 1301.960 1000.000 1303.640 1000.010 ;
        RECT 1304.260 1000.000 1305.940 1000.010 ;
        RECT 1307.780 1000.000 1309.000 1000.010 ;
        RECT 1299.660 999.870 1301.490 1000.000 ;
        RECT 1301.960 999.870 1303.790 1000.000 ;
        RECT 1304.260 999.870 1306.090 1000.000 ;
      LAYER met2 ;
        RECT 1295.330 995.720 1296.790 998.810 ;
      LAYER met2 ;
        RECT 1297.070 996.000 1297.350 999.870 ;
      LAYER met2 ;
        RECT 1297.630 995.720 1298.630 998.810 ;
      LAYER met2 ;
        RECT 1298.910 996.000 1299.190 999.870 ;
      LAYER met2 ;
        RECT 1299.470 995.720 1300.930 998.810 ;
      LAYER met2 ;
        RECT 1301.210 996.000 1301.490 999.870 ;
      LAYER met2 ;
        RECT 1301.770 995.720 1303.230 998.810 ;
      LAYER met2 ;
        RECT 1303.510 996.000 1303.790 999.870 ;
      LAYER met2 ;
        RECT 1304.070 995.720 1305.530 998.810 ;
      LAYER met2 ;
        RECT 1305.810 996.000 1306.090 999.870 ;
        RECT 1307.650 999.870 1309.000 1000.000 ;
        RECT 1309.780 1000.010 1309.920 1010.635 ;
        RECT 1313.400 1008.450 1313.660 1008.770 ;
        RECT 1313.460 1000.010 1313.600 1008.450 ;
        RECT 1309.780 1000.000 1310.080 1000.010 ;
        RECT 1312.380 1000.000 1313.600 1000.010 ;
        RECT 1309.780 999.870 1310.230 1000.000 ;
      LAYER met2 ;
        RECT 1306.370 995.720 1307.370 998.810 ;
      LAYER met2 ;
        RECT 1307.650 996.000 1307.930 999.870 ;
      LAYER met2 ;
        RECT 1308.210 995.720 1309.670 998.810 ;
      LAYER met2 ;
        RECT 1309.950 996.000 1310.230 999.870 ;
        RECT 1312.250 999.870 1313.600 1000.000 ;
        RECT 1313.920 1000.010 1314.060 1018.650 ;
        RECT 1314.780 1018.310 1315.040 1018.630 ;
        RECT 1314.840 1000.010 1314.980 1018.310 ;
        RECT 1327.200 1017.970 1327.460 1018.290 ;
        RECT 1318.000 1013.890 1318.260 1014.210 ;
        RECT 1318.060 1000.010 1318.200 1013.890 ;
        RECT 1319.380 1013.550 1319.640 1013.870 ;
        RECT 1324.440 1013.550 1324.700 1013.870 ;
        RECT 1319.440 1000.010 1319.580 1013.550 ;
        RECT 1324.500 1000.010 1324.640 1013.550 ;
        RECT 1326.740 1009.470 1327.000 1009.790 ;
        RECT 1326.800 1000.010 1326.940 1009.470 ;
        RECT 1313.920 1000.000 1314.220 1000.010 ;
        RECT 1314.840 1000.000 1316.520 1000.010 ;
        RECT 1318.060 1000.000 1318.820 1000.010 ;
        RECT 1319.440 1000.000 1321.120 1000.010 ;
        RECT 1322.960 1000.000 1324.640 1000.010 ;
        RECT 1325.260 1000.000 1326.940 1000.010 ;
        RECT 1313.920 999.870 1314.370 1000.000 ;
        RECT 1314.840 999.870 1316.670 1000.000 ;
        RECT 1318.060 999.870 1318.970 1000.000 ;
        RECT 1319.440 999.870 1321.270 1000.000 ;
      LAYER met2 ;
        RECT 1310.510 995.720 1311.970 998.810 ;
      LAYER met2 ;
        RECT 1312.250 996.000 1312.530 999.870 ;
      LAYER met2 ;
        RECT 1312.810 995.720 1313.810 998.810 ;
      LAYER met2 ;
        RECT 1314.090 996.000 1314.370 999.870 ;
      LAYER met2 ;
        RECT 1314.650 995.720 1316.110 998.810 ;
      LAYER met2 ;
        RECT 1316.390 996.000 1316.670 999.870 ;
      LAYER met2 ;
        RECT 1316.950 995.720 1318.410 998.810 ;
      LAYER met2 ;
        RECT 1318.690 996.000 1318.970 999.870 ;
      LAYER met2 ;
        RECT 1319.250 995.720 1320.710 998.810 ;
      LAYER met2 ;
        RECT 1320.990 996.000 1321.270 999.870 ;
        RECT 1322.830 999.870 1324.640 1000.000 ;
        RECT 1325.130 999.870 1326.940 1000.000 ;
        RECT 1327.260 1000.010 1327.400 1017.970 ;
        RECT 1331.340 1013.890 1331.600 1014.210 ;
        RECT 1331.400 1012.510 1331.540 1013.890 ;
        RECT 1331.340 1012.190 1331.600 1012.510 ;
        RECT 1330.420 1011.510 1330.680 1011.830 ;
        RECT 1330.880 1011.510 1331.140 1011.830 ;
        RECT 1330.480 1009.450 1330.620 1011.510 ;
        RECT 1329.960 1009.130 1330.220 1009.450 ;
        RECT 1330.420 1009.130 1330.680 1009.450 ;
        RECT 1330.020 1008.770 1330.160 1009.130 ;
        RECT 1329.500 1008.450 1329.760 1008.770 ;
        RECT 1329.960 1008.450 1330.220 1008.770 ;
        RECT 1329.560 1007.410 1329.700 1008.450 ;
        RECT 1329.500 1007.090 1329.760 1007.410 ;
        RECT 1330.940 1000.010 1331.080 1011.510 ;
        RECT 1331.860 1008.090 1332.000 2054.970 ;
        RECT 1335.020 2054.630 1335.280 2054.950 ;
        RECT 1332.720 2053.950 1332.980 2054.270 ;
        RECT 1332.260 2052.250 1332.520 2052.570 ;
        RECT 1332.320 1010.130 1332.460 2052.250 ;
        RECT 1332.260 1009.810 1332.520 1010.130 ;
        RECT 1332.780 1009.530 1332.920 2053.950 ;
        RECT 1333.640 2053.270 1333.900 2053.590 ;
        RECT 1333.180 2049.870 1333.440 2050.190 ;
        RECT 1332.320 1009.390 1332.920 1009.530 ;
        RECT 1333.240 1009.530 1333.380 2049.870 ;
        RECT 1333.700 1011.150 1333.840 2053.270 ;
        RECT 1334.090 1997.995 1334.370 1998.365 ;
        RECT 1333.640 1010.830 1333.900 1011.150 ;
        RECT 1334.160 1009.790 1334.300 1997.995 ;
        RECT 1334.550 1913.675 1334.830 1914.045 ;
        RECT 1334.620 1021.350 1334.760 1913.675 ;
        RECT 1334.560 1021.030 1334.820 1021.350 ;
        RECT 1335.080 1009.790 1335.220 2054.630 ;
        RECT 1346.060 2052.590 1346.320 2052.910 ;
        RECT 1336.400 2051.910 1336.660 2052.230 ;
        RECT 1335.470 1787.195 1335.750 1787.565 ;
        RECT 1333.240 1009.390 1333.840 1009.530 ;
        RECT 1334.100 1009.470 1334.360 1009.790 ;
        RECT 1335.020 1009.470 1335.280 1009.790 ;
        RECT 1332.320 1009.110 1332.460 1009.390 ;
        RECT 1332.260 1008.790 1332.520 1009.110 ;
        RECT 1333.700 1008.430 1333.840 1009.390 ;
        RECT 1335.540 1008.680 1335.680 1787.195 ;
        RECT 1335.930 1745.035 1336.210 1745.405 ;
        RECT 1336.000 1019.650 1336.140 1745.035 ;
        RECT 1336.460 1694.210 1336.600 2051.910 ;
        RECT 1336.860 2049.530 1337.120 2049.850 ;
        RECT 1336.400 1693.890 1336.660 1694.210 ;
        RECT 1336.920 1693.870 1337.060 2049.530 ;
        RECT 1343.760 2049.190 1344.020 2049.510 ;
        RECT 1338.690 2018.395 1338.970 2018.765 ;
        RECT 1336.860 1693.550 1337.120 1693.870 ;
        RECT 1335.940 1019.330 1336.200 1019.650 ;
        RECT 1335.940 1017.630 1336.200 1017.950 ;
        RECT 1334.160 1008.540 1335.680 1008.680 ;
        RECT 1333.640 1008.110 1333.900 1008.430 ;
        RECT 1331.800 1007.770 1332.060 1008.090 ;
        RECT 1332.260 1007.490 1332.520 1007.750 ;
        RECT 1333.180 1007.490 1333.440 1007.750 ;
        RECT 1332.260 1007.430 1333.440 1007.490 ;
        RECT 1332.320 1007.350 1333.380 1007.430 ;
        RECT 1334.160 1000.690 1334.300 1008.540 ;
        RECT 1335.480 1007.770 1335.740 1008.090 ;
        RECT 1333.240 1000.550 1334.300 1000.690 ;
        RECT 1333.240 1000.010 1333.380 1000.550 ;
        RECT 1335.540 1000.010 1335.680 1007.770 ;
        RECT 1327.260 1000.000 1327.560 1000.010 ;
        RECT 1329.860 1000.000 1331.080 1000.010 ;
        RECT 1331.700 1000.000 1333.380 1000.010 ;
        RECT 1334.000 1000.000 1335.680 1000.010 ;
        RECT 1327.260 999.870 1327.710 1000.000 ;
      LAYER met2 ;
        RECT 1321.550 995.720 1322.550 998.810 ;
      LAYER met2 ;
        RECT 1322.830 996.000 1323.110 999.870 ;
      LAYER met2 ;
        RECT 1323.390 995.720 1324.850 998.810 ;
      LAYER met2 ;
        RECT 1325.130 996.000 1325.410 999.870 ;
      LAYER met2 ;
        RECT 1325.690 995.720 1327.150 998.810 ;
      LAYER met2 ;
        RECT 1327.430 996.000 1327.710 999.870 ;
        RECT 1329.730 999.870 1331.080 1000.000 ;
        RECT 1331.570 999.870 1333.380 1000.000 ;
        RECT 1333.870 999.870 1335.680 1000.000 ;
        RECT 1336.000 1000.010 1336.140 1017.630 ;
        RECT 1338.240 1012.190 1338.500 1012.510 ;
        RECT 1338.300 1000.010 1338.440 1012.190 ;
        RECT 1338.760 1010.470 1338.900 2018.395 ;
        RECT 1339.150 1976.235 1339.430 1976.605 ;
        RECT 1339.220 1021.010 1339.360 1976.235 ;
        RECT 1339.610 1955.835 1339.890 1956.205 ;
        RECT 1339.160 1020.690 1339.420 1021.010 ;
        RECT 1339.680 1012.850 1339.820 1955.835 ;
        RECT 1340.070 1934.075 1340.350 1934.445 ;
        RECT 1339.620 1012.530 1339.880 1012.850 ;
        RECT 1340.140 1012.170 1340.280 1934.075 ;
        RECT 1340.530 1891.915 1340.810 1892.285 ;
        RECT 1340.600 1013.190 1340.740 1891.915 ;
        RECT 1340.990 1871.515 1341.270 1871.885 ;
        RECT 1340.540 1012.870 1340.800 1013.190 ;
        RECT 1340.080 1011.850 1340.340 1012.170 ;
        RECT 1338.700 1010.150 1338.960 1010.470 ;
        RECT 1341.060 1010.210 1341.200 1871.515 ;
        RECT 1341.450 1849.755 1341.730 1850.125 ;
        RECT 1341.520 1010.810 1341.660 1849.755 ;
        RECT 1341.910 1829.355 1342.190 1829.725 ;
        RECT 1341.980 1020.330 1342.120 1829.355 ;
        RECT 1342.370 1807.595 1342.650 1807.965 ;
        RECT 1342.440 1052.290 1342.580 1807.595 ;
        RECT 1342.830 1766.795 1343.110 1767.165 ;
        RECT 1342.380 1051.970 1342.640 1052.290 ;
        RECT 1341.920 1020.010 1342.180 1020.330 ;
        RECT 1342.900 1017.610 1343.040 1766.795 ;
        RECT 1343.290 1724.635 1343.570 1725.005 ;
        RECT 1343.360 1020.670 1343.500 1724.635 ;
        RECT 1343.820 1693.190 1343.960 2049.190 ;
        RECT 1343.760 1692.870 1344.020 1693.190 ;
        RECT 1344.220 1051.970 1344.480 1052.290 ;
        RECT 1343.300 1020.350 1343.560 1020.670 ;
        RECT 1342.840 1017.290 1343.100 1017.610 ;
        RECT 1341.460 1010.490 1341.720 1010.810 ;
        RECT 1340.140 1010.070 1341.200 1010.210 ;
        RECT 1340.140 1007.750 1340.280 1010.070 ;
        RECT 1341.000 1009.470 1341.260 1009.790 ;
        RECT 1340.540 1008.450 1340.800 1008.770 ;
        RECT 1340.080 1007.430 1340.340 1007.750 ;
        RECT 1340.600 1000.010 1340.740 1008.450 ;
        RECT 1336.000 1000.000 1336.300 1000.010 ;
        RECT 1338.140 1000.000 1338.440 1000.010 ;
        RECT 1340.440 1000.000 1340.740 1000.010 ;
        RECT 1336.000 999.870 1336.450 1000.000 ;
      LAYER met2 ;
        RECT 1327.990 995.720 1329.450 998.810 ;
      LAYER met2 ;
        RECT 1329.730 996.000 1330.010 999.870 ;
      LAYER met2 ;
        RECT 1330.290 995.720 1331.290 998.810 ;
      LAYER met2 ;
        RECT 1331.570 996.000 1331.850 999.870 ;
      LAYER met2 ;
        RECT 1332.130 995.720 1333.590 998.810 ;
      LAYER met2 ;
        RECT 1333.870 996.000 1334.150 999.870 ;
      LAYER met2 ;
        RECT 1334.430 995.720 1335.890 998.810 ;
      LAYER met2 ;
        RECT 1336.170 996.000 1336.450 999.870 ;
        RECT 1338.010 999.870 1338.440 1000.000 ;
        RECT 1340.310 999.870 1340.740 1000.000 ;
        RECT 1341.060 1000.010 1341.200 1009.470 ;
        RECT 1344.280 1000.010 1344.420 1051.970 ;
        RECT 1346.120 1013.530 1346.260 2052.590 ;
        RECT 1346.520 2051.570 1346.780 2051.890 ;
        RECT 1346.060 1013.210 1346.320 1013.530 ;
        RECT 1346.580 1012.510 1346.720 2051.570 ;
        RECT 1346.980 2050.550 1347.240 2050.870 ;
        RECT 1347.040 1014.210 1347.180 2050.550 ;
        RECT 1347.440 2050.210 1347.700 2050.530 ;
        RECT 1346.980 1013.890 1347.240 1014.210 ;
        RECT 1347.500 1013.870 1347.640 2050.210 ;
        RECT 1347.440 1013.550 1347.700 1013.870 ;
        RECT 1346.520 1012.190 1346.780 1012.510 ;
        RECT 1347.960 1011.830 1348.100 2055.310 ;
        RECT 1348.360 1684.030 1348.620 1684.350 ;
        RECT 1347.900 1011.510 1348.160 1011.830 ;
        RECT 1348.420 1000.010 1348.560 1684.030 ;
        RECT 1348.820 1011.170 1349.080 1011.490 ;
        RECT 1341.060 1000.000 1342.740 1000.010 ;
        RECT 1344.280 1000.000 1345.040 1000.010 ;
        RECT 1346.880 1000.000 1348.560 1000.010 ;
        RECT 1341.060 999.870 1342.890 1000.000 ;
        RECT 1344.280 999.870 1345.190 1000.000 ;
      LAYER met2 ;
        RECT 1336.730 995.720 1337.730 998.810 ;
      LAYER met2 ;
        RECT 1338.010 996.000 1338.290 999.870 ;
      LAYER met2 ;
        RECT 1338.570 995.720 1340.030 998.810 ;
      LAYER met2 ;
        RECT 1340.310 996.000 1340.590 999.870 ;
      LAYER met2 ;
        RECT 1340.870 995.720 1342.330 998.810 ;
      LAYER met2 ;
        RECT 1342.610 996.000 1342.890 999.870 ;
      LAYER met2 ;
        RECT 1343.170 995.720 1344.630 998.810 ;
      LAYER met2 ;
        RECT 1344.910 996.000 1345.190 999.870 ;
        RECT 1346.750 999.870 1348.560 1000.000 ;
        RECT 1348.880 1000.010 1349.020 1011.170 ;
        RECT 1352.100 1000.010 1352.240 2917.890 ;
        RECT 1414.140 2917.550 1414.400 2917.870 ;
        RECT 1379.640 2915.510 1379.900 2915.830 ;
        RECT 1372.740 2913.470 1373.000 2913.790 ;
        RECT 1358.940 2849.550 1359.200 2849.870 ;
        RECT 1359.000 2815.725 1359.140 2849.550 ;
        RECT 1358.930 2815.355 1359.210 2815.725 ;
        RECT 1358.470 2814.675 1358.750 2815.045 ;
        RECT 1358.540 2801.445 1358.680 2814.675 ;
        RECT 1357.550 2801.075 1357.830 2801.445 ;
        RECT 1358.470 2801.075 1358.750 2801.445 ;
        RECT 1357.620 2753.310 1357.760 2801.075 ;
        RECT 1365.840 2780.870 1366.100 2781.190 ;
        RECT 1357.560 2752.990 1357.820 2753.310 ;
        RECT 1358.940 2752.990 1359.200 2753.310 ;
        RECT 1359.000 2729.170 1359.140 2752.990 ;
        RECT 1357.560 2728.850 1357.820 2729.170 ;
        RECT 1358.940 2728.850 1359.200 2729.170 ;
        RECT 1357.620 2705.030 1357.760 2728.850 ;
        RECT 1357.560 2704.710 1357.820 2705.030 ;
        RECT 1358.020 2704.770 1358.280 2705.030 ;
        RECT 1358.470 2704.770 1358.750 2704.885 ;
        RECT 1358.020 2704.710 1358.750 2704.770 ;
        RECT 1358.080 2704.630 1358.750 2704.710 ;
        RECT 1358.470 2704.515 1358.750 2704.630 ;
        RECT 1359.850 2704.515 1360.130 2704.885 ;
        RECT 1359.920 2656.750 1360.060 2704.515 ;
        RECT 1358.940 2656.430 1359.200 2656.750 ;
        RECT 1359.860 2656.430 1360.120 2656.750 ;
        RECT 1359.000 2622.750 1359.140 2656.430 ;
        RECT 1358.940 2622.430 1359.200 2622.750 ;
        RECT 1358.940 2621.750 1359.200 2622.070 ;
        RECT 1359.000 2574.130 1359.140 2621.750 ;
        RECT 1358.940 2573.810 1359.200 2574.130 ;
        RECT 1358.480 2573.470 1358.740 2573.790 ;
        RECT 1358.540 2560.190 1358.680 2573.470 ;
        RECT 1358.480 2559.870 1358.740 2560.190 ;
        RECT 1358.940 2559.870 1359.200 2560.190 ;
        RECT 1359.000 2536.050 1359.140 2559.870 ;
        RECT 1357.560 2535.730 1357.820 2536.050 ;
        RECT 1358.940 2535.730 1359.200 2536.050 ;
        RECT 1357.620 2511.910 1357.760 2535.730 ;
        RECT 1357.560 2511.590 1357.820 2511.910 ;
        RECT 1358.020 2511.765 1358.280 2511.910 ;
        RECT 1358.010 2511.395 1358.290 2511.765 ;
        RECT 1358.930 2463.115 1359.210 2463.485 ;
        RECT 1359.000 2439.150 1359.140 2463.115 ;
        RECT 1357.560 2438.830 1357.820 2439.150 ;
        RECT 1358.940 2438.830 1359.200 2439.150 ;
        RECT 1357.620 2415.690 1357.760 2438.830 ;
        RECT 1357.560 2415.370 1357.820 2415.690 ;
        RECT 1358.480 2415.370 1358.740 2415.690 ;
        RECT 1358.540 2415.010 1358.680 2415.370 ;
        RECT 1358.480 2414.690 1358.740 2415.010 ;
        RECT 1358.940 2414.690 1359.200 2415.010 ;
        RECT 1359.000 2380.670 1359.140 2414.690 ;
        RECT 1358.940 2380.350 1359.200 2380.670 ;
        RECT 1358.480 2380.010 1358.740 2380.330 ;
        RECT 1358.540 2366.810 1358.680 2380.010 ;
        RECT 1358.540 2366.670 1359.140 2366.810 ;
        RECT 1359.000 2342.590 1359.140 2366.670 ;
        RECT 1357.560 2342.270 1357.820 2342.590 ;
        RECT 1358.940 2342.270 1359.200 2342.590 ;
        RECT 1357.620 2319.130 1357.760 2342.270 ;
        RECT 1357.560 2318.810 1357.820 2319.130 ;
        RECT 1358.480 2318.810 1358.740 2319.130 ;
        RECT 1358.540 2318.450 1358.680 2318.810 ;
        RECT 1358.480 2318.130 1358.740 2318.450 ;
        RECT 1358.940 2318.130 1359.200 2318.450 ;
        RECT 1359.000 2284.110 1359.140 2318.130 ;
        RECT 1358.940 2283.790 1359.200 2284.110 ;
        RECT 1358.480 2283.450 1358.740 2283.770 ;
        RECT 1358.540 2270.250 1358.680 2283.450 ;
        RECT 1358.540 2270.110 1359.140 2270.250 ;
        RECT 1359.000 2246.030 1359.140 2270.110 ;
        RECT 1357.560 2245.710 1357.820 2246.030 ;
        RECT 1358.940 2245.710 1359.200 2246.030 ;
        RECT 1357.620 2222.570 1357.760 2245.710 ;
        RECT 1357.560 2222.250 1357.820 2222.570 ;
        RECT 1358.480 2222.250 1358.740 2222.570 ;
        RECT 1358.540 2221.890 1358.680 2222.250 ;
        RECT 1358.480 2221.570 1358.740 2221.890 ;
        RECT 1358.940 2221.570 1359.200 2221.890 ;
        RECT 1359.000 2187.550 1359.140 2221.570 ;
        RECT 1358.940 2187.230 1359.200 2187.550 ;
        RECT 1358.480 2186.890 1358.740 2187.210 ;
        RECT 1358.540 2173.690 1358.680 2186.890 ;
        RECT 1358.540 2173.550 1359.140 2173.690 ;
        RECT 1359.000 2149.470 1359.140 2173.550 ;
        RECT 1357.560 2149.150 1357.820 2149.470 ;
        RECT 1358.940 2149.150 1359.200 2149.470 ;
        RECT 1357.620 2126.010 1357.760 2149.150 ;
        RECT 1357.560 2125.690 1357.820 2126.010 ;
        RECT 1358.480 2125.690 1358.740 2126.010 ;
        RECT 1358.540 2125.330 1358.680 2125.690 ;
        RECT 1358.480 2125.010 1358.740 2125.330 ;
        RECT 1358.940 2125.010 1359.200 2125.330 ;
        RECT 1359.000 2097.645 1359.140 2125.010 ;
        RECT 1358.930 2097.275 1359.210 2097.645 ;
        RECT 1359.850 2097.275 1360.130 2097.645 ;
        RECT 1353.880 2054.290 1354.140 2054.610 ;
        RECT 1353.420 2053.610 1353.680 2053.930 ;
        RECT 1352.500 2052.930 1352.760 2053.250 ;
        RECT 1352.560 1008.090 1352.700 2052.930 ;
        RECT 1352.960 2050.890 1353.220 2051.210 ;
        RECT 1353.020 1008.770 1353.160 2050.890 ;
        RECT 1353.480 1009.450 1353.620 2053.610 ;
        RECT 1353.420 1009.130 1353.680 1009.450 ;
        RECT 1352.960 1008.450 1353.220 1008.770 ;
        RECT 1353.940 1008.430 1354.080 2054.290 ;
        RECT 1354.340 2051.230 1354.600 2051.550 ;
        RECT 1354.400 1009.110 1354.540 2051.230 ;
        RECT 1359.920 2042.710 1360.060 2097.275 ;
        RECT 1358.020 2042.390 1358.280 2042.710 ;
        RECT 1359.860 2042.390 1360.120 2042.710 ;
        RECT 1358.080 1994.090 1358.220 2042.390 ;
        RECT 1358.020 1993.770 1358.280 1994.090 ;
        RECT 1358.940 1993.770 1359.200 1994.090 ;
        RECT 1359.000 1946.005 1359.140 1993.770 ;
        RECT 1357.560 1945.490 1357.820 1945.810 ;
        RECT 1358.010 1945.635 1358.290 1946.005 ;
        RECT 1358.930 1945.635 1359.210 1946.005 ;
        RECT 1358.020 1945.490 1358.280 1945.635 ;
        RECT 1357.620 1921.330 1357.760 1945.490 ;
        RECT 1357.560 1921.010 1357.820 1921.330 ;
        RECT 1358.480 1921.010 1358.740 1921.330 ;
        RECT 1358.540 1897.610 1358.680 1921.010 ;
        RECT 1358.540 1897.530 1359.140 1897.610 ;
        RECT 1358.480 1897.470 1359.200 1897.530 ;
        RECT 1358.480 1897.210 1358.740 1897.470 ;
        RECT 1358.940 1897.210 1359.200 1897.470 ;
        RECT 1358.540 1801.310 1358.680 1897.210 ;
        RECT 1359.000 1897.055 1359.140 1897.210 ;
        RECT 1358.480 1800.990 1358.740 1801.310 ;
        RECT 1358.940 1800.990 1359.200 1801.310 ;
        RECT 1359.000 1684.690 1359.140 1800.990 ;
        RECT 1358.940 1684.370 1359.200 1684.690 ;
        RECT 1358.480 1684.030 1358.740 1684.350 ;
        RECT 1358.540 1663.010 1358.680 1684.030 ;
        RECT 1358.080 1662.870 1358.680 1663.010 ;
        RECT 1358.080 1652.730 1358.220 1662.870 ;
        RECT 1357.100 1652.410 1357.360 1652.730 ;
        RECT 1358.020 1652.410 1358.280 1652.730 ;
        RECT 1357.160 1628.590 1357.300 1652.410 ;
        RECT 1357.100 1628.270 1357.360 1628.590 ;
        RECT 1357.560 1628.270 1357.820 1628.590 ;
        RECT 1357.620 1614.650 1357.760 1628.270 ;
        RECT 1357.560 1614.330 1357.820 1614.650 ;
        RECT 1358.480 1614.330 1358.740 1614.650 ;
        RECT 1358.540 1566.450 1358.680 1614.330 ;
        RECT 1358.540 1566.310 1359.140 1566.450 ;
        RECT 1359.000 1518.090 1359.140 1566.310 ;
        RECT 1358.940 1517.770 1359.200 1518.090 ;
        RECT 1359.860 1517.770 1360.120 1518.090 ;
        RECT 1359.920 1470.685 1360.060 1517.770 ;
        RECT 1359.850 1470.315 1360.130 1470.685 ;
        RECT 1358.930 1469.635 1359.210 1470.005 ;
        RECT 1359.000 1421.530 1359.140 1469.635 ;
        RECT 1358.940 1421.210 1359.200 1421.530 ;
        RECT 1359.860 1421.210 1360.120 1421.530 ;
        RECT 1359.920 1374.125 1360.060 1421.210 ;
        RECT 1359.850 1373.755 1360.130 1374.125 ;
        RECT 1358.930 1373.075 1359.210 1373.445 ;
        RECT 1359.000 1324.630 1359.140 1373.075 ;
        RECT 1358.020 1324.310 1358.280 1324.630 ;
        RECT 1358.940 1324.310 1359.200 1324.630 ;
        RECT 1358.080 1276.885 1358.220 1324.310 ;
        RECT 1358.010 1276.515 1358.290 1276.885 ;
        RECT 1358.930 1276.515 1359.210 1276.885 ;
        RECT 1359.000 1276.350 1359.140 1276.515 ;
        RECT 1357.100 1276.030 1357.360 1276.350 ;
        RECT 1358.940 1276.030 1359.200 1276.350 ;
        RECT 1357.160 1228.410 1357.300 1276.030 ;
        RECT 1357.100 1228.090 1357.360 1228.410 ;
        RECT 1357.560 1228.090 1357.820 1228.410 ;
        RECT 1357.620 1211.070 1357.760 1228.090 ;
        RECT 1357.560 1210.750 1357.820 1211.070 ;
        RECT 1358.940 1210.750 1359.200 1211.070 ;
        RECT 1359.000 1138.730 1359.140 1210.750 ;
        RECT 1359.000 1138.650 1359.600 1138.730 ;
        RECT 1358.480 1138.330 1358.740 1138.650 ;
        RECT 1359.000 1138.590 1359.660 1138.650 ;
        RECT 1359.400 1138.330 1359.660 1138.590 ;
        RECT 1358.540 1090.370 1358.680 1138.330 ;
        RECT 1359.460 1138.175 1359.600 1138.330 ;
        RECT 1358.480 1090.050 1358.740 1090.370 ;
        RECT 1359.860 1090.050 1360.120 1090.370 ;
        RECT 1359.920 1062.830 1360.060 1090.050 ;
        RECT 1357.560 1062.510 1357.820 1062.830 ;
        RECT 1359.860 1062.510 1360.120 1062.830 ;
        RECT 1357.620 1028.570 1357.760 1062.510 ;
        RECT 1357.160 1028.430 1357.760 1028.570 ;
        RECT 1354.800 1010.830 1355.060 1011.150 ;
        RECT 1354.340 1008.790 1354.600 1009.110 ;
        RECT 1353.880 1008.110 1354.140 1008.430 ;
        RECT 1352.500 1007.770 1352.760 1008.090 ;
        RECT 1354.860 1000.010 1355.000 1010.830 ;
        RECT 1357.160 1000.010 1357.300 1028.430 ;
        RECT 1358.940 1017.970 1359.200 1018.290 ;
        RECT 1359.000 1000.010 1359.140 1017.970 ;
        RECT 1365.900 1008.770 1366.040 2780.870 ;
        RECT 1372.280 1735.030 1372.540 1735.350 ;
        RECT 1369.980 1012.190 1370.240 1012.510 ;
        RECT 1361.240 1008.450 1361.500 1008.770 ;
        RECT 1365.840 1008.450 1366.100 1008.770 ;
        RECT 1368.140 1008.450 1368.400 1008.770 ;
        RECT 1361.300 1000.010 1361.440 1008.450 ;
        RECT 1368.200 1000.010 1368.340 1008.450 ;
        RECT 1370.040 1000.010 1370.180 1012.190 ;
        RECT 1372.340 1008.770 1372.480 1735.030 ;
        RECT 1372.800 1012.510 1372.940 2913.470 ;
        RECT 1379.180 2485.750 1379.440 2486.070 ;
        RECT 1378.260 1062.510 1378.520 1062.830 ;
        RECT 1372.740 1012.190 1373.000 1012.510 ;
        RECT 1372.280 1008.450 1372.540 1008.770 ;
        RECT 1376.420 1008.450 1376.680 1008.770 ;
        RECT 1376.480 1000.010 1376.620 1008.450 ;
        RECT 1378.320 1000.010 1378.460 1062.510 ;
        RECT 1379.240 1008.770 1379.380 2485.750 ;
        RECT 1379.700 1062.830 1379.840 2915.510 ;
        RECT 1405.860 2915.170 1406.120 2915.490 ;
        RECT 1405.920 2903.330 1406.060 2915.170 ;
        RECT 1405.920 2903.190 1406.520 2903.330 ;
        RECT 1406.380 2863.810 1406.520 2903.190 ;
        RECT 1406.320 2863.490 1406.580 2863.810 ;
        RECT 1406.320 2862.810 1406.580 2863.130 ;
        RECT 1406.380 2849.190 1406.520 2862.810 ;
        RECT 1405.400 2848.870 1405.660 2849.190 ;
        RECT 1406.320 2848.870 1406.580 2849.190 ;
        RECT 1405.460 2801.590 1405.600 2848.870 ;
        RECT 1405.400 2801.270 1405.660 2801.590 ;
        RECT 1406.320 2801.270 1406.580 2801.590 ;
        RECT 1406.380 2767.250 1406.520 2801.270 ;
        RECT 1406.320 2766.930 1406.580 2767.250 ;
        RECT 1406.780 2766.590 1407.040 2766.910 ;
        RECT 1406.840 2753.310 1406.980 2766.590 ;
        RECT 1406.320 2752.990 1406.580 2753.310 ;
        RECT 1406.780 2752.990 1407.040 2753.310 ;
        RECT 1406.380 2752.630 1406.520 2752.990 ;
        RECT 1405.400 2752.310 1405.660 2752.630 ;
        RECT 1406.320 2752.310 1406.580 2752.630 ;
        RECT 1405.460 2705.030 1405.600 2752.310 ;
        RECT 1405.400 2704.710 1405.660 2705.030 ;
        RECT 1406.320 2704.710 1406.580 2705.030 ;
        RECT 1406.380 2670.690 1406.520 2704.710 ;
        RECT 1406.320 2670.370 1406.580 2670.690 ;
        RECT 1406.780 2670.030 1407.040 2670.350 ;
        RECT 1406.840 2656.750 1406.980 2670.030 ;
        RECT 1406.320 2656.430 1406.580 2656.750 ;
        RECT 1406.780 2656.430 1407.040 2656.750 ;
        RECT 1406.380 2622.750 1406.520 2656.430 ;
        RECT 1406.320 2622.430 1406.580 2622.750 ;
        RECT 1406.320 2621.750 1406.580 2622.070 ;
        RECT 1406.380 2609.685 1406.520 2621.750 ;
        RECT 1406.310 2609.315 1406.590 2609.685 ;
        RECT 1400.340 2608.150 1400.600 2608.470 ;
        RECT 1406.770 2608.210 1407.050 2608.495 ;
        RECT 1393.440 2594.550 1393.700 2594.870 ;
        RECT 1386.540 2485.410 1386.800 2485.730 ;
        RECT 1379.640 1062.510 1379.900 1062.830 ;
        RECT 1386.600 1011.570 1386.740 2485.410 ;
        RECT 1384.760 1011.430 1386.740 1011.570 ;
        RECT 1379.180 1008.450 1379.440 1008.770 ;
        RECT 1384.760 1000.010 1384.900 1011.430 ;
        RECT 1386.530 1010.635 1386.810 1011.005 ;
        RECT 1386.600 1000.010 1386.740 1010.635 ;
        RECT 1393.500 1000.010 1393.640 2594.550 ;
        RECT 1400.400 1008.770 1400.540 2608.150 ;
        RECT 1406.380 2608.125 1407.050 2608.210 ;
        RECT 1406.380 2608.070 1406.980 2608.125 ;
        RECT 1406.380 2574.130 1406.520 2608.070 ;
        RECT 1413.680 2580.610 1413.940 2580.930 ;
        RECT 1406.320 2573.810 1406.580 2574.130 ;
        RECT 1406.780 2573.470 1407.040 2573.790 ;
        RECT 1406.840 2560.190 1406.980 2573.470 ;
        RECT 1406.320 2559.870 1406.580 2560.190 ;
        RECT 1406.780 2559.870 1407.040 2560.190 ;
        RECT 1406.380 2559.510 1406.520 2559.870 ;
        RECT 1405.400 2559.190 1405.660 2559.510 ;
        RECT 1406.320 2559.190 1406.580 2559.510 ;
        RECT 1405.460 2511.910 1405.600 2559.190 ;
        RECT 1405.400 2511.590 1405.660 2511.910 ;
        RECT 1406.320 2511.590 1406.580 2511.910 ;
        RECT 1406.380 2488.110 1406.520 2511.590 ;
        RECT 1405.400 2487.790 1405.660 2488.110 ;
        RECT 1406.320 2487.790 1406.580 2488.110 ;
        RECT 1405.460 2463.485 1405.600 2487.790 ;
        RECT 1405.390 2463.115 1405.670 2463.485 ;
        RECT 1406.310 2463.115 1406.590 2463.485 ;
        RECT 1406.380 2429.630 1406.520 2463.115 ;
        RECT 1406.320 2429.310 1406.580 2429.630 ;
        RECT 1406.320 2428.630 1406.580 2428.950 ;
        RECT 1406.380 2380.670 1406.520 2428.630 ;
        RECT 1406.320 2380.350 1406.580 2380.670 ;
        RECT 1406.780 2380.350 1407.040 2380.670 ;
        RECT 1406.840 2367.070 1406.980 2380.350 ;
        RECT 1406.320 2366.750 1406.580 2367.070 ;
        RECT 1406.780 2366.750 1407.040 2367.070 ;
        RECT 1406.380 2332.730 1406.520 2366.750 ;
        RECT 1406.320 2332.410 1406.580 2332.730 ;
        RECT 1406.320 2331.730 1406.580 2332.050 ;
        RECT 1406.380 2294.310 1406.520 2331.730 ;
        RECT 1405.400 2293.990 1405.660 2294.310 ;
        RECT 1406.320 2293.990 1406.580 2294.310 ;
        RECT 1405.460 2270.365 1405.600 2293.990 ;
        RECT 1405.390 2269.995 1405.670 2270.365 ;
        RECT 1406.310 2269.995 1406.590 2270.365 ;
        RECT 1406.380 2236.170 1406.520 2269.995 ;
        RECT 1406.320 2235.850 1406.580 2236.170 ;
        RECT 1406.320 2235.170 1406.580 2235.490 ;
        RECT 1406.380 2197.750 1406.520 2235.170 ;
        RECT 1405.400 2197.430 1405.660 2197.750 ;
        RECT 1406.320 2197.430 1406.580 2197.750 ;
        RECT 1405.460 2173.805 1405.600 2197.430 ;
        RECT 1405.390 2173.435 1405.670 2173.805 ;
        RECT 1406.310 2173.435 1406.590 2173.805 ;
        RECT 1406.380 2139.610 1406.520 2173.435 ;
        RECT 1406.320 2139.290 1406.580 2139.610 ;
        RECT 1406.320 2138.610 1406.580 2138.930 ;
        RECT 1406.380 2118.190 1406.520 2138.610 ;
        RECT 1406.320 2117.870 1406.580 2118.190 ;
        RECT 1407.700 2117.870 1407.960 2118.190 ;
        RECT 1407.760 2070.330 1407.900 2117.870 ;
        RECT 1407.760 2070.190 1408.360 2070.330 ;
        RECT 1408.220 2069.910 1408.360 2070.190 ;
        RECT 1408.160 2069.590 1408.420 2069.910 ;
        RECT 1409.080 2069.590 1409.340 2069.910 ;
        RECT 1409.140 2024.770 1409.280 2069.590 ;
        RECT 1408.220 2024.630 1409.280 2024.770 ;
        RECT 1408.220 1980.685 1408.360 2024.630 ;
        RECT 1408.150 1980.315 1408.430 1980.685 ;
        RECT 1408.150 1979.635 1408.430 1980.005 ;
        RECT 1408.220 1932.290 1408.360 1979.635 ;
        RECT 1406.840 1932.150 1408.360 1932.290 ;
        RECT 1406.840 1931.870 1406.980 1932.150 ;
        RECT 1406.780 1931.550 1407.040 1931.870 ;
        RECT 1407.700 1931.550 1407.960 1931.870 ;
        RECT 1407.760 1884.270 1407.900 1931.550 ;
        RECT 1405.860 1883.950 1406.120 1884.270 ;
        RECT 1407.700 1883.950 1407.960 1884.270 ;
        RECT 1405.920 1883.590 1406.060 1883.950 ;
        RECT 1405.400 1883.270 1405.660 1883.590 ;
        RECT 1405.860 1883.270 1406.120 1883.590 ;
        RECT 1405.460 1835.990 1405.600 1883.270 ;
        RECT 1405.400 1835.670 1405.660 1835.990 ;
        RECT 1406.780 1835.670 1407.040 1835.990 ;
        RECT 1406.840 1835.310 1406.980 1835.670 ;
        RECT 1405.400 1834.990 1405.660 1835.310 ;
        RECT 1406.780 1834.990 1407.040 1835.310 ;
        RECT 1405.460 1787.710 1405.600 1834.990 ;
        RECT 1405.400 1787.390 1405.660 1787.710 ;
        RECT 1405.860 1787.390 1406.120 1787.710 ;
        RECT 1405.920 1787.030 1406.060 1787.390 ;
        RECT 1405.400 1786.710 1405.660 1787.030 ;
        RECT 1405.860 1786.710 1406.120 1787.030 ;
        RECT 1405.460 1739.430 1405.600 1786.710 ;
        RECT 1405.400 1739.110 1405.660 1739.430 ;
        RECT 1406.780 1739.110 1407.040 1739.430 ;
        RECT 1406.840 1738.750 1406.980 1739.110 ;
        RECT 1405.400 1738.430 1405.660 1738.750 ;
        RECT 1406.780 1738.430 1407.040 1738.750 ;
        RECT 1405.460 1690.810 1405.600 1738.430 ;
        RECT 1405.400 1690.490 1405.660 1690.810 ;
        RECT 1406.320 1690.490 1406.580 1690.810 ;
        RECT 1406.380 1690.210 1406.520 1690.490 ;
        RECT 1405.920 1690.070 1406.520 1690.210 ;
        RECT 1405.920 1642.530 1406.060 1690.070 ;
        RECT 1405.860 1642.210 1406.120 1642.530 ;
        RECT 1406.320 1642.210 1406.580 1642.530 ;
        RECT 1406.380 1607.850 1406.520 1642.210 ;
        RECT 1406.320 1607.530 1406.580 1607.850 ;
        RECT 1406.780 1607.530 1407.040 1607.850 ;
        RECT 1406.840 1593.910 1406.980 1607.530 ;
        RECT 1405.400 1593.590 1405.660 1593.910 ;
        RECT 1406.780 1593.590 1407.040 1593.910 ;
        RECT 1405.460 1545.970 1405.600 1593.590 ;
        RECT 1405.400 1545.650 1405.660 1545.970 ;
        RECT 1406.320 1545.650 1406.580 1545.970 ;
        RECT 1406.380 1511.290 1406.520 1545.650 ;
        RECT 1406.320 1510.970 1406.580 1511.290 ;
        RECT 1406.780 1510.630 1407.040 1510.950 ;
        RECT 1406.840 1497.350 1406.980 1510.630 ;
        RECT 1405.400 1497.030 1405.660 1497.350 ;
        RECT 1406.780 1497.030 1407.040 1497.350 ;
        RECT 1405.460 1449.410 1405.600 1497.030 ;
        RECT 1405.400 1449.090 1405.660 1449.410 ;
        RECT 1406.320 1449.090 1406.580 1449.410 ;
        RECT 1406.380 1414.730 1406.520 1449.090 ;
        RECT 1406.320 1414.410 1406.580 1414.730 ;
        RECT 1406.780 1414.070 1407.040 1414.390 ;
        RECT 1406.840 1400.790 1406.980 1414.070 ;
        RECT 1406.780 1400.470 1407.040 1400.790 ;
        RECT 1408.160 1400.470 1408.420 1400.790 ;
        RECT 1408.220 1353.190 1408.360 1400.470 ;
        RECT 1406.780 1352.870 1407.040 1353.190 ;
        RECT 1408.160 1352.870 1408.420 1353.190 ;
        RECT 1406.840 1352.510 1406.980 1352.870 ;
        RECT 1405.400 1352.190 1405.660 1352.510 ;
        RECT 1406.780 1352.190 1407.040 1352.510 ;
        RECT 1405.460 1304.570 1405.600 1352.190 ;
        RECT 1405.400 1304.250 1405.660 1304.570 ;
        RECT 1406.320 1304.250 1406.580 1304.570 ;
        RECT 1405.850 1303.970 1406.130 1304.085 ;
        RECT 1406.380 1303.970 1406.520 1304.250 ;
        RECT 1405.850 1303.830 1406.520 1303.970 ;
        RECT 1405.850 1303.715 1406.130 1303.830 ;
        RECT 1405.390 1255.435 1405.670 1255.805 ;
        RECT 1405.460 1207.670 1405.600 1255.435 ;
        RECT 1405.400 1207.350 1405.660 1207.670 ;
        RECT 1406.320 1207.350 1406.580 1207.670 ;
        RECT 1406.380 1206.990 1406.520 1207.350 ;
        RECT 1405.400 1206.670 1405.660 1206.990 ;
        RECT 1406.320 1206.670 1406.580 1206.990 ;
        RECT 1405.460 1159.390 1405.600 1206.670 ;
        RECT 1405.400 1159.070 1405.660 1159.390 ;
        RECT 1406.320 1159.070 1406.580 1159.390 ;
        RECT 1406.380 1135.330 1406.520 1159.070 ;
        RECT 1405.460 1135.190 1406.520 1135.330 ;
        RECT 1405.460 1111.110 1405.600 1135.190 ;
        RECT 1405.400 1110.790 1405.660 1111.110 ;
        RECT 1405.860 1110.790 1406.120 1111.110 ;
        RECT 1405.920 1076.770 1406.060 1110.790 ;
        RECT 1405.860 1076.450 1406.120 1076.770 ;
        RECT 1406.320 1075.770 1406.580 1076.090 ;
        RECT 1402.640 1017.630 1402.900 1017.950 ;
        RECT 1396.200 1008.450 1396.460 1008.770 ;
        RECT 1400.340 1008.450 1400.600 1008.770 ;
        RECT 1396.260 1000.010 1396.400 1008.450 ;
        RECT 1402.700 1000.010 1402.840 1017.630 ;
        RECT 1406.380 1012.510 1406.520 1075.770 ;
        RECT 1413.740 1012.510 1413.880 2580.610 ;
        RECT 1404.940 1012.190 1405.200 1012.510 ;
        RECT 1406.320 1012.190 1406.580 1012.510 ;
        RECT 1411.380 1012.190 1411.640 1012.510 ;
        RECT 1413.680 1012.190 1413.940 1012.510 ;
        RECT 1405.000 1000.010 1405.140 1012.190 ;
        RECT 1411.440 1000.010 1411.580 1012.190 ;
        RECT 1414.200 1000.690 1414.340 2917.550 ;
        RECT 1448.640 2915.850 1448.900 2916.170 ;
        RECT 1434.840 2691.110 1435.100 2691.430 ;
        RECT 1421.040 2488.470 1421.300 2488.790 ;
        RECT 1420.580 2487.790 1420.840 2488.110 ;
        RECT 1419.660 1012.870 1419.920 1013.190 ;
        RECT 1417.820 1010.490 1418.080 1010.810 ;
        RECT 1413.740 1000.550 1414.340 1000.690 ;
        RECT 1413.740 1000.010 1413.880 1000.550 ;
        RECT 1417.880 1000.010 1418.020 1010.490 ;
        RECT 1419.720 1000.010 1419.860 1012.870 ;
        RECT 1348.880 1000.000 1349.180 1000.010 ;
        RECT 1351.480 1000.000 1352.240 1000.010 ;
        RECT 1353.320 1000.000 1355.000 1000.010 ;
        RECT 1355.620 1000.000 1357.300 1000.010 ;
        RECT 1357.920 1000.000 1359.140 1000.010 ;
        RECT 1360.220 1000.000 1361.440 1000.010 ;
        RECT 1366.660 1000.000 1368.340 1000.010 ;
        RECT 1368.960 1000.000 1370.180 1000.010 ;
        RECT 1375.400 1000.000 1376.620 1000.010 ;
        RECT 1377.240 1000.000 1378.460 1000.010 ;
        RECT 1384.140 1000.000 1384.900 1000.010 ;
        RECT 1385.980 1000.000 1386.740 1000.010 ;
        RECT 1392.880 1000.000 1393.640 1000.010 ;
        RECT 1394.720 1000.000 1396.400 1000.010 ;
        RECT 1401.160 1000.000 1402.840 1000.010 ;
        RECT 1403.460 1000.000 1405.140 1000.010 ;
        RECT 1409.900 1000.000 1411.580 1000.010 ;
        RECT 1412.200 1000.000 1413.880 1000.010 ;
        RECT 1416.800 1000.000 1418.020 1000.010 ;
        RECT 1418.640 1000.000 1419.860 1000.010 ;
        RECT 1348.880 999.870 1349.330 1000.000 ;
      LAYER met2 ;
        RECT 1345.470 995.720 1346.470 998.810 ;
      LAYER met2 ;
        RECT 1346.750 996.000 1347.030 999.870 ;
      LAYER met2 ;
        RECT 1347.310 995.720 1348.770 998.810 ;
      LAYER met2 ;
        RECT 1349.050 996.000 1349.330 999.870 ;
        RECT 1351.350 999.870 1352.240 1000.000 ;
        RECT 1353.190 999.870 1355.000 1000.000 ;
        RECT 1355.490 999.870 1357.300 1000.000 ;
        RECT 1357.790 999.870 1359.140 1000.000 ;
        RECT 1360.090 999.870 1361.440 1000.000 ;
      LAYER met2 ;
        RECT 1349.610 995.720 1351.070 998.810 ;
      LAYER met2 ;
        RECT 1351.350 996.000 1351.630 999.870 ;
      LAYER met2 ;
        RECT 1351.910 995.720 1352.910 998.810 ;
      LAYER met2 ;
        RECT 1353.190 996.000 1353.470 999.870 ;
      LAYER met2 ;
        RECT 1353.750 995.720 1355.210 998.810 ;
      LAYER met2 ;
        RECT 1355.490 996.000 1355.770 999.870 ;
      LAYER met2 ;
        RECT 1356.050 995.720 1357.510 998.810 ;
      LAYER met2 ;
        RECT 1357.790 996.000 1358.070 999.870 ;
      LAYER met2 ;
        RECT 1358.350 995.720 1359.810 998.810 ;
      LAYER met2 ;
        RECT 1360.090 996.000 1360.370 999.870 ;
      LAYER met2 ;
        RECT 1360.650 995.720 1361.650 998.810 ;
      LAYER met2 ;
        RECT 1361.930 996.000 1362.210 1000.000 ;
      LAYER met2 ;
        RECT 1362.490 995.720 1363.950 998.810 ;
      LAYER met2 ;
        RECT 1364.230 996.000 1364.510 1000.000 ;
        RECT 1366.530 999.870 1368.340 1000.000 ;
        RECT 1368.830 999.870 1370.180 1000.000 ;
      LAYER met2 ;
        RECT 1364.790 995.720 1366.250 998.810 ;
      LAYER met2 ;
        RECT 1366.530 996.000 1366.810 999.870 ;
      LAYER met2 ;
        RECT 1367.090 995.720 1368.550 998.810 ;
      LAYER met2 ;
        RECT 1368.830 996.000 1369.110 999.870 ;
      LAYER met2 ;
        RECT 1369.390 995.720 1370.390 998.810 ;
      LAYER met2 ;
        RECT 1370.670 996.000 1370.950 1000.000 ;
      LAYER met2 ;
        RECT 1371.230 995.720 1372.690 998.810 ;
      LAYER met2 ;
        RECT 1372.970 996.000 1373.250 1000.000 ;
        RECT 1375.270 999.870 1376.620 1000.000 ;
        RECT 1377.110 999.870 1378.460 1000.000 ;
      LAYER met2 ;
        RECT 1373.530 995.720 1374.990 998.810 ;
      LAYER met2 ;
        RECT 1375.270 996.000 1375.550 999.870 ;
      LAYER met2 ;
        RECT 1375.830 995.720 1376.830 998.810 ;
      LAYER met2 ;
        RECT 1377.110 996.000 1377.390 999.870 ;
      LAYER met2 ;
        RECT 1377.670 995.720 1379.130 998.810 ;
      LAYER met2 ;
        RECT 1379.410 996.000 1379.690 1000.000 ;
      LAYER met2 ;
        RECT 1379.970 995.720 1381.430 998.810 ;
      LAYER met2 ;
        RECT 1381.710 996.000 1381.990 1000.000 ;
        RECT 1384.010 999.870 1384.900 1000.000 ;
        RECT 1385.850 999.870 1386.740 1000.000 ;
      LAYER met2 ;
        RECT 1382.270 995.720 1383.730 998.810 ;
      LAYER met2 ;
        RECT 1384.010 996.000 1384.290 999.870 ;
      LAYER met2 ;
        RECT 1384.570 995.720 1385.570 998.810 ;
      LAYER met2 ;
        RECT 1385.850 996.000 1386.130 999.870 ;
      LAYER met2 ;
        RECT 1386.410 995.720 1387.870 998.810 ;
      LAYER met2 ;
        RECT 1388.150 996.000 1388.430 1000.000 ;
      LAYER met2 ;
        RECT 1388.710 995.720 1390.170 998.810 ;
      LAYER met2 ;
        RECT 1390.450 996.000 1390.730 1000.000 ;
        RECT 1392.750 999.870 1393.640 1000.000 ;
        RECT 1394.590 999.870 1396.400 1000.000 ;
      LAYER met2 ;
        RECT 1391.010 995.720 1392.470 998.810 ;
      LAYER met2 ;
        RECT 1392.750 996.000 1393.030 999.870 ;
      LAYER met2 ;
        RECT 1393.310 995.720 1394.310 998.810 ;
      LAYER met2 ;
        RECT 1394.590 996.000 1394.870 999.870 ;
      LAYER met2 ;
        RECT 1395.150 995.720 1396.610 998.810 ;
      LAYER met2 ;
        RECT 1396.890 996.000 1397.170 1000.000 ;
      LAYER met2 ;
        RECT 1397.450 995.720 1398.910 998.810 ;
      LAYER met2 ;
        RECT 1399.190 996.000 1399.470 1000.000 ;
        RECT 1401.030 999.870 1402.840 1000.000 ;
        RECT 1403.330 999.870 1405.140 1000.000 ;
      LAYER met2 ;
        RECT 1399.750 995.720 1400.750 998.810 ;
      LAYER met2 ;
        RECT 1401.030 996.000 1401.310 999.870 ;
      LAYER met2 ;
        RECT 1401.590 995.720 1403.050 998.810 ;
      LAYER met2 ;
        RECT 1403.330 996.000 1403.610 999.870 ;
      LAYER met2 ;
        RECT 1403.890 995.720 1405.350 998.810 ;
      LAYER met2 ;
        RECT 1405.630 996.000 1405.910 1000.000 ;
      LAYER met2 ;
        RECT 1406.190 995.720 1407.650 998.810 ;
      LAYER met2 ;
        RECT 1407.930 996.000 1408.210 1000.000 ;
        RECT 1409.770 999.870 1411.580 1000.000 ;
        RECT 1412.070 999.870 1413.880 1000.000 ;
      LAYER met2 ;
        RECT 1408.490 995.720 1409.490 998.810 ;
      LAYER met2 ;
        RECT 1409.770 996.000 1410.050 999.870 ;
      LAYER met2 ;
        RECT 1410.330 995.720 1411.790 998.810 ;
      LAYER met2 ;
        RECT 1412.070 996.000 1412.350 999.870 ;
      LAYER met2 ;
        RECT 1412.630 995.720 1414.090 998.810 ;
      LAYER met2 ;
        RECT 1414.370 996.000 1414.650 1000.000 ;
        RECT 1416.670 999.870 1418.020 1000.000 ;
        RECT 1418.510 999.870 1419.860 1000.000 ;
        RECT 1420.640 1000.010 1420.780 2487.790 ;
        RECT 1421.100 1013.190 1421.240 2488.470 ;
        RECT 1427.940 2486.430 1428.200 2486.750 ;
        RECT 1421.040 1012.870 1421.300 1013.190 ;
        RECT 1428.000 1000.010 1428.140 2486.430 ;
        RECT 1431.160 1024.430 1431.420 1024.750 ;
        RECT 1431.220 1000.010 1431.360 1024.430 ;
        RECT 1434.900 1000.010 1435.040 2691.110 ;
        RECT 1448.180 2486.770 1448.440 2487.090 ;
        RECT 1441.280 2485.070 1441.540 2485.390 ;
        RECT 1441.340 1076.170 1441.480 2485.070 ;
        RECT 1440.420 1076.030 1441.480 1076.170 ;
        RECT 1440.420 1028.570 1440.560 1076.030 ;
        RECT 1439.960 1028.430 1440.560 1028.570 ;
        RECT 1437.600 1018.310 1437.860 1018.630 ;
        RECT 1437.660 1000.010 1437.800 1018.310 ;
        RECT 1439.960 1000.010 1440.100 1028.430 ;
        RECT 1446.340 1013.890 1446.600 1014.210 ;
        RECT 1444.040 1012.190 1444.300 1012.510 ;
        RECT 1444.100 1000.010 1444.240 1012.190 ;
        RECT 1446.400 1000.010 1446.540 1013.890 ;
        RECT 1448.240 1000.010 1448.380 2486.770 ;
        RECT 1448.700 1014.210 1448.840 2915.850 ;
        RECT 1469.340 2914.830 1469.600 2915.150 ;
        RECT 1455.540 2913.810 1455.800 2914.130 ;
        RECT 1455.080 2488.130 1455.340 2488.450 ;
        RECT 1454.620 1051.970 1454.880 1052.290 ;
        RECT 1448.640 1013.890 1448.900 1014.210 ;
        RECT 1452.780 1013.890 1453.040 1014.210 ;
        RECT 1452.840 1000.010 1452.980 1013.890 ;
        RECT 1454.680 1000.690 1454.820 1051.970 ;
        RECT 1455.140 1014.210 1455.280 2488.130 ;
        RECT 1455.600 1052.290 1455.740 2913.810 ;
        RECT 1468.880 2546.270 1469.140 2546.590 ;
        RECT 1461.980 2486.090 1462.240 2486.410 ;
        RECT 1455.540 1051.970 1455.800 1052.290 ;
        RECT 1462.040 1014.210 1462.180 2486.090 ;
        RECT 1462.440 1018.650 1462.700 1018.970 ;
        RECT 1455.080 1013.890 1455.340 1014.210 ;
        RECT 1456.920 1013.890 1457.180 1014.210 ;
        RECT 1461.980 1013.890 1462.240 1014.210 ;
        RECT 1454.680 1000.550 1455.280 1000.690 ;
        RECT 1455.140 1000.010 1455.280 1000.550 ;
        RECT 1456.980 1000.010 1457.120 1013.890 ;
        RECT 1461.520 1011.170 1461.780 1011.490 ;
        RECT 1461.580 1000.010 1461.720 1011.170 ;
        RECT 1462.500 1000.010 1462.640 1018.650 ;
        RECT 1465.660 1013.890 1465.920 1014.210 ;
        RECT 1465.720 1000.010 1465.860 1013.890 ;
        RECT 1468.940 1000.010 1469.080 2546.270 ;
        RECT 1469.400 1014.210 1469.540 2914.830 ;
        RECT 1502.000 2914.490 1502.260 2914.810 ;
        RECT 1494.640 2913.130 1494.900 2913.450 ;
        RECT 1493.720 2912.110 1493.980 2912.430 ;
        RECT 1490.040 2894.090 1490.300 2894.410 ;
        RECT 1483.590 2850.035 1483.870 2850.405 ;
        RECT 1483.660 2849.870 1483.800 2850.035 ;
        RECT 1483.600 2849.550 1483.860 2849.870 ;
        RECT 1482.210 2830.315 1482.490 2830.685 ;
        RECT 1474.400 1024.770 1474.660 1025.090 ;
        RECT 1472.100 1016.950 1472.360 1017.270 ;
        RECT 1469.340 1013.890 1469.600 1014.210 ;
        RECT 1472.160 1000.010 1472.300 1016.950 ;
        RECT 1474.460 1000.010 1474.600 1024.770 ;
        RECT 1480.840 1017.290 1481.100 1017.610 ;
        RECT 1479.000 1013.890 1479.260 1014.210 ;
        RECT 1479.060 1000.010 1479.200 1013.890 ;
        RECT 1480.900 1000.010 1481.040 1017.290 ;
        RECT 1482.280 1014.210 1482.420 2830.315 ;
        RECT 1489.570 2801.755 1489.850 2802.125 ;
        RECT 1489.110 2784.075 1489.390 2784.445 ;
        RECT 1489.180 2781.190 1489.320 2784.075 ;
        RECT 1489.120 2780.870 1489.380 2781.190 ;
        RECT 1489.110 2767.755 1489.390 2768.125 ;
        RECT 1488.650 2753.475 1488.930 2753.845 ;
        RECT 1488.190 2691.595 1488.470 2691.965 ;
        RECT 1488.260 2691.430 1488.400 2691.595 ;
        RECT 1488.200 2691.110 1488.460 2691.430 ;
        RECT 1488.190 2673.915 1488.470 2674.285 ;
        RECT 1482.670 2657.595 1482.950 2657.965 ;
        RECT 1482.220 1013.890 1482.480 1014.210 ;
        RECT 1482.740 1000.010 1482.880 2657.595 ;
        RECT 1487.270 2629.035 1487.550 2629.405 ;
        RECT 1487.340 2607.530 1487.480 2629.035 ;
        RECT 1487.730 2609.995 1488.010 2610.365 ;
        RECT 1487.800 2608.470 1487.940 2609.995 ;
        RECT 1487.740 2608.150 1488.000 2608.470 ;
        RECT 1487.340 2607.390 1487.940 2607.530 ;
        RECT 1487.270 2595.035 1487.550 2595.405 ;
        RECT 1487.340 2594.870 1487.480 2595.035 ;
        RECT 1487.280 2594.550 1487.540 2594.870 ;
        RECT 1487.270 2580.755 1487.550 2581.125 ;
        RECT 1487.280 2580.610 1487.540 2580.755 ;
        RECT 1487.270 2567.155 1487.550 2567.525 ;
        RECT 1483.590 2547.435 1483.870 2547.805 ;
        RECT 1483.660 2546.590 1483.800 2547.435 ;
        RECT 1483.600 2546.270 1483.860 2546.590 ;
        RECT 1485.900 2525.190 1486.160 2525.510 ;
        RECT 1485.960 2477.570 1486.100 2525.190 ;
        RECT 1486.810 2518.875 1487.090 2519.245 ;
        RECT 1485.900 2477.250 1486.160 2477.570 ;
        RECT 1485.900 1945.490 1486.160 1945.810 ;
        RECT 1485.960 1897.870 1486.100 1945.490 ;
        RECT 1485.900 1897.550 1486.160 1897.870 ;
        RECT 1486.360 1076.110 1486.620 1076.430 ;
        RECT 1486.420 1028.490 1486.560 1076.110 ;
        RECT 1486.360 1028.170 1486.620 1028.490 ;
        RECT 1486.360 1009.130 1486.620 1009.450 ;
        RECT 1486.420 1000.010 1486.560 1009.130 ;
        RECT 1486.880 1008.430 1487.020 2518.875 ;
        RECT 1487.340 1010.470 1487.480 2567.155 ;
        RECT 1487.800 1011.830 1487.940 2607.390 ;
        RECT 1487.740 1011.510 1488.000 1011.830 ;
        RECT 1487.280 1010.150 1487.540 1010.470 ;
        RECT 1486.820 1008.110 1487.080 1008.430 ;
        RECT 1488.260 1007.750 1488.400 2673.915 ;
        RECT 1488.720 1052.290 1488.860 2753.475 ;
        RECT 1489.180 1055.690 1489.320 2767.755 ;
        RECT 1489.120 1055.370 1489.380 1055.690 ;
        RECT 1488.660 1051.970 1488.920 1052.290 ;
        RECT 1489.120 1028.170 1489.380 1028.490 ;
        RECT 1488.200 1007.430 1488.460 1007.750 ;
        RECT 1489.180 1000.690 1489.320 1028.170 ;
        RECT 1489.640 1016.590 1489.780 2801.755 ;
        RECT 1490.100 2525.510 1490.240 2894.090 ;
        RECT 1490.040 2525.190 1490.300 2525.510 ;
        RECT 1490.040 2477.250 1490.300 2477.570 ;
        RECT 1490.100 1945.810 1490.240 2477.250 ;
        RECT 1490.040 1945.490 1490.300 1945.810 ;
        RECT 1490.040 1897.550 1490.300 1897.870 ;
        RECT 1490.100 1076.430 1490.240 1897.550 ;
        RECT 1490.040 1076.110 1490.300 1076.430 ;
        RECT 1489.580 1016.270 1489.840 1016.590 ;
        RECT 1491.880 1008.450 1492.140 1008.770 ;
        RECT 1489.180 1000.550 1489.780 1000.690 ;
        RECT 1489.640 1000.010 1489.780 1000.550 ;
        RECT 1491.940 1000.010 1492.080 1008.450 ;
        RECT 1493.780 1008.090 1493.920 2912.110 ;
        RECT 1494.180 2911.770 1494.440 2912.090 ;
        RECT 1494.240 2497.290 1494.380 2911.770 ;
        RECT 1494.180 2496.970 1494.440 2497.290 ;
        RECT 1494.700 2495.250 1494.840 2913.130 ;
        RECT 1501.540 2912.790 1501.800 2913.110 ;
        RECT 1496.480 2912.450 1496.740 2912.770 ;
        RECT 1496.020 2898.170 1496.280 2898.490 ;
        RECT 1495.550 2739.195 1495.830 2739.565 ;
        RECT 1495.090 2720.155 1495.370 2720.525 ;
        RECT 1494.640 2494.930 1494.900 2495.250 ;
        RECT 1495.160 1013.190 1495.300 2720.155 ;
        RECT 1495.620 1013.530 1495.760 2739.195 ;
        RECT 1495.560 1013.210 1495.820 1013.530 ;
        RECT 1495.100 1012.870 1495.360 1013.190 ;
        RECT 1496.080 1012.170 1496.220 2898.170 ;
        RECT 1496.540 1012.850 1496.680 2912.450 ;
        RECT 1497.400 2896.470 1497.660 2896.790 ;
        RECT 1496.940 1018.990 1497.200 1019.310 ;
        RECT 1496.480 1012.530 1496.740 1012.850 ;
        RECT 1496.020 1011.850 1496.280 1012.170 ;
        RECT 1496.020 1009.470 1496.280 1009.790 ;
        RECT 1493.720 1007.770 1493.980 1008.090 ;
        RECT 1496.080 1000.010 1496.220 1009.470 ;
        RECT 1497.000 1000.010 1497.140 1018.990 ;
        RECT 1497.460 1013.870 1497.600 2896.470 ;
        RECT 1501.600 2494.910 1501.740 2912.790 ;
        RECT 1501.540 2494.590 1501.800 2494.910 ;
        RECT 1500.620 1013.890 1500.880 1014.210 ;
        RECT 1497.400 1013.550 1497.660 1013.870 ;
        RECT 1500.680 1000.010 1500.820 1013.890 ;
        RECT 1502.060 1009.110 1502.200 2914.490 ;
        RECT 1502.460 2914.150 1502.720 2914.470 ;
        RECT 1502.520 1010.130 1502.660 2914.150 ;
        RECT 1535.180 2900.055 1535.320 2917.890 ;
        RECT 1567.320 2917.550 1567.580 2917.870 ;
        RECT 1546.160 2911.770 1546.420 2912.090 ;
        RECT 1546.220 2900.055 1546.360 2911.770 ;
        RECT 1567.380 2900.055 1567.520 2917.550 ;
        RECT 1641.840 2915.850 1642.100 2916.170 ;
        RECT 1598.600 2915.510 1598.860 2915.830 ;
        RECT 1598.660 2900.055 1598.800 2915.510 ;
        RECT 1630.800 2915.170 1631.060 2915.490 ;
        RECT 1609.640 2912.110 1609.900 2912.430 ;
        RECT 1609.700 2900.055 1609.840 2912.110 ;
        RECT 1630.860 2900.055 1631.000 2915.170 ;
        RECT 1641.900 2900.055 1642.040 2915.850 ;
        RECT 1694.280 2914.830 1694.540 2915.150 ;
        RECT 1663.000 2912.450 1663.260 2912.770 ;
        RECT 1663.060 2900.055 1663.200 2912.450 ;
        RECT 1694.340 2900.055 1694.480 2914.830 ;
        RECT 1768.800 2914.490 1769.060 2914.810 ;
        RECT 1758.680 2913.810 1758.940 2914.130 ;
        RECT 1705.320 2913.130 1705.580 2913.450 ;
        RECT 1705.380 2900.055 1705.520 2913.130 ;
        RECT 1758.740 2900.055 1758.880 2913.810 ;
        RECT 1768.860 2900.055 1769.000 2914.490 ;
        RECT 1779.840 2914.150 1780.100 2914.470 ;
        RECT 1779.900 2900.055 1780.040 2914.150 ;
        RECT 1843.320 2913.470 1843.580 2913.790 ;
        RECT 1789.960 2913.130 1790.220 2913.450 ;
        RECT 1790.020 2900.055 1790.160 2913.130 ;
        RECT 1812.040 2912.790 1812.300 2913.110 ;
        RECT 1833.200 2912.790 1833.460 2913.110 ;
        RECT 1812.100 2900.055 1812.240 2912.790 ;
        RECT 1833.260 2900.055 1833.400 2912.790 ;
        RECT 1843.380 2900.055 1843.520 2913.470 ;
        RECT 1895.300 2913.130 1895.560 2913.450 ;
        RECT 1887.940 2912.790 1888.200 2913.110 ;
        RECT 1854.360 2912.450 1854.620 2912.770 ;
        RECT 1886.560 2912.450 1886.820 2912.770 ;
        RECT 1854.420 2900.055 1854.560 2912.450 ;
        RECT 1864.480 2912.110 1864.740 2912.430 ;
        RECT 1864.540 2900.055 1864.680 2912.110 ;
        RECT 1502.850 2896.530 1503.130 2900.055 ;
        RECT 1524.930 2898.570 1525.210 2900.055 ;
        RECT 1524.140 2898.490 1525.210 2898.570 ;
        RECT 1524.080 2898.430 1525.210 2898.490 ;
        RECT 1524.080 2898.170 1524.340 2898.430 ;
        RECT 1503.380 2896.530 1503.640 2896.790 ;
        RECT 1502.850 2896.470 1503.640 2896.530 ;
        RECT 1502.850 2896.390 1503.580 2896.470 ;
        RECT 1502.850 2896.055 1503.130 2896.390 ;
        RECT 1524.930 2896.055 1525.210 2898.430 ;
        RECT 1535.050 2896.055 1535.330 2900.055 ;
        RECT 1546.090 2896.055 1546.370 2900.055 ;
        RECT 1567.250 2896.055 1567.530 2900.055 ;
        RECT 1598.530 2896.055 1598.810 2900.055 ;
        RECT 1609.570 2896.055 1609.850 2900.055 ;
        RECT 1630.730 2896.055 1631.010 2900.055 ;
        RECT 1641.770 2896.055 1642.050 2900.055 ;
        RECT 1652.880 2897.150 1653.140 2897.470 ;
        RECT 1652.940 2896.790 1653.080 2897.150 ;
        RECT 1652.880 2896.470 1653.140 2896.790 ;
        RECT 1662.930 2896.055 1663.210 2900.055 ;
        RECT 1693.360 2897.150 1693.620 2897.470 ;
        RECT 1693.420 2896.790 1693.560 2897.150 ;
        RECT 1693.360 2896.470 1693.620 2896.790 ;
        RECT 1694.210 2896.055 1694.490 2900.055 ;
        RECT 1705.250 2896.055 1705.530 2900.055 ;
        RECT 1758.610 2896.055 1758.890 2900.055 ;
        RECT 1768.730 2896.055 1769.010 2900.055 ;
        RECT 1779.770 2896.055 1780.050 2900.055 ;
        RECT 1789.890 2896.055 1790.170 2900.055 ;
        RECT 1800.930 2896.530 1801.210 2900.055 ;
        RECT 1801.920 2896.530 1802.180 2896.790 ;
        RECT 1800.930 2896.470 1802.180 2896.530 ;
        RECT 1800.930 2896.390 1802.120 2896.470 ;
        RECT 1800.930 2896.055 1801.210 2896.390 ;
        RECT 1811.970 2896.055 1812.250 2900.055 ;
        RECT 1833.130 2896.055 1833.410 2900.055 ;
        RECT 1843.250 2896.055 1843.530 2900.055 ;
        RECT 1854.290 2896.055 1854.570 2900.055 ;
        RECT 1864.410 2896.055 1864.690 2900.055 ;
        RECT 1875.450 2896.530 1875.730 2900.055 ;
        RECT 1876.900 2896.530 1877.160 2896.790 ;
        RECT 1875.450 2896.470 1877.160 2896.530 ;
        RECT 1885.570 2896.530 1885.850 2900.055 ;
        RECT 1875.450 2896.390 1877.100 2896.470 ;
        RECT 1885.570 2896.390 1886.300 2896.530 ;
        RECT 1875.450 2896.055 1875.730 2896.390 ;
        RECT 1885.570 2896.055 1885.850 2896.390 ;
      LAYER met2 ;
        RECT 1503.410 2895.775 1513.610 2896.055 ;
        RECT 1514.450 2895.775 1524.650 2896.055 ;
        RECT 1525.490 2895.775 1534.770 2896.055 ;
        RECT 1535.610 2895.775 1545.810 2896.055 ;
        RECT 1546.650 2895.775 1555.930 2896.055 ;
        RECT 1556.770 2895.775 1566.970 2896.055 ;
        RECT 1567.810 2895.775 1577.090 2896.055 ;
        RECT 1577.930 2895.775 1588.130 2896.055 ;
        RECT 1588.970 2895.775 1598.250 2896.055 ;
        RECT 1599.090 2895.775 1609.290 2896.055 ;
        RECT 1610.130 2895.775 1620.330 2896.055 ;
        RECT 1621.170 2895.775 1630.450 2896.055 ;
        RECT 1631.290 2895.775 1641.490 2896.055 ;
        RECT 1642.330 2895.775 1651.610 2896.055 ;
        RECT 1652.450 2895.775 1662.650 2896.055 ;
        RECT 1663.490 2895.775 1672.770 2896.055 ;
        RECT 1673.610 2895.775 1683.810 2896.055 ;
        RECT 1684.650 2895.775 1693.930 2896.055 ;
        RECT 1694.770 2895.775 1704.970 2896.055 ;
        RECT 1705.810 2895.775 1716.010 2896.055 ;
        RECT 1716.850 2895.775 1726.130 2896.055 ;
        RECT 1726.970 2895.775 1737.170 2896.055 ;
        RECT 1738.010 2895.775 1747.290 2896.055 ;
        RECT 1748.130 2895.775 1758.330 2896.055 ;
        RECT 1759.170 2895.775 1768.450 2896.055 ;
        RECT 1769.290 2895.775 1779.490 2896.055 ;
        RECT 1780.330 2895.775 1789.610 2896.055 ;
        RECT 1790.450 2895.775 1800.650 2896.055 ;
        RECT 1801.490 2895.775 1811.690 2896.055 ;
        RECT 1812.530 2895.775 1821.810 2896.055 ;
        RECT 1822.650 2895.775 1832.850 2896.055 ;
        RECT 1833.690 2895.775 1842.970 2896.055 ;
        RECT 1843.810 2895.775 1854.010 2896.055 ;
        RECT 1854.850 2895.775 1864.130 2896.055 ;
        RECT 1864.970 2895.775 1875.170 2896.055 ;
        RECT 1876.010 2895.775 1885.290 2896.055 ;
        RECT 1502.860 2504.280 1885.840 2895.775 ;
        RECT 1503.410 2504.000 1512.690 2504.280 ;
        RECT 1513.530 2504.000 1523.730 2504.280 ;
        RECT 1524.570 2504.000 1533.850 2504.280 ;
        RECT 1534.690 2504.000 1544.890 2504.280 ;
        RECT 1545.730 2504.000 1555.010 2504.280 ;
        RECT 1555.850 2504.000 1566.050 2504.280 ;
        RECT 1566.890 2504.000 1576.170 2504.280 ;
        RECT 1577.010 2504.000 1587.210 2504.280 ;
        RECT 1588.050 2504.000 1598.250 2504.280 ;
        RECT 1599.090 2504.000 1608.370 2504.280 ;
        RECT 1609.210 2504.000 1619.410 2504.280 ;
        RECT 1620.250 2504.000 1629.530 2504.280 ;
        RECT 1630.370 2504.000 1640.570 2504.280 ;
        RECT 1641.410 2504.000 1650.690 2504.280 ;
        RECT 1651.530 2504.000 1661.730 2504.280 ;
        RECT 1662.570 2504.000 1671.850 2504.280 ;
        RECT 1672.690 2504.000 1682.890 2504.280 ;
        RECT 1683.730 2504.000 1693.930 2504.280 ;
        RECT 1694.770 2504.000 1704.050 2504.280 ;
        RECT 1704.890 2504.000 1715.090 2504.280 ;
        RECT 1715.930 2504.000 1725.210 2504.280 ;
        RECT 1726.050 2504.000 1736.250 2504.280 ;
        RECT 1737.090 2504.000 1746.370 2504.280 ;
        RECT 1747.210 2504.000 1757.410 2504.280 ;
        RECT 1758.250 2504.000 1767.530 2504.280 ;
        RECT 1768.370 2504.000 1778.570 2504.280 ;
        RECT 1779.410 2504.000 1789.610 2504.280 ;
        RECT 1790.450 2504.000 1799.730 2504.280 ;
        RECT 1800.570 2504.000 1810.770 2504.280 ;
        RECT 1811.610 2504.000 1820.890 2504.280 ;
        RECT 1821.730 2504.000 1831.930 2504.280 ;
        RECT 1832.770 2504.000 1842.050 2504.280 ;
        RECT 1842.890 2504.000 1853.090 2504.280 ;
        RECT 1853.930 2504.000 1863.210 2504.280 ;
        RECT 1864.050 2504.000 1874.250 2504.280 ;
        RECT 1875.090 2504.000 1885.290 2504.280 ;
      LAYER met2 ;
        RECT 1524.010 2500.000 1524.290 2504.000 ;
        RECT 1534.130 2500.000 1534.410 2504.000 ;
        RECT 1545.170 2500.090 1545.450 2504.000 ;
        RECT 1555.290 2500.090 1555.570 2504.000 ;
        RECT 1576.450 2500.090 1576.730 2504.000 ;
        RECT 1544.840 2500.000 1545.450 2500.090 ;
        RECT 1553.120 2500.000 1555.570 2500.090 ;
        RECT 1575.200 2500.000 1576.730 2500.090 ;
        RECT 1587.490 2500.000 1587.770 2504.000 ;
        RECT 1608.650 2500.000 1608.930 2504.000 ;
        RECT 1619.690 2500.000 1619.970 2504.000 ;
        RECT 1629.810 2500.090 1630.090 2504.000 ;
        RECT 1628.560 2500.000 1630.090 2500.090 ;
        RECT 1640.850 2500.000 1641.130 2504.000 ;
        RECT 1662.010 2500.090 1662.290 2504.000 ;
        RECT 1656.160 2500.000 1662.290 2500.090 ;
        RECT 1683.170 2500.000 1683.450 2504.000 ;
        RECT 1704.330 2500.000 1704.610 2504.000 ;
        RECT 1715.370 2500.000 1715.650 2504.000 ;
        RECT 1725.490 2500.000 1725.770 2504.000 ;
        RECT 1746.650 2500.000 1746.930 2504.000 ;
        RECT 1757.690 2500.000 1757.970 2504.000 ;
        RECT 1767.810 2500.090 1768.090 2504.000 ;
        RECT 1766.560 2500.000 1768.090 2500.090 ;
        RECT 1778.850 2500.000 1779.130 2504.000 ;
        RECT 1789.890 2500.000 1790.170 2504.000 ;
        RECT 1811.050 2500.000 1811.330 2504.000 ;
        RECT 1832.210 2500.000 1832.490 2504.000 ;
        RECT 1842.330 2500.000 1842.610 2504.000 ;
        RECT 1853.370 2500.090 1853.650 2504.000 ;
        RECT 1849.360 2500.000 1853.650 2500.090 ;
        RECT 1874.530 2500.000 1874.810 2504.000 ;
        RECT 1885.570 2500.000 1885.850 2504.000 ;
        RECT 1512.120 2496.970 1512.380 2497.290 ;
        RECT 1503.840 1459.290 1504.100 1459.610 ;
        RECT 1503.380 1458.950 1503.640 1459.270 ;
        RECT 1503.440 1014.210 1503.580 1458.950 ;
        RECT 1503.380 1013.890 1503.640 1014.210 ;
        RECT 1502.460 1009.810 1502.720 1010.130 ;
        RECT 1502.000 1008.790 1502.260 1009.110 ;
        RECT 1503.900 1000.010 1504.040 1459.290 ;
        RECT 1507.060 1019.330 1507.320 1019.650 ;
        RECT 1505.220 1013.550 1505.480 1013.870 ;
        RECT 1505.280 1008.770 1505.420 1013.550 ;
        RECT 1505.220 1008.450 1505.480 1008.770 ;
        RECT 1507.120 1000.010 1507.260 1019.330 ;
        RECT 1511.190 1012.675 1511.470 1013.045 ;
        RECT 1511.200 1012.530 1511.460 1012.675 ;
        RECT 1511.660 1012.530 1511.920 1012.850 ;
        RECT 1511.720 1012.250 1511.860 1012.530 ;
        RECT 1511.260 1012.110 1511.860 1012.250 ;
        RECT 1511.260 1011.830 1511.400 1012.110 ;
        RECT 1511.200 1011.510 1511.460 1011.830 ;
        RECT 1509.360 1008.110 1509.620 1008.430 ;
        RECT 1509.420 1000.010 1509.560 1008.110 ;
        RECT 1512.180 1000.010 1512.320 2496.970 ;
        RECT 1524.140 2484.710 1524.280 2500.000 ;
        RECT 1534.260 2486.070 1534.400 2500.000 ;
        RECT 1544.840 2499.950 1545.370 2500.000 ;
        RECT 1553.120 2499.950 1555.490 2500.000 ;
        RECT 1575.200 2499.950 1576.650 2500.000 ;
        RECT 1534.200 2485.750 1534.460 2486.070 ;
        RECT 1535.120 2485.750 1535.380 2486.070 ;
        RECT 1524.080 2484.390 1524.340 2484.710 ;
        RECT 1535.180 2415.885 1535.320 2485.750 ;
        RECT 1537.880 2484.730 1538.140 2485.050 ;
        RECT 1535.110 2415.515 1535.390 2415.885 ;
        RECT 1535.110 2414.835 1535.390 2415.205 ;
        RECT 1535.180 2319.325 1535.320 2414.835 ;
        RECT 1535.110 2318.955 1535.390 2319.325 ;
        RECT 1534.200 2318.130 1534.460 2318.450 ;
        RECT 1535.110 2318.275 1535.390 2318.645 ;
        RECT 1535.120 2318.130 1535.380 2318.275 ;
        RECT 1534.260 2270.365 1534.400 2318.130 ;
        RECT 1534.190 2269.995 1534.470 2270.365 ;
        RECT 1535.110 2269.995 1535.390 2270.365 ;
        RECT 1535.180 2221.890 1535.320 2269.995 ;
        RECT 1534.200 2221.570 1534.460 2221.890 ;
        RECT 1535.120 2221.570 1535.380 2221.890 ;
        RECT 1534.260 2173.950 1534.400 2221.570 ;
        RECT 1534.200 2173.630 1534.460 2173.950 ;
        RECT 1535.120 2173.630 1535.380 2173.950 ;
        RECT 1535.180 1931.870 1535.320 2173.630 ;
        RECT 1534.200 1931.550 1534.460 1931.870 ;
        RECT 1535.120 1931.550 1535.380 1931.870 ;
        RECT 1534.260 1883.930 1534.400 1931.550 ;
        RECT 1534.200 1883.610 1534.460 1883.930 ;
        RECT 1535.120 1883.610 1535.380 1883.930 ;
        RECT 1535.180 1835.310 1535.320 1883.610 ;
        RECT 1534.200 1834.990 1534.460 1835.310 ;
        RECT 1535.120 1834.990 1535.380 1835.310 ;
        RECT 1534.260 1787.370 1534.400 1834.990 ;
        RECT 1534.200 1787.050 1534.460 1787.370 ;
        RECT 1535.120 1787.050 1535.380 1787.370 ;
        RECT 1535.180 1739.850 1535.320 1787.050 ;
        RECT 1534.720 1739.710 1535.320 1739.850 ;
        RECT 1534.720 1738.750 1534.860 1739.710 ;
        RECT 1534.200 1738.430 1534.460 1738.750 ;
        RECT 1534.660 1738.430 1534.920 1738.750 ;
        RECT 1534.260 1690.810 1534.400 1738.430 ;
        RECT 1534.200 1690.490 1534.460 1690.810 ;
        RECT 1535.120 1690.490 1535.380 1690.810 ;
        RECT 1535.180 1642.190 1535.320 1690.490 ;
        RECT 1535.120 1641.870 1535.380 1642.190 ;
        RECT 1535.120 1641.190 1535.380 1641.510 ;
        RECT 1535.180 1545.970 1535.320 1641.190 ;
        RECT 1535.120 1545.650 1535.380 1545.970 ;
        RECT 1535.580 1545.310 1535.840 1545.630 ;
        RECT 1535.640 1539.170 1535.780 1545.310 ;
        RECT 1535.580 1538.850 1535.840 1539.170 ;
        RECT 1536.040 1538.850 1536.300 1539.170 ;
        RECT 1536.100 1497.690 1536.240 1538.850 ;
        RECT 1535.120 1497.370 1535.380 1497.690 ;
        RECT 1536.040 1497.370 1536.300 1497.690 ;
        RECT 1535.180 1352.850 1535.320 1497.370 ;
        RECT 1535.120 1352.530 1535.380 1352.850 ;
        RECT 1534.660 1352.190 1534.920 1352.510 ;
        RECT 1534.720 1345.370 1534.860 1352.190 ;
        RECT 1533.740 1345.050 1534.000 1345.370 ;
        RECT 1534.660 1345.050 1534.920 1345.370 ;
        RECT 1533.800 1297.430 1533.940 1345.050 ;
        RECT 1533.740 1297.110 1534.000 1297.430 ;
        RECT 1535.120 1297.110 1535.380 1297.430 ;
        RECT 1535.180 1257.650 1535.320 1297.110 ;
        RECT 1535.120 1257.330 1535.380 1257.650 ;
        RECT 1535.120 1256.650 1535.380 1256.970 ;
        RECT 1535.180 1255.010 1535.320 1256.650 ;
        RECT 1535.180 1254.870 1536.240 1255.010 ;
        RECT 1536.100 1208.010 1536.240 1254.870 ;
        RECT 1535.120 1207.690 1535.380 1208.010 ;
        RECT 1536.040 1207.690 1536.300 1208.010 ;
        RECT 1535.180 1200.610 1535.320 1207.690 ;
        RECT 1534.720 1200.470 1535.320 1200.610 ;
        RECT 1534.720 1159.390 1534.860 1200.470 ;
        RECT 1534.660 1159.070 1534.920 1159.390 ;
        RECT 1535.120 1158.730 1535.380 1159.050 ;
        RECT 1535.180 1152.590 1535.320 1158.730 ;
        RECT 1534.660 1152.270 1534.920 1152.590 ;
        RECT 1535.120 1152.270 1535.380 1152.590 ;
        RECT 1534.720 1124.450 1534.860 1152.270 ;
        RECT 1534.720 1124.310 1535.780 1124.450 ;
        RECT 1535.640 1110.770 1535.780 1124.310 ;
        RECT 1535.120 1110.450 1535.380 1110.770 ;
        RECT 1535.580 1110.450 1535.840 1110.770 ;
        RECT 1535.180 1062.830 1535.320 1110.450 ;
        RECT 1535.120 1062.510 1535.380 1062.830 ;
        RECT 1536.040 1062.510 1536.300 1062.830 ;
        RECT 1519.480 1055.370 1519.740 1055.690 ;
        RECT 1514.420 1016.610 1514.680 1016.930 ;
        RECT 1514.480 1000.010 1514.620 1016.610 ;
        RECT 1514.880 1012.530 1515.140 1012.850 ;
        RECT 1420.640 1000.000 1420.940 1000.010 ;
        RECT 1427.380 1000.000 1428.140 1000.010 ;
        RECT 1429.680 1000.000 1431.360 1000.010 ;
        RECT 1433.820 1000.000 1435.040 1000.010 ;
        RECT 1436.120 1000.000 1437.800 1000.010 ;
        RECT 1438.420 1000.000 1440.100 1000.010 ;
        RECT 1442.560 1000.000 1444.240 1000.010 ;
        RECT 1444.860 1000.000 1446.540 1000.010 ;
        RECT 1447.160 1000.000 1448.380 1000.010 ;
        RECT 1451.300 1000.000 1452.980 1000.010 ;
        RECT 1453.600 1000.000 1455.280 1000.010 ;
        RECT 1455.900 1000.000 1457.120 1000.010 ;
        RECT 1460.040 1000.000 1461.720 1000.010 ;
        RECT 1462.340 1000.000 1462.640 1000.010 ;
        RECT 1464.640 1000.000 1465.860 1000.010 ;
        RECT 1468.780 1000.000 1469.080 1000.010 ;
        RECT 1471.080 1000.000 1472.300 1000.010 ;
        RECT 1472.920 1000.000 1474.600 1000.010 ;
        RECT 1477.520 1000.000 1479.200 1000.010 ;
        RECT 1479.820 1000.000 1481.040 1000.010 ;
        RECT 1481.660 1000.000 1482.880 1000.010 ;
        RECT 1486.260 1000.000 1486.560 1000.010 ;
        RECT 1488.560 1000.000 1489.780 1000.010 ;
        RECT 1490.400 1000.000 1492.080 1000.010 ;
        RECT 1495.000 1000.000 1496.220 1000.010 ;
        RECT 1496.840 1000.000 1497.140 1000.010 ;
        RECT 1499.140 1000.000 1500.820 1000.010 ;
        RECT 1503.740 1000.000 1504.040 1000.010 ;
        RECT 1505.580 1000.000 1507.260 1000.010 ;
        RECT 1507.880 1000.000 1509.560 1000.010 ;
        RECT 1512.020 1000.000 1512.320 1000.010 ;
        RECT 1514.320 1000.000 1514.620 1000.010 ;
        RECT 1420.640 999.870 1421.090 1000.000 ;
      LAYER met2 ;
        RECT 1414.930 995.720 1416.390 998.810 ;
      LAYER met2 ;
        RECT 1416.670 996.000 1416.950 999.870 ;
      LAYER met2 ;
        RECT 1417.230 995.720 1418.230 998.810 ;
      LAYER met2 ;
        RECT 1418.510 996.000 1418.790 999.870 ;
      LAYER met2 ;
        RECT 1419.070 995.720 1420.530 998.810 ;
      LAYER met2 ;
        RECT 1420.810 996.000 1421.090 999.870 ;
      LAYER met2 ;
        RECT 1421.370 995.720 1422.830 998.810 ;
      LAYER met2 ;
        RECT 1423.110 996.000 1423.390 1000.000 ;
      LAYER met2 ;
        RECT 1423.670 995.720 1424.670 998.810 ;
      LAYER met2 ;
        RECT 1424.950 996.000 1425.230 1000.000 ;
        RECT 1427.250 999.870 1428.140 1000.000 ;
        RECT 1429.550 999.870 1431.360 1000.000 ;
      LAYER met2 ;
        RECT 1425.510 995.720 1426.970 998.810 ;
      LAYER met2 ;
        RECT 1427.250 996.000 1427.530 999.870 ;
      LAYER met2 ;
        RECT 1427.810 995.720 1429.270 998.810 ;
      LAYER met2 ;
        RECT 1429.550 996.000 1429.830 999.870 ;
      LAYER met2 ;
        RECT 1430.110 995.720 1431.570 998.810 ;
      LAYER met2 ;
        RECT 1431.850 996.000 1432.130 1000.000 ;
        RECT 1433.690 999.870 1435.040 1000.000 ;
        RECT 1435.990 999.870 1437.800 1000.000 ;
        RECT 1438.290 999.870 1440.100 1000.000 ;
      LAYER met2 ;
        RECT 1432.410 995.720 1433.410 998.810 ;
      LAYER met2 ;
        RECT 1433.690 996.000 1433.970 999.870 ;
      LAYER met2 ;
        RECT 1434.250 995.720 1435.710 998.810 ;
      LAYER met2 ;
        RECT 1435.990 996.000 1436.270 999.870 ;
      LAYER met2 ;
        RECT 1436.550 995.720 1438.010 998.810 ;
      LAYER met2 ;
        RECT 1438.290 996.000 1438.570 999.870 ;
      LAYER met2 ;
        RECT 1438.850 995.720 1440.310 998.810 ;
      LAYER met2 ;
        RECT 1440.590 996.000 1440.870 1000.000 ;
        RECT 1442.430 999.870 1444.240 1000.000 ;
        RECT 1444.730 999.870 1446.540 1000.000 ;
        RECT 1447.030 999.870 1448.380 1000.000 ;
      LAYER met2 ;
        RECT 1441.150 995.720 1442.150 998.810 ;
      LAYER met2 ;
        RECT 1442.430 996.000 1442.710 999.870 ;
      LAYER met2 ;
        RECT 1442.990 995.720 1444.450 998.810 ;
      LAYER met2 ;
        RECT 1444.730 996.000 1445.010 999.870 ;
      LAYER met2 ;
        RECT 1445.290 995.720 1446.750 998.810 ;
      LAYER met2 ;
        RECT 1447.030 996.000 1447.310 999.870 ;
      LAYER met2 ;
        RECT 1447.590 995.720 1448.590 998.810 ;
      LAYER met2 ;
        RECT 1448.870 996.000 1449.150 1000.000 ;
        RECT 1451.170 999.870 1452.980 1000.000 ;
        RECT 1453.470 999.870 1455.280 1000.000 ;
        RECT 1455.770 999.870 1457.120 1000.000 ;
      LAYER met2 ;
        RECT 1449.430 995.720 1450.890 998.810 ;
      LAYER met2 ;
        RECT 1451.170 996.000 1451.450 999.870 ;
      LAYER met2 ;
        RECT 1451.730 995.720 1453.190 998.810 ;
      LAYER met2 ;
        RECT 1453.470 996.000 1453.750 999.870 ;
      LAYER met2 ;
        RECT 1454.030 995.720 1455.490 998.810 ;
      LAYER met2 ;
        RECT 1455.770 996.000 1456.050 999.870 ;
      LAYER met2 ;
        RECT 1456.330 995.720 1457.330 998.810 ;
      LAYER met2 ;
        RECT 1457.610 996.000 1457.890 1000.000 ;
        RECT 1459.910 999.870 1461.720 1000.000 ;
        RECT 1462.210 999.870 1462.640 1000.000 ;
        RECT 1464.510 999.870 1465.860 1000.000 ;
      LAYER met2 ;
        RECT 1458.170 995.720 1459.630 998.810 ;
      LAYER met2 ;
        RECT 1459.910 996.000 1460.190 999.870 ;
      LAYER met2 ;
        RECT 1460.470 995.720 1461.930 998.810 ;
      LAYER met2 ;
        RECT 1462.210 996.000 1462.490 999.870 ;
      LAYER met2 ;
        RECT 1462.770 995.720 1464.230 998.810 ;
      LAYER met2 ;
        RECT 1464.510 996.000 1464.790 999.870 ;
      LAYER met2 ;
        RECT 1465.070 995.720 1466.070 998.810 ;
      LAYER met2 ;
        RECT 1466.350 996.000 1466.630 1000.000 ;
        RECT 1468.650 999.870 1469.080 1000.000 ;
        RECT 1470.950 999.870 1472.300 1000.000 ;
        RECT 1472.790 999.870 1474.600 1000.000 ;
      LAYER met2 ;
        RECT 1466.910 995.720 1468.370 998.810 ;
      LAYER met2 ;
        RECT 1468.650 996.000 1468.930 999.870 ;
      LAYER met2 ;
        RECT 1469.210 995.720 1470.670 998.810 ;
      LAYER met2 ;
        RECT 1470.950 996.000 1471.230 999.870 ;
      LAYER met2 ;
        RECT 1471.510 995.720 1472.510 998.810 ;
      LAYER met2 ;
        RECT 1472.790 996.000 1473.070 999.870 ;
      LAYER met2 ;
        RECT 1473.350 995.720 1474.810 998.810 ;
      LAYER met2 ;
        RECT 1475.090 996.000 1475.370 1000.000 ;
        RECT 1477.390 999.870 1479.200 1000.000 ;
        RECT 1479.690 999.870 1481.040 1000.000 ;
        RECT 1481.530 999.870 1482.880 1000.000 ;
      LAYER met2 ;
        RECT 1475.650 995.720 1477.110 998.810 ;
      LAYER met2 ;
        RECT 1477.390 996.000 1477.670 999.870 ;
      LAYER met2 ;
        RECT 1477.950 995.720 1479.410 998.810 ;
      LAYER met2 ;
        RECT 1479.690 996.000 1479.970 999.870 ;
      LAYER met2 ;
        RECT 1480.250 995.720 1481.250 998.810 ;
      LAYER met2 ;
        RECT 1481.530 996.000 1481.810 999.870 ;
      LAYER met2 ;
        RECT 1482.090 995.720 1483.550 998.810 ;
      LAYER met2 ;
        RECT 1483.830 996.000 1484.110 1000.000 ;
        RECT 1486.130 999.870 1486.560 1000.000 ;
        RECT 1488.430 999.870 1489.780 1000.000 ;
        RECT 1490.270 999.870 1492.080 1000.000 ;
      LAYER met2 ;
        RECT 1484.390 995.720 1485.850 998.810 ;
      LAYER met2 ;
        RECT 1486.130 996.000 1486.410 999.870 ;
      LAYER met2 ;
        RECT 1486.690 995.720 1488.150 998.810 ;
      LAYER met2 ;
        RECT 1488.430 996.000 1488.710 999.870 ;
      LAYER met2 ;
        RECT 1488.990 995.720 1489.990 998.810 ;
      LAYER met2 ;
        RECT 1490.270 996.000 1490.550 999.870 ;
      LAYER met2 ;
        RECT 1490.830 995.720 1492.290 998.810 ;
      LAYER met2 ;
        RECT 1492.570 996.000 1492.850 1000.000 ;
        RECT 1494.870 999.870 1496.220 1000.000 ;
        RECT 1496.710 999.870 1497.140 1000.000 ;
        RECT 1499.010 999.870 1500.820 1000.000 ;
      LAYER met2 ;
        RECT 1493.130 995.720 1494.590 998.810 ;
      LAYER met2 ;
        RECT 1494.870 996.000 1495.150 999.870 ;
      LAYER met2 ;
        RECT 1495.430 995.720 1496.430 998.810 ;
      LAYER met2 ;
        RECT 1496.710 996.000 1496.990 999.870 ;
      LAYER met2 ;
        RECT 1497.270 995.720 1498.730 998.810 ;
      LAYER met2 ;
        RECT 1499.010 996.000 1499.290 999.870 ;
      LAYER met2 ;
        RECT 1499.570 995.720 1501.030 998.810 ;
      LAYER met2 ;
        RECT 1501.310 996.000 1501.590 1000.000 ;
        RECT 1503.610 999.870 1504.040 1000.000 ;
        RECT 1505.450 999.870 1507.260 1000.000 ;
        RECT 1507.750 999.870 1509.560 1000.000 ;
      LAYER met2 ;
        RECT 1501.870 995.720 1503.330 998.810 ;
      LAYER met2 ;
        RECT 1503.610 996.000 1503.890 999.870 ;
      LAYER met2 ;
        RECT 1504.170 995.720 1505.170 998.810 ;
      LAYER met2 ;
        RECT 1505.450 996.000 1505.730 999.870 ;
      LAYER met2 ;
        RECT 1506.010 995.720 1507.470 998.810 ;
      LAYER met2 ;
        RECT 1507.750 996.000 1508.030 999.870 ;
      LAYER met2 ;
        RECT 1508.310 995.720 1509.770 998.810 ;
      LAYER met2 ;
        RECT 1510.050 996.000 1510.330 1000.000 ;
        RECT 1511.890 999.870 1512.320 1000.000 ;
        RECT 1514.190 999.870 1514.620 1000.000 ;
        RECT 1514.940 1000.010 1515.080 1012.530 ;
        RECT 1519.540 1010.890 1519.680 1055.370 ;
        RECT 1533.280 1019.670 1533.540 1019.990 ;
        RECT 1525.000 1013.210 1525.260 1013.530 ;
        RECT 1519.540 1010.750 1522.440 1010.890 ;
        RECT 1519.480 1010.150 1519.740 1010.470 ;
        RECT 1519.540 1000.010 1519.680 1010.150 ;
        RECT 1521.310 1009.955 1521.590 1010.325 ;
        RECT 1521.380 1009.790 1521.520 1009.955 ;
        RECT 1521.320 1009.470 1521.580 1009.790 ;
        RECT 1522.300 1000.010 1522.440 1010.750 ;
        RECT 1525.060 1000.010 1525.200 1013.210 ;
        RECT 1528.220 1012.870 1528.480 1013.190 ;
        RECT 1527.760 1011.510 1528.020 1011.830 ;
        RECT 1527.820 1009.450 1527.960 1011.510 ;
        RECT 1527.760 1009.130 1528.020 1009.450 ;
        RECT 1528.280 1000.010 1528.420 1012.870 ;
        RECT 1533.340 1000.010 1533.480 1019.670 ;
        RECT 1535.580 1013.890 1535.840 1014.210 ;
        RECT 1534.660 1013.210 1534.920 1013.530 ;
        RECT 1534.720 1012.170 1534.860 1013.210 ;
        RECT 1534.660 1011.850 1534.920 1012.170 ;
        RECT 1535.120 1011.850 1535.380 1012.170 ;
        RECT 1534.660 1010.150 1534.920 1010.470 ;
        RECT 1534.720 1007.750 1534.860 1010.150 ;
        RECT 1534.660 1007.430 1534.920 1007.750 ;
        RECT 1535.180 1000.010 1535.320 1011.850 ;
        RECT 1535.640 1009.110 1535.780 1013.890 ;
        RECT 1536.100 1013.870 1536.240 1062.510 ;
        RECT 1536.040 1013.550 1536.300 1013.870 ;
        RECT 1536.040 1013.045 1536.300 1013.190 ;
        RECT 1536.030 1012.675 1536.310 1013.045 ;
        RECT 1536.500 1012.530 1536.760 1012.850 ;
        RECT 1536.560 1010.325 1536.700 1012.530 ;
        RECT 1537.940 1012.170 1538.080 2484.730 ;
        RECT 1544.320 2463.650 1544.580 2463.970 ;
        RECT 1544.380 2432.090 1544.520 2463.650 ;
        RECT 1543.920 2431.950 1544.520 2432.090 ;
        RECT 1543.920 2408.210 1544.060 2431.950 ;
        RECT 1543.860 2407.890 1544.120 2408.210 ;
        RECT 1544.320 2407.890 1544.580 2408.210 ;
        RECT 1544.380 2367.070 1544.520 2407.890 ;
        RECT 1544.320 2366.750 1544.580 2367.070 ;
        RECT 1543.860 2366.410 1544.120 2366.730 ;
        RECT 1543.920 2360.010 1544.060 2366.410 ;
        RECT 1543.920 2359.870 1544.520 2360.010 ;
        RECT 1544.380 2262.770 1544.520 2359.870 ;
        RECT 1543.920 2262.630 1544.520 2262.770 ;
        RECT 1543.920 2215.090 1544.060 2262.630 ;
        RECT 1543.860 2214.770 1544.120 2215.090 ;
        RECT 1544.320 2214.770 1544.580 2215.090 ;
        RECT 1544.380 2166.210 1544.520 2214.770 ;
        RECT 1543.920 2166.070 1544.520 2166.210 ;
        RECT 1543.920 2118.530 1544.060 2166.070 ;
        RECT 1543.860 2118.210 1544.120 2118.530 ;
        RECT 1544.320 2118.210 1544.580 2118.530 ;
        RECT 1544.380 2069.650 1544.520 2118.210 ;
        RECT 1543.920 2069.510 1544.520 2069.650 ;
        RECT 1543.920 2021.970 1544.060 2069.510 ;
        RECT 1543.860 2021.650 1544.120 2021.970 ;
        RECT 1544.320 2021.650 1544.580 2021.970 ;
        RECT 1544.380 1973.010 1544.520 2021.650 ;
        RECT 1542.940 1972.690 1543.200 1973.010 ;
        RECT 1544.320 1972.690 1544.580 1973.010 ;
        RECT 1543.000 1883.930 1543.140 1972.690 ;
        RECT 1542.940 1883.610 1543.200 1883.930 ;
        RECT 1543.400 1883.610 1543.660 1883.930 ;
        RECT 1543.460 1829.190 1543.600 1883.610 ;
        RECT 1543.400 1828.870 1543.660 1829.190 ;
        RECT 1544.320 1828.870 1544.580 1829.190 ;
        RECT 1544.380 1828.510 1544.520 1828.870 ;
        RECT 1543.400 1828.190 1543.660 1828.510 ;
        RECT 1544.320 1828.190 1544.580 1828.510 ;
        RECT 1543.460 1787.370 1543.600 1828.190 ;
        RECT 1543.400 1787.050 1543.660 1787.370 ;
        RECT 1544.320 1786.710 1544.580 1787.030 ;
        RECT 1544.380 1756.170 1544.520 1786.710 ;
        RECT 1543.460 1756.030 1544.520 1756.170 ;
        RECT 1543.460 1732.290 1543.600 1756.030 ;
        RECT 1543.400 1731.970 1543.660 1732.290 ;
        RECT 1543.860 1731.970 1544.120 1732.290 ;
        RECT 1543.920 1690.810 1544.060 1731.970 ;
        RECT 1543.860 1690.490 1544.120 1690.810 ;
        RECT 1544.320 1689.810 1544.580 1690.130 ;
        RECT 1544.380 1683.410 1544.520 1689.810 ;
        RECT 1543.920 1683.270 1544.520 1683.410 ;
        RECT 1543.920 1636.070 1544.060 1683.270 ;
        RECT 1543.860 1635.750 1544.120 1636.070 ;
        RECT 1544.320 1635.410 1544.580 1635.730 ;
        RECT 1544.380 1586.850 1544.520 1635.410 ;
        RECT 1543.920 1586.710 1544.520 1586.850 ;
        RECT 1543.920 1497.690 1544.060 1586.710 ;
        RECT 1543.400 1497.370 1543.660 1497.690 ;
        RECT 1543.860 1497.370 1544.120 1497.690 ;
        RECT 1543.460 1463.010 1543.600 1497.370 ;
        RECT 1543.400 1462.690 1543.660 1463.010 ;
        RECT 1544.320 1462.690 1544.580 1463.010 ;
        RECT 1544.380 1418.130 1544.520 1462.690 ;
        RECT 1542.940 1417.810 1543.200 1418.130 ;
        RECT 1544.320 1417.810 1544.580 1418.130 ;
        RECT 1543.000 1393.990 1543.140 1417.810 ;
        RECT 1542.940 1393.670 1543.200 1393.990 ;
        RECT 1543.400 1393.670 1543.660 1393.990 ;
        RECT 1543.460 1345.710 1543.600 1393.670 ;
        RECT 1543.400 1345.390 1543.660 1345.710 ;
        RECT 1544.320 1345.390 1544.580 1345.710 ;
        RECT 1544.380 1257.165 1544.520 1345.390 ;
        RECT 1544.310 1256.795 1544.590 1257.165 ;
        RECT 1544.310 1256.115 1544.590 1256.485 ;
        RECT 1544.380 1227.050 1544.520 1256.115 ;
        RECT 1542.940 1226.730 1543.200 1227.050 ;
        RECT 1544.320 1226.730 1544.580 1227.050 ;
        RECT 1543.000 1176.730 1543.140 1226.730 ;
        RECT 1542.940 1176.410 1543.200 1176.730 ;
        RECT 1543.860 1176.410 1544.120 1176.730 ;
        RECT 1543.920 1152.330 1544.060 1176.410 ;
        RECT 1543.460 1152.190 1544.060 1152.330 ;
        RECT 1543.460 1111.110 1543.600 1152.190 ;
        RECT 1543.400 1110.790 1543.660 1111.110 ;
        RECT 1543.860 1110.450 1544.120 1110.770 ;
        RECT 1543.920 1104.310 1544.060 1110.450 ;
        RECT 1543.400 1103.990 1543.660 1104.310 ;
        RECT 1543.860 1103.990 1544.120 1104.310 ;
        RECT 1543.460 1080.170 1543.600 1103.990 ;
        RECT 1541.560 1079.850 1541.820 1080.170 ;
        RECT 1543.400 1079.850 1543.660 1080.170 ;
        RECT 1541.620 1061.890 1541.760 1079.850 ;
        RECT 1541.620 1061.750 1542.220 1061.890 ;
        RECT 1542.080 1028.150 1542.220 1061.750 ;
        RECT 1542.020 1027.830 1542.280 1028.150 ;
        RECT 1542.940 1027.830 1543.200 1028.150 ;
        RECT 1542.020 1020.010 1542.280 1020.330 ;
        RECT 1537.880 1011.850 1538.140 1012.170 ;
        RECT 1536.490 1009.955 1536.770 1010.325 ;
        RECT 1535.580 1008.790 1535.840 1009.110 ;
        RECT 1536.500 1007.770 1536.760 1008.090 ;
        RECT 1514.940 1000.000 1516.620 1000.010 ;
        RECT 1519.540 1000.000 1520.760 1000.010 ;
        RECT 1522.300 1000.000 1523.060 1000.010 ;
        RECT 1525.060 1000.000 1525.360 1000.010 ;
        RECT 1528.280 1000.000 1529.500 1000.010 ;
        RECT 1531.800 1000.000 1533.480 1000.010 ;
        RECT 1534.100 1000.000 1535.320 1000.010 ;
        RECT 1536.560 1000.010 1536.700 1007.770 ;
        RECT 1542.080 1000.010 1542.220 1020.010 ;
        RECT 1543.000 1014.290 1543.140 1027.830 ;
        RECT 1544.840 1015.910 1544.980 2499.950 ;
        RECT 1552.600 2494.930 1552.860 2495.250 ;
        RECT 1545.240 2494.250 1545.500 2494.570 ;
        RECT 1545.300 2463.970 1545.440 2494.250 ;
        RECT 1546.620 2484.390 1546.880 2484.710 ;
        RECT 1545.240 2463.650 1545.500 2463.970 ;
        RECT 1544.780 1015.590 1545.040 1015.910 ;
        RECT 1543.000 1014.150 1544.060 1014.290 ;
        RECT 1543.920 1001.290 1544.060 1014.150 ;
        RECT 1542.710 1000.970 1542.970 1001.290 ;
        RECT 1543.860 1000.970 1544.120 1001.290 ;
        RECT 1536.560 1000.000 1538.240 1000.010 ;
        RECT 1540.540 1000.000 1542.220 1000.010 ;
        RECT 1542.770 1000.000 1542.910 1000.970 ;
        RECT 1546.680 1000.010 1546.820 2484.390 ;
        RECT 1552.140 1013.550 1552.400 1013.870 ;
        RECT 1547.540 1012.870 1547.800 1013.190 ;
        RECT 1547.600 1000.010 1547.740 1012.870 ;
        RECT 1552.200 1000.010 1552.340 1013.550 ;
        RECT 1552.660 1012.170 1552.800 2494.930 ;
        RECT 1553.120 1735.350 1553.260 2499.950 ;
        RECT 1559.500 2494.590 1559.760 2494.910 ;
        RECT 1553.060 1735.030 1553.320 1735.350 ;
        RECT 1559.560 1014.210 1559.700 2494.590 ;
        RECT 1575.200 2485.050 1575.340 2499.950 ;
        RECT 1586.640 2494.590 1586.900 2494.910 ;
        RECT 1575.140 2484.730 1575.400 2485.050 ;
        RECT 1576.520 2484.730 1576.780 2485.050 ;
        RECT 1559.960 1051.970 1560.220 1052.290 ;
        RECT 1559.500 1013.890 1559.760 1014.210 ;
        RECT 1555.820 1012.870 1556.080 1013.190 ;
        RECT 1552.600 1011.850 1552.860 1012.170 ;
        RECT 1555.880 1000.010 1556.020 1012.870 ;
        RECT 1556.280 1011.850 1556.540 1012.170 ;
        RECT 1556.740 1011.850 1557.000 1012.170 ;
        RECT 1546.680 1000.000 1546.980 1000.010 ;
        RECT 1547.600 1000.000 1549.280 1000.010 ;
        RECT 1551.580 1000.000 1552.340 1000.010 ;
        RECT 1555.720 1000.000 1556.020 1000.010 ;
        RECT 1514.940 999.870 1516.770 1000.000 ;
      LAYER met2 ;
        RECT 1510.610 995.720 1511.610 998.810 ;
      LAYER met2 ;
        RECT 1511.890 996.000 1512.170 999.870 ;
      LAYER met2 ;
        RECT 1512.450 995.720 1513.910 998.810 ;
      LAYER met2 ;
        RECT 1514.190 996.000 1514.470 999.870 ;
      LAYER met2 ;
        RECT 1514.750 995.720 1516.210 998.810 ;
      LAYER met2 ;
        RECT 1516.490 996.000 1516.770 999.870 ;
      LAYER met2 ;
        RECT 1517.050 995.720 1518.510 998.810 ;
      LAYER met2 ;
        RECT 1518.790 996.000 1519.070 1000.000 ;
        RECT 1519.540 999.870 1520.910 1000.000 ;
        RECT 1522.300 999.870 1523.210 1000.000 ;
        RECT 1525.060 999.870 1525.510 1000.000 ;
      LAYER met2 ;
        RECT 1519.350 995.720 1520.350 998.810 ;
      LAYER met2 ;
        RECT 1520.630 996.000 1520.910 999.870 ;
      LAYER met2 ;
        RECT 1521.190 995.720 1522.650 998.810 ;
      LAYER met2 ;
        RECT 1522.930 996.000 1523.210 999.870 ;
      LAYER met2 ;
        RECT 1523.490 995.720 1524.950 998.810 ;
      LAYER met2 ;
        RECT 1525.230 996.000 1525.510 999.870 ;
      LAYER met2 ;
        RECT 1525.790 995.720 1527.250 998.810 ;
      LAYER met2 ;
        RECT 1527.530 996.000 1527.810 1000.000 ;
        RECT 1528.280 999.870 1529.650 1000.000 ;
      LAYER met2 ;
        RECT 1528.090 995.720 1529.090 998.810 ;
      LAYER met2 ;
        RECT 1529.370 996.000 1529.650 999.870 ;
        RECT 1531.670 999.870 1533.480 1000.000 ;
        RECT 1533.970 999.870 1535.320 1000.000 ;
      LAYER met2 ;
        RECT 1529.930 995.720 1531.390 998.810 ;
      LAYER met2 ;
        RECT 1531.670 996.000 1531.950 999.870 ;
      LAYER met2 ;
        RECT 1532.230 995.720 1533.690 998.810 ;
      LAYER met2 ;
        RECT 1533.970 996.000 1534.250 999.870 ;
      LAYER met2 ;
        RECT 1534.530 995.720 1535.530 998.810 ;
      LAYER met2 ;
        RECT 1535.810 996.000 1536.090 1000.000 ;
        RECT 1536.560 999.870 1538.390 1000.000 ;
      LAYER met2 ;
        RECT 1536.370 995.720 1537.830 998.810 ;
      LAYER met2 ;
        RECT 1538.110 996.000 1538.390 999.870 ;
        RECT 1540.410 999.870 1542.220 1000.000 ;
      LAYER met2 ;
        RECT 1538.670 995.720 1540.130 998.810 ;
      LAYER met2 ;
        RECT 1540.410 996.000 1540.690 999.870 ;
      LAYER met2 ;
        RECT 1540.970 995.720 1542.430 998.810 ;
      LAYER met2 ;
        RECT 1542.710 996.000 1542.990 1000.000 ;
      LAYER met2 ;
        RECT 1543.270 995.720 1544.270 998.810 ;
      LAYER met2 ;
        RECT 1544.550 996.000 1544.830 1000.000 ;
        RECT 1546.680 999.870 1547.130 1000.000 ;
        RECT 1547.600 999.870 1549.430 1000.000 ;
      LAYER met2 ;
        RECT 1545.110 995.720 1546.570 998.810 ;
      LAYER met2 ;
        RECT 1546.850 996.000 1547.130 999.870 ;
      LAYER met2 ;
        RECT 1547.410 995.720 1548.870 998.810 ;
      LAYER met2 ;
        RECT 1549.150 996.000 1549.430 999.870 ;
        RECT 1551.450 999.870 1552.340 1000.000 ;
      LAYER met2 ;
        RECT 1549.710 995.720 1551.170 998.810 ;
      LAYER met2 ;
        RECT 1551.450 996.000 1551.730 999.870 ;
      LAYER met2 ;
        RECT 1552.010 995.720 1553.010 998.810 ;
      LAYER met2 ;
        RECT 1553.290 996.000 1553.570 1000.000 ;
        RECT 1555.590 999.870 1556.020 1000.000 ;
        RECT 1556.340 1000.010 1556.480 1011.850 ;
        RECT 1556.800 1008.770 1556.940 1011.850 ;
        RECT 1556.740 1008.450 1557.000 1008.770 ;
        RECT 1560.020 1000.010 1560.160 1051.970 ;
        RECT 1567.780 1020.690 1568.040 1021.010 ;
        RECT 1562.720 1013.890 1562.980 1014.210 ;
        RECT 1563.180 1013.890 1563.440 1014.210 ;
        RECT 1556.340 1000.000 1558.020 1000.010 ;
        RECT 1559.860 1000.000 1560.160 1000.010 ;
        RECT 1562.780 1000.010 1562.920 1013.890 ;
        RECT 1563.240 1008.430 1563.380 1013.890 ;
        RECT 1563.180 1008.110 1563.440 1008.430 ;
        RECT 1567.840 1000.010 1567.980 1020.690 ;
        RECT 1574.680 1020.350 1574.940 1020.670 ;
        RECT 1568.240 1008.790 1568.500 1009.110 ;
        RECT 1562.780 1000.000 1564.460 1000.010 ;
        RECT 1566.760 1000.000 1567.980 1000.010 ;
        RECT 1556.340 999.870 1558.170 1000.000 ;
      LAYER met2 ;
        RECT 1553.850 995.720 1555.310 998.810 ;
      LAYER met2 ;
        RECT 1555.590 996.000 1555.870 999.870 ;
      LAYER met2 ;
        RECT 1556.150 995.720 1557.610 998.810 ;
      LAYER met2 ;
        RECT 1557.890 996.000 1558.170 999.870 ;
        RECT 1559.730 999.870 1560.160 1000.000 ;
      LAYER met2 ;
        RECT 1558.450 995.720 1559.450 998.810 ;
      LAYER met2 ;
        RECT 1559.730 996.000 1560.010 999.870 ;
      LAYER met2 ;
        RECT 1560.290 995.720 1561.750 998.810 ;
      LAYER met2 ;
        RECT 1562.030 996.000 1562.310 1000.000 ;
        RECT 1562.780 999.870 1564.610 1000.000 ;
      LAYER met2 ;
        RECT 1562.590 995.720 1564.050 998.810 ;
      LAYER met2 ;
        RECT 1564.330 996.000 1564.610 999.870 ;
        RECT 1566.630 999.870 1567.980 1000.000 ;
        RECT 1568.300 1000.010 1568.440 1008.790 ;
        RECT 1574.740 1000.010 1574.880 1020.350 ;
        RECT 1576.060 1015.930 1576.320 1016.250 ;
        RECT 1576.120 1000.010 1576.260 1015.930 ;
        RECT 1576.580 1012.510 1576.720 2484.730 ;
        RECT 1586.700 1023.810 1586.840 2494.590 ;
        RECT 1587.620 2485.730 1587.760 2500.000 ;
        RECT 1607.340 2494.930 1607.600 2495.250 ;
        RECT 1593.540 2489.150 1593.800 2489.470 ;
        RECT 1587.560 2485.410 1587.820 2485.730 ;
        RECT 1585.320 1023.670 1586.840 1023.810 ;
        RECT 1576.520 1012.190 1576.780 1012.510 ;
        RECT 1576.520 1010.150 1576.780 1010.470 ;
        RECT 1568.300 1000.000 1568.600 1000.010 ;
        RECT 1573.200 1000.000 1574.880 1000.010 ;
        RECT 1575.500 1000.000 1576.260 1000.010 ;
        RECT 1568.300 999.870 1568.750 1000.000 ;
      LAYER met2 ;
        RECT 1564.890 995.720 1566.350 998.810 ;
      LAYER met2 ;
        RECT 1566.630 996.000 1566.910 999.870 ;
      LAYER met2 ;
        RECT 1567.190 995.720 1568.190 998.810 ;
      LAYER met2 ;
        RECT 1568.470 996.000 1568.750 999.870 ;
      LAYER met2 ;
        RECT 1569.030 995.720 1570.490 998.810 ;
      LAYER met2 ;
        RECT 1570.770 996.000 1571.050 1000.000 ;
        RECT 1573.070 999.870 1574.880 1000.000 ;
        RECT 1575.370 999.870 1576.260 1000.000 ;
        RECT 1576.580 1000.010 1576.720 1010.150 ;
        RECT 1577.900 1009.470 1578.160 1009.790 ;
        RECT 1577.960 1000.010 1578.100 1009.470 ;
        RECT 1585.320 1000.010 1585.460 1023.670 ;
        RECT 1585.720 1009.810 1585.980 1010.130 ;
        RECT 1576.580 1000.000 1577.340 1000.010 ;
        RECT 1577.960 1000.000 1579.640 1000.010 ;
        RECT 1583.780 1000.000 1585.460 1000.010 ;
        RECT 1576.580 999.870 1577.490 1000.000 ;
        RECT 1577.960 999.870 1579.790 1000.000 ;
      LAYER met2 ;
        RECT 1571.330 995.720 1572.790 998.810 ;
      LAYER met2 ;
        RECT 1573.070 996.000 1573.350 999.870 ;
      LAYER met2 ;
        RECT 1573.630 995.720 1575.090 998.810 ;
      LAYER met2 ;
        RECT 1575.370 996.000 1575.650 999.870 ;
      LAYER met2 ;
        RECT 1575.930 995.720 1576.930 998.810 ;
      LAYER met2 ;
        RECT 1577.210 996.000 1577.490 999.870 ;
      LAYER met2 ;
        RECT 1577.770 995.720 1579.230 998.810 ;
      LAYER met2 ;
        RECT 1579.510 996.000 1579.790 999.870 ;
      LAYER met2 ;
        RECT 1580.070 995.720 1581.530 998.810 ;
      LAYER met2 ;
        RECT 1581.810 996.000 1582.090 1000.000 ;
        RECT 1583.650 999.870 1585.460 1000.000 ;
        RECT 1585.780 1000.010 1585.920 1009.810 ;
        RECT 1593.600 1000.010 1593.740 2489.150 ;
        RECT 1600.440 2488.810 1600.700 2489.130 ;
        RECT 1595.840 1021.030 1596.100 1021.350 ;
        RECT 1595.900 1014.210 1596.040 1021.030 ;
        RECT 1600.500 1014.210 1600.640 2488.810 ;
        RECT 1595.840 1013.890 1596.100 1014.210 ;
        RECT 1596.300 1013.890 1596.560 1014.210 ;
        RECT 1600.440 1013.890 1600.700 1014.210 ;
        RECT 1596.360 1000.010 1596.500 1013.890 ;
        RECT 1603.200 1013.210 1603.460 1013.530 ;
        RECT 1602.740 1009.810 1603.000 1010.130 ;
        RECT 1602.800 1000.010 1602.940 1009.810 ;
        RECT 1585.780 1000.000 1586.080 1000.010 ;
        RECT 1592.520 1000.000 1593.740 1000.010 ;
        RECT 1594.820 1000.000 1596.500 1000.010 ;
        RECT 1601.260 1000.000 1602.940 1000.010 ;
        RECT 1585.780 999.870 1586.230 1000.000 ;
      LAYER met2 ;
        RECT 1582.370 995.720 1583.370 998.810 ;
      LAYER met2 ;
        RECT 1583.650 996.000 1583.930 999.870 ;
      LAYER met2 ;
        RECT 1584.210 995.720 1585.670 998.810 ;
      LAYER met2 ;
        RECT 1585.950 996.000 1586.230 999.870 ;
      LAYER met2 ;
        RECT 1586.510 995.720 1587.970 998.810 ;
      LAYER met2 ;
        RECT 1588.250 996.000 1588.530 1000.000 ;
      LAYER met2 ;
        RECT 1588.810 995.720 1590.270 998.810 ;
      LAYER met2 ;
        RECT 1590.550 996.000 1590.830 1000.000 ;
        RECT 1592.390 999.870 1593.740 1000.000 ;
        RECT 1594.690 999.870 1596.500 1000.000 ;
      LAYER met2 ;
        RECT 1591.110 995.720 1592.110 998.810 ;
      LAYER met2 ;
        RECT 1592.390 996.000 1592.670 999.870 ;
      LAYER met2 ;
        RECT 1592.950 995.720 1594.410 998.810 ;
      LAYER met2 ;
        RECT 1594.690 996.000 1594.970 999.870 ;
      LAYER met2 ;
        RECT 1595.250 995.720 1596.710 998.810 ;
      LAYER met2 ;
        RECT 1596.990 996.000 1597.270 1000.000 ;
      LAYER met2 ;
        RECT 1597.550 995.720 1599.010 998.810 ;
      LAYER met2 ;
        RECT 1599.290 996.000 1599.570 1000.000 ;
        RECT 1601.130 999.870 1602.940 1000.000 ;
        RECT 1603.260 1000.010 1603.400 1013.210 ;
        RECT 1607.400 1010.130 1607.540 2494.930 ;
        RECT 1608.780 2485.390 1608.920 2500.000 ;
        RECT 1608.720 2485.070 1608.980 2485.390 ;
        RECT 1619.820 2485.050 1619.960 2500.000 ;
        RECT 1628.560 2499.950 1630.010 2500.000 ;
        RECT 1621.140 2495.270 1621.400 2495.590 ;
        RECT 1619.760 2484.730 1620.020 2485.050 ;
        RECT 1614.240 1459.630 1614.500 1459.950 ;
        RECT 1608.720 1015.590 1608.980 1015.910 ;
        RECT 1607.340 1009.810 1607.600 1010.130 ;
        RECT 1608.780 1000.010 1608.920 1015.590 ;
        RECT 1614.300 1000.690 1614.440 1459.630 ;
        RECT 1620.220 1009.810 1620.480 1010.130 ;
        RECT 1613.380 1000.550 1614.440 1000.690 ;
        RECT 1613.380 1000.010 1613.520 1000.550 ;
        RECT 1620.280 1000.010 1620.420 1009.810 ;
        RECT 1621.200 1000.010 1621.340 2495.270 ;
        RECT 1624.820 2484.390 1625.080 2484.710 ;
        RECT 1624.880 1010.130 1625.020 2484.390 ;
        RECT 1625.740 1016.270 1626.000 1016.590 ;
        RECT 1624.820 1009.810 1625.080 1010.130 ;
        RECT 1603.260 1000.000 1603.560 1000.010 ;
        RECT 1608.780 1000.000 1610.000 1000.010 ;
        RECT 1612.300 1000.000 1613.520 1000.010 ;
        RECT 1618.740 1000.000 1620.420 1000.010 ;
        RECT 1621.040 1000.000 1621.340 1000.010 ;
        RECT 1625.800 1000.010 1625.940 1016.270 ;
        RECT 1628.560 1012.850 1628.700 2499.950 ;
        RECT 1640.980 2484.710 1641.120 2500.000 ;
        RECT 1656.160 2499.950 1662.210 2500.000 ;
        RECT 1640.920 2484.390 1641.180 2484.710 ;
        RECT 1656.160 1016.930 1656.300 2499.950 ;
        RECT 1680.020 2489.490 1680.280 2489.810 ;
        RECT 1673.120 2485.410 1673.380 2485.730 ;
        RECT 1659.320 2484.390 1659.580 2484.710 ;
        RECT 1656.100 1016.610 1656.360 1016.930 ;
        RECT 1659.380 1013.190 1659.520 2484.390 ;
        RECT 1669.440 1814.590 1669.700 1814.910 ;
        RECT 1668.980 1735.030 1669.240 1735.350 ;
        RECT 1659.320 1012.870 1659.580 1013.190 ;
        RECT 1628.500 1012.530 1628.760 1012.850 ;
        RECT 1665.760 1012.190 1666.020 1012.510 ;
        RECT 1628.500 1011.850 1628.760 1012.170 ;
        RECT 1662.540 1011.850 1662.800 1012.170 ;
        RECT 1628.560 1000.010 1628.700 1011.850 ;
        RECT 1662.600 1000.010 1662.740 1011.850 ;
        RECT 1665.820 1000.010 1665.960 1012.190 ;
        RECT 1669.040 1000.690 1669.180 1735.030 ;
        RECT 1669.500 1012.510 1669.640 1814.590 ;
        RECT 1669.440 1012.190 1669.700 1012.510 ;
        RECT 1673.180 1010.130 1673.320 2485.410 ;
        RECT 1680.080 1016.250 1680.220 2489.490 ;
        RECT 1683.300 2484.710 1683.440 2500.000 ;
        RECT 1683.240 2484.390 1683.500 2484.710 ;
        RECT 1704.460 1017.270 1704.600 2500.000 ;
        RECT 1715.500 2485.730 1715.640 2500.000 ;
        RECT 1725.620 2486.750 1725.760 2500.000 ;
        RECT 1746.780 2489.810 1746.920 2500.000 ;
        RECT 1746.720 2489.490 1746.980 2489.810 ;
        RECT 1725.560 2486.430 1725.820 2486.750 ;
        RECT 1757.820 2486.410 1757.960 2500.000 ;
        RECT 1766.560 2499.950 1768.010 2500.000 ;
        RECT 1757.760 2486.090 1758.020 2486.410 ;
        RECT 1715.440 2485.410 1715.700 2485.730 ;
        RECT 1724.640 1928.490 1724.900 1928.810 ;
        RECT 1717.740 1925.770 1718.000 1926.090 ;
        RECT 1710.840 1736.390 1711.100 1736.710 ;
        RECT 1704.400 1016.950 1704.660 1017.270 ;
        RECT 1680.020 1015.930 1680.280 1016.250 ;
        RECT 1710.380 1012.870 1710.640 1013.190 ;
        RECT 1707.160 1012.190 1707.420 1012.510 ;
        RECT 1673.120 1009.810 1673.380 1010.130 ;
        RECT 1667.660 1000.550 1669.180 1000.690 ;
        RECT 1667.660 1000.010 1667.800 1000.550 ;
        RECT 1707.220 1000.010 1707.360 1012.190 ;
        RECT 1710.440 1000.010 1710.580 1012.870 ;
        RECT 1710.900 1012.510 1711.040 1736.390 ;
        RECT 1717.800 1012.510 1717.940 1925.770 ;
        RECT 1720.040 1013.210 1720.300 1013.530 ;
        RECT 1710.840 1012.190 1711.100 1012.510 ;
        RECT 1715.900 1012.190 1716.160 1012.510 ;
        RECT 1717.740 1012.190 1718.000 1012.510 ;
        RECT 1715.960 1000.010 1716.100 1012.190 ;
        RECT 1720.100 1000.010 1720.240 1013.210 ;
        RECT 1724.700 1000.010 1724.840 1928.490 ;
        RECT 1745.340 1927.470 1745.600 1927.790 ;
        RECT 1738.440 1926.110 1738.700 1926.430 ;
        RECT 1737.980 1849.270 1738.240 1849.590 ;
        RECT 1738.040 1012.510 1738.180 1849.270 ;
        RECT 1733.380 1012.190 1733.640 1012.510 ;
        RECT 1737.980 1012.190 1738.240 1012.510 ;
        RECT 1728.780 1010.490 1729.040 1010.810 ;
        RECT 1728.840 1000.010 1728.980 1010.490 ;
        RECT 1733.440 1000.010 1733.580 1012.190 ;
        RECT 1738.500 1000.690 1738.640 1926.110 ;
        RECT 1741.660 1012.870 1741.920 1013.190 ;
        RECT 1737.580 1000.550 1738.640 1000.690 ;
        RECT 1737.580 1000.010 1737.720 1000.550 ;
        RECT 1741.720 1000.010 1741.860 1012.870 ;
        RECT 1745.400 1000.010 1745.540 1927.470 ;
        RECT 1766.040 1926.790 1766.300 1927.110 ;
        RECT 1759.140 1883.610 1759.400 1883.930 ;
        RECT 1752.700 1736.730 1752.960 1737.050 ;
        RECT 1752.760 1690.810 1752.900 1736.730 ;
        RECT 1751.320 1690.490 1751.580 1690.810 ;
        RECT 1752.700 1690.490 1752.960 1690.810 ;
        RECT 1751.380 1656.210 1751.520 1690.490 ;
        RECT 1751.380 1656.070 1752.440 1656.210 ;
        RECT 1752.300 1013.530 1752.440 1656.070 ;
        RECT 1759.200 1014.210 1759.340 1883.610 ;
        RECT 1766.100 1014.210 1766.240 1926.790 ;
        RECT 1766.560 1017.610 1766.700 2499.950 ;
        RECT 1778.980 2489.470 1779.120 2500.000 ;
        RECT 1778.920 2489.150 1779.180 2489.470 ;
        RECT 1790.020 2489.130 1790.160 2500.000 ;
        RECT 1789.960 2488.810 1790.220 2489.130 ;
        RECT 1811.180 2486.070 1811.320 2500.000 ;
        RECT 1832.340 2487.090 1832.480 2500.000 ;
        RECT 1842.460 2488.790 1842.600 2500.000 ;
        RECT 1849.360 2499.950 1853.570 2500.000 ;
        RECT 1842.400 2488.470 1842.660 2488.790 ;
        RECT 1832.280 2486.770 1832.540 2487.090 ;
        RECT 1811.120 2485.750 1811.380 2486.070 ;
        RECT 1828.140 1927.810 1828.400 1928.130 ;
        RECT 1779.380 1927.130 1779.640 1927.450 ;
        RECT 1772.940 1766.310 1773.200 1766.630 ;
        RECT 1772.480 1735.710 1772.740 1736.030 ;
        RECT 1766.500 1017.290 1766.760 1017.610 ;
        RECT 1755.000 1013.890 1755.260 1014.210 ;
        RECT 1759.140 1013.890 1759.400 1014.210 ;
        RECT 1763.740 1013.890 1764.000 1014.210 ;
        RECT 1766.040 1013.890 1766.300 1014.210 ;
        RECT 1766.500 1013.890 1766.760 1014.210 ;
        RECT 1749.940 1013.210 1750.200 1013.530 ;
        RECT 1752.240 1013.210 1752.500 1013.530 ;
        RECT 1750.000 1000.010 1750.140 1013.210 ;
        RECT 1755.060 1000.010 1755.200 1013.890 ;
        RECT 1758.680 1013.210 1758.940 1013.530 ;
        RECT 1758.740 1000.010 1758.880 1013.210 ;
        RECT 1763.800 1000.010 1763.940 1013.890 ;
        RECT 1766.560 1013.530 1766.700 1013.890 ;
        RECT 1766.500 1013.210 1766.760 1013.530 ;
        RECT 1767.420 1012.870 1767.680 1013.190 ;
        RECT 1767.480 1010.810 1767.620 1012.870 ;
        RECT 1767.420 1010.490 1767.680 1010.810 ;
        RECT 1767.880 1010.490 1768.140 1010.810 ;
        RECT 1767.940 1000.010 1768.080 1010.490 ;
        RECT 1772.540 1000.010 1772.680 1735.710 ;
        RECT 1773.000 1010.810 1773.140 1766.310 ;
        RECT 1772.940 1010.490 1773.200 1010.810 ;
        RECT 1776.620 1007.430 1776.880 1007.750 ;
        RECT 1776.680 1000.010 1776.820 1007.430 ;
        RECT 1625.800 1000.000 1627.480 1000.010 ;
        RECT 1628.560 1000.000 1629.780 1000.010 ;
        RECT 1662.440 1000.000 1662.740 1000.010 ;
        RECT 1664.280 1000.000 1665.960 1000.010 ;
        RECT 1666.580 1000.000 1667.800 1000.010 ;
        RECT 1705.680 1000.000 1707.360 1000.010 ;
        RECT 1710.280 1000.000 1710.580 1000.010 ;
        RECT 1714.420 1000.000 1716.100 1000.010 ;
        RECT 1718.560 1000.000 1720.240 1000.010 ;
        RECT 1723.160 1000.000 1724.840 1000.010 ;
        RECT 1727.300 1000.000 1728.980 1000.010 ;
        RECT 1731.900 1000.000 1733.580 1000.010 ;
        RECT 1736.040 1000.000 1737.720 1000.010 ;
        RECT 1740.640 1000.000 1741.860 1000.010 ;
        RECT 1744.780 1000.000 1745.540 1000.010 ;
        RECT 1749.380 1000.000 1750.140 1000.010 ;
        RECT 1753.520 1000.000 1755.200 1000.010 ;
        RECT 1758.120 1000.000 1758.880 1000.010 ;
        RECT 1762.260 1000.000 1763.940 1000.010 ;
        RECT 1766.400 1000.000 1768.080 1000.010 ;
        RECT 1771.000 1000.000 1772.680 1000.010 ;
        RECT 1775.140 1000.000 1776.820 1000.010 ;
        RECT 1779.440 1000.010 1779.580 1927.130 ;
        RECT 1786.740 1926.450 1787.000 1926.770 ;
        RECT 1779.840 1925.430 1780.100 1925.750 ;
        RECT 1779.900 1007.750 1780.040 1925.430 ;
        RECT 1779.840 1007.430 1780.100 1007.750 ;
        RECT 1786.800 1000.690 1786.940 1926.450 ;
        RECT 1821.240 1870.010 1821.500 1870.330 ;
        RECT 1800.540 1738.090 1800.800 1738.410 ;
        RECT 1793.640 1737.750 1793.900 1738.070 ;
        RECT 1789.500 1010.150 1789.760 1010.470 ;
        RECT 1785.420 1000.550 1786.940 1000.690 ;
        RECT 1785.420 1000.010 1785.560 1000.550 ;
        RECT 1789.560 1000.010 1789.700 1010.150 ;
        RECT 1793.700 1000.010 1793.840 1737.750 ;
        RECT 1800.600 1007.750 1800.740 1738.090 ;
        RECT 1814.340 1737.410 1814.600 1737.730 ;
        RECT 1813.880 1737.070 1814.140 1737.390 ;
        RECT 1807.440 1736.050 1807.700 1736.370 ;
        RECT 1806.980 1735.370 1807.240 1735.690 ;
        RECT 1807.040 1007.750 1807.180 1735.370 ;
        RECT 1798.240 1007.430 1798.500 1007.750 ;
        RECT 1800.540 1007.430 1800.800 1007.750 ;
        RECT 1802.840 1007.430 1803.100 1007.750 ;
        RECT 1806.980 1007.430 1807.240 1007.750 ;
        RECT 1798.300 1000.010 1798.440 1007.430 ;
        RECT 1802.900 1000.010 1803.040 1007.430 ;
        RECT 1807.500 1000.690 1807.640 1736.050 ;
        RECT 1813.940 1007.750 1814.080 1737.070 ;
        RECT 1811.580 1007.430 1811.840 1007.750 ;
        RECT 1813.880 1007.430 1814.140 1007.750 ;
        RECT 1807.040 1000.550 1807.640 1000.690 ;
        RECT 1807.040 1000.010 1807.180 1000.550 ;
        RECT 1811.640 1000.010 1811.780 1007.430 ;
        RECT 1814.400 1000.010 1814.540 1737.410 ;
        RECT 1821.300 1000.690 1821.440 1870.010 ;
        RECT 1827.680 1738.430 1827.940 1738.750 ;
        RECT 1827.740 1010.810 1827.880 1738.430 ;
        RECT 1824.460 1010.490 1824.720 1010.810 ;
        RECT 1827.680 1010.490 1827.940 1010.810 ;
        RECT 1820.380 1000.550 1821.440 1000.690 ;
        RECT 1820.380 1000.010 1820.520 1000.550 ;
        RECT 1824.520 1000.010 1824.660 1010.490 ;
        RECT 1828.200 1010.210 1828.340 1927.810 ;
        RECT 1835.040 1925.090 1835.300 1925.410 ;
        RECT 1835.100 1010.810 1835.240 1925.090 ;
        RECT 1849.360 1018.290 1849.500 2499.950 ;
        RECT 1874.660 2488.110 1874.800 2500.000 ;
        RECT 1876.440 2493.910 1876.700 2494.230 ;
        RECT 1874.600 2487.790 1874.860 2488.110 ;
        RECT 1849.300 1017.970 1849.560 1018.290 ;
        RECT 1876.500 1011.150 1876.640 2493.910 ;
        RECT 1885.700 2488.450 1885.840 2500.000 ;
        RECT 1885.640 2488.130 1885.900 2488.450 ;
        RECT 1886.160 1020.330 1886.300 2896.390 ;
        RECT 1886.100 1020.010 1886.360 1020.330 ;
        RECT 1878.280 1013.550 1878.540 1013.870 ;
        RECT 1878.740 1013.550 1879.000 1013.870 ;
        RECT 1878.340 1011.830 1878.480 1013.550 ;
        RECT 1878.280 1011.510 1878.540 1011.830 ;
        RECT 1871.840 1010.830 1872.100 1011.150 ;
        RECT 1872.300 1010.830 1872.560 1011.150 ;
        RECT 1876.440 1010.830 1876.700 1011.150 ;
        RECT 1830.900 1010.490 1831.160 1010.810 ;
        RECT 1835.040 1010.490 1835.300 1010.810 ;
        RECT 1826.820 1010.070 1828.340 1010.210 ;
        RECT 1826.820 1000.010 1826.960 1010.070 ;
        RECT 1830.960 1000.010 1831.100 1010.490 ;
        RECT 1834.580 1009.810 1834.840 1010.130 ;
        RECT 1834.640 1000.010 1834.780 1009.810 ;
        RECT 1871.900 1009.790 1872.040 1010.830 ;
        RECT 1871.840 1009.470 1872.100 1009.790 ;
        RECT 1872.360 1000.010 1872.500 1010.830 ;
        RECT 1878.800 1000.010 1878.940 1013.550 ;
        RECT 1886.620 1011.830 1886.760 2912.450 ;
        RECT 1887.480 2912.110 1887.740 2912.430 ;
        RECT 1887.540 2494.570 1887.680 2912.110 ;
        RECT 1888.000 2494.910 1888.140 2912.790 ;
        RECT 1894.840 2896.470 1895.100 2896.790 ;
        RECT 1890.690 2848.335 1890.970 2848.705 ;
        RECT 1887.940 2494.590 1888.200 2494.910 ;
        RECT 1887.480 2494.250 1887.740 2494.570 ;
        RECT 1890.760 1021.010 1890.900 2848.335 ;
        RECT 1891.150 2832.015 1891.430 2832.385 ;
        RECT 1891.220 1024.750 1891.360 2832.015 ;
        RECT 1891.610 2817.055 1891.890 2817.425 ;
        RECT 1891.680 1025.090 1891.820 2817.055 ;
        RECT 1892.070 2797.675 1892.350 2798.045 ;
        RECT 1891.620 1024.770 1891.880 1025.090 ;
        RECT 1891.160 1024.430 1891.420 1024.750 ;
        RECT 1890.700 1020.690 1890.960 1021.010 ;
        RECT 1886.560 1011.510 1886.820 1011.830 ;
        RECT 1892.140 1011.005 1892.280 2797.675 ;
        RECT 1892.990 2782.715 1893.270 2783.085 ;
        RECT 1892.530 2608.635 1892.810 2609.005 ;
        RECT 1892.600 1011.490 1892.740 2608.635 ;
        RECT 1893.060 1459.610 1893.200 2782.715 ;
        RECT 1893.920 2780.870 1894.180 2781.190 ;
        RECT 1893.450 2753.475 1893.730 2753.845 ;
        RECT 1893.520 1459.950 1893.660 2753.475 ;
        RECT 1893.460 1459.630 1893.720 1459.950 ;
        RECT 1893.000 1459.290 1893.260 1459.610 ;
        RECT 1893.980 1013.870 1894.120 2780.870 ;
        RECT 1894.370 2735.115 1894.650 2735.485 ;
        RECT 1894.440 1459.270 1894.580 2735.115 ;
        RECT 1894.900 2495.250 1895.040 2896.470 ;
        RECT 1895.360 2495.590 1895.500 2913.130 ;
        RECT 2094.020 2781.210 2094.280 2781.530 ;
        RECT 2556.320 2781.210 2556.580 2781.530 ;
        RECT 1897.590 2767.075 1897.870 2767.445 ;
        RECT 1895.300 2495.270 1895.560 2495.590 ;
        RECT 1894.840 2494.930 1895.100 2495.250 ;
        RECT 1894.380 1458.950 1894.640 1459.270 ;
        RECT 1897.660 1019.650 1897.800 2767.075 ;
        RECT 1898.050 2718.795 1898.330 2719.165 ;
        RECT 1897.600 1019.330 1897.860 1019.650 ;
        RECT 1898.120 1018.630 1898.260 2718.795 ;
        RECT 1898.510 2687.515 1898.790 2687.885 ;
        RECT 1898.060 1018.310 1898.320 1018.630 ;
        RECT 1893.920 1013.550 1894.180 1013.870 ;
        RECT 1892.540 1011.170 1892.800 1011.490 ;
        RECT 1898.580 1011.150 1898.720 2687.515 ;
        RECT 1898.970 2672.555 1899.250 2672.925 ;
        RECT 1899.040 1018.970 1899.180 2672.555 ;
        RECT 1899.430 2656.915 1899.710 2657.285 ;
        RECT 1898.980 1018.650 1899.240 1018.970 ;
        RECT 1899.500 1017.950 1899.640 2656.915 ;
        RECT 1899.890 2624.955 1900.170 2625.325 ;
        RECT 1899.440 1017.630 1899.700 1017.950 ;
        RECT 1882.420 1010.490 1882.680 1010.810 ;
        RECT 1892.070 1010.635 1892.350 1011.005 ;
        RECT 1898.520 1010.830 1898.780 1011.150 ;
        RECT 1882.480 1000.010 1882.620 1010.490 ;
        RECT 1899.960 1009.790 1900.100 2624.955 ;
        RECT 1900.350 2577.355 1900.630 2577.725 ;
        RECT 1900.420 1021.350 1900.560 2577.355 ;
        RECT 1900.810 2562.395 1901.090 2562.765 ;
        RECT 1900.360 1021.030 1900.620 1021.350 ;
        RECT 1900.880 1020.670 1901.020 2562.395 ;
        RECT 1901.270 2547.435 1901.550 2547.805 ;
        RECT 1900.820 1020.350 1901.080 1020.670 ;
        RECT 1901.340 1019.310 1901.480 2547.435 ;
        RECT 1903.570 2514.795 1903.850 2515.165 ;
        RECT 1903.640 1019.990 1903.780 2514.795 ;
        RECT 2083.440 1946.510 2083.700 1946.830 ;
        RECT 2082.980 1945.830 2083.240 1946.150 ;
        RECT 2044.340 1928.490 2044.600 1928.810 ;
        RECT 1964.300 1927.810 1964.560 1928.130 ;
        RECT 1929.340 1927.470 1929.600 1927.790 ;
        RECT 1929.400 1917.095 1929.540 1927.470 ;
        RECT 1952.340 1925.090 1952.600 1925.410 ;
        RECT 1952.400 1917.095 1952.540 1925.090 ;
        RECT 1964.360 1917.095 1964.500 1927.810 ;
        RECT 1998.340 1927.130 1998.600 1927.450 ;
        RECT 1987.300 1926.110 1987.560 1926.430 ;
        RECT 1975.340 1925.770 1975.600 1926.090 ;
        RECT 1975.400 1917.095 1975.540 1925.770 ;
        RECT 1987.360 1917.095 1987.500 1926.110 ;
        RECT 1998.400 1917.095 1998.540 1927.130 ;
        RECT 2010.300 1926.790 2010.560 1927.110 ;
        RECT 2010.360 1917.095 2010.500 1926.790 ;
        RECT 2033.300 1926.450 2033.560 1926.770 ;
        RECT 2033.360 1917.095 2033.500 1926.450 ;
        RECT 2044.400 1917.095 2044.540 1928.490 ;
        RECT 2067.340 1925.430 2067.600 1925.750 ;
        RECT 2067.400 1917.095 2067.540 1925.430 ;
        RECT 1929.290 1913.095 1929.570 1917.095 ;
        RECT 1952.290 1913.095 1952.570 1917.095 ;
        RECT 1964.250 1913.095 1964.530 1917.095 ;
        RECT 1975.290 1913.095 1975.570 1917.095 ;
        RECT 1987.250 1913.095 1987.530 1917.095 ;
        RECT 1998.290 1913.095 1998.570 1917.095 ;
        RECT 2010.250 1913.095 2010.530 1917.095 ;
        RECT 2033.250 1913.095 2033.530 1917.095 ;
        RECT 2044.290 1913.095 2044.570 1917.095 ;
        RECT 2067.290 1913.095 2067.570 1917.095 ;
      LAYER met2 ;
        RECT 1922.860 1912.815 1929.010 1913.095 ;
        RECT 1929.850 1912.815 1940.970 1913.095 ;
        RECT 1941.810 1912.815 1952.010 1913.095 ;
        RECT 1952.850 1912.815 1963.970 1913.095 ;
        RECT 1964.810 1912.815 1975.010 1913.095 ;
        RECT 1975.850 1912.815 1986.970 1913.095 ;
        RECT 1987.810 1912.815 1998.010 1913.095 ;
        RECT 1998.850 1912.815 2009.970 1913.095 ;
        RECT 2010.810 1912.815 2021.010 1913.095 ;
        RECT 2021.850 1912.815 2032.970 1913.095 ;
        RECT 2033.810 1912.815 2044.010 1913.095 ;
        RECT 2044.850 1912.815 2055.970 1913.095 ;
        RECT 2056.810 1912.815 2067.010 1913.095 ;
        RECT 2067.850 1912.815 2072.160 1913.095 ;
      LAYER met2 ;
        RECT 1904.490 1885.795 1904.770 1886.165 ;
        RECT 1904.560 1883.930 1904.700 1885.795 ;
        RECT 1904.500 1883.610 1904.760 1883.930 ;
        RECT 1904.490 1870.155 1904.770 1870.525 ;
        RECT 1904.500 1870.010 1904.760 1870.155 ;
        RECT 1904.490 1851.795 1904.770 1852.165 ;
        RECT 1904.560 1849.590 1904.700 1851.795 ;
        RECT 1904.500 1849.270 1904.760 1849.590 ;
        RECT 1904.490 1817.795 1904.770 1818.165 ;
        RECT 1904.560 1814.910 1904.700 1817.795 ;
        RECT 1904.500 1814.590 1904.760 1814.910 ;
        RECT 1904.490 1767.475 1904.770 1767.845 ;
        RECT 1904.560 1766.630 1904.700 1767.475 ;
        RECT 1904.500 1766.310 1904.760 1766.630 ;
      LAYER met2 ;
        RECT 1922.860 1754.280 2072.160 1912.815 ;
      LAYER met2 ;
        RECT 2073.320 1870.010 2073.580 1870.330 ;
      LAYER met2 ;
        RECT 1923.410 1754.000 1933.610 1754.280 ;
        RECT 1934.450 1754.000 1944.650 1754.280 ;
        RECT 1945.490 1754.000 1956.610 1754.280 ;
        RECT 1957.450 1754.000 1967.650 1754.280 ;
        RECT 1968.490 1754.000 1979.610 1754.280 ;
        RECT 1980.450 1754.000 1990.650 1754.280 ;
        RECT 1991.490 1754.000 2002.610 1754.280 ;
        RECT 2003.450 1754.000 2013.650 1754.280 ;
        RECT 2014.490 1754.000 2025.610 1754.280 ;
        RECT 2026.450 1754.000 2036.650 1754.280 ;
        RECT 2037.490 1754.000 2048.610 1754.280 ;
        RECT 2049.450 1754.000 2059.650 1754.280 ;
        RECT 2060.490 1754.000 2071.610 1754.280 ;
      LAYER met2 ;
        RECT 1933.890 1750.000 1934.170 1754.000 ;
        RECT 1944.930 1750.000 1945.210 1754.000 ;
        RECT 1956.890 1750.000 1957.170 1754.000 ;
        RECT 1967.930 1750.000 1968.210 1754.000 ;
        RECT 1979.890 1750.000 1980.170 1754.000 ;
        RECT 1990.930 1750.000 1991.210 1754.000 ;
        RECT 2002.890 1750.000 2003.170 1754.000 ;
        RECT 2013.930 1750.000 2014.210 1754.000 ;
        RECT 2036.930 1750.000 2037.210 1754.000 ;
        RECT 2059.930 1750.000 2060.210 1754.000 ;
        RECT 2071.890 1750.000 2072.170 1754.000 ;
        RECT 1934.000 1738.750 1934.140 1750.000 ;
        RECT 1933.940 1738.430 1934.200 1738.750 ;
        RECT 1945.040 1736.710 1945.180 1750.000 ;
        RECT 1957.000 1738.410 1957.140 1750.000 ;
        RECT 1956.940 1738.090 1957.200 1738.410 ;
        RECT 1968.040 1738.070 1968.180 1750.000 ;
        RECT 1967.980 1737.750 1968.240 1738.070 ;
        RECT 1980.000 1737.050 1980.140 1750.000 ;
        RECT 1991.040 1737.730 1991.180 1750.000 ;
        RECT 1990.980 1737.410 1991.240 1737.730 ;
        RECT 1979.940 1736.730 1980.200 1737.050 ;
        RECT 1944.980 1736.390 1945.240 1736.710 ;
        RECT 2003.000 1736.030 2003.140 1750.000 ;
        RECT 2014.040 1737.390 2014.180 1750.000 ;
        RECT 2013.980 1737.070 2014.240 1737.390 ;
        RECT 2037.040 1736.370 2037.180 1750.000 ;
        RECT 2036.980 1736.050 2037.240 1736.370 ;
        RECT 2002.940 1735.710 2003.200 1736.030 ;
        RECT 2060.040 1735.350 2060.180 1750.000 ;
        RECT 2072.000 1735.690 2072.140 1750.000 ;
        RECT 2071.940 1735.370 2072.200 1735.690 ;
        RECT 2059.980 1735.030 2060.240 1735.350 ;
        RECT 2007.540 1687.770 2007.800 1688.090 ;
        RECT 1903.580 1019.670 1903.840 1019.990 ;
        RECT 1901.280 1018.990 1901.540 1019.310 ;
        RECT 2007.600 1013.870 2007.740 1687.770 ;
        RECT 2055.840 1687.430 2056.100 1687.750 ;
        RECT 2042.040 1687.090 2042.300 1687.410 ;
        RECT 2002.940 1013.550 2003.200 1013.870 ;
        RECT 2007.540 1013.550 2007.800 1013.870 ;
        RECT 2008.000 1013.550 2008.260 1013.870 ;
        RECT 1899.900 1009.470 1900.160 1009.790 ;
        RECT 2003.000 1000.010 2003.140 1013.550 ;
        RECT 2008.060 1012.930 2008.200 1013.550 ;
        RECT 2007.600 1012.790 2008.200 1012.930 ;
        RECT 2007.600 1007.750 2007.740 1012.790 ;
        RECT 2004.780 1007.430 2005.040 1007.750 ;
        RECT 2007.540 1007.430 2007.800 1007.750 ;
        RECT 2004.840 1000.010 2004.980 1007.430 ;
        RECT 2042.100 1000.010 2042.240 1687.090 ;
        RECT 2055.900 1011.830 2056.040 1687.430 ;
        RECT 2069.640 1686.750 2069.900 1687.070 ;
        RECT 2065.040 1013.890 2065.300 1014.210 ;
        RECT 2065.500 1013.890 2065.760 1014.210 ;
        RECT 2065.100 1013.530 2065.240 1013.890 ;
        RECT 2064.580 1013.210 2064.840 1013.530 ;
        RECT 2065.040 1013.210 2065.300 1013.530 ;
        RECT 2064.640 1012.510 2064.780 1013.210 ;
        RECT 2064.120 1012.190 2064.380 1012.510 ;
        RECT 2064.580 1012.190 2064.840 1012.510 ;
        RECT 2050.780 1011.510 2051.040 1011.830 ;
        RECT 2055.840 1011.510 2056.100 1011.830 ;
        RECT 2046.180 1010.830 2046.440 1011.150 ;
        RECT 2046.240 1000.010 2046.380 1010.830 ;
        RECT 2050.840 1000.010 2050.980 1011.510 ;
        RECT 2055.380 1011.170 2055.640 1011.490 ;
        RECT 1779.440 1000.000 1779.740 1000.010 ;
        RECT 1783.880 1000.000 1785.560 1000.010 ;
        RECT 1788.480 1000.000 1789.700 1000.010 ;
        RECT 1792.620 1000.000 1793.840 1000.010 ;
        RECT 1797.220 1000.000 1798.440 1000.010 ;
        RECT 1801.360 1000.000 1803.040 1000.010 ;
        RECT 1805.960 1000.000 1807.180 1000.010 ;
        RECT 1810.100 1000.000 1811.780 1000.010 ;
        RECT 1814.240 1000.000 1814.540 1000.010 ;
        RECT 1818.840 1000.000 1820.520 1000.010 ;
        RECT 1822.980 1000.000 1824.660 1000.010 ;
        RECT 1825.280 1000.000 1826.960 1000.010 ;
        RECT 1829.880 1000.000 1831.100 1000.010 ;
        RECT 1834.020 1000.000 1834.780 1000.010 ;
        RECT 1870.820 1000.000 1872.500 1000.010 ;
        RECT 1877.260 1000.000 1878.940 1000.010 ;
        RECT 1881.860 1000.000 1882.620 1000.010 ;
        RECT 2001.460 1000.000 2003.140 1000.010 ;
        RECT 2003.760 1000.000 2004.980 1000.010 ;
        RECT 2040.560 1000.000 2042.240 1000.010 ;
        RECT 2044.700 1000.000 2046.380 1000.010 ;
        RECT 2049.300 1000.000 2050.980 1000.010 ;
        RECT 2055.440 1000.010 2055.580 1011.170 ;
        RECT 2061.360 1009.470 2061.620 1009.790 ;
        RECT 2061.420 1000.010 2061.560 1009.470 ;
        RECT 2064.180 1009.450 2064.320 1012.190 ;
        RECT 2064.120 1009.130 2064.380 1009.450 ;
        RECT 2065.560 1000.010 2065.700 1013.890 ;
        RECT 2069.700 1000.010 2069.840 1686.750 ;
        RECT 2073.380 1014.210 2073.520 1870.010 ;
        RECT 2073.320 1013.890 2073.580 1014.210 ;
        RECT 2075.160 1013.890 2075.420 1014.210 ;
        RECT 2075.220 1012.170 2075.360 1013.890 ;
        RECT 2075.160 1011.850 2075.420 1012.170 ;
        RECT 2078.840 1011.850 2079.100 1012.170 ;
        RECT 2074.700 1010.150 2074.960 1010.470 ;
        RECT 2073.320 1009.810 2073.580 1010.130 ;
        RECT 2073.380 1009.110 2073.520 1009.810 ;
        RECT 2073.320 1008.790 2073.580 1009.110 ;
        RECT 2074.760 1000.010 2074.900 1010.150 ;
        RECT 2078.900 1000.010 2079.040 1011.850 ;
        RECT 2083.040 1000.010 2083.180 1945.830 ;
        RECT 2083.500 1012.170 2083.640 1946.510 ;
        RECT 2090.340 1946.170 2090.600 1946.490 ;
        RECT 2087.110 1884.435 2087.390 1884.805 ;
        RECT 2084.350 1850.435 2084.630 1850.805 ;
        RECT 2084.420 1012.850 2084.560 1850.435 ;
        RECT 2084.810 1835.475 2085.090 1835.845 ;
        RECT 2084.360 1012.530 2084.620 1012.850 ;
        RECT 2083.440 1011.850 2083.700 1012.170 ;
        RECT 2084.880 1010.130 2085.020 1835.475 ;
        RECT 2085.270 1816.435 2085.550 1816.805 ;
        RECT 2084.820 1009.810 2085.080 1010.130 ;
        RECT 2085.340 1009.450 2085.480 1816.435 ;
        RECT 2085.730 1800.795 2086.010 1801.165 ;
        RECT 2085.800 1013.190 2085.940 1800.795 ;
        RECT 2086.190 1782.435 2086.470 1782.805 ;
        RECT 2085.740 1012.870 2086.000 1013.190 ;
        RECT 2086.260 1012.510 2086.400 1782.435 ;
        RECT 2086.650 1766.795 2086.930 1767.165 ;
        RECT 2086.720 1013.530 2086.860 1766.795 ;
        RECT 2087.180 1014.210 2087.320 1884.435 ;
        RECT 2090.400 1014.210 2090.540 1946.170 ;
        RECT 2087.120 1013.890 2087.380 1014.210 ;
        RECT 2087.580 1013.890 2087.840 1014.210 ;
        RECT 2090.340 1013.890 2090.600 1014.210 ;
        RECT 2086.660 1013.210 2086.920 1013.530 ;
        RECT 2086.200 1012.190 2086.460 1012.510 ;
        RECT 2085.740 1011.510 2086.000 1011.830 ;
        RECT 2085.800 1010.470 2085.940 1011.510 ;
        RECT 2085.740 1010.150 2086.000 1010.470 ;
        RECT 2085.280 1009.130 2085.540 1009.450 ;
        RECT 2087.640 1000.010 2087.780 1013.890 ;
        RECT 2094.080 1009.110 2094.220 2781.210 ;
        RECT 2422.000 2780.870 2422.260 2781.190 ;
        RECT 2422.060 2773.820 2422.200 2780.870 ;
        RECT 2556.380 2773.820 2556.520 2781.210 ;
        RECT 2422.060 2773.380 2422.380 2773.820 ;
        RECT 2556.380 2773.380 2556.700 2773.820 ;
        RECT 2422.100 2769.820 2422.380 2773.380 ;
        RECT 2556.420 2769.820 2556.700 2773.380 ;
      LAYER met2 ;
        RECT 2400.030 2769.540 2421.820 2769.820 ;
        RECT 2422.660 2769.540 2556.140 2769.820 ;
        RECT 2400.030 2604.280 2556.690 2769.540 ;
        RECT 2400.580 2604.000 2534.060 2604.280 ;
        RECT 2534.900 2604.000 2556.690 2604.280 ;
      LAYER met2 ;
        RECT 2400.020 2600.730 2400.300 2604.000 ;
        RECT 2394.460 2600.590 2400.300 2600.730 ;
        RECT 2534.340 2600.660 2534.620 2604.000 ;
        RECT 2394.460 2494.230 2394.600 2600.590 ;
        RECT 2400.020 2600.000 2400.300 2600.590 ;
        RECT 2534.300 2600.000 2534.620 2600.660 ;
        RECT 2534.300 2587.730 2534.440 2600.000 ;
        RECT 2528.720 2587.410 2528.980 2587.730 ;
        RECT 2534.240 2587.410 2534.500 2587.730 ;
        RECT 2394.400 2493.910 2394.660 2494.230 ;
        RECT 2294.120 1946.850 2294.380 1947.170 ;
        RECT 2379.220 1946.850 2379.480 1947.170 ;
        RECT 2283.990 1875.595 2284.270 1875.965 ;
        RECT 2284.060 1870.330 2284.200 1875.595 ;
        RECT 2284.000 1870.010 2284.260 1870.330 ;
        RECT 2287.210 1789.915 2287.490 1790.285 ;
        RECT 2287.280 1009.790 2287.420 1789.915 ;
        RECT 2294.180 1013.870 2294.320 1946.850 ;
        RECT 2321.260 1946.510 2321.520 1946.830 ;
        RECT 2321.320 1937.745 2321.460 1946.510 ;
        RECT 2379.280 1937.745 2379.420 1946.850 ;
        RECT 2437.180 1946.170 2437.440 1946.490 ;
        RECT 2437.240 1937.745 2437.380 1946.170 ;
        RECT 2495.140 1945.830 2495.400 1946.150 ;
        RECT 2495.200 1937.745 2495.340 1945.830 ;
        RECT 2321.250 1933.745 2321.530 1937.745 ;
        RECT 2379.210 1933.745 2379.490 1937.745 ;
        RECT 2437.170 1933.745 2437.450 1937.745 ;
        RECT 2495.130 1933.745 2495.410 1937.745 ;
      LAYER met2 ;
        RECT 2302.860 1933.465 2320.970 1933.745 ;
        RECT 2321.810 1933.465 2378.930 1933.745 ;
        RECT 2379.770 1933.465 2436.890 1933.745 ;
        RECT 2437.730 1933.465 2494.850 1933.745 ;
        RECT 2495.690 1933.465 2514.720 1933.745 ;
        RECT 2302.860 1704.280 2514.720 1933.465 ;
      LAYER met2 ;
        RECT 2523.650 1892.170 2523.930 1892.285 ;
        RECT 2518.660 1892.030 2523.930 1892.170 ;
        RECT 2518.660 1807.170 2518.800 1892.030 ;
        RECT 2523.650 1891.915 2523.930 1892.030 ;
        RECT 2518.200 1807.030 2518.800 1807.170 ;
        RECT 2518.200 1800.370 2518.340 1807.030 ;
        RECT 2523.650 1802.410 2523.930 1802.525 ;
        RECT 2521.880 1802.270 2523.930 1802.410 ;
        RECT 2518.200 1800.230 2518.800 1800.370 ;
        RECT 2518.660 1799.690 2518.800 1800.230 ;
        RECT 2518.660 1799.550 2519.260 1799.690 ;
        RECT 2519.120 1752.770 2519.260 1799.550 ;
        RECT 2521.880 1759.570 2522.020 1802.270 ;
        RECT 2523.650 1802.155 2523.930 1802.270 ;
        RECT 2520.500 1759.430 2522.020 1759.570 ;
        RECT 2520.500 1752.770 2520.640 1759.430 ;
        RECT 2519.120 1752.630 2520.180 1752.770 ;
        RECT 2520.500 1752.630 2521.100 1752.770 ;
        RECT 2520.040 1724.890 2520.180 1752.630 ;
        RECT 2519.580 1724.750 2520.180 1724.890 ;
        RECT 2519.060 1709.870 2519.320 1710.190 ;
      LAYER met2 ;
        RECT 2303.410 1704.000 2360.530 1704.280 ;
        RECT 2361.370 1704.000 2418.490 1704.280 ;
        RECT 2419.330 1704.000 2476.450 1704.280 ;
        RECT 2477.290 1704.000 2514.720 1704.280 ;
      LAYER met2 ;
        RECT 2518.590 1704.235 2518.870 1704.605 ;
        RECT 2302.850 1700.000 2303.130 1704.000 ;
        RECT 2360.810 1700.000 2361.090 1704.000 ;
        RECT 2418.770 1700.000 2419.050 1704.000 ;
        RECT 2476.730 1700.000 2477.010 1704.000 ;
        RECT 2302.920 1688.090 2303.060 1700.000 ;
        RECT 2302.860 1687.770 2303.120 1688.090 ;
        RECT 2360.880 1687.750 2361.020 1700.000 ;
        RECT 2360.820 1687.430 2361.080 1687.750 ;
        RECT 2418.840 1687.410 2418.980 1700.000 ;
        RECT 2418.780 1687.090 2419.040 1687.410 ;
        RECT 2476.800 1687.070 2476.940 1700.000 ;
        RECT 2476.740 1686.750 2477.000 1687.070 ;
        RECT 2518.660 1656.890 2518.800 1704.235 ;
        RECT 2518.200 1656.750 2518.800 1656.890 ;
        RECT 2518.200 1656.130 2518.340 1656.750 ;
        RECT 2518.140 1655.810 2518.400 1656.130 ;
        RECT 2519.120 1655.530 2519.260 1709.870 ;
        RECT 2519.580 1704.605 2519.720 1724.750 ;
        RECT 2520.960 1710.190 2521.100 1752.630 ;
        RECT 2523.650 1717.835 2523.930 1718.205 ;
        RECT 2520.900 1709.870 2521.160 1710.190 ;
        RECT 2519.510 1704.235 2519.790 1704.605 ;
        RECT 2523.720 1704.410 2523.860 1717.835 ;
        RECT 2523.660 1704.090 2523.920 1704.410 ;
        RECT 2519.520 1703.750 2519.780 1704.070 ;
        RECT 2518.660 1655.390 2519.260 1655.530 ;
        RECT 2518.660 1642.190 2518.800 1655.390 ;
        RECT 2517.680 1641.870 2517.940 1642.190 ;
        RECT 2518.600 1641.870 2518.860 1642.190 ;
        RECT 2517.740 1594.250 2517.880 1641.870 ;
        RECT 2519.580 1608.725 2519.720 1703.750 ;
        RECT 2519.980 1655.810 2520.240 1656.130 ;
        RECT 2520.040 1618.050 2520.180 1655.810 ;
        RECT 2519.980 1617.730 2520.240 1618.050 ;
        RECT 2520.900 1617.730 2521.160 1618.050 ;
        RECT 2519.510 1608.355 2519.790 1608.725 ;
        RECT 2519.510 1606.995 2519.790 1607.365 ;
        RECT 2517.680 1593.930 2517.940 1594.250 ;
        RECT 2518.600 1593.930 2518.860 1594.250 ;
        RECT 2518.660 1569.770 2518.800 1593.930 ;
        RECT 2517.220 1569.450 2517.480 1569.770 ;
        RECT 2518.600 1569.450 2518.860 1569.770 ;
        RECT 2517.280 1545.970 2517.420 1569.450 ;
        RECT 2518.140 1559.250 2518.400 1559.570 ;
        RECT 2518.200 1558.890 2518.340 1559.250 ;
        RECT 2518.140 1558.570 2518.400 1558.890 ;
        RECT 2517.220 1545.650 2517.480 1545.970 ;
        RECT 2519.060 1545.650 2519.320 1545.970 ;
        RECT 2519.120 1462.410 2519.260 1545.650 ;
        RECT 2518.660 1462.270 2519.260 1462.410 ;
        RECT 2518.660 1415.410 2518.800 1462.270 ;
        RECT 2518.600 1415.090 2518.860 1415.410 ;
        RECT 2519.060 1414.750 2519.320 1415.070 ;
        RECT 2518.140 1366.470 2518.400 1366.790 ;
        RECT 2518.200 1366.110 2518.340 1366.470 ;
        RECT 2518.140 1365.790 2518.400 1366.110 ;
        RECT 2518.600 1318.190 2518.860 1318.510 ;
        RECT 2518.660 1317.830 2518.800 1318.190 ;
        RECT 2518.600 1317.510 2518.860 1317.830 ;
        RECT 2518.140 1269.910 2518.400 1270.230 ;
        RECT 2518.200 1269.550 2518.340 1269.910 ;
        RECT 2518.140 1269.230 2518.400 1269.550 ;
        RECT 2519.120 1269.290 2519.260 1414.750 ;
        RECT 2518.660 1269.150 2519.260 1269.290 ;
        RECT 2518.660 1222.290 2518.800 1269.150 ;
        RECT 2518.600 1221.970 2518.860 1222.290 ;
        RECT 2519.060 1221.630 2519.320 1221.950 ;
        RECT 2518.140 1173.350 2518.400 1173.670 ;
        RECT 2518.200 1172.990 2518.340 1173.350 ;
        RECT 2518.140 1172.670 2518.400 1172.990 ;
        RECT 2519.120 1172.730 2519.260 1221.630 ;
        RECT 2518.660 1172.590 2519.260 1172.730 ;
        RECT 2518.660 1125.730 2518.800 1172.590 ;
        RECT 2518.600 1125.410 2518.860 1125.730 ;
        RECT 2519.060 1125.070 2519.320 1125.390 ;
        RECT 2518.140 1076.790 2518.400 1077.110 ;
        RECT 2518.200 1076.430 2518.340 1076.790 ;
        RECT 2518.140 1076.110 2518.400 1076.430 ;
        RECT 2519.120 1076.170 2519.260 1125.070 ;
        RECT 2518.660 1076.030 2519.260 1076.170 ;
        RECT 2518.660 1029.170 2518.800 1076.030 ;
        RECT 2518.600 1028.850 2518.860 1029.170 ;
        RECT 2519.060 1028.510 2519.320 1028.830 ;
        RECT 2518.600 1028.170 2518.860 1028.490 ;
        RECT 2294.120 1013.550 2294.380 1013.870 ;
        RECT 2518.660 1011.150 2518.800 1028.170 ;
        RECT 2519.120 1011.490 2519.260 1028.510 ;
        RECT 2519.580 1011.830 2519.720 1606.995 ;
        RECT 2520.960 1594.250 2521.100 1617.730 ;
        RECT 2519.980 1593.930 2520.240 1594.250 ;
        RECT 2520.900 1593.930 2521.160 1594.250 ;
        RECT 2520.040 1559.570 2520.180 1593.930 ;
        RECT 2519.980 1559.250 2520.240 1559.570 ;
        RECT 2519.980 1558.570 2520.240 1558.890 ;
        RECT 2520.040 1366.790 2520.180 1558.570 ;
        RECT 2519.980 1366.470 2520.240 1366.790 ;
        RECT 2519.980 1365.790 2520.240 1366.110 ;
        RECT 2520.040 1318.510 2520.180 1365.790 ;
        RECT 2519.980 1318.190 2520.240 1318.510 ;
        RECT 2519.980 1317.510 2520.240 1317.830 ;
        RECT 2520.040 1270.230 2520.180 1317.510 ;
        RECT 2519.980 1269.910 2520.240 1270.230 ;
        RECT 2519.980 1269.230 2520.240 1269.550 ;
        RECT 2520.040 1173.670 2520.180 1269.230 ;
        RECT 2519.980 1173.350 2520.240 1173.670 ;
        RECT 2519.980 1172.670 2520.240 1172.990 ;
        RECT 2520.040 1077.110 2520.180 1172.670 ;
        RECT 2519.980 1076.790 2520.240 1077.110 ;
        RECT 2519.980 1076.110 2520.240 1076.430 ;
        RECT 2520.040 1028.490 2520.180 1076.110 ;
        RECT 2519.980 1028.170 2520.240 1028.490 ;
        RECT 2519.520 1011.510 2519.780 1011.830 ;
        RECT 2519.060 1011.170 2519.320 1011.490 ;
        RECT 2518.600 1010.830 2518.860 1011.150 ;
        RECT 2528.780 1010.810 2528.920 2587.410 ;
        RECT 2528.720 1010.490 2528.980 1010.810 ;
        RECT 2287.220 1009.470 2287.480 1009.790 ;
        RECT 2094.020 1008.790 2094.280 1009.110 ;
        RECT 2055.440 1000.000 2055.740 1000.010 ;
        RECT 2059.880 1000.000 2061.560 1000.010 ;
        RECT 2064.480 1000.000 2065.700 1000.010 ;
        RECT 2068.620 1000.000 2069.840 1000.010 ;
        RECT 2073.220 1000.000 2074.900 1000.010 ;
        RECT 2077.360 1000.000 2079.040 1000.010 ;
        RECT 2081.960 1000.000 2083.180 1000.010 ;
        RECT 2086.100 1000.000 2087.780 1000.010 ;
        RECT 1603.260 999.870 1603.710 1000.000 ;
      LAYER met2 ;
        RECT 1599.850 995.720 1600.850 998.810 ;
      LAYER met2 ;
        RECT 1601.130 996.000 1601.410 999.870 ;
      LAYER met2 ;
        RECT 1601.690 995.720 1603.150 998.810 ;
      LAYER met2 ;
        RECT 1603.430 996.000 1603.710 999.870 ;
      LAYER met2 ;
        RECT 1603.990 995.720 1605.450 998.810 ;
      LAYER met2 ;
        RECT 1605.730 996.000 1606.010 1000.000 ;
      LAYER met2 ;
        RECT 1606.290 995.720 1607.290 998.810 ;
      LAYER met2 ;
        RECT 1607.570 996.000 1607.850 1000.000 ;
        RECT 1608.780 999.870 1610.150 1000.000 ;
      LAYER met2 ;
        RECT 1608.130 995.720 1609.590 998.810 ;
      LAYER met2 ;
        RECT 1609.870 996.000 1610.150 999.870 ;
        RECT 1612.170 999.870 1613.520 1000.000 ;
      LAYER met2 ;
        RECT 1610.430 995.720 1611.890 998.810 ;
      LAYER met2 ;
        RECT 1612.170 996.000 1612.450 999.870 ;
      LAYER met2 ;
        RECT 1612.730 995.720 1614.190 998.810 ;
      LAYER met2 ;
        RECT 1614.470 996.000 1614.750 1000.000 ;
      LAYER met2 ;
        RECT 1615.030 995.720 1616.030 998.810 ;
      LAYER met2 ;
        RECT 1616.310 996.000 1616.590 1000.000 ;
        RECT 1618.610 999.870 1620.420 1000.000 ;
        RECT 1620.910 999.870 1621.340 1000.000 ;
      LAYER met2 ;
        RECT 1616.870 995.720 1618.330 998.810 ;
      LAYER met2 ;
        RECT 1618.610 996.000 1618.890 999.870 ;
      LAYER met2 ;
        RECT 1619.170 995.720 1620.630 998.810 ;
      LAYER met2 ;
        RECT 1620.910 996.000 1621.190 999.870 ;
      LAYER met2 ;
        RECT 1621.470 995.720 1622.930 998.810 ;
      LAYER met2 ;
        RECT 1623.210 996.000 1623.490 1000.000 ;
      LAYER met2 ;
        RECT 1623.770 995.720 1624.770 998.810 ;
      LAYER met2 ;
        RECT 1625.050 996.000 1625.330 1000.000 ;
        RECT 1625.800 999.870 1627.630 1000.000 ;
        RECT 1628.560 999.870 1629.930 1000.000 ;
      LAYER met2 ;
        RECT 1625.610 995.720 1627.070 998.810 ;
      LAYER met2 ;
        RECT 1627.350 996.000 1627.630 999.870 ;
      LAYER met2 ;
        RECT 1627.910 995.720 1629.370 998.810 ;
      LAYER met2 ;
        RECT 1629.650 996.000 1629.930 999.870 ;
      LAYER met2 ;
        RECT 1630.210 995.720 1631.210 998.810 ;
      LAYER met2 ;
        RECT 1631.490 996.000 1631.770 1000.000 ;
      LAYER met2 ;
        RECT 1632.050 995.720 1633.510 998.810 ;
      LAYER met2 ;
        RECT 1633.790 996.000 1634.070 1000.000 ;
      LAYER met2 ;
        RECT 1634.350 995.720 1635.810 998.810 ;
      LAYER met2 ;
        RECT 1636.090 996.000 1636.370 1000.000 ;
      LAYER met2 ;
        RECT 1636.650 995.720 1638.110 998.810 ;
      LAYER met2 ;
        RECT 1638.390 996.000 1638.670 1000.000 ;
      LAYER met2 ;
        RECT 1638.950 995.720 1639.950 998.810 ;
      LAYER met2 ;
        RECT 1640.230 996.000 1640.510 1000.000 ;
      LAYER met2 ;
        RECT 1640.790 995.720 1642.250 998.810 ;
      LAYER met2 ;
        RECT 1642.530 996.000 1642.810 1000.000 ;
      LAYER met2 ;
        RECT 1643.090 995.720 1644.550 998.810 ;
      LAYER met2 ;
        RECT 1644.830 996.000 1645.110 1000.000 ;
      LAYER met2 ;
        RECT 1645.390 995.720 1646.850 998.810 ;
      LAYER met2 ;
        RECT 1647.130 996.000 1647.410 1000.000 ;
      LAYER met2 ;
        RECT 1647.690 995.720 1648.690 998.810 ;
      LAYER met2 ;
        RECT 1648.970 996.000 1649.250 1000.000 ;
      LAYER met2 ;
        RECT 1649.530 995.720 1650.990 998.810 ;
      LAYER met2 ;
        RECT 1651.270 996.000 1651.550 1000.000 ;
      LAYER met2 ;
        RECT 1651.830 995.720 1653.290 998.810 ;
      LAYER met2 ;
        RECT 1653.570 996.000 1653.850 1000.000 ;
      LAYER met2 ;
        RECT 1654.130 995.720 1655.130 998.810 ;
      LAYER met2 ;
        RECT 1655.410 996.000 1655.690 1000.000 ;
      LAYER met2 ;
        RECT 1655.970 995.720 1657.430 998.810 ;
      LAYER met2 ;
        RECT 1657.710 996.000 1657.990 1000.000 ;
      LAYER met2 ;
        RECT 1658.270 995.720 1659.730 998.810 ;
      LAYER met2 ;
        RECT 1660.010 996.000 1660.290 1000.000 ;
        RECT 1662.310 999.870 1662.740 1000.000 ;
        RECT 1664.150 999.870 1665.960 1000.000 ;
        RECT 1666.450 999.870 1667.800 1000.000 ;
      LAYER met2 ;
        RECT 1660.570 995.720 1662.030 998.810 ;
      LAYER met2 ;
        RECT 1662.310 996.000 1662.590 999.870 ;
      LAYER met2 ;
        RECT 1662.870 995.720 1663.870 998.810 ;
      LAYER met2 ;
        RECT 1664.150 996.000 1664.430 999.870 ;
      LAYER met2 ;
        RECT 1664.710 995.720 1666.170 998.810 ;
      LAYER met2 ;
        RECT 1666.450 996.000 1666.730 999.870 ;
      LAYER met2 ;
        RECT 1667.010 995.720 1668.470 998.810 ;
      LAYER met2 ;
        RECT 1668.750 996.000 1669.030 1000.000 ;
      LAYER met2 ;
        RECT 1669.310 995.720 1670.770 998.810 ;
      LAYER met2 ;
        RECT 1671.050 996.000 1671.330 1000.000 ;
      LAYER met2 ;
        RECT 1671.610 995.720 1672.610 998.810 ;
      LAYER met2 ;
        RECT 1672.890 996.000 1673.170 1000.000 ;
      LAYER met2 ;
        RECT 1673.450 995.720 1674.910 998.810 ;
      LAYER met2 ;
        RECT 1675.190 996.000 1675.470 1000.000 ;
      LAYER met2 ;
        RECT 1675.750 995.720 1677.210 998.810 ;
      LAYER met2 ;
        RECT 1677.490 996.000 1677.770 1000.000 ;
      LAYER met2 ;
        RECT 1678.050 995.720 1679.050 998.810 ;
      LAYER met2 ;
        RECT 1679.330 996.000 1679.610 1000.000 ;
      LAYER met2 ;
        RECT 1679.890 995.720 1681.350 998.810 ;
      LAYER met2 ;
        RECT 1681.630 996.000 1681.910 1000.000 ;
      LAYER met2 ;
        RECT 1682.190 995.720 1683.650 998.810 ;
      LAYER met2 ;
        RECT 1683.930 996.000 1684.210 1000.000 ;
      LAYER met2 ;
        RECT 1684.490 995.720 1685.950 998.810 ;
      LAYER met2 ;
        RECT 1686.230 996.000 1686.510 1000.000 ;
      LAYER met2 ;
        RECT 1686.790 995.720 1687.790 998.810 ;
      LAYER met2 ;
        RECT 1688.070 996.000 1688.350 1000.000 ;
      LAYER met2 ;
        RECT 1688.630 995.720 1690.090 998.810 ;
      LAYER met2 ;
        RECT 1690.370 996.000 1690.650 1000.000 ;
      LAYER met2 ;
        RECT 1690.930 995.720 1692.390 998.810 ;
      LAYER met2 ;
        RECT 1692.670 996.000 1692.950 1000.000 ;
      LAYER met2 ;
        RECT 1693.230 995.720 1694.230 998.810 ;
      LAYER met2 ;
        RECT 1694.510 996.000 1694.790 1000.000 ;
      LAYER met2 ;
        RECT 1695.070 995.720 1696.530 998.810 ;
      LAYER met2 ;
        RECT 1696.810 996.000 1697.090 1000.000 ;
      LAYER met2 ;
        RECT 1697.370 995.720 1698.830 998.810 ;
      LAYER met2 ;
        RECT 1699.110 996.000 1699.390 1000.000 ;
      LAYER met2 ;
        RECT 1699.670 995.720 1701.130 998.810 ;
      LAYER met2 ;
        RECT 1701.410 996.000 1701.690 1000.000 ;
      LAYER met2 ;
        RECT 1701.970 995.720 1702.970 998.810 ;
      LAYER met2 ;
        RECT 1703.250 996.000 1703.530 1000.000 ;
        RECT 1705.550 999.870 1707.360 1000.000 ;
      LAYER met2 ;
        RECT 1703.810 995.720 1705.270 998.810 ;
      LAYER met2 ;
        RECT 1705.550 996.000 1705.830 999.870 ;
      LAYER met2 ;
        RECT 1706.110 995.720 1707.570 998.810 ;
      LAYER met2 ;
        RECT 1707.850 996.000 1708.130 1000.000 ;
        RECT 1710.150 999.870 1710.580 1000.000 ;
      LAYER met2 ;
        RECT 1708.410 995.720 1709.870 998.810 ;
      LAYER met2 ;
        RECT 1710.150 996.000 1710.430 999.870 ;
      LAYER met2 ;
        RECT 1710.710 995.720 1711.710 998.810 ;
      LAYER met2 ;
        RECT 1711.990 996.000 1712.270 1000.000 ;
        RECT 1714.290 999.870 1716.100 1000.000 ;
      LAYER met2 ;
        RECT 1712.550 995.720 1714.010 998.810 ;
      LAYER met2 ;
        RECT 1714.290 996.000 1714.570 999.870 ;
      LAYER met2 ;
        RECT 1714.850 995.720 1716.310 998.810 ;
      LAYER met2 ;
        RECT 1716.590 996.000 1716.870 1000.000 ;
        RECT 1718.430 999.870 1720.240 1000.000 ;
      LAYER met2 ;
        RECT 1717.150 995.720 1718.150 998.810 ;
      LAYER met2 ;
        RECT 1718.430 996.000 1718.710 999.870 ;
      LAYER met2 ;
        RECT 1718.990 995.720 1720.450 998.810 ;
      LAYER met2 ;
        RECT 1720.730 996.000 1721.010 1000.000 ;
        RECT 1723.030 999.870 1724.840 1000.000 ;
      LAYER met2 ;
        RECT 1721.290 995.720 1722.750 998.810 ;
      LAYER met2 ;
        RECT 1723.030 996.000 1723.310 999.870 ;
      LAYER met2 ;
        RECT 1723.590 995.720 1725.050 998.810 ;
      LAYER met2 ;
        RECT 1725.330 996.000 1725.610 1000.000 ;
        RECT 1727.170 999.870 1728.980 1000.000 ;
      LAYER met2 ;
        RECT 1725.890 995.720 1726.890 998.810 ;
      LAYER met2 ;
        RECT 1727.170 996.000 1727.450 999.870 ;
      LAYER met2 ;
        RECT 1727.730 995.720 1729.190 998.810 ;
      LAYER met2 ;
        RECT 1729.470 996.000 1729.750 1000.000 ;
        RECT 1731.770 999.870 1733.580 1000.000 ;
      LAYER met2 ;
        RECT 1730.030 995.720 1731.490 998.810 ;
      LAYER met2 ;
        RECT 1731.770 996.000 1732.050 999.870 ;
      LAYER met2 ;
        RECT 1732.330 995.720 1733.790 998.810 ;
      LAYER met2 ;
        RECT 1734.070 996.000 1734.350 1000.000 ;
        RECT 1735.910 999.870 1737.720 1000.000 ;
      LAYER met2 ;
        RECT 1734.630 995.720 1735.630 998.810 ;
      LAYER met2 ;
        RECT 1735.910 996.000 1736.190 999.870 ;
      LAYER met2 ;
        RECT 1736.470 995.720 1737.930 998.810 ;
      LAYER met2 ;
        RECT 1738.210 996.000 1738.490 1000.000 ;
        RECT 1740.510 999.870 1741.860 1000.000 ;
      LAYER met2 ;
        RECT 1738.770 995.720 1740.230 998.810 ;
      LAYER met2 ;
        RECT 1740.510 996.000 1740.790 999.870 ;
      LAYER met2 ;
        RECT 1741.070 995.720 1742.070 998.810 ;
      LAYER met2 ;
        RECT 1742.350 996.000 1742.630 1000.000 ;
        RECT 1744.650 999.870 1745.540 1000.000 ;
      LAYER met2 ;
        RECT 1742.910 995.720 1744.370 998.810 ;
      LAYER met2 ;
        RECT 1744.650 996.000 1744.930 999.870 ;
      LAYER met2 ;
        RECT 1745.210 995.720 1746.670 998.810 ;
      LAYER met2 ;
        RECT 1746.950 996.000 1747.230 1000.000 ;
        RECT 1749.250 999.870 1750.140 1000.000 ;
      LAYER met2 ;
        RECT 1747.510 995.720 1748.970 998.810 ;
      LAYER met2 ;
        RECT 1749.250 996.000 1749.530 999.870 ;
      LAYER met2 ;
        RECT 1749.810 995.720 1750.810 998.810 ;
      LAYER met2 ;
        RECT 1751.090 996.000 1751.370 1000.000 ;
        RECT 1753.390 999.870 1755.200 1000.000 ;
      LAYER met2 ;
        RECT 1751.650 995.720 1753.110 998.810 ;
      LAYER met2 ;
        RECT 1753.390 996.000 1753.670 999.870 ;
      LAYER met2 ;
        RECT 1753.950 995.720 1755.410 998.810 ;
      LAYER met2 ;
        RECT 1755.690 996.000 1755.970 1000.000 ;
        RECT 1757.990 999.870 1758.880 1000.000 ;
      LAYER met2 ;
        RECT 1756.250 995.720 1757.710 998.810 ;
      LAYER met2 ;
        RECT 1757.990 996.000 1758.270 999.870 ;
      LAYER met2 ;
        RECT 1758.550 995.720 1759.550 998.810 ;
      LAYER met2 ;
        RECT 1759.830 996.000 1760.110 1000.000 ;
        RECT 1762.130 999.870 1763.940 1000.000 ;
      LAYER met2 ;
        RECT 1760.390 995.720 1761.850 998.810 ;
      LAYER met2 ;
        RECT 1762.130 996.000 1762.410 999.870 ;
      LAYER met2 ;
        RECT 1762.690 995.720 1764.150 998.810 ;
      LAYER met2 ;
        RECT 1764.430 996.000 1764.710 1000.000 ;
        RECT 1766.270 999.870 1768.080 1000.000 ;
      LAYER met2 ;
        RECT 1764.990 995.720 1765.990 998.810 ;
      LAYER met2 ;
        RECT 1766.270 996.000 1766.550 999.870 ;
      LAYER met2 ;
        RECT 1766.830 995.720 1768.290 998.810 ;
      LAYER met2 ;
        RECT 1768.570 996.000 1768.850 1000.000 ;
        RECT 1770.870 999.870 1772.680 1000.000 ;
      LAYER met2 ;
        RECT 1769.130 995.720 1770.590 998.810 ;
      LAYER met2 ;
        RECT 1770.870 996.000 1771.150 999.870 ;
      LAYER met2 ;
        RECT 1771.430 995.720 1772.890 998.810 ;
      LAYER met2 ;
        RECT 1773.170 996.000 1773.450 1000.000 ;
        RECT 1775.010 999.870 1776.820 1000.000 ;
      LAYER met2 ;
        RECT 1773.730 995.720 1774.730 998.810 ;
      LAYER met2 ;
        RECT 1775.010 996.000 1775.290 999.870 ;
      LAYER met2 ;
        RECT 1775.570 995.720 1777.030 998.810 ;
      LAYER met2 ;
        RECT 1777.310 996.000 1777.590 1000.000 ;
        RECT 1779.440 999.870 1779.890 1000.000 ;
      LAYER met2 ;
        RECT 1777.870 995.720 1779.330 998.810 ;
      LAYER met2 ;
        RECT 1779.610 996.000 1779.890 999.870 ;
      LAYER met2 ;
        RECT 1780.170 995.720 1781.630 998.810 ;
      LAYER met2 ;
        RECT 1781.910 996.000 1782.190 1000.000 ;
        RECT 1783.750 999.870 1785.560 1000.000 ;
      LAYER met2 ;
        RECT 1782.470 995.720 1783.470 998.810 ;
      LAYER met2 ;
        RECT 1783.750 996.000 1784.030 999.870 ;
      LAYER met2 ;
        RECT 1784.310 995.720 1785.770 998.810 ;
      LAYER met2 ;
        RECT 1786.050 996.000 1786.330 1000.000 ;
        RECT 1788.350 999.870 1789.700 1000.000 ;
      LAYER met2 ;
        RECT 1786.610 995.720 1788.070 998.810 ;
      LAYER met2 ;
        RECT 1788.350 996.000 1788.630 999.870 ;
      LAYER met2 ;
        RECT 1788.910 995.720 1789.910 998.810 ;
      LAYER met2 ;
        RECT 1790.190 996.000 1790.470 1000.000 ;
        RECT 1792.490 999.870 1793.840 1000.000 ;
      LAYER met2 ;
        RECT 1790.750 995.720 1792.210 998.810 ;
      LAYER met2 ;
        RECT 1792.490 996.000 1792.770 999.870 ;
      LAYER met2 ;
        RECT 1793.050 995.720 1794.510 998.810 ;
      LAYER met2 ;
        RECT 1794.790 996.000 1795.070 1000.000 ;
        RECT 1797.090 999.870 1798.440 1000.000 ;
      LAYER met2 ;
        RECT 1795.350 995.720 1796.810 998.810 ;
      LAYER met2 ;
        RECT 1797.090 996.000 1797.370 999.870 ;
      LAYER met2 ;
        RECT 1797.650 995.720 1798.650 998.810 ;
      LAYER met2 ;
        RECT 1798.930 996.000 1799.210 1000.000 ;
        RECT 1801.230 999.870 1803.040 1000.000 ;
      LAYER met2 ;
        RECT 1799.490 995.720 1800.950 998.810 ;
      LAYER met2 ;
        RECT 1801.230 996.000 1801.510 999.870 ;
      LAYER met2 ;
        RECT 1801.790 995.720 1803.250 998.810 ;
      LAYER met2 ;
        RECT 1803.530 996.000 1803.810 1000.000 ;
        RECT 1805.830 999.870 1807.180 1000.000 ;
      LAYER met2 ;
        RECT 1804.090 995.720 1805.550 998.810 ;
      LAYER met2 ;
        RECT 1805.830 996.000 1806.110 999.870 ;
      LAYER met2 ;
        RECT 1806.390 995.720 1807.390 998.810 ;
      LAYER met2 ;
        RECT 1807.670 996.000 1807.950 1000.000 ;
        RECT 1809.970 999.870 1811.780 1000.000 ;
      LAYER met2 ;
        RECT 1808.230 995.720 1809.690 998.810 ;
      LAYER met2 ;
        RECT 1809.970 996.000 1810.250 999.870 ;
      LAYER met2 ;
        RECT 1810.530 995.720 1811.990 998.810 ;
      LAYER met2 ;
        RECT 1812.270 996.000 1812.550 1000.000 ;
        RECT 1814.110 999.870 1814.540 1000.000 ;
      LAYER met2 ;
        RECT 1812.830 995.720 1813.830 998.810 ;
      LAYER met2 ;
        RECT 1814.110 996.000 1814.390 999.870 ;
      LAYER met2 ;
        RECT 1814.670 995.720 1816.130 998.810 ;
      LAYER met2 ;
        RECT 1816.410 996.000 1816.690 1000.000 ;
        RECT 1818.710 999.870 1820.520 1000.000 ;
      LAYER met2 ;
        RECT 1816.970 995.720 1818.430 998.810 ;
      LAYER met2 ;
        RECT 1818.710 996.000 1818.990 999.870 ;
      LAYER met2 ;
        RECT 1819.270 995.720 1820.730 998.810 ;
      LAYER met2 ;
        RECT 1821.010 996.000 1821.290 1000.000 ;
        RECT 1822.850 999.870 1824.660 1000.000 ;
        RECT 1825.150 999.870 1826.960 1000.000 ;
      LAYER met2 ;
        RECT 1821.570 995.720 1822.570 998.810 ;
      LAYER met2 ;
        RECT 1822.850 996.000 1823.130 999.870 ;
      LAYER met2 ;
        RECT 1823.410 995.720 1824.870 998.810 ;
      LAYER met2 ;
        RECT 1825.150 996.000 1825.430 999.870 ;
      LAYER met2 ;
        RECT 1825.710 995.720 1827.170 998.810 ;
      LAYER met2 ;
        RECT 1827.450 996.000 1827.730 1000.000 ;
        RECT 1829.750 999.870 1831.100 1000.000 ;
      LAYER met2 ;
        RECT 1828.010 995.720 1829.470 998.810 ;
      LAYER met2 ;
        RECT 1829.750 996.000 1830.030 999.870 ;
      LAYER met2 ;
        RECT 1830.310 995.720 1831.310 998.810 ;
      LAYER met2 ;
        RECT 1831.590 996.000 1831.870 1000.000 ;
        RECT 1833.890 999.870 1834.780 1000.000 ;
      LAYER met2 ;
        RECT 1832.150 995.720 1833.610 998.810 ;
      LAYER met2 ;
        RECT 1833.890 996.000 1834.170 999.870 ;
      LAYER met2 ;
        RECT 1834.450 995.720 1835.910 998.810 ;
      LAYER met2 ;
        RECT 1836.190 996.000 1836.470 1000.000 ;
      LAYER met2 ;
        RECT 1836.750 995.720 1837.750 998.810 ;
      LAYER met2 ;
        RECT 1838.030 996.000 1838.310 1000.000 ;
      LAYER met2 ;
        RECT 1838.590 995.720 1840.050 998.810 ;
      LAYER met2 ;
        RECT 1840.330 996.000 1840.610 1000.000 ;
      LAYER met2 ;
        RECT 1840.890 995.720 1842.350 998.810 ;
      LAYER met2 ;
        RECT 1842.630 996.000 1842.910 1000.000 ;
      LAYER met2 ;
        RECT 1843.190 995.720 1844.650 998.810 ;
      LAYER met2 ;
        RECT 1844.930 996.000 1845.210 1000.000 ;
      LAYER met2 ;
        RECT 1845.490 995.720 1846.490 998.810 ;
      LAYER met2 ;
        RECT 1846.770 996.000 1847.050 1000.000 ;
      LAYER met2 ;
        RECT 1847.330 995.720 1848.790 998.810 ;
      LAYER met2 ;
        RECT 1849.070 996.000 1849.350 1000.000 ;
      LAYER met2 ;
        RECT 1849.630 995.720 1851.090 998.810 ;
      LAYER met2 ;
        RECT 1851.370 996.000 1851.650 1000.000 ;
      LAYER met2 ;
        RECT 1851.930 995.720 1852.930 998.810 ;
      LAYER met2 ;
        RECT 1853.210 996.000 1853.490 1000.000 ;
      LAYER met2 ;
        RECT 1853.770 995.720 1855.230 998.810 ;
      LAYER met2 ;
        RECT 1855.510 996.000 1855.790 1000.000 ;
      LAYER met2 ;
        RECT 1856.070 995.720 1857.530 998.810 ;
      LAYER met2 ;
        RECT 1857.810 996.000 1858.090 1000.000 ;
      LAYER met2 ;
        RECT 1858.370 995.720 1859.830 998.810 ;
      LAYER met2 ;
        RECT 1860.110 996.000 1860.390 1000.000 ;
      LAYER met2 ;
        RECT 1860.670 995.720 1861.670 998.810 ;
      LAYER met2 ;
        RECT 1861.950 996.000 1862.230 1000.000 ;
      LAYER met2 ;
        RECT 1862.510 995.720 1863.970 998.810 ;
      LAYER met2 ;
        RECT 1864.250 996.000 1864.530 1000.000 ;
      LAYER met2 ;
        RECT 1864.810 995.720 1866.270 998.810 ;
      LAYER met2 ;
        RECT 1866.550 996.000 1866.830 1000.000 ;
      LAYER met2 ;
        RECT 1867.110 995.720 1868.570 998.810 ;
      LAYER met2 ;
        RECT 1868.850 996.000 1869.130 1000.000 ;
        RECT 1870.690 999.870 1872.500 1000.000 ;
      LAYER met2 ;
        RECT 1869.410 995.720 1870.410 998.810 ;
      LAYER met2 ;
        RECT 1870.690 996.000 1870.970 999.870 ;
      LAYER met2 ;
        RECT 1871.250 995.720 1872.710 998.810 ;
      LAYER met2 ;
        RECT 1872.990 996.000 1873.270 1000.000 ;
      LAYER met2 ;
        RECT 1873.550 995.720 1875.010 998.810 ;
      LAYER met2 ;
        RECT 1875.290 996.000 1875.570 1000.000 ;
        RECT 1877.130 999.870 1878.940 1000.000 ;
      LAYER met2 ;
        RECT 1875.850 995.720 1876.850 998.810 ;
      LAYER met2 ;
        RECT 1877.130 996.000 1877.410 999.870 ;
      LAYER met2 ;
        RECT 1877.690 995.720 1879.150 998.810 ;
      LAYER met2 ;
        RECT 1879.430 996.000 1879.710 1000.000 ;
        RECT 1881.730 999.870 1882.620 1000.000 ;
      LAYER met2 ;
        RECT 1879.990 995.720 1881.450 998.810 ;
      LAYER met2 ;
        RECT 1881.730 996.000 1882.010 999.870 ;
      LAYER met2 ;
        RECT 1882.290 995.720 1883.750 998.810 ;
      LAYER met2 ;
        RECT 1884.030 996.000 1884.310 1000.000 ;
      LAYER met2 ;
        RECT 1884.590 995.720 1885.590 998.810 ;
      LAYER met2 ;
        RECT 1885.870 996.000 1886.150 1000.000 ;
      LAYER met2 ;
        RECT 1886.430 995.720 1887.890 998.810 ;
      LAYER met2 ;
        RECT 1888.170 996.000 1888.450 1000.000 ;
      LAYER met2 ;
        RECT 1888.730 995.720 1890.190 998.810 ;
      LAYER met2 ;
        RECT 1890.470 996.000 1890.750 1000.000 ;
      LAYER met2 ;
        RECT 1891.030 995.720 1892.490 998.810 ;
      LAYER met2 ;
        RECT 1892.770 996.000 1893.050 1000.000 ;
      LAYER met2 ;
        RECT 1893.330 995.720 1894.330 998.810 ;
      LAYER met2 ;
        RECT 1894.610 996.000 1894.890 1000.000 ;
      LAYER met2 ;
        RECT 1895.170 995.720 1896.630 998.810 ;
      LAYER met2 ;
        RECT 1896.910 996.000 1897.190 1000.000 ;
      LAYER met2 ;
        RECT 1897.470 995.720 1898.930 998.810 ;
      LAYER met2 ;
        RECT 1899.210 996.000 1899.490 1000.000 ;
      LAYER met2 ;
        RECT 1899.770 995.720 1900.770 998.810 ;
      LAYER met2 ;
        RECT 1901.050 996.000 1901.330 1000.000 ;
      LAYER met2 ;
        RECT 1901.610 995.720 1903.070 998.810 ;
      LAYER met2 ;
        RECT 1903.350 996.000 1903.630 1000.000 ;
      LAYER met2 ;
        RECT 1903.910 995.720 1905.370 998.810 ;
      LAYER met2 ;
        RECT 1905.650 996.000 1905.930 1000.000 ;
      LAYER met2 ;
        RECT 1906.210 995.720 1907.670 998.810 ;
      LAYER met2 ;
        RECT 1907.950 996.000 1908.230 1000.000 ;
      LAYER met2 ;
        RECT 1908.510 995.720 1909.510 998.810 ;
      LAYER met2 ;
        RECT 1909.790 996.000 1910.070 1000.000 ;
      LAYER met2 ;
        RECT 1910.350 995.720 1911.810 998.810 ;
      LAYER met2 ;
        RECT 1912.090 996.000 1912.370 1000.000 ;
      LAYER met2 ;
        RECT 1912.650 995.720 1914.110 998.810 ;
      LAYER met2 ;
        RECT 1914.390 996.000 1914.670 1000.000 ;
      LAYER met2 ;
        RECT 1914.950 995.720 1916.410 998.810 ;
      LAYER met2 ;
        RECT 1916.690 996.000 1916.970 1000.000 ;
      LAYER met2 ;
        RECT 1917.250 995.720 1918.250 998.810 ;
      LAYER met2 ;
        RECT 1918.530 996.000 1918.810 1000.000 ;
      LAYER met2 ;
        RECT 1919.090 995.720 1920.550 998.810 ;
      LAYER met2 ;
        RECT 1920.830 996.000 1921.110 1000.000 ;
      LAYER met2 ;
        RECT 1921.390 995.720 1922.850 998.810 ;
      LAYER met2 ;
        RECT 1923.130 996.000 1923.410 1000.000 ;
      LAYER met2 ;
        RECT 1923.690 995.720 1924.690 998.810 ;
      LAYER met2 ;
        RECT 1924.970 996.000 1925.250 1000.000 ;
      LAYER met2 ;
        RECT 1925.530 995.720 1926.990 998.810 ;
      LAYER met2 ;
        RECT 1927.270 996.000 1927.550 1000.000 ;
      LAYER met2 ;
        RECT 1927.830 995.720 1929.290 998.810 ;
      LAYER met2 ;
        RECT 1929.570 996.000 1929.850 1000.000 ;
      LAYER met2 ;
        RECT 1930.130 995.720 1931.590 998.810 ;
      LAYER met2 ;
        RECT 1931.870 996.000 1932.150 1000.000 ;
      LAYER met2 ;
        RECT 1932.430 995.720 1933.430 998.810 ;
      LAYER met2 ;
        RECT 1933.710 996.000 1933.990 1000.000 ;
      LAYER met2 ;
        RECT 1934.270 995.720 1935.730 998.810 ;
      LAYER met2 ;
        RECT 1936.010 996.000 1936.290 1000.000 ;
      LAYER met2 ;
        RECT 1936.570 995.720 1938.030 998.810 ;
      LAYER met2 ;
        RECT 1938.310 996.000 1938.590 1000.000 ;
      LAYER met2 ;
        RECT 1938.870 995.720 1940.330 998.810 ;
      LAYER met2 ;
        RECT 1940.610 996.000 1940.890 1000.000 ;
      LAYER met2 ;
        RECT 1941.170 995.720 1942.170 998.810 ;
      LAYER met2 ;
        RECT 1942.450 996.000 1942.730 1000.000 ;
      LAYER met2 ;
        RECT 1943.010 995.720 1944.470 998.810 ;
      LAYER met2 ;
        RECT 1944.750 996.000 1945.030 1000.000 ;
      LAYER met2 ;
        RECT 1945.310 995.720 1946.770 998.810 ;
      LAYER met2 ;
        RECT 1947.050 996.000 1947.330 1000.000 ;
      LAYER met2 ;
        RECT 1947.610 995.720 1948.610 998.810 ;
      LAYER met2 ;
        RECT 1948.890 996.000 1949.170 1000.000 ;
      LAYER met2 ;
        RECT 1949.450 995.720 1950.910 998.810 ;
      LAYER met2 ;
        RECT 1951.190 996.000 1951.470 1000.000 ;
      LAYER met2 ;
        RECT 1951.750 995.720 1953.210 998.810 ;
      LAYER met2 ;
        RECT 1953.490 996.000 1953.770 1000.000 ;
      LAYER met2 ;
        RECT 1954.050 995.720 1955.510 998.810 ;
      LAYER met2 ;
        RECT 1955.790 996.000 1956.070 1000.000 ;
      LAYER met2 ;
        RECT 1956.350 995.720 1957.350 998.810 ;
      LAYER met2 ;
        RECT 1957.630 996.000 1957.910 1000.000 ;
      LAYER met2 ;
        RECT 1958.190 995.720 1959.650 998.810 ;
      LAYER met2 ;
        RECT 1959.930 996.000 1960.210 1000.000 ;
      LAYER met2 ;
        RECT 1960.490 995.720 1961.950 998.810 ;
      LAYER met2 ;
        RECT 1962.230 996.000 1962.510 1000.000 ;
      LAYER met2 ;
        RECT 1962.790 995.720 1964.250 998.810 ;
      LAYER met2 ;
        RECT 1964.530 996.000 1964.810 1000.000 ;
      LAYER met2 ;
        RECT 1965.090 995.720 1966.090 998.810 ;
      LAYER met2 ;
        RECT 1966.370 996.000 1966.650 1000.000 ;
      LAYER met2 ;
        RECT 1966.930 995.720 1968.390 998.810 ;
      LAYER met2 ;
        RECT 1968.670 996.000 1968.950 1000.000 ;
      LAYER met2 ;
        RECT 1969.230 995.720 1970.690 998.810 ;
      LAYER met2 ;
        RECT 1970.970 996.000 1971.250 1000.000 ;
      LAYER met2 ;
        RECT 1971.530 995.720 1972.530 998.810 ;
      LAYER met2 ;
        RECT 1972.810 996.000 1973.090 1000.000 ;
      LAYER met2 ;
        RECT 1973.370 995.720 1974.830 998.810 ;
      LAYER met2 ;
        RECT 1975.110 996.000 1975.390 1000.000 ;
      LAYER met2 ;
        RECT 1975.670 995.720 1977.130 998.810 ;
      LAYER met2 ;
        RECT 1977.410 996.000 1977.690 1000.000 ;
      LAYER met2 ;
        RECT 1977.970 995.720 1979.430 998.810 ;
      LAYER met2 ;
        RECT 1979.710 996.000 1979.990 1000.000 ;
      LAYER met2 ;
        RECT 1980.270 995.720 1981.270 998.810 ;
      LAYER met2 ;
        RECT 1981.550 996.000 1981.830 1000.000 ;
      LAYER met2 ;
        RECT 1982.110 995.720 1983.570 998.810 ;
      LAYER met2 ;
        RECT 1983.850 996.000 1984.130 1000.000 ;
      LAYER met2 ;
        RECT 1984.410 995.720 1985.870 998.810 ;
      LAYER met2 ;
        RECT 1986.150 996.000 1986.430 1000.000 ;
      LAYER met2 ;
        RECT 1986.710 995.720 1988.170 998.810 ;
      LAYER met2 ;
        RECT 1988.450 996.000 1988.730 1000.000 ;
      LAYER met2 ;
        RECT 1989.010 995.720 1990.010 998.810 ;
      LAYER met2 ;
        RECT 1990.290 996.000 1990.570 1000.000 ;
      LAYER met2 ;
        RECT 1990.850 995.720 1992.310 998.810 ;
      LAYER met2 ;
        RECT 1992.590 996.000 1992.870 1000.000 ;
      LAYER met2 ;
        RECT 1993.150 995.720 1994.610 998.810 ;
      LAYER met2 ;
        RECT 1994.890 996.000 1995.170 1000.000 ;
      LAYER met2 ;
        RECT 1995.450 995.720 1996.450 998.810 ;
      LAYER met2 ;
        RECT 1996.730 996.000 1997.010 1000.000 ;
      LAYER met2 ;
        RECT 1997.290 995.720 1998.750 998.810 ;
      LAYER met2 ;
        RECT 1999.030 996.000 1999.310 1000.000 ;
        RECT 2001.330 999.870 2003.140 1000.000 ;
        RECT 2003.630 999.870 2004.980 1000.000 ;
      LAYER met2 ;
        RECT 1999.590 995.720 2001.050 998.810 ;
      LAYER met2 ;
        RECT 2001.330 996.000 2001.610 999.870 ;
      LAYER met2 ;
        RECT 2001.890 995.720 2003.350 998.810 ;
      LAYER met2 ;
        RECT 2003.630 996.000 2003.910 999.870 ;
      LAYER met2 ;
        RECT 2004.190 995.720 2005.190 998.810 ;
      LAYER met2 ;
        RECT 2005.470 996.000 2005.750 1000.000 ;
      LAYER met2 ;
        RECT 2006.030 995.720 2007.490 998.810 ;
      LAYER met2 ;
        RECT 2007.770 996.000 2008.050 1000.000 ;
      LAYER met2 ;
        RECT 2008.330 995.720 2009.790 998.810 ;
      LAYER met2 ;
        RECT 2010.070 996.000 2010.350 1000.000 ;
      LAYER met2 ;
        RECT 2010.630 995.720 2011.630 998.810 ;
      LAYER met2 ;
        RECT 2011.910 996.000 2012.190 1000.000 ;
      LAYER met2 ;
        RECT 2012.470 995.720 2013.930 998.810 ;
      LAYER met2 ;
        RECT 2014.210 996.000 2014.490 1000.000 ;
      LAYER met2 ;
        RECT 2014.770 995.720 2016.230 998.810 ;
      LAYER met2 ;
        RECT 2016.510 996.000 2016.790 1000.000 ;
      LAYER met2 ;
        RECT 2017.070 995.720 2018.530 998.810 ;
      LAYER met2 ;
        RECT 2018.810 996.000 2019.090 1000.000 ;
      LAYER met2 ;
        RECT 2019.370 995.720 2020.370 998.810 ;
      LAYER met2 ;
        RECT 2020.650 996.000 2020.930 1000.000 ;
      LAYER met2 ;
        RECT 2021.210 995.720 2022.670 998.810 ;
      LAYER met2 ;
        RECT 2022.950 996.000 2023.230 1000.000 ;
      LAYER met2 ;
        RECT 2023.510 995.720 2024.970 998.810 ;
      LAYER met2 ;
        RECT 2025.250 996.000 2025.530 1000.000 ;
      LAYER met2 ;
        RECT 2025.810 995.720 2027.270 998.810 ;
      LAYER met2 ;
        RECT 2027.550 996.000 2027.830 1000.000 ;
      LAYER met2 ;
        RECT 2028.110 995.720 2029.110 998.810 ;
      LAYER met2 ;
        RECT 2029.390 996.000 2029.670 1000.000 ;
      LAYER met2 ;
        RECT 2029.950 995.720 2031.410 998.810 ;
      LAYER met2 ;
        RECT 2031.690 996.000 2031.970 1000.000 ;
      LAYER met2 ;
        RECT 2032.250 995.720 2033.710 998.810 ;
      LAYER met2 ;
        RECT 2033.990 996.000 2034.270 1000.000 ;
      LAYER met2 ;
        RECT 2034.550 995.720 2035.550 998.810 ;
      LAYER met2 ;
        RECT 2035.830 996.000 2036.110 1000.000 ;
      LAYER met2 ;
        RECT 2036.390 995.720 2037.850 998.810 ;
      LAYER met2 ;
        RECT 2038.130 996.000 2038.410 1000.000 ;
        RECT 2040.430 999.870 2042.240 1000.000 ;
      LAYER met2 ;
        RECT 2038.690 995.720 2040.150 998.810 ;
      LAYER met2 ;
        RECT 2040.430 996.000 2040.710 999.870 ;
      LAYER met2 ;
        RECT 2040.990 995.720 2042.450 998.810 ;
      LAYER met2 ;
        RECT 2042.730 996.000 2043.010 1000.000 ;
        RECT 2044.570 999.870 2046.380 1000.000 ;
      LAYER met2 ;
        RECT 2043.290 995.720 2044.290 998.810 ;
      LAYER met2 ;
        RECT 2044.570 996.000 2044.850 999.870 ;
      LAYER met2 ;
        RECT 2045.130 995.720 2046.590 998.810 ;
      LAYER met2 ;
        RECT 2046.870 996.000 2047.150 1000.000 ;
        RECT 2049.170 999.870 2050.980 1000.000 ;
      LAYER met2 ;
        RECT 2047.430 995.720 2048.890 998.810 ;
      LAYER met2 ;
        RECT 2049.170 996.000 2049.450 999.870 ;
      LAYER met2 ;
        RECT 2049.730 995.720 2051.190 998.810 ;
      LAYER met2 ;
        RECT 2051.470 996.000 2051.750 1000.000 ;
      LAYER met2 ;
        RECT 2052.030 995.720 2053.030 998.810 ;
      LAYER met2 ;
        RECT 2053.310 996.000 2053.590 1000.000 ;
        RECT 2055.440 999.870 2055.890 1000.000 ;
      LAYER met2 ;
        RECT 2053.870 995.720 2055.330 998.810 ;
      LAYER met2 ;
        RECT 2055.610 996.000 2055.890 999.870 ;
      LAYER met2 ;
        RECT 2056.170 995.720 2057.630 998.810 ;
      LAYER met2 ;
        RECT 2057.910 996.000 2058.190 1000.000 ;
        RECT 2059.750 999.870 2061.560 1000.000 ;
      LAYER met2 ;
        RECT 2058.470 995.720 2059.470 998.810 ;
      LAYER met2 ;
        RECT 2059.750 996.000 2060.030 999.870 ;
      LAYER met2 ;
        RECT 2060.310 995.720 2061.770 998.810 ;
      LAYER met2 ;
        RECT 2062.050 996.000 2062.330 1000.000 ;
        RECT 2064.350 999.870 2065.700 1000.000 ;
      LAYER met2 ;
        RECT 2062.610 995.720 2064.070 998.810 ;
      LAYER met2 ;
        RECT 2064.350 996.000 2064.630 999.870 ;
      LAYER met2 ;
        RECT 2064.910 995.720 2066.370 998.810 ;
      LAYER met2 ;
        RECT 2066.650 996.000 2066.930 1000.000 ;
        RECT 2068.490 999.870 2069.840 1000.000 ;
      LAYER met2 ;
        RECT 2067.210 995.720 2068.210 998.810 ;
      LAYER met2 ;
        RECT 2068.490 996.000 2068.770 999.870 ;
      LAYER met2 ;
        RECT 2069.050 995.720 2070.510 998.810 ;
      LAYER met2 ;
        RECT 2070.790 996.000 2071.070 1000.000 ;
        RECT 2073.090 999.870 2074.900 1000.000 ;
      LAYER met2 ;
        RECT 2071.350 995.720 2072.810 998.810 ;
      LAYER met2 ;
        RECT 2073.090 996.000 2073.370 999.870 ;
      LAYER met2 ;
        RECT 2073.650 995.720 2075.110 998.810 ;
      LAYER met2 ;
        RECT 2075.390 996.000 2075.670 1000.000 ;
        RECT 2077.230 999.870 2079.040 1000.000 ;
      LAYER met2 ;
        RECT 2075.950 995.720 2076.950 998.810 ;
      LAYER met2 ;
        RECT 2077.230 996.000 2077.510 999.870 ;
      LAYER met2 ;
        RECT 2077.790 995.720 2079.250 998.810 ;
      LAYER met2 ;
        RECT 2079.530 996.000 2079.810 1000.000 ;
        RECT 2081.830 999.870 2083.180 1000.000 ;
      LAYER met2 ;
        RECT 2080.090 995.720 2081.550 998.810 ;
      LAYER met2 ;
        RECT 2081.830 996.000 2082.110 999.870 ;
      LAYER met2 ;
        RECT 2082.390 995.720 2083.390 998.810 ;
      LAYER met2 ;
        RECT 2083.670 996.000 2083.950 1000.000 ;
        RECT 2085.970 999.870 2087.780 1000.000 ;
      LAYER met2 ;
        RECT 2084.230 995.720 2085.690 998.810 ;
      LAYER met2 ;
        RECT 2085.970 996.000 2086.250 999.870 ;
      LAYER met2 ;
        RECT 2086.530 995.720 2087.990 998.810 ;
      LAYER met2 ;
        RECT 2088.270 996.000 2088.550 1000.000 ;
      LAYER met2 ;
        RECT 2088.830 995.720 2090.290 998.810 ;
      LAYER met2 ;
        RECT 2090.570 996.000 2090.850 1000.000 ;
      LAYER met2 ;
        RECT 2091.130 995.720 2092.130 998.810 ;
      LAYER met2 ;
        RECT 2092.410 996.000 2092.690 1000.000 ;
      LAYER met2 ;
        RECT 2092.970 995.720 2094.430 998.810 ;
      LAYER met2 ;
        RECT 2094.710 996.000 2094.990 1000.000 ;
      LAYER met2 ;
        RECT 2095.270 995.720 2096.730 998.810 ;
      LAYER met2 ;
        RECT 2097.010 996.000 2097.290 1000.000 ;
      LAYER met2 ;
        RECT 2097.570 995.720 2099.030 998.810 ;
      LAYER met2 ;
        RECT 2099.310 996.000 2099.590 1000.000 ;
      LAYER met2 ;
        RECT 2099.870 995.720 2100.870 998.810 ;
      LAYER met2 ;
        RECT 2101.150 996.000 2101.430 1000.000 ;
      LAYER met2 ;
        RECT 2101.710 995.720 2103.170 998.810 ;
      LAYER met2 ;
        RECT 2103.450 996.000 2103.730 1000.000 ;
      LAYER met2 ;
        RECT 2104.010 995.720 2105.470 998.810 ;
      LAYER met2 ;
        RECT 2105.750 996.000 2106.030 1000.000 ;
      LAYER met2 ;
        RECT 2106.310 995.720 2107.310 998.810 ;
      LAYER met2 ;
        RECT 2107.590 996.000 2107.870 1000.000 ;
      LAYER met2 ;
        RECT 2108.150 995.720 2109.610 998.810 ;
      LAYER met2 ;
        RECT 2109.890 996.000 2110.170 1000.000 ;
      LAYER met2 ;
        RECT 2110.450 995.720 2111.910 998.810 ;
      LAYER met2 ;
        RECT 2112.190 996.000 2112.470 1000.000 ;
      LAYER met2 ;
        RECT 2112.750 995.720 2114.210 998.810 ;
      LAYER met2 ;
        RECT 2114.490 996.000 2114.770 1000.000 ;
      LAYER met2 ;
        RECT 2115.050 995.720 2116.050 998.810 ;
      LAYER met2 ;
        RECT 2116.330 996.000 2116.610 1000.000 ;
      LAYER met2 ;
        RECT 2116.890 995.720 2118.350 998.810 ;
      LAYER met2 ;
        RECT 2118.630 996.000 2118.910 1000.000 ;
      LAYER met2 ;
        RECT 2119.190 995.720 2120.650 998.810 ;
      LAYER met2 ;
        RECT 2120.930 996.000 2121.210 1000.000 ;
      LAYER met2 ;
        RECT 2121.490 995.720 2122.950 998.810 ;
      LAYER met2 ;
        RECT 2123.230 996.000 2123.510 1000.000 ;
      LAYER met2 ;
        RECT 2123.790 995.720 2124.790 998.810 ;
      LAYER met2 ;
        RECT 2125.070 996.000 2125.350 1000.000 ;
      LAYER met2 ;
        RECT 2125.630 995.720 2127.090 998.810 ;
      LAYER met2 ;
        RECT 2127.370 996.000 2127.650 1000.000 ;
      LAYER met2 ;
        RECT 2127.930 995.720 2129.390 998.810 ;
      LAYER met2 ;
        RECT 2129.670 996.000 2129.950 1000.000 ;
      LAYER met2 ;
        RECT 2130.230 995.720 2131.230 998.810 ;
      LAYER met2 ;
        RECT 2131.510 996.000 2131.790 1000.000 ;
      LAYER met2 ;
        RECT 2132.070 995.720 2133.530 998.810 ;
      LAYER met2 ;
        RECT 2133.810 996.000 2134.090 1000.000 ;
      LAYER met2 ;
        RECT 2134.370 995.720 2135.830 998.810 ;
      LAYER met2 ;
        RECT 2136.110 996.000 2136.390 1000.000 ;
      LAYER met2 ;
        RECT 2136.670 995.720 2138.130 998.810 ;
      LAYER met2 ;
        RECT 2138.410 996.000 2138.690 1000.000 ;
      LAYER met2 ;
        RECT 2138.970 995.720 2139.970 998.810 ;
      LAYER met2 ;
        RECT 2140.250 996.000 2140.530 1000.000 ;
      LAYER met2 ;
        RECT 2140.810 995.720 2142.270 998.810 ;
      LAYER met2 ;
        RECT 2142.550 996.000 2142.830 1000.000 ;
      LAYER met2 ;
        RECT 2143.110 995.720 2144.570 998.810 ;
      LAYER met2 ;
        RECT 2144.850 996.000 2145.130 1000.000 ;
      LAYER met2 ;
        RECT 2145.410 995.720 2146.870 998.810 ;
      LAYER met2 ;
        RECT 2147.150 996.000 2147.430 1000.000 ;
      LAYER met2 ;
        RECT 2147.710 995.720 2148.710 998.810 ;
      LAYER met2 ;
        RECT 2148.990 996.000 2149.270 1000.000 ;
      LAYER met2 ;
        RECT 2149.550 995.720 2151.010 998.810 ;
      LAYER met2 ;
        RECT 2151.290 996.000 2151.570 1000.000 ;
      LAYER met2 ;
        RECT 2151.850 995.720 2153.310 998.810 ;
      LAYER met2 ;
        RECT 2153.590 996.000 2153.870 1000.000 ;
      LAYER met2 ;
        RECT 2154.150 995.720 2155.150 998.810 ;
      LAYER met2 ;
        RECT 2155.430 996.000 2155.710 1000.000 ;
      LAYER met2 ;
        RECT 2155.990 995.720 2157.450 998.810 ;
      LAYER met2 ;
        RECT 2157.730 996.000 2158.010 1000.000 ;
      LAYER met2 ;
        RECT 2158.290 995.720 2159.750 998.810 ;
      LAYER met2 ;
        RECT 2160.030 996.000 2160.310 1000.000 ;
      LAYER met2 ;
        RECT 2160.590 995.720 2162.050 998.810 ;
      LAYER met2 ;
        RECT 2162.330 996.000 2162.610 1000.000 ;
      LAYER met2 ;
        RECT 2162.890 995.720 2163.890 998.810 ;
      LAYER met2 ;
        RECT 2164.170 996.000 2164.450 1000.000 ;
      LAYER met2 ;
        RECT 2164.730 995.720 2166.190 998.810 ;
      LAYER met2 ;
        RECT 2166.470 996.000 2166.750 1000.000 ;
      LAYER met2 ;
        RECT 2167.030 995.720 2168.490 998.810 ;
      LAYER met2 ;
        RECT 2168.770 996.000 2169.050 1000.000 ;
      LAYER met2 ;
        RECT 671.020 604.280 2169.040 995.720 ;
        RECT 671.020 602.195 671.190 604.280 ;
        RECT 672.030 602.195 673.950 604.280 ;
        RECT 674.790 602.195 677.170 604.280 ;
        RECT 678.010 602.195 679.930 604.280 ;
        RECT 680.770 602.195 683.150 604.280 ;
        RECT 683.990 602.195 686.370 604.280 ;
        RECT 687.210 602.195 689.130 604.280 ;
        RECT 689.970 602.195 692.350 604.280 ;
        RECT 693.190 602.195 695.570 604.280 ;
        RECT 696.410 602.195 698.330 604.280 ;
        RECT 699.170 602.195 701.550 604.280 ;
        RECT 702.390 602.195 704.770 604.280 ;
        RECT 705.610 602.195 707.530 604.280 ;
        RECT 708.370 602.195 710.750 604.280 ;
        RECT 711.590 602.195 713.970 604.280 ;
        RECT 714.810 602.195 716.730 604.280 ;
        RECT 717.570 602.195 719.950 604.280 ;
        RECT 720.790 602.195 723.170 604.280 ;
        RECT 724.010 602.195 725.930 604.280 ;
        RECT 726.770 602.195 729.150 604.280 ;
        RECT 729.990 602.195 732.370 604.280 ;
        RECT 733.210 602.195 735.130 604.280 ;
        RECT 735.970 602.195 738.350 604.280 ;
        RECT 739.190 602.195 741.570 604.280 ;
        RECT 742.410 602.195 744.330 604.280 ;
        RECT 745.170 602.195 747.550 604.280 ;
        RECT 748.390 602.195 750.770 604.280 ;
        RECT 751.610 602.195 753.530 604.280 ;
        RECT 754.370 602.195 756.750 604.280 ;
        RECT 757.590 602.195 759.510 604.280 ;
        RECT 760.350 602.195 762.730 604.280 ;
        RECT 763.570 602.195 765.950 604.280 ;
        RECT 766.790 602.195 768.710 604.280 ;
        RECT 769.550 602.195 771.930 604.280 ;
        RECT 772.770 602.195 775.150 604.280 ;
        RECT 775.990 602.195 777.910 604.280 ;
        RECT 778.750 602.195 781.130 604.280 ;
        RECT 781.970 602.195 784.350 604.280 ;
        RECT 785.190 602.195 787.110 604.280 ;
        RECT 787.950 602.195 790.330 604.280 ;
        RECT 791.170 602.195 793.550 604.280 ;
        RECT 794.390 602.195 796.310 604.280 ;
        RECT 797.150 602.195 799.530 604.280 ;
        RECT 800.370 602.195 802.750 604.280 ;
        RECT 803.590 602.195 805.510 604.280 ;
        RECT 806.350 602.195 808.730 604.280 ;
        RECT 809.570 602.195 811.950 604.280 ;
        RECT 812.790 602.195 814.710 604.280 ;
        RECT 815.550 602.195 817.930 604.280 ;
        RECT 818.770 602.195 821.150 604.280 ;
        RECT 821.990 602.195 823.910 604.280 ;
        RECT 824.750 602.195 827.130 604.280 ;
        RECT 827.970 602.195 830.350 604.280 ;
        RECT 831.190 602.195 833.110 604.280 ;
        RECT 833.950 602.195 836.330 604.280 ;
        RECT 837.170 602.195 839.550 604.280 ;
        RECT 840.390 602.195 842.310 604.280 ;
        RECT 843.150 602.195 845.530 604.280 ;
        RECT 846.370 602.195 848.290 604.280 ;
        RECT 849.130 602.195 851.510 604.280 ;
        RECT 852.350 602.195 854.730 604.280 ;
        RECT 855.570 602.195 857.490 604.280 ;
        RECT 858.330 602.195 860.710 604.280 ;
        RECT 861.550 602.195 863.930 604.280 ;
        RECT 864.770 602.195 866.690 604.280 ;
        RECT 867.530 602.195 869.910 604.280 ;
        RECT 870.750 602.195 873.130 604.280 ;
        RECT 873.970 602.195 875.890 604.280 ;
        RECT 876.730 602.195 879.110 604.280 ;
        RECT 879.950 602.195 882.330 604.280 ;
        RECT 883.170 602.195 885.090 604.280 ;
        RECT 885.930 602.195 888.310 604.280 ;
        RECT 889.150 602.195 891.530 604.280 ;
        RECT 892.370 602.195 894.290 604.280 ;
        RECT 895.130 602.195 897.510 604.280 ;
        RECT 898.350 602.195 900.730 604.280 ;
        RECT 901.570 602.195 903.490 604.280 ;
        RECT 904.330 602.195 906.710 604.280 ;
        RECT 907.550 602.195 909.930 604.280 ;
        RECT 910.770 602.195 912.690 604.280 ;
        RECT 913.530 602.195 915.910 604.280 ;
        RECT 916.750 602.195 919.130 604.280 ;
        RECT 919.970 602.195 921.890 604.280 ;
        RECT 922.730 602.195 925.110 604.280 ;
        RECT 925.950 602.195 928.330 604.280 ;
        RECT 929.170 602.195 931.090 604.280 ;
        RECT 931.930 602.195 934.310 604.280 ;
        RECT 935.150 602.195 937.070 604.280 ;
        RECT 937.910 602.195 940.290 604.280 ;
        RECT 941.130 602.195 943.510 604.280 ;
        RECT 944.350 602.195 946.270 604.280 ;
        RECT 947.110 602.195 949.490 604.280 ;
        RECT 950.330 602.195 952.710 604.280 ;
        RECT 953.550 602.195 955.470 604.280 ;
        RECT 956.310 602.195 958.690 604.280 ;
        RECT 959.530 602.195 961.910 604.280 ;
        RECT 962.750 602.195 964.670 604.280 ;
        RECT 965.510 602.195 967.890 604.280 ;
        RECT 968.730 602.195 971.110 604.280 ;
        RECT 971.950 602.195 973.870 604.280 ;
        RECT 974.710 602.195 977.090 604.280 ;
        RECT 977.930 602.195 980.310 604.280 ;
        RECT 981.150 602.195 983.070 604.280 ;
        RECT 983.910 602.195 986.290 604.280 ;
        RECT 987.130 602.195 989.510 604.280 ;
        RECT 990.350 602.195 992.270 604.280 ;
        RECT 993.110 602.195 995.490 604.280 ;
        RECT 996.330 602.195 998.710 604.280 ;
        RECT 999.550 602.195 1001.470 604.280 ;
        RECT 1002.310 602.195 1004.690 604.280 ;
        RECT 1005.530 602.195 1007.910 604.280 ;
        RECT 1008.750 602.195 1010.670 604.280 ;
        RECT 1011.510 602.195 1013.890 604.280 ;
        RECT 1014.730 602.195 1017.110 604.280 ;
        RECT 1017.950 602.195 1019.870 604.280 ;
        RECT 1020.710 602.195 1023.090 604.280 ;
        RECT 1023.930 602.195 1025.850 604.280 ;
        RECT 1026.690 602.195 1029.070 604.280 ;
        RECT 1029.910 602.195 1032.290 604.280 ;
        RECT 1033.130 602.195 1035.050 604.280 ;
        RECT 1035.890 602.195 1038.270 604.280 ;
        RECT 1039.110 602.195 1041.490 604.280 ;
        RECT 1042.330 602.195 1044.250 604.280 ;
        RECT 1045.090 602.195 1047.470 604.280 ;
        RECT 1048.310 602.195 1050.690 604.280 ;
        RECT 1051.530 602.195 1053.450 604.280 ;
        RECT 1054.290 602.195 1056.670 604.280 ;
        RECT 1057.510 602.195 1059.890 604.280 ;
        RECT 1060.730 602.195 1062.650 604.280 ;
        RECT 1063.490 602.195 1065.870 604.280 ;
        RECT 1066.710 602.195 1069.090 604.280 ;
        RECT 1069.930 602.195 1071.850 604.280 ;
        RECT 1072.690 602.195 1075.070 604.280 ;
        RECT 1075.910 602.195 1078.290 604.280 ;
        RECT 1079.130 602.195 1081.050 604.280 ;
        RECT 1081.890 602.195 1084.270 604.280 ;
        RECT 1085.110 602.195 1087.490 604.280 ;
        RECT 1088.330 602.195 1090.250 604.280 ;
        RECT 1091.090 602.195 1093.470 604.280 ;
        RECT 1094.310 602.195 1096.690 604.280 ;
        RECT 1097.530 602.195 1099.450 604.280 ;
        RECT 1100.290 602.195 1102.670 604.280 ;
        RECT 1103.510 602.195 1105.890 604.280 ;
        RECT 1106.730 602.195 1108.650 604.280 ;
        RECT 1109.490 602.195 1111.870 604.280 ;
        RECT 1112.710 602.195 1114.630 604.280 ;
        RECT 1115.470 602.195 1117.850 604.280 ;
        RECT 1118.690 602.195 1121.070 604.280 ;
        RECT 1121.910 602.195 1123.830 604.280 ;
        RECT 1124.670 602.195 1127.050 604.280 ;
        RECT 1127.890 602.195 1130.270 604.280 ;
        RECT 1131.110 602.195 1133.030 604.280 ;
        RECT 1133.870 602.195 1136.250 604.280 ;
        RECT 1137.090 602.195 1139.470 604.280 ;
        RECT 1140.310 602.195 1142.230 604.280 ;
        RECT 1143.070 602.195 1145.450 604.280 ;
        RECT 1146.290 602.195 1148.670 604.280 ;
        RECT 1149.510 602.195 1151.430 604.280 ;
        RECT 1152.270 602.195 1154.650 604.280 ;
        RECT 1155.490 602.195 1157.870 604.280 ;
        RECT 1158.710 602.195 1160.630 604.280 ;
        RECT 1161.470 602.195 1163.850 604.280 ;
        RECT 1164.690 602.195 1167.070 604.280 ;
        RECT 1167.910 602.195 1169.830 604.280 ;
        RECT 1170.670 602.195 1173.050 604.280 ;
        RECT 1173.890 602.195 1176.270 604.280 ;
        RECT 1177.110 602.195 1179.030 604.280 ;
        RECT 1179.870 602.195 1182.250 604.280 ;
        RECT 1183.090 602.195 1185.470 604.280 ;
        RECT 1186.310 602.195 1188.230 604.280 ;
        RECT 1189.070 602.195 1191.450 604.280 ;
        RECT 1192.290 602.195 1194.670 604.280 ;
        RECT 1195.510 602.195 1197.430 604.280 ;
        RECT 1198.270 602.195 1200.650 604.280 ;
        RECT 1201.490 602.195 1203.410 604.280 ;
        RECT 1204.250 602.195 1206.630 604.280 ;
        RECT 1207.470 602.195 1209.850 604.280 ;
        RECT 1210.690 602.195 1212.610 604.280 ;
        RECT 1213.450 602.195 1215.830 604.280 ;
        RECT 1216.670 602.195 1219.050 604.280 ;
        RECT 1219.890 602.195 1221.810 604.280 ;
        RECT 1222.650 602.195 1225.030 604.280 ;
        RECT 1225.870 602.195 1228.250 604.280 ;
        RECT 1229.090 602.195 1231.010 604.280 ;
        RECT 1231.850 602.195 1234.230 604.280 ;
        RECT 1235.070 602.195 1237.450 604.280 ;
        RECT 1238.290 602.195 1240.210 604.280 ;
        RECT 1241.050 602.195 1243.430 604.280 ;
        RECT 1244.270 602.195 1246.650 604.280 ;
        RECT 1247.490 602.195 1249.410 604.280 ;
        RECT 1250.250 602.195 1252.630 604.280 ;
        RECT 1253.470 602.195 1255.850 604.280 ;
        RECT 1256.690 602.195 1258.610 604.280 ;
        RECT 1259.450 602.195 1261.830 604.280 ;
        RECT 1262.670 602.195 1265.050 604.280 ;
        RECT 1265.890 602.195 1267.810 604.280 ;
        RECT 1268.650 602.195 1271.030 604.280 ;
        RECT 1271.870 602.195 1274.250 604.280 ;
        RECT 1275.090 602.195 1277.010 604.280 ;
        RECT 1277.850 602.195 1280.230 604.280 ;
        RECT 1281.070 602.195 1283.450 604.280 ;
        RECT 1284.290 602.195 1286.210 604.280 ;
        RECT 1287.050 602.195 1289.430 604.280 ;
        RECT 1290.270 602.195 1292.190 604.280 ;
        RECT 1293.030 602.195 1295.410 604.280 ;
        RECT 1296.250 602.195 1298.630 604.280 ;
        RECT 1299.470 602.195 1301.390 604.280 ;
        RECT 1302.230 602.195 1304.610 604.280 ;
        RECT 1305.450 602.195 1307.830 604.280 ;
        RECT 1308.670 602.195 1310.590 604.280 ;
        RECT 1311.430 602.195 1313.810 604.280 ;
        RECT 1314.650 602.195 1317.030 604.280 ;
        RECT 1317.870 602.195 1319.790 604.280 ;
        RECT 1320.630 602.195 1323.010 604.280 ;
        RECT 1323.850 602.195 1326.230 604.280 ;
        RECT 1327.070 602.195 1328.990 604.280 ;
        RECT 1329.830 602.195 1332.210 604.280 ;
        RECT 1333.050 602.195 1335.430 604.280 ;
        RECT 1336.270 602.195 1338.190 604.280 ;
        RECT 1339.030 602.195 1341.410 604.280 ;
        RECT 1342.250 602.195 1344.630 604.280 ;
        RECT 1345.470 602.195 1347.390 604.280 ;
        RECT 1348.230 602.195 1350.610 604.280 ;
        RECT 1351.450 602.195 1353.830 604.280 ;
        RECT 1354.670 602.195 1356.590 604.280 ;
        RECT 1357.430 602.195 1359.810 604.280 ;
        RECT 1360.650 602.195 1363.030 604.280 ;
        RECT 1363.870 602.195 1365.790 604.280 ;
        RECT 1366.630 602.195 1369.010 604.280 ;
        RECT 1369.850 602.195 1372.230 604.280 ;
        RECT 1373.070 602.195 1374.990 604.280 ;
        RECT 1375.830 602.195 1378.210 604.280 ;
        RECT 1379.050 602.195 1380.970 604.280 ;
        RECT 1381.810 602.195 1384.190 604.280 ;
        RECT 1385.030 602.195 1387.410 604.280 ;
        RECT 1388.250 602.195 1390.170 604.280 ;
        RECT 1391.010 602.195 1393.390 604.280 ;
        RECT 1394.230 602.195 1396.610 604.280 ;
        RECT 1397.450 602.195 1399.370 604.280 ;
        RECT 1400.210 602.195 1402.590 604.280 ;
        RECT 1403.430 602.195 1405.810 604.280 ;
        RECT 1406.650 602.195 1408.570 604.280 ;
        RECT 1409.410 602.195 1411.790 604.280 ;
        RECT 1412.630 602.195 1415.010 604.280 ;
        RECT 1415.850 602.195 1417.770 604.280 ;
        RECT 1418.610 602.195 1420.990 604.280 ;
        RECT 1421.830 602.195 1424.210 604.280 ;
        RECT 1425.050 602.195 1426.970 604.280 ;
        RECT 1427.810 602.195 1430.190 604.280 ;
        RECT 1431.030 602.195 1433.410 604.280 ;
        RECT 1434.250 602.195 1436.170 604.280 ;
        RECT 1437.010 602.195 1439.390 604.280 ;
        RECT 1440.230 602.195 1442.610 604.280 ;
        RECT 1443.450 602.195 1445.370 604.280 ;
        RECT 1446.210 602.195 1448.590 604.280 ;
        RECT 1449.430 602.195 1451.810 604.280 ;
        RECT 1452.650 602.195 1454.570 604.280 ;
        RECT 1455.410 602.195 1457.790 604.280 ;
        RECT 1458.630 602.195 1461.010 604.280 ;
        RECT 1461.850 602.195 1463.770 604.280 ;
        RECT 1464.610 602.195 1466.990 604.280 ;
        RECT 1467.830 602.195 1469.750 604.280 ;
        RECT 1470.590 602.195 1472.970 604.280 ;
        RECT 1473.810 602.195 1476.190 604.280 ;
        RECT 1477.030 602.195 1478.950 604.280 ;
        RECT 1479.790 602.195 1482.170 604.280 ;
        RECT 1483.010 602.195 1485.390 604.280 ;
        RECT 1486.230 602.195 1488.150 604.280 ;
        RECT 1488.990 602.195 1491.370 604.280 ;
        RECT 1492.210 602.195 1494.590 604.280 ;
        RECT 1495.430 602.195 1497.350 604.280 ;
        RECT 1498.190 602.195 1500.570 604.280 ;
        RECT 1501.410 602.195 1503.790 604.280 ;
        RECT 1504.630 602.195 1506.550 604.280 ;
        RECT 1507.390 602.195 1509.770 604.280 ;
        RECT 1510.610 602.195 1512.990 604.280 ;
        RECT 1513.830 602.195 1515.750 604.280 ;
        RECT 1516.590 602.195 1518.970 604.280 ;
        RECT 1519.810 602.195 1522.190 604.280 ;
        RECT 1523.030 602.195 1524.950 604.280 ;
        RECT 1525.790 602.195 1528.170 604.280 ;
        RECT 1529.010 602.195 1531.390 604.280 ;
        RECT 1532.230 602.195 1534.150 604.280 ;
        RECT 1534.990 602.195 1537.370 604.280 ;
        RECT 1538.210 602.195 1540.590 604.280 ;
        RECT 1541.430 602.195 1543.350 604.280 ;
        RECT 1544.190 602.195 1546.570 604.280 ;
        RECT 1547.410 602.195 1549.790 604.280 ;
        RECT 1550.630 602.195 1552.550 604.280 ;
        RECT 1553.390 602.195 1555.770 604.280 ;
        RECT 1556.610 602.195 1558.530 604.280 ;
        RECT 1559.370 602.195 1561.750 604.280 ;
        RECT 1562.590 602.195 1564.970 604.280 ;
        RECT 1565.810 602.195 1567.730 604.280 ;
        RECT 1568.570 602.195 1570.950 604.280 ;
        RECT 1571.790 602.195 1574.170 604.280 ;
        RECT 1575.010 602.195 1576.930 604.280 ;
        RECT 1577.770 602.195 1580.150 604.280 ;
        RECT 1580.990 602.195 1583.370 604.280 ;
        RECT 1584.210 602.195 1586.130 604.280 ;
        RECT 1586.970 602.195 1589.350 604.280 ;
        RECT 1590.190 602.195 1592.570 604.280 ;
        RECT 1593.410 602.195 1595.330 604.280 ;
        RECT 1596.170 602.195 1598.550 604.280 ;
        RECT 1599.390 602.195 1601.770 604.280 ;
        RECT 1602.610 602.195 1604.530 604.280 ;
        RECT 1605.370 602.195 1607.750 604.280 ;
        RECT 1608.590 602.195 1610.970 604.280 ;
        RECT 1611.810 602.195 1613.730 604.280 ;
        RECT 1614.570 602.195 1616.950 604.280 ;
        RECT 1617.790 602.195 1620.170 604.280 ;
        RECT 1621.010 602.195 1622.930 604.280 ;
        RECT 1623.770 602.195 1626.150 604.280 ;
        RECT 1626.990 602.195 1629.370 604.280 ;
        RECT 1630.210 602.195 1632.130 604.280 ;
        RECT 1632.970 602.195 1635.350 604.280 ;
        RECT 1636.190 602.195 1638.570 604.280 ;
        RECT 1639.410 602.195 1641.330 604.280 ;
        RECT 1642.170 602.195 1644.550 604.280 ;
        RECT 1645.390 602.195 1647.310 604.280 ;
        RECT 1648.150 602.195 1650.530 604.280 ;
        RECT 1651.370 602.195 1653.750 604.280 ;
        RECT 1654.590 602.195 1656.510 604.280 ;
        RECT 1657.350 602.195 1659.730 604.280 ;
        RECT 1660.570 602.195 1662.950 604.280 ;
        RECT 1663.790 602.195 1665.710 604.280 ;
        RECT 1666.550 602.195 1668.930 604.280 ;
        RECT 1669.770 602.195 1672.150 604.280 ;
        RECT 1672.990 602.195 1674.910 604.280 ;
        RECT 1675.750 602.195 1678.130 604.280 ;
        RECT 1678.970 602.195 1681.350 604.280 ;
        RECT 1682.190 602.195 1684.110 604.280 ;
        RECT 1684.950 602.195 1687.330 604.280 ;
        RECT 1688.170 602.195 1690.550 604.280 ;
        RECT 1691.390 602.195 1693.310 604.280 ;
        RECT 1694.150 602.195 1696.530 604.280 ;
        RECT 1697.370 602.195 1699.750 604.280 ;
        RECT 1700.590 602.195 1702.510 604.280 ;
        RECT 1703.350 602.195 1705.730 604.280 ;
        RECT 1706.570 602.195 1708.950 604.280 ;
        RECT 1709.790 602.195 1711.710 604.280 ;
        RECT 1712.550 602.195 1714.930 604.280 ;
        RECT 1715.770 602.195 1718.150 604.280 ;
        RECT 1718.990 602.195 1720.910 604.280 ;
        RECT 1721.750 602.195 1724.130 604.280 ;
        RECT 1724.970 602.195 1727.350 604.280 ;
        RECT 1728.190 602.195 1730.110 604.280 ;
        RECT 1730.950 602.195 1733.330 604.280 ;
        RECT 1734.170 602.195 1736.090 604.280 ;
        RECT 1736.930 602.195 1739.310 604.280 ;
        RECT 1740.150 602.195 1742.530 604.280 ;
        RECT 1743.370 602.195 1745.290 604.280 ;
        RECT 1746.130 602.195 1748.510 604.280 ;
        RECT 1749.350 602.195 1751.730 604.280 ;
        RECT 1752.570 602.195 1754.490 604.280 ;
        RECT 1755.330 602.195 1757.710 604.280 ;
        RECT 1758.550 602.195 1760.930 604.280 ;
        RECT 1761.770 602.195 1763.690 604.280 ;
        RECT 1764.530 602.195 1766.910 604.280 ;
        RECT 1767.750 602.195 1770.130 604.280 ;
        RECT 1770.970 602.195 1772.890 604.280 ;
        RECT 1773.730 602.195 1776.110 604.280 ;
        RECT 1776.950 602.195 1779.330 604.280 ;
        RECT 1780.170 602.195 1782.090 604.280 ;
        RECT 1782.930 602.195 1785.310 604.280 ;
        RECT 1786.150 602.195 1788.530 604.280 ;
        RECT 1789.370 602.195 1791.290 604.280 ;
        RECT 1792.130 602.195 1794.510 604.280 ;
        RECT 1795.350 602.195 1797.730 604.280 ;
        RECT 1798.570 602.195 1800.490 604.280 ;
        RECT 1801.330 602.195 1803.710 604.280 ;
        RECT 1804.550 602.195 1806.930 604.280 ;
        RECT 1807.770 602.195 1809.690 604.280 ;
        RECT 1810.530 602.195 1812.910 604.280 ;
        RECT 1813.750 602.195 1816.130 604.280 ;
        RECT 1816.970 602.195 1818.890 604.280 ;
        RECT 1819.730 602.195 1822.110 604.280 ;
        RECT 1822.950 602.195 1824.870 604.280 ;
        RECT 1825.710 602.195 1828.090 604.280 ;
        RECT 1828.930 602.195 1831.310 604.280 ;
        RECT 1832.150 602.195 1834.070 604.280 ;
        RECT 1834.910 602.195 1837.290 604.280 ;
        RECT 1838.130 602.195 1840.510 604.280 ;
        RECT 1841.350 602.195 1843.270 604.280 ;
        RECT 1844.110 602.195 1846.490 604.280 ;
        RECT 1847.330 602.195 1849.710 604.280 ;
        RECT 1850.550 602.195 1852.470 604.280 ;
        RECT 1853.310 602.195 1855.690 604.280 ;
        RECT 1856.530 602.195 1858.910 604.280 ;
        RECT 1859.750 602.195 1861.670 604.280 ;
        RECT 1862.510 602.195 1864.890 604.280 ;
        RECT 1865.730 602.195 1868.110 604.280 ;
        RECT 1868.950 602.195 1870.870 604.280 ;
        RECT 1871.710 602.195 1874.090 604.280 ;
        RECT 1874.930 602.195 1877.310 604.280 ;
        RECT 1878.150 602.195 1880.070 604.280 ;
        RECT 1880.910 602.195 1883.290 604.280 ;
        RECT 1884.130 602.195 1886.510 604.280 ;
        RECT 1887.350 602.195 1889.270 604.280 ;
        RECT 1890.110 602.195 1892.490 604.280 ;
        RECT 1893.330 602.195 1895.710 604.280 ;
        RECT 1896.550 602.195 1898.470 604.280 ;
        RECT 1899.310 602.195 1901.690 604.280 ;
        RECT 1902.530 602.195 1904.910 604.280 ;
        RECT 1905.750 602.195 1907.670 604.280 ;
        RECT 1908.510 602.195 1910.890 604.280 ;
        RECT 1911.730 602.195 1913.650 604.280 ;
        RECT 1914.490 602.195 1916.870 604.280 ;
        RECT 1917.710 602.195 1920.090 604.280 ;
        RECT 1920.930 602.195 1922.850 604.280 ;
        RECT 1923.690 602.195 1926.070 604.280 ;
        RECT 1926.910 602.195 1929.290 604.280 ;
        RECT 1930.130 602.195 1932.050 604.280 ;
        RECT 1932.890 602.195 1935.270 604.280 ;
        RECT 1936.110 602.195 1938.490 604.280 ;
        RECT 1939.330 602.195 1941.250 604.280 ;
        RECT 1942.090 602.195 1944.470 604.280 ;
        RECT 1945.310 602.195 1947.690 604.280 ;
        RECT 1948.530 602.195 1950.450 604.280 ;
        RECT 1951.290 602.195 1953.670 604.280 ;
        RECT 1954.510 602.195 1956.890 604.280 ;
        RECT 1957.730 602.195 1959.650 604.280 ;
        RECT 1960.490 602.195 1962.870 604.280 ;
        RECT 1963.710 602.195 1966.090 604.280 ;
        RECT 1966.930 602.195 1968.850 604.280 ;
        RECT 1969.690 602.195 1972.070 604.280 ;
        RECT 1972.910 602.195 1975.290 604.280 ;
        RECT 1976.130 602.195 1978.050 604.280 ;
        RECT 1978.890 602.195 1981.270 604.280 ;
        RECT 1982.110 602.195 1984.490 604.280 ;
        RECT 1985.330 602.195 1987.250 604.280 ;
        RECT 1988.090 602.195 1990.470 604.280 ;
        RECT 1991.310 602.195 1993.690 604.280 ;
        RECT 1994.530 602.195 1996.450 604.280 ;
        RECT 1997.290 602.195 1999.670 604.280 ;
        RECT 2000.510 602.195 2002.430 604.280 ;
        RECT 2003.270 602.195 2005.650 604.280 ;
        RECT 2006.490 602.195 2008.870 604.280 ;
        RECT 2009.710 602.195 2011.630 604.280 ;
        RECT 2012.470 602.195 2014.850 604.280 ;
        RECT 2015.690 602.195 2018.070 604.280 ;
        RECT 2018.910 602.195 2020.830 604.280 ;
        RECT 2021.670 602.195 2024.050 604.280 ;
        RECT 2024.890 602.195 2027.270 604.280 ;
        RECT 2028.110 602.195 2030.030 604.280 ;
        RECT 2030.870 602.195 2033.250 604.280 ;
        RECT 2034.090 602.195 2036.470 604.280 ;
        RECT 2037.310 602.195 2039.230 604.280 ;
        RECT 2040.070 602.195 2042.450 604.280 ;
        RECT 2043.290 602.195 2045.670 604.280 ;
        RECT 2046.510 602.195 2048.430 604.280 ;
        RECT 2049.270 602.195 2051.650 604.280 ;
        RECT 2052.490 602.195 2054.870 604.280 ;
        RECT 2055.710 602.195 2057.630 604.280 ;
        RECT 2058.470 602.195 2060.850 604.280 ;
        RECT 2061.690 602.195 2064.070 604.280 ;
        RECT 2064.910 602.195 2066.830 604.280 ;
        RECT 2067.670 602.195 2070.050 604.280 ;
        RECT 2070.890 602.195 2073.270 604.280 ;
        RECT 2074.110 602.195 2076.030 604.280 ;
        RECT 2076.870 602.195 2079.250 604.280 ;
        RECT 2080.090 602.195 2082.470 604.280 ;
        RECT 2083.310 602.195 2085.230 604.280 ;
        RECT 2086.070 602.195 2088.450 604.280 ;
        RECT 2089.290 602.195 2091.210 604.280 ;
        RECT 2092.050 602.195 2094.430 604.280 ;
        RECT 2095.270 602.195 2097.650 604.280 ;
        RECT 2098.490 602.195 2100.410 604.280 ;
        RECT 2101.250 602.195 2103.630 604.280 ;
        RECT 2104.470 602.195 2106.850 604.280 ;
        RECT 2107.690 602.195 2109.610 604.280 ;
        RECT 2110.450 602.195 2112.830 604.280 ;
        RECT 2113.670 602.195 2116.050 604.280 ;
        RECT 2116.890 602.195 2118.810 604.280 ;
        RECT 2119.650 602.195 2122.030 604.280 ;
        RECT 2122.870 602.195 2125.250 604.280 ;
        RECT 2126.090 602.195 2128.010 604.280 ;
        RECT 2128.850 602.195 2131.230 604.280 ;
        RECT 2132.070 602.195 2134.450 604.280 ;
        RECT 2135.290 602.195 2137.210 604.280 ;
        RECT 2138.050 602.195 2140.430 604.280 ;
        RECT 2141.270 602.195 2143.650 604.280 ;
        RECT 2144.490 602.195 2146.410 604.280 ;
        RECT 2147.250 602.195 2149.630 604.280 ;
        RECT 2150.470 602.195 2152.850 604.280 ;
        RECT 2153.690 602.195 2155.610 604.280 ;
        RECT 2156.450 602.195 2158.830 604.280 ;
        RECT 2159.670 602.195 2162.050 604.280 ;
        RECT 2162.890 602.195 2164.810 604.280 ;
        RECT 2165.650 602.195 2168.030 604.280 ;
        RECT 2168.870 602.195 2169.040 604.280 ;
      LAYER via2 ;
        RECT 420.530 2729.040 420.810 2729.320 ;
        RECT 420.070 2707.280 420.350 2707.560 ;
        RECT 588.890 2686.880 589.170 2687.160 ;
        RECT 588.890 2666.480 589.170 2666.760 ;
        RECT 978.510 1013.400 978.790 1013.680 ;
        RECT 978.970 1012.720 979.250 1013.000 ;
        RECT 993.230 2783.440 993.510 2783.720 ;
        RECT 992.770 2760.320 993.050 2760.600 ;
        RECT 992.310 2718.840 992.590 2719.120 ;
        RECT 991.850 2692.320 992.130 2692.600 ;
        RECT 991.390 2622.960 991.670 2623.240 ;
        RECT 990.930 1998.040 991.210 1998.320 ;
        RECT 990.470 1955.880 990.750 1956.160 ;
        RECT 990.010 1935.480 990.290 1935.760 ;
        RECT 989.550 1893.320 989.830 1893.600 ;
        RECT 989.090 1851.160 989.370 1851.440 ;
        RECT 988.630 1809.000 988.910 1809.280 ;
        RECT 988.170 1787.240 988.450 1787.520 ;
        RECT 987.710 1766.840 987.990 1767.120 ;
        RECT 987.250 1745.080 987.530 1745.360 ;
        RECT 986.330 1014.080 986.610 1014.360 ;
        RECT 985.870 1012.040 986.150 1012.320 ;
        RECT 985.410 1011.360 985.690 1011.640 ;
        RECT 994.610 2739.240 994.890 2739.520 ;
        RECT 993.690 2670.560 993.970 2670.840 ;
        RECT 993.230 1010.000 993.510 1010.280 ;
        RECT 994.150 2646.080 994.430 2646.360 ;
        RECT 995.070 2018.440 995.350 2018.720 ;
        RECT 995.530 1976.280 995.810 1976.560 ;
        RECT 995.990 1913.720 996.270 1914.000 ;
        RECT 996.450 1871.560 996.730 1871.840 ;
        RECT 995.070 1010.680 995.350 1010.960 ;
        RECT 996.910 1829.400 997.190 1829.680 ;
        RECT 997.370 1724.680 997.650 1724.960 ;
        RECT 1110.990 2780.720 1111.270 2781.000 ;
        RECT 1097.190 2644.720 1097.470 2645.000 ;
        RECT 1097.650 2622.280 1097.930 2622.560 ;
        RECT 1111.450 2760.320 1111.730 2760.600 ;
        RECT 1111.910 2734.480 1112.190 2734.760 ;
        RECT 1112.370 2712.720 1112.650 2713.000 ;
        RECT 1112.830 2691.640 1113.110 2691.920 ;
        RECT 1113.290 2666.480 1113.570 2666.760 ;
        RECT 1067.290 1010.000 1067.570 1010.280 ;
        RECT 1101.790 1014.080 1102.070 1014.360 ;
        RECT 1119.270 1013.400 1119.550 1013.680 ;
        RECT 1131.690 1012.720 1131.970 1013.000 ;
        RECT 1143.190 1012.040 1143.470 1012.320 ;
        RECT 1167.110 1011.360 1167.390 1011.640 ;
        RECT 1263.250 1012.040 1263.530 1012.320 ;
        RECT 1267.390 1011.360 1267.670 1011.640 ;
        RECT 1290.850 1634.920 1291.130 1635.200 ;
        RECT 1291.770 1634.920 1292.050 1635.200 ;
        RECT 1277.970 1545.840 1278.250 1546.120 ;
        RECT 1279.350 1545.840 1279.630 1546.120 ;
        RECT 1291.770 1545.840 1292.050 1546.120 ;
        RECT 1293.150 1545.840 1293.430 1546.120 ;
        RECT 1289.930 1207.200 1290.210 1207.480 ;
        RECT 1290.850 1207.200 1291.130 1207.480 ;
        RECT 1269.690 1011.360 1269.970 1011.640 ;
        RECT 1270.610 1012.040 1270.890 1012.320 ;
        RECT 1292.690 1011.360 1292.970 1011.640 ;
        RECT 1297.290 1011.360 1297.570 1011.640 ;
        RECT 1309.710 1010.680 1309.990 1010.960 ;
        RECT 1334.090 1998.040 1334.370 1998.320 ;
        RECT 1334.550 1913.720 1334.830 1914.000 ;
        RECT 1335.470 1787.240 1335.750 1787.520 ;
        RECT 1335.930 1745.080 1336.210 1745.360 ;
        RECT 1338.690 2018.440 1338.970 2018.720 ;
        RECT 1339.150 1976.280 1339.430 1976.560 ;
        RECT 1339.610 1955.880 1339.890 1956.160 ;
        RECT 1340.070 1934.120 1340.350 1934.400 ;
        RECT 1340.530 1891.960 1340.810 1892.240 ;
        RECT 1340.990 1871.560 1341.270 1871.840 ;
        RECT 1341.450 1849.800 1341.730 1850.080 ;
        RECT 1341.910 1829.400 1342.190 1829.680 ;
        RECT 1342.370 1807.640 1342.650 1807.920 ;
        RECT 1342.830 1766.840 1343.110 1767.120 ;
        RECT 1343.290 1724.680 1343.570 1724.960 ;
        RECT 1358.930 2815.400 1359.210 2815.680 ;
        RECT 1358.470 2814.720 1358.750 2815.000 ;
        RECT 1357.550 2801.120 1357.830 2801.400 ;
        RECT 1358.470 2801.120 1358.750 2801.400 ;
        RECT 1358.470 2704.560 1358.750 2704.840 ;
        RECT 1359.850 2704.560 1360.130 2704.840 ;
        RECT 1358.010 2511.440 1358.290 2511.720 ;
        RECT 1358.930 2463.160 1359.210 2463.440 ;
        RECT 1358.930 2097.320 1359.210 2097.600 ;
        RECT 1359.850 2097.320 1360.130 2097.600 ;
        RECT 1358.010 1945.680 1358.290 1945.960 ;
        RECT 1358.930 1945.680 1359.210 1945.960 ;
        RECT 1359.850 1470.360 1360.130 1470.640 ;
        RECT 1358.930 1469.680 1359.210 1469.960 ;
        RECT 1359.850 1373.800 1360.130 1374.080 ;
        RECT 1358.930 1373.120 1359.210 1373.400 ;
        RECT 1358.010 1276.560 1358.290 1276.840 ;
        RECT 1358.930 1276.560 1359.210 1276.840 ;
        RECT 1406.310 2609.360 1406.590 2609.640 ;
        RECT 1406.770 2608.170 1407.050 2608.450 ;
        RECT 1386.530 1010.680 1386.810 1010.960 ;
        RECT 1405.390 2463.160 1405.670 2463.440 ;
        RECT 1406.310 2463.160 1406.590 2463.440 ;
        RECT 1405.390 2270.040 1405.670 2270.320 ;
        RECT 1406.310 2270.040 1406.590 2270.320 ;
        RECT 1405.390 2173.480 1405.670 2173.760 ;
        RECT 1406.310 2173.480 1406.590 2173.760 ;
        RECT 1408.150 1980.360 1408.430 1980.640 ;
        RECT 1408.150 1979.680 1408.430 1979.960 ;
        RECT 1405.850 1303.760 1406.130 1304.040 ;
        RECT 1405.390 1255.480 1405.670 1255.760 ;
        RECT 1483.590 2850.080 1483.870 2850.360 ;
        RECT 1482.210 2830.360 1482.490 2830.640 ;
        RECT 1489.570 2801.800 1489.850 2802.080 ;
        RECT 1489.110 2784.120 1489.390 2784.400 ;
        RECT 1489.110 2767.800 1489.390 2768.080 ;
        RECT 1488.650 2753.520 1488.930 2753.800 ;
        RECT 1488.190 2691.640 1488.470 2691.920 ;
        RECT 1488.190 2673.960 1488.470 2674.240 ;
        RECT 1482.670 2657.640 1482.950 2657.920 ;
        RECT 1487.270 2629.080 1487.550 2629.360 ;
        RECT 1487.730 2610.040 1488.010 2610.320 ;
        RECT 1487.270 2595.080 1487.550 2595.360 ;
        RECT 1487.270 2580.800 1487.550 2581.080 ;
        RECT 1487.270 2567.200 1487.550 2567.480 ;
        RECT 1483.590 2547.480 1483.870 2547.760 ;
        RECT 1486.810 2518.920 1487.090 2519.200 ;
        RECT 1495.550 2739.240 1495.830 2739.520 ;
        RECT 1495.090 2720.200 1495.370 2720.480 ;
        RECT 1511.190 1012.720 1511.470 1013.000 ;
        RECT 1535.110 2415.560 1535.390 2415.840 ;
        RECT 1535.110 2414.880 1535.390 2415.160 ;
        RECT 1535.110 2319.000 1535.390 2319.280 ;
        RECT 1535.110 2318.320 1535.390 2318.600 ;
        RECT 1534.190 2270.040 1534.470 2270.320 ;
        RECT 1535.110 2270.040 1535.390 2270.320 ;
        RECT 1521.310 1010.000 1521.590 1010.280 ;
        RECT 1536.030 1012.720 1536.310 1013.000 ;
        RECT 1544.310 1256.840 1544.590 1257.120 ;
        RECT 1544.310 1256.160 1544.590 1256.440 ;
        RECT 1536.490 1010.000 1536.770 1010.280 ;
        RECT 1890.690 2848.380 1890.970 2848.660 ;
        RECT 1891.150 2832.060 1891.430 2832.340 ;
        RECT 1891.610 2817.100 1891.890 2817.380 ;
        RECT 1892.070 2797.720 1892.350 2798.000 ;
        RECT 1892.990 2782.760 1893.270 2783.040 ;
        RECT 1892.530 2608.680 1892.810 2608.960 ;
        RECT 1893.450 2753.520 1893.730 2753.800 ;
        RECT 1894.370 2735.160 1894.650 2735.440 ;
        RECT 1897.590 2767.120 1897.870 2767.400 ;
        RECT 1898.050 2718.840 1898.330 2719.120 ;
        RECT 1898.510 2687.560 1898.790 2687.840 ;
        RECT 1898.970 2672.600 1899.250 2672.880 ;
        RECT 1899.430 2656.960 1899.710 2657.240 ;
        RECT 1899.890 2625.000 1900.170 2625.280 ;
        RECT 1892.070 1010.680 1892.350 1010.960 ;
        RECT 1900.350 2577.400 1900.630 2577.680 ;
        RECT 1900.810 2562.440 1901.090 2562.720 ;
        RECT 1901.270 2547.480 1901.550 2547.760 ;
        RECT 1903.570 2514.840 1903.850 2515.120 ;
        RECT 1904.490 1885.840 1904.770 1886.120 ;
        RECT 1904.490 1870.200 1904.770 1870.480 ;
        RECT 1904.490 1851.840 1904.770 1852.120 ;
        RECT 1904.490 1817.840 1904.770 1818.120 ;
        RECT 1904.490 1767.520 1904.770 1767.800 ;
        RECT 2087.110 1884.480 2087.390 1884.760 ;
        RECT 2084.350 1850.480 2084.630 1850.760 ;
        RECT 2084.810 1835.520 2085.090 1835.800 ;
        RECT 2085.270 1816.480 2085.550 1816.760 ;
        RECT 2085.730 1800.840 2086.010 1801.120 ;
        RECT 2086.190 1782.480 2086.470 1782.760 ;
        RECT 2086.650 1766.840 2086.930 1767.120 ;
        RECT 2283.990 1875.640 2284.270 1875.920 ;
        RECT 2287.210 1789.960 2287.490 1790.240 ;
        RECT 2523.650 1891.960 2523.930 1892.240 ;
        RECT 2523.650 1802.200 2523.930 1802.480 ;
        RECT 2518.590 1704.280 2518.870 1704.560 ;
        RECT 2523.650 1717.880 2523.930 1718.160 ;
        RECT 2519.510 1704.280 2519.790 1704.560 ;
        RECT 2519.510 1608.400 2519.790 1608.680 ;
        RECT 2519.510 1607.040 2519.790 1607.320 ;
      LAYER met3 ;
        RECT 1504.000 2881.840 1885.335 2889.125 ;
        RECT 1504.400 2880.480 1885.335 2881.840 ;
        RECT 1504.400 2880.440 1884.935 2880.480 ;
        RECT 1504.000 2879.080 1884.935 2880.440 ;
        RECT 1504.000 2865.520 1885.335 2879.080 ;
        RECT 1504.400 2864.160 1885.335 2865.520 ;
        RECT 1504.400 2864.120 1884.935 2864.160 ;
        RECT 1504.000 2862.760 1884.935 2864.120 ;
        RECT 1504.000 2850.560 1885.335 2862.760 ;
      LAYER met3 ;
        RECT 1483.565 2850.370 1483.895 2850.385 ;
        RECT 1483.565 2850.160 1500.210 2850.370 ;
        RECT 1483.565 2850.070 1504.000 2850.160 ;
        RECT 1483.565 2850.055 1483.895 2850.070 ;
        RECT 1499.910 2849.880 1504.000 2850.070 ;
        RECT 1500.000 2849.560 1504.000 2849.880 ;
      LAYER met3 ;
        RECT 1504.400 2849.200 1885.335 2850.560 ;
        RECT 1504.400 2849.160 1884.935 2849.200 ;
        RECT 1504.000 2847.800 1884.935 2849.160 ;
      LAYER met3 ;
        RECT 1885.335 2848.670 1889.335 2848.800 ;
        RECT 1890.665 2848.670 1890.995 2848.685 ;
        RECT 1885.335 2848.370 1890.995 2848.670 ;
        RECT 1885.335 2848.200 1889.335 2848.370 ;
        RECT 1890.665 2848.355 1890.995 2848.370 ;
      LAYER met3 ;
        RECT 1504.000 2834.240 1885.335 2847.800 ;
      LAYER met3 ;
        RECT 1500.000 2833.560 1504.000 2833.840 ;
        RECT 1499.910 2833.240 1504.000 2833.560 ;
        RECT 1482.185 2830.650 1482.515 2830.665 ;
        RECT 1499.910 2830.650 1500.210 2833.240 ;
      LAYER met3 ;
        RECT 1504.400 2832.880 1885.335 2834.240 ;
        RECT 1504.400 2832.840 1884.935 2832.880 ;
      LAYER met3 ;
        RECT 1482.185 2830.350 1500.210 2830.650 ;
      LAYER met3 ;
        RECT 1504.000 2831.480 1884.935 2832.840 ;
      LAYER met3 ;
        RECT 1885.335 2832.350 1889.335 2832.480 ;
        RECT 1891.125 2832.350 1891.455 2832.365 ;
        RECT 1885.335 2832.050 1891.455 2832.350 ;
        RECT 1885.335 2831.880 1889.335 2832.050 ;
        RECT 1891.125 2832.035 1891.455 2832.050 ;
        RECT 1482.185 2830.335 1482.515 2830.350 ;
      LAYER met3 ;
        RECT 1504.000 2819.280 1885.335 2831.480 ;
        RECT 1504.400 2817.920 1885.335 2819.280 ;
        RECT 1504.400 2817.880 1884.935 2817.920 ;
        RECT 1504.000 2816.520 1884.935 2817.880 ;
      LAYER met3 ;
        RECT 1885.335 2817.390 1889.335 2817.520 ;
        RECT 1891.585 2817.390 1891.915 2817.405 ;
        RECT 1885.335 2817.090 1891.915 2817.390 ;
        RECT 1885.335 2816.920 1889.335 2817.090 ;
        RECT 1891.585 2817.075 1891.915 2817.090 ;
        RECT 1358.905 2815.690 1359.235 2815.705 ;
        RECT 1358.230 2815.390 1359.235 2815.690 ;
        RECT 1358.230 2815.025 1358.530 2815.390 ;
        RECT 1358.905 2815.375 1359.235 2815.390 ;
        RECT 1358.230 2814.710 1358.775 2815.025 ;
        RECT 1358.445 2814.695 1358.775 2814.710 ;
      LAYER met3 ;
        RECT 1504.000 2802.960 1885.335 2816.520 ;
      LAYER met3 ;
        RECT 1500.000 2802.280 1504.000 2802.560 ;
        RECT 1489.545 2802.090 1489.875 2802.105 ;
        RECT 1499.910 2802.090 1504.000 2802.280 ;
        RECT 1489.545 2801.960 1504.000 2802.090 ;
        RECT 1489.545 2801.790 1500.210 2801.960 ;
        RECT 1489.545 2801.775 1489.875 2801.790 ;
      LAYER met3 ;
        RECT 1504.400 2801.600 1885.335 2802.960 ;
        RECT 1504.400 2801.560 1884.935 2801.600 ;
      LAYER met3 ;
        RECT 1357.525 2801.410 1357.855 2801.425 ;
        RECT 1358.445 2801.410 1358.775 2801.425 ;
        RECT 1357.525 2801.110 1358.775 2801.410 ;
        RECT 1357.525 2801.095 1357.855 2801.110 ;
        RECT 1358.445 2801.095 1358.775 2801.110 ;
      LAYER met3 ;
        RECT 1504.000 2800.200 1884.935 2801.560 ;
      LAYER met3 ;
        RECT 1885.335 2800.920 1889.335 2801.200 ;
        RECT 1885.335 2800.600 1889.370 2800.920 ;
      LAYER met3 ;
        RECT 1504.000 2788.000 1885.335 2800.200 ;
      LAYER met3 ;
        RECT 1889.070 2798.010 1889.370 2800.600 ;
        RECT 1892.045 2798.010 1892.375 2798.025 ;
        RECT 1889.070 2797.710 1892.375 2798.010 ;
        RECT 1892.045 2797.695 1892.375 2797.710 ;
      LAYER met3 ;
        RECT 1004.000 2787.360 1096.000 2787.845 ;
      LAYER met3 ;
        RECT 1000.000 2786.360 1004.000 2786.960 ;
        RECT 993.205 2783.730 993.535 2783.745 ;
        RECT 1000.350 2783.730 1000.650 2786.360 ;
      LAYER met3 ;
        RECT 1004.400 2785.960 1096.000 2787.360 ;
      LAYER met3 ;
        RECT 1500.000 2787.320 1504.000 2787.600 ;
        RECT 993.205 2783.430 1000.650 2783.730 ;
      LAYER met3 ;
        RECT 1004.000 2784.640 1096.000 2785.960 ;
      LAYER met3 ;
        RECT 1499.910 2787.000 1504.000 2787.320 ;
        RECT 993.205 2783.415 993.535 2783.430 ;
      LAYER met3 ;
        RECT 1004.000 2783.240 1095.600 2784.640 ;
      LAYER met3 ;
        RECT 1489.085 2784.410 1489.415 2784.425 ;
        RECT 1499.910 2784.410 1500.210 2787.000 ;
      LAYER met3 ;
        RECT 1504.400 2786.640 1885.335 2788.000 ;
        RECT 1504.400 2786.600 1884.935 2786.640 ;
      LAYER met3 ;
        RECT 1096.000 2783.920 1100.000 2784.240 ;
        RECT 1489.085 2784.110 1500.210 2784.410 ;
      LAYER met3 ;
        RECT 1504.000 2785.240 1884.935 2786.600 ;
      LAYER met3 ;
        RECT 1885.335 2785.960 1889.335 2786.240 ;
        RECT 1885.335 2785.640 1889.370 2785.960 ;
        RECT 1489.085 2784.095 1489.415 2784.110 ;
        RECT 1096.000 2783.640 1100.010 2783.920 ;
      LAYER met3 ;
        RECT 1004.000 2764.240 1096.000 2783.240 ;
      LAYER met3 ;
        RECT 1099.710 2781.010 1100.010 2783.640 ;
        RECT 1110.965 2781.010 1111.295 2781.025 ;
        RECT 1099.710 2780.710 1111.295 2781.010 ;
        RECT 1110.965 2780.695 1111.295 2780.710 ;
      LAYER met3 ;
        RECT 1504.000 2771.680 1885.335 2785.240 ;
      LAYER met3 ;
        RECT 1889.070 2783.050 1889.370 2785.640 ;
        RECT 1892.965 2783.050 1893.295 2783.065 ;
        RECT 1889.070 2782.750 1893.295 2783.050 ;
        RECT 1892.965 2782.735 1893.295 2782.750 ;
        RECT 1500.000 2771.000 1504.000 2771.280 ;
        RECT 1499.910 2770.680 1504.000 2771.000 ;
        RECT 1489.085 2768.090 1489.415 2768.105 ;
        RECT 1499.910 2768.090 1500.210 2770.680 ;
      LAYER met3 ;
        RECT 1504.400 2770.320 1885.335 2771.680 ;
        RECT 1504.400 2770.280 1884.935 2770.320 ;
      LAYER met3 ;
        RECT 1489.085 2767.790 1500.210 2768.090 ;
      LAYER met3 ;
        RECT 1504.000 2768.920 1884.935 2770.280 ;
      LAYER met3 ;
        RECT 1885.335 2769.640 1889.335 2769.920 ;
        RECT 1885.335 2769.320 1889.370 2769.640 ;
        RECT 1489.085 2767.775 1489.415 2767.790 ;
        RECT 1000.000 2763.240 1004.000 2763.840 ;
        RECT 992.745 2760.610 993.075 2760.625 ;
        RECT 1000.350 2760.610 1000.650 2763.240 ;
      LAYER met3 ;
        RECT 1004.400 2762.840 1096.000 2764.240 ;
      LAYER met3 ;
        RECT 992.745 2760.310 1000.650 2760.610 ;
      LAYER met3 ;
        RECT 1004.000 2761.520 1096.000 2762.840 ;
      LAYER met3 ;
        RECT 992.745 2760.295 993.075 2760.310 ;
      LAYER met3 ;
        RECT 1004.000 2760.120 1095.600 2761.520 ;
      LAYER met3 ;
        RECT 1096.000 2760.800 1100.000 2761.120 ;
        RECT 1096.000 2760.610 1100.010 2760.800 ;
        RECT 1111.425 2760.610 1111.755 2760.625 ;
        RECT 1096.000 2760.520 1111.755 2760.610 ;
        RECT 1099.710 2760.310 1111.755 2760.520 ;
        RECT 1111.425 2760.295 1111.755 2760.310 ;
      LAYER met3 ;
        RECT 434.400 2751.960 574.800 2752.825 ;
        RECT 434.000 2734.320 574.800 2751.960 ;
        RECT 1004.000 2741.120 1096.000 2760.120 ;
        RECT 1504.000 2755.360 1885.335 2768.920 ;
      LAYER met3 ;
        RECT 1889.070 2767.410 1889.370 2769.320 ;
        RECT 1897.565 2767.410 1897.895 2767.425 ;
        RECT 1889.070 2767.110 1897.895 2767.410 ;
        RECT 1897.565 2767.095 1897.895 2767.110 ;
        RECT 1500.000 2754.680 1504.000 2754.960 ;
        RECT 1499.910 2754.360 1504.000 2754.680 ;
        RECT 1488.625 2753.810 1488.955 2753.825 ;
        RECT 1499.910 2753.810 1500.210 2754.360 ;
      LAYER met3 ;
        RECT 1504.400 2754.000 1885.335 2755.360 ;
        RECT 1504.400 2753.960 1884.935 2754.000 ;
      LAYER met3 ;
        RECT 1488.625 2753.510 1500.210 2753.810 ;
        RECT 1488.625 2753.495 1488.955 2753.510 ;
        RECT 1000.000 2740.120 1004.000 2740.720 ;
        RECT 994.585 2739.530 994.915 2739.545 ;
        RECT 1000.350 2739.530 1000.650 2740.120 ;
      LAYER met3 ;
        RECT 1004.400 2739.720 1096.000 2741.120 ;
        RECT 1504.000 2752.600 1884.935 2753.960 ;
      LAYER met3 ;
        RECT 1893.425 2753.810 1893.755 2753.825 ;
        RECT 1889.070 2753.600 1893.755 2753.810 ;
        RECT 1885.335 2753.510 1893.755 2753.600 ;
        RECT 1885.335 2753.320 1889.370 2753.510 ;
        RECT 1893.425 2753.495 1893.755 2753.510 ;
        RECT 1885.335 2753.000 1889.335 2753.320 ;
      LAYER met3 ;
        RECT 1504.000 2740.400 1885.335 2752.600 ;
      LAYER met3 ;
        RECT 1500.000 2739.720 1504.000 2740.000 ;
        RECT 994.585 2739.230 1000.650 2739.530 ;
        RECT 994.585 2739.215 994.915 2739.230 ;
      LAYER met3 ;
        RECT 1004.000 2738.400 1096.000 2739.720 ;
      LAYER met3 ;
        RECT 1495.525 2739.530 1495.855 2739.545 ;
        RECT 1499.910 2739.530 1504.000 2739.720 ;
        RECT 1495.525 2739.400 1504.000 2739.530 ;
        RECT 1495.525 2739.230 1500.210 2739.400 ;
        RECT 1495.525 2739.215 1495.855 2739.230 ;
      LAYER met3 ;
        RECT 1504.400 2739.040 1885.335 2740.400 ;
        RECT 1504.400 2739.000 1884.935 2739.040 ;
        RECT 1004.000 2737.000 1095.600 2738.400 ;
      LAYER met3 ;
        RECT 1096.000 2737.680 1100.000 2738.000 ;
        RECT 1096.000 2737.400 1100.010 2737.680 ;
      LAYER met3 ;
        RECT 434.000 2732.960 574.400 2734.320 ;
        RECT 434.400 2732.920 574.400 2732.960 ;
      LAYER met3 ;
        RECT 430.000 2732.240 434.000 2732.560 ;
        RECT 429.950 2731.960 434.000 2732.240 ;
        RECT 420.505 2729.330 420.835 2729.345 ;
        RECT 429.950 2729.330 430.250 2731.960 ;
      LAYER met3 ;
        RECT 434.400 2731.560 574.800 2732.920 ;
      LAYER met3 ;
        RECT 420.505 2729.030 430.250 2729.330 ;
        RECT 420.505 2729.015 420.835 2729.030 ;
      LAYER met3 ;
        RECT 434.000 2712.560 574.800 2731.560 ;
        RECT 1004.000 2719.360 1096.000 2737.000 ;
      LAYER met3 ;
        RECT 1099.710 2734.770 1100.010 2737.400 ;
      LAYER met3 ;
        RECT 1504.000 2737.640 1884.935 2739.000 ;
      LAYER met3 ;
        RECT 1885.335 2738.360 1889.335 2738.640 ;
        RECT 1885.335 2738.040 1889.370 2738.360 ;
        RECT 1111.885 2734.770 1112.215 2734.785 ;
        RECT 1099.710 2734.470 1112.215 2734.770 ;
        RECT 1111.885 2734.455 1112.215 2734.470 ;
      LAYER met3 ;
        RECT 1504.000 2724.080 1885.335 2737.640 ;
      LAYER met3 ;
        RECT 1889.070 2735.450 1889.370 2738.040 ;
        RECT 1894.345 2735.450 1894.675 2735.465 ;
        RECT 1889.070 2735.150 1894.675 2735.450 ;
        RECT 1894.345 2735.135 1894.675 2735.150 ;
        RECT 1500.000 2723.400 1504.000 2723.680 ;
        RECT 1499.910 2723.080 1504.000 2723.400 ;
        RECT 1495.065 2720.490 1495.395 2720.505 ;
        RECT 1499.910 2720.490 1500.210 2723.080 ;
      LAYER met3 ;
        RECT 1504.400 2722.720 1885.335 2724.080 ;
        RECT 1504.400 2722.680 1884.935 2722.720 ;
      LAYER met3 ;
        RECT 1495.065 2720.190 1500.210 2720.490 ;
      LAYER met3 ;
        RECT 1504.000 2721.320 1884.935 2722.680 ;
      LAYER met3 ;
        RECT 1885.335 2722.040 1889.335 2722.320 ;
        RECT 1885.335 2721.720 1889.370 2722.040 ;
        RECT 1495.065 2720.175 1495.395 2720.190 ;
        RECT 992.285 2719.130 992.615 2719.145 ;
        RECT 992.285 2718.960 1000.650 2719.130 ;
        RECT 992.285 2718.830 1004.000 2718.960 ;
        RECT 992.285 2718.815 992.615 2718.830 ;
        RECT 1000.000 2718.360 1004.000 2718.830 ;
      LAYER met3 ;
        RECT 1004.400 2717.960 1096.000 2719.360 ;
        RECT 1004.000 2716.640 1096.000 2717.960 ;
        RECT 1004.000 2715.240 1095.600 2716.640 ;
      LAYER met3 ;
        RECT 1096.000 2715.920 1100.000 2716.240 ;
        RECT 1096.000 2715.640 1100.010 2715.920 ;
      LAYER met3 ;
        RECT 434.000 2711.200 574.400 2712.560 ;
        RECT 434.400 2711.160 574.400 2711.200 ;
      LAYER met3 ;
        RECT 430.000 2710.480 434.000 2710.800 ;
        RECT 429.950 2710.200 434.000 2710.480 ;
        RECT 420.045 2707.570 420.375 2707.585 ;
        RECT 429.950 2707.570 430.250 2710.200 ;
      LAYER met3 ;
        RECT 434.400 2709.800 574.800 2711.160 ;
      LAYER met3 ;
        RECT 420.045 2707.270 430.250 2707.570 ;
        RECT 420.045 2707.255 420.375 2707.270 ;
      LAYER met3 ;
        RECT 434.000 2690.800 574.800 2709.800 ;
        RECT 1004.000 2696.240 1096.000 2715.240 ;
      LAYER met3 ;
        RECT 1099.710 2713.010 1100.010 2715.640 ;
        RECT 1112.345 2713.010 1112.675 2713.025 ;
        RECT 1099.710 2712.710 1112.675 2713.010 ;
        RECT 1112.345 2712.695 1112.675 2712.710 ;
      LAYER met3 ;
        RECT 1504.000 2709.120 1885.335 2721.320 ;
      LAYER met3 ;
        RECT 1889.070 2719.130 1889.370 2721.720 ;
        RECT 1898.025 2719.130 1898.355 2719.145 ;
        RECT 1889.070 2718.830 1898.355 2719.130 ;
        RECT 1898.025 2718.815 1898.355 2718.830 ;
      LAYER met3 ;
        RECT 1504.400 2707.760 1885.335 2709.120 ;
        RECT 1504.400 2707.720 1884.935 2707.760 ;
        RECT 1504.000 2706.360 1884.935 2707.720 ;
      LAYER met3 ;
        RECT 1358.445 2704.850 1358.775 2704.865 ;
        RECT 1359.825 2704.850 1360.155 2704.865 ;
        RECT 1358.445 2704.550 1360.155 2704.850 ;
        RECT 1358.445 2704.535 1358.775 2704.550 ;
        RECT 1359.825 2704.535 1360.155 2704.550 ;
        RECT 1000.000 2695.240 1004.000 2695.840 ;
        RECT 991.825 2692.610 992.155 2692.625 ;
        RECT 1000.350 2692.610 1000.650 2695.240 ;
      LAYER met3 ;
        RECT 1004.400 2694.840 1096.000 2696.240 ;
      LAYER met3 ;
        RECT 991.825 2692.310 1000.650 2692.610 ;
      LAYER met3 ;
        RECT 1004.000 2693.520 1096.000 2694.840 ;
      LAYER met3 ;
        RECT 991.825 2692.295 992.155 2692.310 ;
      LAYER met3 ;
        RECT 1004.000 2692.120 1095.600 2693.520 ;
      LAYER met3 ;
        RECT 1096.000 2692.800 1100.000 2693.120 ;
      LAYER met3 ;
        RECT 1504.000 2692.800 1885.335 2706.360 ;
      LAYER met3 ;
        RECT 1096.000 2692.520 1100.010 2692.800 ;
      LAYER met3 ;
        RECT 434.000 2689.440 574.400 2690.800 ;
      LAYER met3 ;
        RECT 574.800 2689.800 578.800 2690.400 ;
      LAYER met3 ;
        RECT 434.400 2689.400 574.400 2689.440 ;
        RECT 434.400 2688.040 574.800 2689.400 ;
        RECT 434.000 2670.400 574.800 2688.040 ;
      LAYER met3 ;
        RECT 578.070 2687.170 578.370 2689.800 ;
        RECT 588.865 2687.170 589.195 2687.185 ;
        RECT 578.070 2686.870 589.195 2687.170 ;
        RECT 588.865 2686.855 589.195 2686.870 ;
      LAYER met3 ;
        RECT 1004.000 2673.120 1096.000 2692.120 ;
      LAYER met3 ;
        RECT 1099.710 2691.930 1100.010 2692.520 ;
        RECT 1500.000 2692.120 1504.000 2692.400 ;
        RECT 1112.805 2691.930 1113.135 2691.945 ;
        RECT 1099.710 2691.630 1113.135 2691.930 ;
        RECT 1112.805 2691.615 1113.135 2691.630 ;
        RECT 1488.165 2691.930 1488.495 2691.945 ;
        RECT 1499.910 2691.930 1504.000 2692.120 ;
        RECT 1488.165 2691.800 1504.000 2691.930 ;
        RECT 1488.165 2691.630 1500.210 2691.800 ;
        RECT 1488.165 2691.615 1488.495 2691.630 ;
      LAYER met3 ;
        RECT 1504.400 2691.440 1885.335 2692.800 ;
        RECT 1504.400 2691.400 1884.935 2691.440 ;
        RECT 1504.000 2690.040 1884.935 2691.400 ;
      LAYER met3 ;
        RECT 1885.335 2690.760 1889.335 2691.040 ;
        RECT 1885.335 2690.440 1889.370 2690.760 ;
      LAYER met3 ;
        RECT 1504.000 2677.840 1885.335 2690.040 ;
      LAYER met3 ;
        RECT 1889.070 2687.850 1889.370 2690.440 ;
        RECT 1898.485 2687.850 1898.815 2687.865 ;
        RECT 1889.070 2687.550 1898.815 2687.850 ;
        RECT 1898.485 2687.535 1898.815 2687.550 ;
        RECT 1500.000 2677.160 1504.000 2677.440 ;
        RECT 1499.910 2676.840 1504.000 2677.160 ;
        RECT 1488.165 2674.250 1488.495 2674.265 ;
        RECT 1499.910 2674.250 1500.210 2676.840 ;
      LAYER met3 ;
        RECT 1504.400 2676.480 1885.335 2677.840 ;
        RECT 1504.400 2676.440 1884.935 2676.480 ;
      LAYER met3 ;
        RECT 1488.165 2673.950 1500.210 2674.250 ;
      LAYER met3 ;
        RECT 1504.000 2675.080 1884.935 2676.440 ;
      LAYER met3 ;
        RECT 1885.335 2675.800 1889.335 2676.080 ;
        RECT 1885.335 2675.480 1889.370 2675.800 ;
        RECT 1488.165 2673.935 1488.495 2673.950 ;
        RECT 1000.000 2672.120 1004.000 2672.720 ;
        RECT 993.665 2670.850 993.995 2670.865 ;
        RECT 1000.350 2670.850 1000.650 2672.120 ;
      LAYER met3 ;
        RECT 1004.400 2671.720 1096.000 2673.120 ;
      LAYER met3 ;
        RECT 993.665 2670.550 1000.650 2670.850 ;
        RECT 993.665 2670.535 993.995 2670.550 ;
      LAYER met3 ;
        RECT 1004.000 2670.400 1096.000 2671.720 ;
        RECT 434.000 2669.040 574.400 2670.400 ;
      LAYER met3 ;
        RECT 574.800 2669.400 578.800 2670.000 ;
      LAYER met3 ;
        RECT 434.400 2669.000 574.400 2669.040 ;
        RECT 434.400 2667.640 574.800 2669.000 ;
        RECT 434.000 2648.640 574.800 2667.640 ;
      LAYER met3 ;
        RECT 578.070 2666.770 578.370 2669.400 ;
      LAYER met3 ;
        RECT 1004.000 2669.000 1095.600 2670.400 ;
      LAYER met3 ;
        RECT 1096.000 2669.680 1100.000 2670.000 ;
        RECT 1096.000 2669.400 1100.010 2669.680 ;
        RECT 588.865 2666.770 589.195 2666.785 ;
        RECT 578.070 2666.470 589.195 2666.770 ;
        RECT 588.865 2666.455 589.195 2666.470 ;
      LAYER met3 ;
        RECT 1004.000 2650.000 1096.000 2669.000 ;
      LAYER met3 ;
        RECT 1099.710 2666.770 1100.010 2669.400 ;
        RECT 1113.265 2666.770 1113.595 2666.785 ;
        RECT 1099.710 2666.470 1113.595 2666.770 ;
        RECT 1113.265 2666.455 1113.595 2666.470 ;
      LAYER met3 ;
        RECT 1504.000 2661.520 1885.335 2675.080 ;
      LAYER met3 ;
        RECT 1889.070 2672.890 1889.370 2675.480 ;
        RECT 1898.945 2672.890 1899.275 2672.905 ;
        RECT 1889.070 2672.590 1899.275 2672.890 ;
        RECT 1898.945 2672.575 1899.275 2672.590 ;
        RECT 1500.000 2660.840 1504.000 2661.120 ;
        RECT 1499.910 2660.520 1504.000 2660.840 ;
        RECT 1482.645 2657.930 1482.975 2657.945 ;
        RECT 1499.910 2657.930 1500.210 2660.520 ;
      LAYER met3 ;
        RECT 1504.400 2660.160 1885.335 2661.520 ;
        RECT 1504.400 2660.120 1884.935 2660.160 ;
      LAYER met3 ;
        RECT 1482.645 2657.630 1500.210 2657.930 ;
      LAYER met3 ;
        RECT 1504.000 2658.760 1884.935 2660.120 ;
      LAYER met3 ;
        RECT 1885.335 2659.480 1889.335 2659.760 ;
        RECT 1885.335 2659.160 1889.370 2659.480 ;
        RECT 1482.645 2657.615 1482.975 2657.630 ;
        RECT 1000.000 2649.000 1004.000 2649.600 ;
      LAYER met3 ;
        RECT 434.000 2647.280 574.400 2648.640 ;
        RECT 434.400 2647.240 574.400 2647.280 ;
        RECT 434.400 2645.880 574.800 2647.240 ;
      LAYER met3 ;
        RECT 994.125 2646.370 994.455 2646.385 ;
        RECT 1000.350 2646.370 1000.650 2649.000 ;
      LAYER met3 ;
        RECT 1004.400 2648.600 1096.000 2650.000 ;
      LAYER met3 ;
        RECT 994.125 2646.070 1000.650 2646.370 ;
      LAYER met3 ;
        RECT 1004.000 2647.280 1096.000 2648.600 ;
      LAYER met3 ;
        RECT 994.125 2646.055 994.455 2646.070 ;
      LAYER met3 ;
        RECT 434.000 2626.880 574.800 2645.880 ;
        RECT 1004.000 2645.880 1095.600 2647.280 ;
      LAYER met3 ;
        RECT 1096.000 2646.280 1100.000 2646.880 ;
      LAYER met3 ;
        RECT 1504.000 2646.560 1885.335 2658.760 ;
      LAYER met3 ;
        RECT 1889.070 2657.250 1889.370 2659.160 ;
        RECT 1899.405 2657.250 1899.735 2657.265 ;
        RECT 1889.070 2656.950 1899.735 2657.250 ;
        RECT 1899.405 2656.935 1899.735 2656.950 ;
      LAYER met3 ;
        RECT 1004.000 2626.880 1096.000 2645.880 ;
      LAYER met3 ;
        RECT 1096.950 2645.025 1097.250 2646.280 ;
      LAYER met3 ;
        RECT 1504.400 2645.200 1885.335 2646.560 ;
        RECT 1504.400 2645.160 1884.935 2645.200 ;
      LAYER met3 ;
        RECT 1096.950 2644.710 1097.495 2645.025 ;
        RECT 1097.165 2644.695 1097.495 2644.710 ;
      LAYER met3 ;
        RECT 1504.000 2643.800 1884.935 2645.160 ;
        RECT 1504.000 2630.240 1885.335 2643.800 ;
      LAYER met3 ;
        RECT 1500.000 2629.560 1504.000 2629.840 ;
        RECT 1487.245 2629.370 1487.575 2629.385 ;
        RECT 1499.910 2629.370 1504.000 2629.560 ;
        RECT 1487.245 2629.240 1504.000 2629.370 ;
        RECT 1487.245 2629.070 1500.210 2629.240 ;
        RECT 1487.245 2629.055 1487.575 2629.070 ;
      LAYER met3 ;
        RECT 1504.400 2628.880 1885.335 2630.240 ;
        RECT 1504.400 2628.840 1884.935 2628.880 ;
        RECT 434.000 2625.520 574.400 2626.880 ;
      LAYER met3 ;
        RECT 1000.000 2625.880 1004.000 2626.480 ;
      LAYER met3 ;
        RECT 434.400 2625.480 574.400 2625.520 ;
        RECT 434.400 2624.120 574.800 2625.480 ;
        RECT 434.000 2606.480 574.800 2624.120 ;
      LAYER met3 ;
        RECT 991.365 2623.250 991.695 2623.265 ;
        RECT 1000.350 2623.250 1000.650 2625.880 ;
      LAYER met3 ;
        RECT 1004.400 2625.480 1096.000 2626.880 ;
      LAYER met3 ;
        RECT 991.365 2622.950 1000.650 2623.250 ;
      LAYER met3 ;
        RECT 1004.000 2624.160 1096.000 2625.480 ;
        RECT 1504.000 2627.480 1884.935 2628.840 ;
      LAYER met3 ;
        RECT 1885.335 2628.200 1889.335 2628.480 ;
        RECT 1885.335 2627.880 1889.370 2628.200 ;
        RECT 991.365 2622.935 991.695 2622.950 ;
      LAYER met3 ;
        RECT 1004.000 2622.760 1095.600 2624.160 ;
      LAYER met3 ;
        RECT 1096.000 2623.160 1100.000 2623.760 ;
      LAYER met3 ;
        RECT 1004.000 2610.715 1096.000 2622.760 ;
      LAYER met3 ;
        RECT 1097.870 2622.585 1098.170 2623.160 ;
        RECT 1097.625 2622.270 1098.170 2622.585 ;
        RECT 1097.625 2622.255 1097.955 2622.270 ;
      LAYER met3 ;
        RECT 1504.000 2613.920 1885.335 2627.480 ;
      LAYER met3 ;
        RECT 1889.070 2625.290 1889.370 2627.880 ;
        RECT 1899.865 2625.290 1900.195 2625.305 ;
        RECT 1889.070 2624.990 1900.195 2625.290 ;
        RECT 1899.865 2624.975 1900.195 2624.990 ;
        RECT 1500.000 2613.240 1504.000 2613.520 ;
        RECT 1499.910 2612.920 1504.000 2613.240 ;
        RECT 1487.705 2610.330 1488.035 2610.345 ;
        RECT 1499.910 2610.330 1500.210 2612.920 ;
      LAYER met3 ;
        RECT 1504.400 2612.560 1885.335 2613.920 ;
        RECT 1504.400 2612.520 1884.935 2612.560 ;
      LAYER met3 ;
        RECT 1487.705 2610.030 1500.210 2610.330 ;
      LAYER met3 ;
        RECT 1504.000 2611.160 1884.935 2612.520 ;
      LAYER met3 ;
        RECT 1885.335 2611.880 1889.335 2612.160 ;
        RECT 1885.335 2611.560 1889.370 2611.880 ;
        RECT 1487.705 2610.015 1488.035 2610.030 ;
        RECT 1406.285 2609.650 1406.615 2609.665 ;
        RECT 1406.070 2609.335 1406.615 2609.650 ;
        RECT 1406.070 2608.460 1406.370 2609.335 ;
        RECT 1406.745 2608.460 1407.075 2608.475 ;
        RECT 1406.070 2608.160 1407.075 2608.460 ;
        RECT 1406.745 2608.145 1407.075 2608.160 ;
      LAYER met3 ;
        RECT 434.000 2605.615 574.400 2606.480 ;
        RECT 1504.000 2598.960 1885.335 2611.160 ;
      LAYER met3 ;
        RECT 1889.070 2608.970 1889.370 2611.560 ;
      LAYER met3 ;
        RECT 2427.190 2610.715 2529.990 2760.645 ;
      LAYER met3 ;
        RECT 1892.505 2608.970 1892.835 2608.985 ;
        RECT 1889.070 2608.670 1892.835 2608.970 ;
        RECT 1892.505 2608.655 1892.835 2608.670 ;
        RECT 1500.000 2598.280 1504.000 2598.560 ;
        RECT 1499.910 2597.960 1504.000 2598.280 ;
        RECT 1487.245 2595.370 1487.575 2595.385 ;
        RECT 1499.910 2595.370 1500.210 2597.960 ;
      LAYER met3 ;
        RECT 1504.400 2597.600 1885.335 2598.960 ;
        RECT 1504.400 2597.560 1884.935 2597.600 ;
      LAYER met3 ;
        RECT 1487.245 2595.070 1500.210 2595.370 ;
      LAYER met3 ;
        RECT 1504.000 2596.200 1884.935 2597.560 ;
      LAYER met3 ;
        RECT 1487.245 2595.055 1487.575 2595.070 ;
      LAYER met3 ;
        RECT 1504.000 2582.640 1885.335 2596.200 ;
      LAYER met3 ;
        RECT 1500.000 2581.960 1504.000 2582.240 ;
        RECT 1499.910 2581.640 1504.000 2581.960 ;
        RECT 1487.245 2581.090 1487.575 2581.105 ;
        RECT 1499.910 2581.090 1500.210 2581.640 ;
      LAYER met3 ;
        RECT 1504.400 2581.280 1885.335 2582.640 ;
        RECT 1504.400 2581.240 1884.935 2581.280 ;
      LAYER met3 ;
        RECT 1487.245 2580.790 1500.210 2581.090 ;
        RECT 1487.245 2580.775 1487.575 2580.790 ;
      LAYER met3 ;
        RECT 1504.000 2579.880 1884.935 2581.240 ;
      LAYER met3 ;
        RECT 1885.335 2580.600 1889.335 2580.880 ;
        RECT 1885.335 2580.280 1889.370 2580.600 ;
      LAYER met3 ;
        RECT 1504.000 2567.680 1885.335 2579.880 ;
      LAYER met3 ;
        RECT 1889.070 2577.690 1889.370 2580.280 ;
        RECT 1900.325 2577.690 1900.655 2577.705 ;
        RECT 1889.070 2577.390 1900.655 2577.690 ;
        RECT 1900.325 2577.375 1900.655 2577.390 ;
        RECT 1487.245 2567.490 1487.575 2567.505 ;
        RECT 1487.245 2567.280 1500.210 2567.490 ;
        RECT 1487.245 2567.190 1504.000 2567.280 ;
        RECT 1487.245 2567.175 1487.575 2567.190 ;
        RECT 1499.910 2567.000 1504.000 2567.190 ;
        RECT 1500.000 2566.680 1504.000 2567.000 ;
      LAYER met3 ;
        RECT 1504.400 2566.320 1885.335 2567.680 ;
        RECT 1504.400 2566.280 1884.935 2566.320 ;
        RECT 1504.000 2564.920 1884.935 2566.280 ;
      LAYER met3 ;
        RECT 1885.335 2565.640 1889.335 2565.920 ;
        RECT 1885.335 2565.320 1889.370 2565.640 ;
      LAYER met3 ;
        RECT 1504.000 2551.360 1885.335 2564.920 ;
      LAYER met3 ;
        RECT 1889.070 2562.730 1889.370 2565.320 ;
        RECT 1900.785 2562.730 1901.115 2562.745 ;
        RECT 1889.070 2562.430 1901.115 2562.730 ;
        RECT 1900.785 2562.415 1901.115 2562.430 ;
        RECT 1500.000 2550.680 1504.000 2550.960 ;
        RECT 1499.910 2550.360 1504.000 2550.680 ;
        RECT 1483.565 2547.770 1483.895 2547.785 ;
        RECT 1499.910 2547.770 1500.210 2550.360 ;
      LAYER met3 ;
        RECT 1504.400 2550.000 1885.335 2551.360 ;
        RECT 1504.400 2549.960 1884.935 2550.000 ;
      LAYER met3 ;
        RECT 1483.565 2547.470 1500.210 2547.770 ;
      LAYER met3 ;
        RECT 1504.000 2548.600 1884.935 2549.960 ;
      LAYER met3 ;
        RECT 1885.335 2549.320 1889.335 2549.600 ;
        RECT 1885.335 2549.000 1889.370 2549.320 ;
        RECT 1483.565 2547.455 1483.895 2547.470 ;
      LAYER met3 ;
        RECT 1504.000 2536.400 1885.335 2548.600 ;
      LAYER met3 ;
        RECT 1889.070 2547.770 1889.370 2549.000 ;
        RECT 1901.245 2547.770 1901.575 2547.785 ;
        RECT 1889.070 2547.470 1901.575 2547.770 ;
        RECT 1901.245 2547.455 1901.575 2547.470 ;
      LAYER met3 ;
        RECT 1504.400 2535.040 1885.335 2536.400 ;
        RECT 1504.400 2535.000 1884.935 2535.040 ;
        RECT 1504.000 2533.640 1884.935 2535.000 ;
        RECT 1504.000 2520.080 1885.335 2533.640 ;
      LAYER met3 ;
        RECT 1500.000 2519.400 1504.000 2519.680 ;
        RECT 1486.785 2519.210 1487.115 2519.225 ;
        RECT 1499.910 2519.210 1504.000 2519.400 ;
        RECT 1486.785 2519.080 1504.000 2519.210 ;
        RECT 1486.785 2518.910 1500.210 2519.080 ;
        RECT 1486.785 2518.895 1487.115 2518.910 ;
      LAYER met3 ;
        RECT 1504.400 2518.720 1885.335 2520.080 ;
        RECT 1504.400 2518.680 1884.935 2518.720 ;
        RECT 1504.000 2517.320 1884.935 2518.680 ;
      LAYER met3 ;
        RECT 1885.335 2518.040 1889.335 2518.320 ;
        RECT 1885.335 2517.720 1889.370 2518.040 ;
        RECT 1357.985 2511.740 1358.315 2511.745 ;
        RECT 1357.985 2511.730 1358.570 2511.740 ;
        RECT 1357.985 2511.430 1358.770 2511.730 ;
        RECT 1357.985 2511.420 1358.570 2511.430 ;
        RECT 1357.985 2511.415 1358.315 2511.420 ;
      LAYER met3 ;
        RECT 1504.000 2504.255 1885.335 2517.320 ;
      LAYER met3 ;
        RECT 1889.070 2515.130 1889.370 2517.720 ;
        RECT 1903.545 2515.130 1903.875 2515.145 ;
        RECT 1889.070 2514.830 1903.875 2515.130 ;
        RECT 1903.545 2514.815 1903.875 2514.830 ;
        RECT 1358.190 2463.450 1358.570 2463.460 ;
        RECT 1358.905 2463.450 1359.235 2463.465 ;
        RECT 1358.190 2463.150 1359.235 2463.450 ;
        RECT 1358.190 2463.140 1358.570 2463.150 ;
        RECT 1358.905 2463.135 1359.235 2463.150 ;
        RECT 1405.365 2463.450 1405.695 2463.465 ;
        RECT 1406.285 2463.450 1406.615 2463.465 ;
        RECT 1405.365 2463.150 1406.615 2463.450 ;
        RECT 1405.365 2463.135 1405.695 2463.150 ;
        RECT 1406.285 2463.135 1406.615 2463.150 ;
        RECT 1535.085 2415.850 1535.415 2415.865 ;
        RECT 1535.085 2415.550 1536.090 2415.850 ;
        RECT 1535.085 2415.535 1535.415 2415.550 ;
        RECT 1535.085 2415.170 1535.415 2415.185 ;
        RECT 1535.790 2415.170 1536.090 2415.550 ;
        RECT 1535.085 2414.870 1536.090 2415.170 ;
        RECT 1535.085 2414.855 1535.415 2414.870 ;
        RECT 1535.085 2319.290 1535.415 2319.305 ;
        RECT 1535.085 2318.990 1536.090 2319.290 ;
        RECT 1535.085 2318.975 1535.415 2318.990 ;
        RECT 1535.085 2318.610 1535.415 2318.625 ;
        RECT 1535.790 2318.610 1536.090 2318.990 ;
        RECT 1535.085 2318.310 1536.090 2318.610 ;
        RECT 1535.085 2318.295 1535.415 2318.310 ;
        RECT 1405.365 2270.330 1405.695 2270.345 ;
        RECT 1406.285 2270.330 1406.615 2270.345 ;
        RECT 1405.365 2270.030 1406.615 2270.330 ;
        RECT 1405.365 2270.015 1405.695 2270.030 ;
        RECT 1406.285 2270.015 1406.615 2270.030 ;
        RECT 1534.165 2270.330 1534.495 2270.345 ;
        RECT 1535.085 2270.330 1535.415 2270.345 ;
        RECT 1534.165 2270.030 1535.415 2270.330 ;
        RECT 1534.165 2270.015 1534.495 2270.030 ;
        RECT 1535.085 2270.015 1535.415 2270.030 ;
        RECT 1405.365 2173.770 1405.695 2173.785 ;
        RECT 1406.285 2173.770 1406.615 2173.785 ;
        RECT 1405.365 2173.470 1406.615 2173.770 ;
        RECT 1405.365 2173.455 1405.695 2173.470 ;
        RECT 1406.285 2173.455 1406.615 2173.470 ;
        RECT 1358.905 2097.610 1359.235 2097.625 ;
        RECT 1359.825 2097.610 1360.155 2097.625 ;
        RECT 1358.905 2097.310 1360.155 2097.610 ;
        RECT 1358.905 2097.295 1359.235 2097.310 ;
        RECT 1359.825 2097.295 1360.155 2097.310 ;
      LAYER met3 ;
        RECT 1004.000 2019.280 1329.390 2032.005 ;
      LAYER met3 ;
        RECT 995.045 2018.730 995.375 2018.745 ;
        RECT 1000.000 2018.730 1004.000 2018.880 ;
        RECT 995.045 2018.430 1004.000 2018.730 ;
        RECT 995.045 2018.415 995.375 2018.430 ;
        RECT 1000.000 2018.280 1004.000 2018.430 ;
      LAYER met3 ;
        RECT 1004.400 2017.880 1328.990 2019.280 ;
      LAYER met3 ;
        RECT 1329.390 2018.730 1333.390 2018.880 ;
        RECT 1338.665 2018.730 1338.995 2018.745 ;
        RECT 1329.390 2018.430 1338.995 2018.730 ;
        RECT 1329.390 2018.280 1333.390 2018.430 ;
        RECT 1338.665 2018.415 1338.995 2018.430 ;
      LAYER met3 ;
        RECT 1004.000 1998.880 1329.390 2017.880 ;
      LAYER met3 ;
        RECT 990.905 1998.330 991.235 1998.345 ;
        RECT 1000.000 1998.330 1004.000 1998.480 ;
        RECT 990.905 1998.030 1004.000 1998.330 ;
        RECT 990.905 1998.015 991.235 1998.030 ;
        RECT 1000.000 1997.880 1004.000 1998.030 ;
      LAYER met3 ;
        RECT 1004.400 1997.480 1328.990 1998.880 ;
      LAYER met3 ;
        RECT 1329.390 1998.330 1333.390 1998.480 ;
        RECT 1334.065 1998.330 1334.395 1998.345 ;
        RECT 1329.390 1998.030 1334.395 1998.330 ;
        RECT 1329.390 1997.880 1333.390 1998.030 ;
        RECT 1334.065 1998.015 1334.395 1998.030 ;
      LAYER met3 ;
        RECT 1004.000 1977.120 1329.390 1997.480 ;
      LAYER met3 ;
        RECT 1408.125 1980.650 1408.455 1980.665 ;
        RECT 1406.990 1980.350 1408.455 1980.650 ;
        RECT 1406.990 1979.970 1407.290 1980.350 ;
        RECT 1408.125 1980.335 1408.455 1980.350 ;
        RECT 1408.125 1979.970 1408.455 1979.985 ;
        RECT 1406.990 1979.670 1408.455 1979.970 ;
        RECT 1408.125 1979.655 1408.455 1979.670 ;
        RECT 995.505 1976.570 995.835 1976.585 ;
        RECT 1000.000 1976.570 1004.000 1976.720 ;
        RECT 995.505 1976.270 1004.000 1976.570 ;
        RECT 995.505 1976.255 995.835 1976.270 ;
        RECT 1000.000 1976.120 1004.000 1976.270 ;
      LAYER met3 ;
        RECT 1004.400 1975.720 1328.990 1977.120 ;
      LAYER met3 ;
        RECT 1329.390 1976.570 1333.390 1976.720 ;
        RECT 1339.125 1976.570 1339.455 1976.585 ;
        RECT 1329.390 1976.270 1339.455 1976.570 ;
        RECT 1329.390 1976.120 1333.390 1976.270 ;
        RECT 1339.125 1976.255 1339.455 1976.270 ;
      LAYER met3 ;
        RECT 364.000 1963.520 627.030 1969.445 ;
        RECT 364.400 1962.120 627.030 1963.520 ;
        RECT 364.000 1940.400 627.030 1962.120 ;
        RECT 1004.000 1956.720 1329.390 1975.720 ;
      LAYER met3 ;
        RECT 990.445 1956.170 990.775 1956.185 ;
        RECT 1000.000 1956.170 1004.000 1956.320 ;
        RECT 990.445 1955.870 1004.000 1956.170 ;
        RECT 990.445 1955.855 990.775 1955.870 ;
        RECT 1000.000 1955.720 1004.000 1955.870 ;
      LAYER met3 ;
        RECT 1004.400 1955.320 1328.990 1956.720 ;
      LAYER met3 ;
        RECT 1329.390 1956.170 1333.390 1956.320 ;
        RECT 1339.585 1956.170 1339.915 1956.185 ;
        RECT 1329.390 1955.870 1339.915 1956.170 ;
        RECT 1329.390 1955.720 1333.390 1955.870 ;
        RECT 1339.585 1955.855 1339.915 1955.870 ;
      LAYER met3 ;
        RECT 364.000 1939.000 626.630 1940.400 ;
        RECT 364.000 1926.800 627.030 1939.000 ;
        RECT 1004.000 1936.320 1329.390 1955.320 ;
      LAYER met3 ;
        RECT 1357.985 1945.970 1358.315 1945.985 ;
        RECT 1358.905 1945.970 1359.235 1945.985 ;
        RECT 1357.985 1945.670 1359.235 1945.970 ;
        RECT 1357.985 1945.655 1358.315 1945.670 ;
        RECT 1358.905 1945.655 1359.235 1945.670 ;
        RECT 989.985 1935.770 990.315 1935.785 ;
        RECT 1000.000 1935.770 1004.000 1935.920 ;
        RECT 989.985 1935.470 1004.000 1935.770 ;
        RECT 989.985 1935.455 990.315 1935.470 ;
        RECT 1000.000 1935.320 1004.000 1935.470 ;
      LAYER met3 ;
        RECT 1004.400 1934.960 1329.390 1936.320 ;
        RECT 1004.400 1934.920 1328.990 1934.960 ;
        RECT 364.400 1925.400 627.030 1926.800 ;
        RECT 364.000 1903.680 627.030 1925.400 ;
        RECT 1004.000 1933.560 1328.990 1934.920 ;
      LAYER met3 ;
        RECT 1329.390 1934.410 1333.390 1934.560 ;
        RECT 1340.045 1934.410 1340.375 1934.425 ;
        RECT 1329.390 1934.110 1340.375 1934.410 ;
        RECT 1329.390 1933.960 1333.390 1934.110 ;
        RECT 1340.045 1934.095 1340.375 1934.110 ;
      LAYER met3 ;
        RECT 1004.000 1914.560 1329.390 1933.560 ;
      LAYER met3 ;
        RECT 995.965 1914.010 996.295 1914.025 ;
        RECT 1000.000 1914.010 1004.000 1914.160 ;
        RECT 995.965 1913.710 1004.000 1914.010 ;
        RECT 995.965 1913.695 996.295 1913.710 ;
        RECT 1000.000 1913.560 1004.000 1913.710 ;
      LAYER met3 ;
        RECT 1004.400 1913.160 1328.990 1914.560 ;
      LAYER met3 ;
        RECT 1329.390 1914.010 1333.390 1914.160 ;
        RECT 1334.525 1914.010 1334.855 1914.025 ;
        RECT 1329.390 1913.710 1334.855 1914.010 ;
        RECT 1329.390 1913.560 1333.390 1913.710 ;
        RECT 1334.525 1913.695 1334.855 1913.710 ;
      LAYER met3 ;
        RECT 364.000 1902.280 626.630 1903.680 ;
        RECT 364.000 1890.080 627.030 1902.280 ;
        RECT 1004.000 1894.160 1329.390 1913.160 ;
        RECT 1924.400 1906.040 2072.375 1906.905 ;
      LAYER met3 ;
        RECT 989.525 1893.610 989.855 1893.625 ;
        RECT 1000.000 1893.610 1004.000 1893.760 ;
        RECT 989.525 1893.310 1004.000 1893.610 ;
        RECT 989.525 1893.295 989.855 1893.310 ;
        RECT 1000.000 1893.160 1004.000 1893.310 ;
      LAYER met3 ;
        RECT 1004.400 1892.800 1329.390 1894.160 ;
        RECT 1924.000 1904.720 2072.375 1906.040 ;
        RECT 1924.000 1903.320 2071.975 1904.720 ;
        RECT 1004.400 1892.760 1328.990 1892.800 ;
        RECT 364.400 1888.680 627.030 1890.080 ;
        RECT 364.000 1866.960 627.030 1888.680 ;
        RECT 1004.000 1891.400 1328.990 1892.760 ;
      LAYER met3 ;
        RECT 1329.390 1892.250 1333.390 1892.400 ;
        RECT 1340.505 1892.250 1340.835 1892.265 ;
        RECT 1329.390 1891.950 1340.835 1892.250 ;
        RECT 1329.390 1891.800 1333.390 1891.950 ;
        RECT 1340.505 1891.935 1340.835 1891.950 ;
      LAYER met3 ;
        RECT 1004.000 1872.400 1329.390 1891.400 ;
        RECT 1924.000 1889.760 2072.375 1903.320 ;
      LAYER met3 ;
        RECT 1920.000 1888.760 1924.000 1889.360 ;
        RECT 1904.465 1886.130 1904.795 1886.145 ;
        RECT 1920.350 1886.130 1920.650 1888.760 ;
      LAYER met3 ;
        RECT 1924.400 1888.400 2072.375 1889.760 ;
        RECT 2304.000 1891.440 2523.025 1925.925 ;
      LAYER met3 ;
        RECT 2523.625 1892.250 2523.955 1892.265 ;
        RECT 2523.625 1891.935 2524.170 1892.250 ;
      LAYER met3 ;
        RECT 2304.000 1890.040 2522.625 1891.440 ;
      LAYER met3 ;
        RECT 2523.870 1891.040 2524.170 1891.935 ;
        RECT 2523.025 1890.440 2527.025 1891.040 ;
      LAYER met3 ;
        RECT 1924.400 1888.360 2071.975 1888.400 ;
      LAYER met3 ;
        RECT 1904.465 1885.830 1920.650 1886.130 ;
      LAYER met3 ;
        RECT 1924.000 1887.000 2071.975 1888.360 ;
      LAYER met3 ;
        RECT 2072.375 1887.400 2076.375 1888.000 ;
        RECT 1904.465 1885.815 1904.795 1885.830 ;
      LAYER met3 ;
        RECT 1924.000 1873.440 2072.375 1887.000 ;
      LAYER met3 ;
        RECT 2075.830 1884.770 2076.130 1887.400 ;
        RECT 2087.085 1884.770 2087.415 1884.785 ;
        RECT 2075.830 1884.470 2087.415 1884.770 ;
        RECT 2087.085 1884.455 2087.415 1884.470 ;
      LAYER met3 ;
        RECT 2304.000 1876.480 2523.025 1890.040 ;
      LAYER met3 ;
        RECT 2283.965 1875.930 2284.295 1875.945 ;
        RECT 2300.000 1875.930 2304.000 1876.080 ;
        RECT 2283.965 1875.630 2304.000 1875.930 ;
        RECT 2283.965 1875.615 2284.295 1875.630 ;
        RECT 2300.000 1875.480 2304.000 1875.630 ;
      LAYER met3 ;
        RECT 2304.400 1875.080 2523.025 1876.480 ;
      LAYER met3 ;
        RECT 1920.000 1872.440 1924.000 1873.040 ;
        RECT 996.425 1871.850 996.755 1871.865 ;
        RECT 1000.000 1871.850 1004.000 1872.000 ;
        RECT 996.425 1871.550 1004.000 1871.850 ;
        RECT 996.425 1871.535 996.755 1871.550 ;
        RECT 1000.000 1871.400 1004.000 1871.550 ;
      LAYER met3 ;
        RECT 1004.400 1871.000 1328.990 1872.400 ;
      LAYER met3 ;
        RECT 1329.390 1871.850 1333.390 1872.000 ;
        RECT 1340.965 1871.850 1341.295 1871.865 ;
        RECT 1329.390 1871.550 1341.295 1871.850 ;
        RECT 1329.390 1871.400 1333.390 1871.550 ;
        RECT 1340.965 1871.535 1341.295 1871.550 ;
      LAYER met3 ;
        RECT 364.000 1865.560 626.630 1866.960 ;
        RECT 364.000 1852.000 627.030 1865.560 ;
        RECT 1004.000 1852.000 1329.390 1871.000 ;
      LAYER met3 ;
        RECT 1904.465 1870.490 1904.795 1870.505 ;
        RECT 1920.350 1870.490 1920.650 1872.440 ;
      LAYER met3 ;
        RECT 1924.400 1872.040 2072.375 1873.440 ;
      LAYER met3 ;
        RECT 1904.465 1870.190 1920.650 1870.490 ;
      LAYER met3 ;
        RECT 1924.000 1870.720 2072.375 1872.040 ;
      LAYER met3 ;
        RECT 1904.465 1870.175 1904.795 1870.190 ;
      LAYER met3 ;
        RECT 1924.000 1869.320 2071.975 1870.720 ;
        RECT 1924.000 1855.760 2072.375 1869.320 ;
      LAYER met3 ;
        RECT 1920.000 1854.760 1924.000 1855.360 ;
      LAYER met3 ;
        RECT 364.400 1850.600 627.030 1852.000 ;
      LAYER met3 ;
        RECT 989.065 1851.450 989.395 1851.465 ;
        RECT 1000.000 1851.450 1004.000 1851.600 ;
        RECT 989.065 1851.150 1004.000 1851.450 ;
        RECT 989.065 1851.135 989.395 1851.150 ;
        RECT 1000.000 1851.000 1004.000 1851.150 ;
      LAYER met3 ;
        RECT 1004.400 1850.640 1329.390 1852.000 ;
      LAYER met3 ;
        RECT 1904.465 1852.130 1904.795 1852.145 ;
        RECT 1920.350 1852.130 1920.650 1854.760 ;
      LAYER met3 ;
        RECT 1924.400 1854.400 2072.375 1855.760 ;
        RECT 1924.400 1854.360 2071.975 1854.400 ;
      LAYER met3 ;
        RECT 1904.465 1851.830 1920.650 1852.130 ;
      LAYER met3 ;
        RECT 1924.000 1853.000 2071.975 1854.360 ;
      LAYER met3 ;
        RECT 2072.375 1853.400 2076.375 1854.000 ;
        RECT 1904.465 1851.815 1904.795 1851.830 ;
      LAYER met3 ;
        RECT 1004.400 1850.600 1328.990 1850.640 ;
        RECT 364.000 1830.240 627.030 1850.600 ;
        RECT 1004.000 1849.240 1328.990 1850.600 ;
      LAYER met3 ;
        RECT 1329.390 1850.090 1333.390 1850.240 ;
        RECT 1341.425 1850.090 1341.755 1850.105 ;
        RECT 1329.390 1849.790 1341.755 1850.090 ;
        RECT 1329.390 1849.640 1333.390 1849.790 ;
        RECT 1341.425 1849.775 1341.755 1849.790 ;
      LAYER met3 ;
        RECT 1004.000 1830.240 1329.390 1849.240 ;
        RECT 1924.000 1839.440 2072.375 1853.000 ;
      LAYER met3 ;
        RECT 2075.830 1850.770 2076.130 1853.400 ;
        RECT 2084.325 1850.770 2084.655 1850.785 ;
        RECT 2075.830 1850.470 2084.655 1850.770 ;
        RECT 2084.325 1850.455 2084.655 1850.470 ;
      LAYER met3 ;
        RECT 1924.400 1838.040 2072.375 1839.440 ;
        RECT 1924.000 1836.720 2072.375 1838.040 ;
        RECT 1924.000 1835.320 2071.975 1836.720 ;
      LAYER met3 ;
        RECT 2072.375 1835.810 2076.375 1836.320 ;
        RECT 2084.785 1835.810 2085.115 1835.825 ;
        RECT 2072.375 1835.720 2085.115 1835.810 ;
        RECT 2075.830 1835.510 2085.115 1835.720 ;
        RECT 2084.785 1835.495 2085.115 1835.510 ;
      LAYER met3 ;
        RECT 364.000 1828.840 626.630 1830.240 ;
      LAYER met3 ;
        RECT 996.885 1829.690 997.215 1829.705 ;
        RECT 1000.000 1829.690 1004.000 1829.840 ;
        RECT 996.885 1829.390 1004.000 1829.690 ;
        RECT 996.885 1829.375 997.215 1829.390 ;
        RECT 1000.000 1829.240 1004.000 1829.390 ;
      LAYER met3 ;
        RECT 1004.400 1828.840 1328.990 1830.240 ;
      LAYER met3 ;
        RECT 1329.390 1829.690 1333.390 1829.840 ;
        RECT 1341.885 1829.690 1342.215 1829.705 ;
        RECT 1329.390 1829.390 1342.215 1829.690 ;
        RECT 1329.390 1829.240 1333.390 1829.390 ;
        RECT 1341.885 1829.375 1342.215 1829.390 ;
      LAYER met3 ;
        RECT 364.000 1815.280 627.030 1828.840 ;
        RECT 364.400 1813.880 627.030 1815.280 ;
        RECT 364.000 1792.160 627.030 1813.880 ;
        RECT 1004.000 1809.840 1329.390 1828.840 ;
        RECT 1924.000 1821.760 2072.375 1835.320 ;
      LAYER met3 ;
        RECT 1920.000 1820.760 1924.000 1821.360 ;
        RECT 1904.465 1818.130 1904.795 1818.145 ;
        RECT 1920.350 1818.130 1920.650 1820.760 ;
      LAYER met3 ;
        RECT 1924.400 1820.400 2072.375 1821.760 ;
        RECT 1924.400 1820.360 2071.975 1820.400 ;
      LAYER met3 ;
        RECT 1904.465 1817.830 1920.650 1818.130 ;
      LAYER met3 ;
        RECT 1924.000 1819.000 2071.975 1820.360 ;
      LAYER met3 ;
        RECT 2072.375 1819.400 2076.375 1820.000 ;
        RECT 1904.465 1817.815 1904.795 1817.830 ;
        RECT 988.605 1809.290 988.935 1809.305 ;
        RECT 1000.000 1809.290 1004.000 1809.440 ;
        RECT 988.605 1808.990 1004.000 1809.290 ;
        RECT 988.605 1808.975 988.935 1808.990 ;
        RECT 1000.000 1808.840 1004.000 1808.990 ;
      LAYER met3 ;
        RECT 1004.400 1808.480 1329.390 1809.840 ;
        RECT 1004.400 1808.440 1328.990 1808.480 ;
        RECT 1004.000 1807.080 1328.990 1808.440 ;
      LAYER met3 ;
        RECT 1329.390 1807.930 1333.390 1808.080 ;
        RECT 1342.345 1807.930 1342.675 1807.945 ;
        RECT 1329.390 1807.630 1342.675 1807.930 ;
        RECT 1329.390 1807.480 1333.390 1807.630 ;
        RECT 1342.345 1807.615 1342.675 1807.630 ;
      LAYER met3 ;
        RECT 364.000 1790.760 626.630 1792.160 ;
        RECT 364.000 1778.560 627.030 1790.760 ;
        RECT 1004.000 1788.080 1329.390 1807.080 ;
        RECT 1924.000 1805.440 2072.375 1819.000 ;
      LAYER met3 ;
        RECT 2075.830 1816.770 2076.130 1819.400 ;
        RECT 2085.245 1816.770 2085.575 1816.785 ;
        RECT 2075.830 1816.470 2085.575 1816.770 ;
        RECT 2085.245 1816.455 2085.575 1816.470 ;
      LAYER met3 ;
        RECT 1924.400 1804.040 2072.375 1805.440 ;
        RECT 1924.000 1802.720 2072.375 1804.040 ;
        RECT 2304.000 1805.760 2523.025 1875.080 ;
        RECT 2304.000 1804.360 2522.625 1805.760 ;
      LAYER met3 ;
        RECT 2523.025 1804.760 2527.025 1805.360 ;
      LAYER met3 ;
        RECT 1924.000 1801.320 2071.975 1802.720 ;
      LAYER met3 ;
        RECT 2072.375 1801.720 2076.375 1802.320 ;
        RECT 988.145 1787.530 988.475 1787.545 ;
        RECT 1000.000 1787.530 1004.000 1787.680 ;
        RECT 988.145 1787.230 1004.000 1787.530 ;
        RECT 988.145 1787.215 988.475 1787.230 ;
        RECT 1000.000 1787.080 1004.000 1787.230 ;
      LAYER met3 ;
        RECT 1004.400 1786.680 1328.990 1788.080 ;
        RECT 1924.000 1787.760 2072.375 1801.320 ;
      LAYER met3 ;
        RECT 2075.830 1801.130 2076.130 1801.720 ;
        RECT 2085.705 1801.130 2086.035 1801.145 ;
        RECT 2075.830 1800.830 2086.035 1801.130 ;
        RECT 2085.705 1800.815 2086.035 1800.830 ;
      LAYER met3 ;
        RECT 2304.000 1790.800 2523.025 1804.360 ;
      LAYER met3 ;
        RECT 2523.870 1802.505 2524.170 1804.760 ;
        RECT 2523.625 1802.190 2524.170 1802.505 ;
        RECT 2523.625 1802.175 2523.955 1802.190 ;
        RECT 2287.185 1790.250 2287.515 1790.265 ;
        RECT 2300.000 1790.250 2304.000 1790.400 ;
        RECT 2287.185 1789.950 2304.000 1790.250 ;
        RECT 2287.185 1789.935 2287.515 1789.950 ;
        RECT 2300.000 1789.800 2304.000 1789.950 ;
      LAYER met3 ;
        RECT 2304.400 1789.400 2523.025 1790.800 ;
      LAYER met3 ;
        RECT 1329.390 1787.530 1333.390 1787.680 ;
        RECT 1335.445 1787.530 1335.775 1787.545 ;
        RECT 1329.390 1787.230 1335.775 1787.530 ;
        RECT 1329.390 1787.080 1333.390 1787.230 ;
        RECT 1335.445 1787.215 1335.775 1787.230 ;
      LAYER met3 ;
        RECT 364.400 1777.160 627.030 1778.560 ;
        RECT 364.000 1755.440 627.030 1777.160 ;
        RECT 1004.000 1767.680 1329.390 1786.680 ;
        RECT 1924.400 1786.400 2072.375 1787.760 ;
        RECT 1924.400 1786.360 2071.975 1786.400 ;
        RECT 1924.000 1785.000 2071.975 1786.360 ;
      LAYER met3 ;
        RECT 2072.375 1785.400 2076.375 1786.000 ;
      LAYER met3 ;
        RECT 1924.000 1771.440 2072.375 1785.000 ;
      LAYER met3 ;
        RECT 2075.830 1782.770 2076.130 1785.400 ;
        RECT 2086.165 1782.770 2086.495 1782.785 ;
        RECT 2075.830 1782.470 2086.495 1782.770 ;
        RECT 2086.165 1782.455 2086.495 1782.470 ;
        RECT 1920.000 1770.440 1924.000 1771.040 ;
        RECT 1904.465 1767.810 1904.795 1767.825 ;
        RECT 1920.350 1767.810 1920.650 1770.440 ;
      LAYER met3 ;
        RECT 1924.400 1770.040 2072.375 1771.440 ;
      LAYER met3 ;
        RECT 987.685 1767.130 988.015 1767.145 ;
        RECT 1000.000 1767.130 1004.000 1767.280 ;
        RECT 987.685 1766.830 1004.000 1767.130 ;
        RECT 987.685 1766.815 988.015 1766.830 ;
        RECT 1000.000 1766.680 1004.000 1766.830 ;
      LAYER met3 ;
        RECT 1004.400 1766.280 1328.990 1767.680 ;
      LAYER met3 ;
        RECT 1904.465 1767.510 1920.650 1767.810 ;
      LAYER met3 ;
        RECT 1924.000 1768.720 2072.375 1770.040 ;
      LAYER met3 ;
        RECT 1904.465 1767.495 1904.795 1767.510 ;
      LAYER met3 ;
        RECT 1924.000 1767.320 2071.975 1768.720 ;
      LAYER met3 ;
        RECT 2072.375 1767.720 2076.375 1768.320 ;
        RECT 1329.390 1767.130 1333.390 1767.280 ;
        RECT 1342.805 1767.130 1343.135 1767.145 ;
        RECT 1329.390 1766.830 1343.135 1767.130 ;
        RECT 1329.390 1766.680 1333.390 1766.830 ;
        RECT 1342.805 1766.815 1343.135 1766.830 ;
      LAYER met3 ;
        RECT 364.000 1754.040 626.630 1755.440 ;
        RECT 364.000 1741.840 627.030 1754.040 ;
        RECT 1004.000 1745.920 1329.390 1766.280 ;
        RECT 1924.000 1760.715 2072.375 1767.320 ;
      LAYER met3 ;
        RECT 2075.830 1767.130 2076.130 1767.720 ;
        RECT 2086.625 1767.130 2086.955 1767.145 ;
        RECT 2075.830 1766.830 2086.955 1767.130 ;
        RECT 2086.625 1766.815 2086.955 1766.830 ;
        RECT 987.225 1745.370 987.555 1745.385 ;
        RECT 1000.000 1745.370 1004.000 1745.520 ;
        RECT 987.225 1745.070 1004.000 1745.370 ;
        RECT 987.225 1745.055 987.555 1745.070 ;
        RECT 1000.000 1744.920 1004.000 1745.070 ;
      LAYER met3 ;
        RECT 1004.400 1744.520 1328.990 1745.920 ;
      LAYER met3 ;
        RECT 1329.390 1745.370 1333.390 1745.520 ;
        RECT 1335.905 1745.370 1336.235 1745.385 ;
        RECT 1329.390 1745.070 1336.235 1745.370 ;
        RECT 1329.390 1744.920 1333.390 1745.070 ;
        RECT 1335.905 1745.055 1336.235 1745.070 ;
      LAYER met3 ;
        RECT 364.400 1740.440 627.030 1741.840 ;
        RECT 364.000 1718.720 627.030 1740.440 ;
        RECT 1004.000 1725.520 1329.390 1744.520 ;
      LAYER met3 ;
        RECT 997.345 1724.970 997.675 1724.985 ;
        RECT 1000.000 1724.970 1004.000 1725.120 ;
        RECT 997.345 1724.670 1004.000 1724.970 ;
        RECT 997.345 1724.655 997.675 1724.670 ;
        RECT 1000.000 1724.520 1004.000 1724.670 ;
      LAYER met3 ;
        RECT 1004.400 1724.120 1328.990 1725.520 ;
      LAYER met3 ;
        RECT 1329.390 1724.970 1333.390 1725.120 ;
        RECT 1343.265 1724.970 1343.595 1724.985 ;
        RECT 1329.390 1724.670 1343.595 1724.970 ;
        RECT 1329.390 1724.520 1333.390 1724.670 ;
        RECT 1343.265 1724.655 1343.595 1724.670 ;
      LAYER met3 ;
        RECT 364.000 1717.320 626.630 1718.720 ;
        RECT 364.000 1710.715 627.030 1717.320 ;
        RECT 1004.000 1710.715 1329.390 1724.120 ;
        RECT 2304.000 1720.080 2523.025 1789.400 ;
        RECT 2304.000 1718.680 2522.625 1720.080 ;
      LAYER met3 ;
        RECT 2523.025 1719.080 2527.025 1719.680 ;
      LAYER met3 ;
        RECT 2304.000 1710.715 2523.025 1718.680 ;
      LAYER met3 ;
        RECT 2523.870 1718.185 2524.170 1719.080 ;
        RECT 2523.625 1717.870 2524.170 1718.185 ;
        RECT 2523.625 1717.855 2523.955 1717.870 ;
        RECT 2518.565 1704.570 2518.895 1704.585 ;
        RECT 2519.485 1704.570 2519.815 1704.585 ;
        RECT 2518.565 1704.270 2519.815 1704.570 ;
        RECT 2518.565 1704.255 2518.895 1704.270 ;
        RECT 2519.485 1704.255 2519.815 1704.270 ;
        RECT 1290.825 1635.210 1291.155 1635.225 ;
        RECT 1291.745 1635.210 1292.075 1635.225 ;
        RECT 1290.825 1634.910 1292.075 1635.210 ;
        RECT 1290.825 1634.895 1291.155 1634.910 ;
        RECT 1291.745 1634.895 1292.075 1634.910 ;
        RECT 2519.485 1608.690 2519.815 1608.705 ;
        RECT 2519.270 1608.375 2519.815 1608.690 ;
        RECT 2519.270 1607.345 2519.570 1608.375 ;
        RECT 2519.270 1607.030 2519.815 1607.345 ;
        RECT 2519.485 1607.015 2519.815 1607.030 ;
        RECT 1277.945 1546.130 1278.275 1546.145 ;
        RECT 1279.325 1546.130 1279.655 1546.145 ;
        RECT 1277.945 1545.830 1279.655 1546.130 ;
        RECT 1277.945 1545.815 1278.275 1545.830 ;
        RECT 1279.325 1545.815 1279.655 1545.830 ;
        RECT 1291.745 1546.130 1292.075 1546.145 ;
        RECT 1293.125 1546.130 1293.455 1546.145 ;
        RECT 1291.745 1545.830 1293.455 1546.130 ;
        RECT 1291.745 1545.815 1292.075 1545.830 ;
        RECT 1293.125 1545.815 1293.455 1545.830 ;
        RECT 1359.825 1470.650 1360.155 1470.665 ;
        RECT 1359.150 1470.350 1360.155 1470.650 ;
        RECT 1359.150 1469.985 1359.450 1470.350 ;
        RECT 1359.825 1470.335 1360.155 1470.350 ;
        RECT 1358.905 1469.670 1359.450 1469.985 ;
        RECT 1358.905 1469.655 1359.235 1469.670 ;
        RECT 1359.825 1374.090 1360.155 1374.105 ;
        RECT 1359.150 1373.790 1360.155 1374.090 ;
        RECT 1359.150 1373.425 1359.450 1373.790 ;
        RECT 1359.825 1373.775 1360.155 1373.790 ;
        RECT 1358.905 1373.110 1359.450 1373.425 ;
        RECT 1358.905 1373.095 1359.235 1373.110 ;
        RECT 1405.825 1304.060 1406.155 1304.065 ;
        RECT 1405.825 1304.050 1406.410 1304.060 ;
        RECT 1405.600 1303.750 1406.410 1304.050 ;
        RECT 1405.825 1303.740 1406.410 1303.750 ;
        RECT 1405.825 1303.735 1406.155 1303.740 ;
        RECT 1357.985 1276.850 1358.315 1276.865 ;
        RECT 1358.905 1276.850 1359.235 1276.865 ;
        RECT 1357.985 1276.550 1359.235 1276.850 ;
        RECT 1357.985 1276.535 1358.315 1276.550 ;
        RECT 1358.905 1276.535 1359.235 1276.550 ;
        RECT 1544.285 1257.130 1544.615 1257.145 ;
        RECT 1544.285 1256.830 1545.290 1257.130 ;
        RECT 1544.285 1256.815 1544.615 1256.830 ;
        RECT 1406.030 1256.140 1406.410 1256.460 ;
        RECT 1544.285 1256.450 1544.615 1256.465 ;
        RECT 1544.990 1256.450 1545.290 1256.830 ;
        RECT 1544.285 1256.150 1545.290 1256.450 ;
        RECT 1405.365 1255.770 1405.695 1255.785 ;
        RECT 1406.070 1255.770 1406.370 1256.140 ;
        RECT 1544.285 1256.135 1544.615 1256.150 ;
        RECT 1405.365 1255.470 1406.370 1255.770 ;
        RECT 1405.365 1255.455 1405.695 1255.470 ;
        RECT 1289.905 1207.490 1290.235 1207.505 ;
        RECT 1290.825 1207.490 1291.155 1207.505 ;
        RECT 1289.905 1207.190 1291.155 1207.490 ;
        RECT 1289.905 1207.175 1290.235 1207.190 ;
        RECT 1290.825 1207.175 1291.155 1207.190 ;
        RECT 986.305 1014.370 986.635 1014.385 ;
        RECT 1101.765 1014.370 1102.095 1014.385 ;
        RECT 986.305 1014.070 1102.095 1014.370 ;
        RECT 986.305 1014.055 986.635 1014.070 ;
        RECT 1101.765 1014.055 1102.095 1014.070 ;
        RECT 978.485 1013.690 978.815 1013.705 ;
        RECT 1119.245 1013.690 1119.575 1013.705 ;
        RECT 978.485 1013.390 1119.575 1013.690 ;
        RECT 978.485 1013.375 978.815 1013.390 ;
        RECT 1119.245 1013.375 1119.575 1013.390 ;
        RECT 978.945 1013.010 979.275 1013.025 ;
        RECT 1131.665 1013.010 1131.995 1013.025 ;
        RECT 978.945 1012.710 1131.995 1013.010 ;
        RECT 978.945 1012.695 979.275 1012.710 ;
        RECT 1131.665 1012.695 1131.995 1012.710 ;
        RECT 1511.165 1013.010 1511.495 1013.025 ;
        RECT 1536.005 1013.010 1536.335 1013.025 ;
        RECT 1511.165 1012.710 1536.335 1013.010 ;
        RECT 1511.165 1012.695 1511.495 1012.710 ;
        RECT 1536.005 1012.695 1536.335 1012.710 ;
        RECT 985.845 1012.330 986.175 1012.345 ;
        RECT 1143.165 1012.330 1143.495 1012.345 ;
        RECT 985.845 1012.030 1143.495 1012.330 ;
        RECT 985.845 1012.015 986.175 1012.030 ;
        RECT 1143.165 1012.015 1143.495 1012.030 ;
        RECT 1263.225 1012.330 1263.555 1012.345 ;
        RECT 1270.585 1012.330 1270.915 1012.345 ;
        RECT 1263.225 1012.030 1270.915 1012.330 ;
        RECT 1263.225 1012.015 1263.555 1012.030 ;
        RECT 1270.585 1012.015 1270.915 1012.030 ;
        RECT 985.385 1011.650 985.715 1011.665 ;
        RECT 1167.085 1011.650 1167.415 1011.665 ;
        RECT 985.385 1011.350 1167.415 1011.650 ;
        RECT 985.385 1011.335 985.715 1011.350 ;
        RECT 1167.085 1011.335 1167.415 1011.350 ;
        RECT 1267.365 1011.650 1267.695 1011.665 ;
        RECT 1269.665 1011.650 1269.995 1011.665 ;
        RECT 1267.365 1011.350 1269.995 1011.650 ;
        RECT 1267.365 1011.335 1267.695 1011.350 ;
        RECT 1269.665 1011.335 1269.995 1011.350 ;
        RECT 1292.665 1011.650 1292.995 1011.665 ;
        RECT 1297.265 1011.650 1297.595 1011.665 ;
        RECT 1292.665 1011.350 1297.595 1011.650 ;
        RECT 1292.665 1011.335 1292.995 1011.350 ;
        RECT 1297.265 1011.335 1297.595 1011.350 ;
        RECT 995.045 1010.970 995.375 1010.985 ;
        RECT 1309.685 1010.970 1310.015 1010.985 ;
        RECT 995.045 1010.670 1310.015 1010.970 ;
        RECT 995.045 1010.655 995.375 1010.670 ;
        RECT 1309.685 1010.655 1310.015 1010.670 ;
        RECT 1386.505 1010.970 1386.835 1010.985 ;
        RECT 1892.045 1010.970 1892.375 1010.985 ;
        RECT 1386.505 1010.670 1892.375 1010.970 ;
        RECT 1386.505 1010.655 1386.835 1010.670 ;
        RECT 1892.045 1010.655 1892.375 1010.670 ;
        RECT 993.205 1010.290 993.535 1010.305 ;
        RECT 1067.265 1010.290 1067.595 1010.305 ;
        RECT 993.205 1009.990 1067.595 1010.290 ;
        RECT 993.205 1009.975 993.535 1009.990 ;
        RECT 1067.265 1009.975 1067.595 1009.990 ;
        RECT 1521.285 1010.290 1521.615 1010.305 ;
        RECT 1536.465 1010.290 1536.795 1010.305 ;
        RECT 1521.285 1009.990 1536.795 1010.290 ;
        RECT 1521.285 1009.975 1521.615 1009.990 ;
        RECT 1536.465 1009.975 1536.795 1009.990 ;
      LAYER met3 ;
        RECT 674.400 996.080 2166.000 996.945 ;
        RECT 674.000 994.760 2166.000 996.080 ;
        RECT 674.000 993.360 2165.600 994.760 ;
        RECT 674.000 992.040 2166.000 993.360 ;
        RECT 674.400 990.640 2166.000 992.040 ;
        RECT 674.000 986.600 2166.000 990.640 ;
        RECT 674.400 985.200 2166.000 986.600 ;
        RECT 674.000 984.560 2166.000 985.200 ;
        RECT 674.000 983.160 2165.600 984.560 ;
        RECT 674.000 981.840 2166.000 983.160 ;
        RECT 674.400 980.440 2166.000 981.840 ;
        RECT 674.000 976.400 2166.000 980.440 ;
        RECT 674.400 975.000 2166.000 976.400 ;
        RECT 674.000 973.680 2166.000 975.000 ;
        RECT 674.000 972.280 2165.600 973.680 ;
        RECT 674.000 970.960 2166.000 972.280 ;
        RECT 674.400 969.560 2166.000 970.960 ;
        RECT 674.000 965.520 2166.000 969.560 ;
        RECT 674.400 964.120 2166.000 965.520 ;
        RECT 674.000 963.480 2166.000 964.120 ;
        RECT 674.000 962.080 2165.600 963.480 ;
        RECT 674.000 960.760 2166.000 962.080 ;
        RECT 674.400 959.360 2166.000 960.760 ;
        RECT 674.000 955.320 2166.000 959.360 ;
        RECT 674.400 953.920 2166.000 955.320 ;
        RECT 674.000 952.600 2166.000 953.920 ;
        RECT 674.000 951.200 2165.600 952.600 ;
        RECT 674.000 949.880 2166.000 951.200 ;
        RECT 674.400 948.480 2166.000 949.880 ;
        RECT 674.000 944.440 2166.000 948.480 ;
        RECT 674.400 943.040 2166.000 944.440 ;
        RECT 674.000 942.400 2166.000 943.040 ;
        RECT 674.000 941.000 2165.600 942.400 ;
        RECT 674.000 939.680 2166.000 941.000 ;
        RECT 674.400 938.280 2166.000 939.680 ;
        RECT 674.000 934.240 2166.000 938.280 ;
        RECT 674.400 932.840 2166.000 934.240 ;
        RECT 674.000 931.520 2166.000 932.840 ;
        RECT 674.000 930.120 2165.600 931.520 ;
        RECT 674.000 928.800 2166.000 930.120 ;
        RECT 674.400 927.400 2166.000 928.800 ;
        RECT 674.000 923.360 2166.000 927.400 ;
        RECT 674.400 921.960 2166.000 923.360 ;
        RECT 674.000 921.320 2166.000 921.960 ;
        RECT 674.000 919.920 2165.600 921.320 ;
        RECT 674.000 918.600 2166.000 919.920 ;
        RECT 674.400 917.200 2166.000 918.600 ;
        RECT 674.000 913.160 2166.000 917.200 ;
        RECT 674.400 911.760 2166.000 913.160 ;
        RECT 674.000 910.440 2166.000 911.760 ;
        RECT 674.000 909.040 2165.600 910.440 ;
        RECT 674.000 907.720 2166.000 909.040 ;
        RECT 674.400 906.320 2166.000 907.720 ;
        RECT 674.000 902.960 2166.000 906.320 ;
        RECT 674.400 901.560 2166.000 902.960 ;
        RECT 674.000 900.240 2166.000 901.560 ;
        RECT 674.000 898.840 2165.600 900.240 ;
        RECT 674.000 897.520 2166.000 898.840 ;
        RECT 674.400 896.120 2166.000 897.520 ;
        RECT 674.000 892.080 2166.000 896.120 ;
        RECT 674.400 890.680 2166.000 892.080 ;
        RECT 674.000 889.360 2166.000 890.680 ;
        RECT 674.000 887.960 2165.600 889.360 ;
        RECT 674.000 886.640 2166.000 887.960 ;
        RECT 674.400 885.240 2166.000 886.640 ;
        RECT 674.000 881.880 2166.000 885.240 ;
        RECT 674.400 880.480 2166.000 881.880 ;
        RECT 674.000 879.160 2166.000 880.480 ;
        RECT 674.000 877.760 2165.600 879.160 ;
        RECT 674.000 876.440 2166.000 877.760 ;
        RECT 674.400 875.040 2166.000 876.440 ;
        RECT 674.000 871.000 2166.000 875.040 ;
        RECT 674.400 869.600 2166.000 871.000 ;
        RECT 674.000 868.280 2166.000 869.600 ;
        RECT 674.000 866.880 2165.600 868.280 ;
        RECT 674.000 865.560 2166.000 866.880 ;
        RECT 674.400 864.160 2166.000 865.560 ;
        RECT 674.000 860.800 2166.000 864.160 ;
        RECT 674.400 859.400 2166.000 860.800 ;
        RECT 674.000 858.080 2166.000 859.400 ;
        RECT 674.000 856.680 2165.600 858.080 ;
        RECT 674.000 855.360 2166.000 856.680 ;
        RECT 674.400 853.960 2166.000 855.360 ;
        RECT 674.000 849.920 2166.000 853.960 ;
        RECT 674.400 848.520 2166.000 849.920 ;
        RECT 674.000 847.200 2166.000 848.520 ;
        RECT 674.000 845.800 2165.600 847.200 ;
        RECT 674.000 844.480 2166.000 845.800 ;
        RECT 674.400 843.080 2166.000 844.480 ;
        RECT 674.000 839.720 2166.000 843.080 ;
        RECT 674.400 838.320 2166.000 839.720 ;
        RECT 674.000 837.000 2166.000 838.320 ;
        RECT 674.000 835.600 2165.600 837.000 ;
        RECT 674.000 834.280 2166.000 835.600 ;
        RECT 674.400 832.880 2166.000 834.280 ;
        RECT 674.000 828.840 2166.000 832.880 ;
        RECT 674.400 827.440 2166.000 828.840 ;
        RECT 674.000 826.120 2166.000 827.440 ;
        RECT 674.000 824.720 2165.600 826.120 ;
        RECT 674.000 823.400 2166.000 824.720 ;
        RECT 674.400 822.000 2166.000 823.400 ;
        RECT 674.000 818.640 2166.000 822.000 ;
        RECT 674.400 817.240 2166.000 818.640 ;
        RECT 674.000 815.920 2166.000 817.240 ;
        RECT 674.000 814.520 2165.600 815.920 ;
        RECT 674.000 813.200 2166.000 814.520 ;
        RECT 674.400 811.800 2166.000 813.200 ;
        RECT 674.000 807.760 2166.000 811.800 ;
        RECT 674.400 806.360 2166.000 807.760 ;
        RECT 674.000 805.720 2166.000 806.360 ;
        RECT 674.000 804.320 2165.600 805.720 ;
        RECT 674.000 803.000 2166.000 804.320 ;
        RECT 674.400 801.600 2166.000 803.000 ;
        RECT 674.000 797.560 2166.000 801.600 ;
        RECT 674.400 796.160 2166.000 797.560 ;
        RECT 674.000 794.840 2166.000 796.160 ;
        RECT 674.000 793.440 2165.600 794.840 ;
        RECT 674.000 792.120 2166.000 793.440 ;
        RECT 674.400 790.720 2166.000 792.120 ;
        RECT 674.000 786.680 2166.000 790.720 ;
        RECT 674.400 785.280 2166.000 786.680 ;
        RECT 674.000 784.640 2166.000 785.280 ;
        RECT 674.000 783.240 2165.600 784.640 ;
        RECT 674.000 781.920 2166.000 783.240 ;
        RECT 674.400 780.520 2166.000 781.920 ;
        RECT 674.000 776.480 2166.000 780.520 ;
        RECT 674.400 775.080 2166.000 776.480 ;
        RECT 674.000 773.760 2166.000 775.080 ;
        RECT 674.000 772.360 2165.600 773.760 ;
        RECT 674.000 771.040 2166.000 772.360 ;
        RECT 674.400 769.640 2166.000 771.040 ;
        RECT 674.000 765.600 2166.000 769.640 ;
        RECT 674.400 764.200 2166.000 765.600 ;
        RECT 674.000 763.560 2166.000 764.200 ;
        RECT 674.000 762.160 2165.600 763.560 ;
        RECT 674.000 760.840 2166.000 762.160 ;
        RECT 674.400 759.440 2166.000 760.840 ;
        RECT 674.000 755.400 2166.000 759.440 ;
        RECT 674.400 754.000 2166.000 755.400 ;
        RECT 674.000 752.680 2166.000 754.000 ;
        RECT 674.000 751.280 2165.600 752.680 ;
        RECT 674.000 749.960 2166.000 751.280 ;
        RECT 674.400 748.560 2166.000 749.960 ;
        RECT 674.000 744.520 2166.000 748.560 ;
        RECT 674.400 743.120 2166.000 744.520 ;
        RECT 674.000 742.480 2166.000 743.120 ;
        RECT 674.000 741.080 2165.600 742.480 ;
        RECT 674.000 739.760 2166.000 741.080 ;
        RECT 674.400 738.360 2166.000 739.760 ;
        RECT 674.000 734.320 2166.000 738.360 ;
        RECT 674.400 732.920 2166.000 734.320 ;
        RECT 674.000 731.600 2166.000 732.920 ;
        RECT 674.000 730.200 2165.600 731.600 ;
        RECT 674.000 728.880 2166.000 730.200 ;
        RECT 674.400 727.480 2166.000 728.880 ;
        RECT 674.000 723.440 2166.000 727.480 ;
        RECT 674.400 722.040 2166.000 723.440 ;
        RECT 674.000 721.400 2166.000 722.040 ;
        RECT 674.000 720.000 2165.600 721.400 ;
        RECT 674.000 718.680 2166.000 720.000 ;
        RECT 674.400 717.280 2166.000 718.680 ;
        RECT 674.000 713.240 2166.000 717.280 ;
        RECT 674.400 711.840 2166.000 713.240 ;
        RECT 674.000 710.520 2166.000 711.840 ;
        RECT 674.000 709.120 2165.600 710.520 ;
        RECT 674.000 707.800 2166.000 709.120 ;
        RECT 674.400 706.400 2166.000 707.800 ;
        RECT 674.000 703.040 2166.000 706.400 ;
        RECT 674.400 701.640 2166.000 703.040 ;
        RECT 674.000 700.320 2166.000 701.640 ;
        RECT 674.000 698.920 2165.600 700.320 ;
        RECT 674.000 697.600 2166.000 698.920 ;
        RECT 674.400 696.200 2166.000 697.600 ;
        RECT 674.000 692.160 2166.000 696.200 ;
        RECT 674.400 690.760 2166.000 692.160 ;
        RECT 674.000 689.440 2166.000 690.760 ;
        RECT 674.000 688.040 2165.600 689.440 ;
        RECT 674.000 686.720 2166.000 688.040 ;
        RECT 674.400 685.320 2166.000 686.720 ;
        RECT 674.000 681.960 2166.000 685.320 ;
        RECT 674.400 680.560 2166.000 681.960 ;
        RECT 674.000 679.240 2166.000 680.560 ;
        RECT 674.000 677.840 2165.600 679.240 ;
        RECT 674.000 676.520 2166.000 677.840 ;
        RECT 674.400 675.120 2166.000 676.520 ;
        RECT 674.000 671.080 2166.000 675.120 ;
        RECT 674.400 669.680 2166.000 671.080 ;
        RECT 674.000 668.360 2166.000 669.680 ;
        RECT 674.000 666.960 2165.600 668.360 ;
        RECT 674.000 665.640 2166.000 666.960 ;
        RECT 674.400 664.240 2166.000 665.640 ;
        RECT 674.000 660.880 2166.000 664.240 ;
        RECT 674.400 659.480 2166.000 660.880 ;
        RECT 674.000 658.160 2166.000 659.480 ;
        RECT 674.000 656.760 2165.600 658.160 ;
        RECT 674.000 655.440 2166.000 656.760 ;
        RECT 674.400 654.040 2166.000 655.440 ;
        RECT 674.000 650.000 2166.000 654.040 ;
        RECT 674.400 648.600 2166.000 650.000 ;
        RECT 674.000 647.280 2166.000 648.600 ;
        RECT 674.000 645.880 2165.600 647.280 ;
        RECT 674.000 644.560 2166.000 645.880 ;
        RECT 674.400 643.160 2166.000 644.560 ;
        RECT 674.000 639.800 2166.000 643.160 ;
        RECT 674.400 638.400 2166.000 639.800 ;
        RECT 674.000 637.080 2166.000 638.400 ;
        RECT 674.000 635.680 2165.600 637.080 ;
        RECT 674.000 634.360 2166.000 635.680 ;
        RECT 674.400 632.960 2166.000 634.360 ;
        RECT 674.000 628.920 2166.000 632.960 ;
        RECT 674.400 627.520 2166.000 628.920 ;
        RECT 674.000 626.200 2166.000 627.520 ;
        RECT 674.000 624.800 2165.600 626.200 ;
        RECT 674.000 623.480 2166.000 624.800 ;
        RECT 674.400 622.080 2166.000 623.480 ;
        RECT 674.000 618.720 2166.000 622.080 ;
        RECT 674.400 617.320 2166.000 618.720 ;
        RECT 674.000 616.000 2166.000 617.320 ;
        RECT 674.000 614.600 2165.600 616.000 ;
        RECT 674.000 613.280 2166.000 614.600 ;
        RECT 674.400 611.880 2166.000 613.280 ;
        RECT 674.000 607.840 2166.000 611.880 ;
        RECT 674.400 606.440 2166.000 607.840 ;
        RECT 674.000 605.800 2166.000 606.440 ;
        RECT 674.000 604.400 2165.600 605.800 ;
        RECT 674.000 603.080 2166.000 604.400 ;
        RECT 674.400 602.215 2166.000 603.080 ;
      LAYER via3 ;
        RECT 1358.220 2511.420 1358.540 2511.740 ;
        RECT 1358.220 2463.140 1358.540 2463.460 ;
        RECT 1406.060 1303.740 1406.380 1304.060 ;
        RECT 1406.060 1256.140 1406.380 1256.460 ;
      LAYER met4 ;
        RECT 459.645 2610.640 480.165 2747.120 ;
        RECT 482.565 2610.640 550.935 2747.120 ;
        RECT 1036.375 2610.640 1080.450 2787.920 ;
      LAYER met4 ;
        RECT 1358.215 2511.415 1358.545 2511.745 ;
        RECT 1358.230 2463.465 1358.530 2511.415 ;
      LAYER met4 ;
        RECT 1674.640 2510.640 1829.840 2889.200 ;
        RECT 2477.790 2610.640 2529.990 2760.720 ;
      LAYER met4 ;
        RECT 1358.215 2463.135 1358.545 2463.465 ;
      LAYER met4 ;
        RECT 531.415 1710.640 613.040 1969.520 ;
        RECT 1174.640 1710.640 1253.040 2032.080 ;
        RECT 1997.170 1760.640 2047.070 1905.280 ;
        RECT 2474.640 1710.640 2476.240 1926.000 ;
      LAYER met4 ;
        RECT 1406.055 1303.735 1406.385 1304.065 ;
        RECT 1406.070 1256.465 1406.370 1303.735 ;
        RECT 1406.055 1256.135 1406.385 1256.465 ;
      LAYER met4 ;
        RECT 718.135 989.600 2151.840 995.585 ;
        RECT 718.135 610.640 767.440 989.600 ;
        RECT 769.840 610.640 2151.840 989.600 ;
      LAYER met5 ;
        RECT 855.500 966.380 1861.740 983.300 ;
        RECT 855.500 948.380 1861.740 963.380 ;
        RECT 855.500 944.300 1861.740 945.380 ;
  END
END user_project_wrapper
END LIBRARY

